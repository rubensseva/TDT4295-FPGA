module DotProd(
  input        clock,
  input        reset,
  input  [7:0] io_dataInA,
  input  [7:0] io_dataInB,
  output [8:0] io_dataOut,
  output       io_outputValid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] countVal; // @[Counter.scala 29:33]
  wire  countReset = countVal == 4'h8; // @[Counter.scala 38:24]
  wire [3:0] _T_2 = countVal + 4'h1; // @[Counter.scala 39:22]
  reg [8:0] accumulator; // @[DotProd.scala 19:28]
  wire [15:0] product = $signed(io_dataInA) * $signed(io_dataInB); // @[DotProd.scala 20:35]
  wire [15:0] _GEN_5 = {{7{accumulator[8]}},accumulator}; // @[DotProd.scala 21:30]
  wire [15:0] _T_6 = $signed(_GEN_5) + $signed(product); // @[DotProd.scala 21:30]
  wire [15:0] _GEN_4 = countReset ? $signed(16'sh0) : $signed(_T_6); // @[DotProd.scala 25:20]
  assign io_dataOut = _T_6[8:0]; // @[DotProd.scala 23:14]
  assign io_outputValid = countVal == 4'h8; // @[DotProd.scala 26:20 DotProd.scala 29:20]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  countVal = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  accumulator = _RAND_1[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      countVal <= 4'h0;
    end else if (countReset) begin
      countVal <= 4'h0;
    end else begin
      countVal <= _T_2;
    end
    if (reset) begin
      accumulator <= 9'sh0;
    end else begin
      accumulator <= _GEN_4[8:0];
    end
  end
endmodule
module KernelConvolution(
  input        clock,
  input        reset,
  input  [4:0] io_kernelVal_in,
  input  [3:0] io_pixelVal_in_0,
  input  [3:0] io_pixelVal_in_1,
  input  [3:0] io_pixelVal_in_2,
  input  [3:0] io_pixelVal_in_3,
  input  [3:0] io_pixelVal_in_4,
  input  [3:0] io_pixelVal_in_5,
  input  [3:0] io_pixelVal_in_6,
  input  [3:0] io_pixelVal_in_7,
  output [8:0] io_pixelVal_out_0,
  output [8:0] io_pixelVal_out_1,
  output [8:0] io_pixelVal_out_2,
  output [8:0] io_pixelVal_out_3,
  output [8:0] io_pixelVal_out_4,
  output [8:0] io_pixelVal_out_5,
  output [8:0] io_pixelVal_out_6,
  output [8:0] io_pixelVal_out_7,
  output       io_valid_out
);
  wire  DotProd_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_1_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_1_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_1_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_1_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_1_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_1_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_2_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_2_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_2_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_2_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_2_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_2_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_3_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_3_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_3_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_3_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_3_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_3_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_4_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_4_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_4_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_4_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_4_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_4_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_5_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_5_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_5_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_5_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_5_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_5_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_6_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_6_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_6_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_6_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_6_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_6_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_7_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_7_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_7_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_7_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_7_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_7_io_outputValid; // @[KernelConvolution.scala 21:58]
  DotProd DotProd ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_clock),
    .reset(DotProd_reset),
    .io_dataInA(DotProd_io_dataInA),
    .io_dataInB(DotProd_io_dataInB),
    .io_dataOut(DotProd_io_dataOut),
    .io_outputValid(DotProd_io_outputValid)
  );
  DotProd DotProd_1 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_1_clock),
    .reset(DotProd_1_reset),
    .io_dataInA(DotProd_1_io_dataInA),
    .io_dataInB(DotProd_1_io_dataInB),
    .io_dataOut(DotProd_1_io_dataOut),
    .io_outputValid(DotProd_1_io_outputValid)
  );
  DotProd DotProd_2 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_2_clock),
    .reset(DotProd_2_reset),
    .io_dataInA(DotProd_2_io_dataInA),
    .io_dataInB(DotProd_2_io_dataInB),
    .io_dataOut(DotProd_2_io_dataOut),
    .io_outputValid(DotProd_2_io_outputValid)
  );
  DotProd DotProd_3 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_3_clock),
    .reset(DotProd_3_reset),
    .io_dataInA(DotProd_3_io_dataInA),
    .io_dataInB(DotProd_3_io_dataInB),
    .io_dataOut(DotProd_3_io_dataOut),
    .io_outputValid(DotProd_3_io_outputValid)
  );
  DotProd DotProd_4 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_4_clock),
    .reset(DotProd_4_reset),
    .io_dataInA(DotProd_4_io_dataInA),
    .io_dataInB(DotProd_4_io_dataInB),
    .io_dataOut(DotProd_4_io_dataOut),
    .io_outputValid(DotProd_4_io_outputValid)
  );
  DotProd DotProd_5 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_5_clock),
    .reset(DotProd_5_reset),
    .io_dataInA(DotProd_5_io_dataInA),
    .io_dataInB(DotProd_5_io_dataInB),
    .io_dataOut(DotProd_5_io_dataOut),
    .io_outputValid(DotProd_5_io_outputValid)
  );
  DotProd DotProd_6 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_6_clock),
    .reset(DotProd_6_reset),
    .io_dataInA(DotProd_6_io_dataInA),
    .io_dataInB(DotProd_6_io_dataInB),
    .io_dataOut(DotProd_6_io_dataOut),
    .io_outputValid(DotProd_6_io_outputValid)
  );
  DotProd DotProd_7 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_7_clock),
    .reset(DotProd_7_reset),
    .io_dataInA(DotProd_7_io_dataInA),
    .io_dataInB(DotProd_7_io_dataInB),
    .io_dataOut(DotProd_7_io_dataOut),
    .io_outputValid(DotProd_7_io_outputValid)
  );
  assign io_pixelVal_out_0 = DotProd_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_1 = DotProd_1_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_2 = DotProd_2_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_3 = DotProd_3_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_4 = DotProd_4_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_5 = DotProd_5_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_6 = DotProd_6_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_7 = DotProd_7_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_valid_out = DotProd_io_outputValid; // @[KernelConvolution.scala 35:30]
  assign DotProd_clock = clock;
  assign DotProd_reset = reset;
  assign DotProd_io_dataInA = {{4'd0}, io_pixelVal_in_0}; // @[KernelConvolution.scala 21:32]
  assign DotProd_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_1_clock = clock;
  assign DotProd_1_reset = reset;
  assign DotProd_1_io_dataInA = {{4'd0}, io_pixelVal_in_1}; // @[KernelConvolution.scala 21:32]
  assign DotProd_1_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_2_clock = clock;
  assign DotProd_2_reset = reset;
  assign DotProd_2_io_dataInA = {{4'd0}, io_pixelVal_in_2}; // @[KernelConvolution.scala 21:32]
  assign DotProd_2_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_3_clock = clock;
  assign DotProd_3_reset = reset;
  assign DotProd_3_io_dataInA = {{4'd0}, io_pixelVal_in_3}; // @[KernelConvolution.scala 21:32]
  assign DotProd_3_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_4_clock = clock;
  assign DotProd_4_reset = reset;
  assign DotProd_4_io_dataInA = {{4'd0}, io_pixelVal_in_4}; // @[KernelConvolution.scala 21:32]
  assign DotProd_4_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_5_clock = clock;
  assign DotProd_5_reset = reset;
  assign DotProd_5_io_dataInA = {{4'd0}, io_pixelVal_in_5}; // @[KernelConvolution.scala 21:32]
  assign DotProd_5_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_6_clock = clock;
  assign DotProd_6_reset = reset;
  assign DotProd_6_io_dataInA = {{4'd0}, io_pixelVal_in_6}; // @[KernelConvolution.scala 21:32]
  assign DotProd_6_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_7_clock = clock;
  assign DotProd_7_reset = reset;
  assign DotProd_7_io_dataInA = {{4'd0}, io_pixelVal_in_7}; // @[KernelConvolution.scala 21:32]
  assign DotProd_7_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
endmodule
module Filter(
  input        clock,
  input        reset,
  input  [5:0] io_SPI_filterIndex,
  input        io_SPI_distort,
  output [3:0] io_pixelVal_out_0_0,
  output [3:0] io_pixelVal_out_0_1,
  output [3:0] io_pixelVal_out_0_2,
  output [3:0] io_pixelVal_out_0_3,
  output [3:0] io_pixelVal_out_0_4,
  output [3:0] io_pixelVal_out_0_5,
  output [3:0] io_pixelVal_out_0_6,
  output [3:0] io_pixelVal_out_0_7,
  output [3:0] io_pixelVal_out_1_0,
  output [3:0] io_pixelVal_out_1_1,
  output [3:0] io_pixelVal_out_1_2,
  output [3:0] io_pixelVal_out_1_3,
  output [3:0] io_pixelVal_out_1_4,
  output [3:0] io_pixelVal_out_1_5,
  output [3:0] io_pixelVal_out_1_6,
  output [3:0] io_pixelVal_out_1_7,
  output [3:0] io_pixelVal_out_2_0,
  output [3:0] io_pixelVal_out_2_1,
  output [3:0] io_pixelVal_out_2_2,
  output [3:0] io_pixelVal_out_2_3,
  output [3:0] io_pixelVal_out_2_4,
  output [3:0] io_pixelVal_out_2_5,
  output [3:0] io_pixelVal_out_2_6,
  output [3:0] io_pixelVal_out_2_7,
  output       io_valid_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
`endif // RANDOMIZE_REG_INIT
  wire  KernelConvolution_clock; // @[Filter.scala 178:36]
  wire  KernelConvolution_reset; // @[Filter.scala 178:36]
  wire [4:0] KernelConvolution_io_kernelVal_in; // @[Filter.scala 178:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_0; // @[Filter.scala 178:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_1; // @[Filter.scala 178:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_2; // @[Filter.scala 178:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_3; // @[Filter.scala 178:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_4; // @[Filter.scala 178:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_5; // @[Filter.scala 178:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_6; // @[Filter.scala 178:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_7; // @[Filter.scala 178:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_0; // @[Filter.scala 178:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_1; // @[Filter.scala 178:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_2; // @[Filter.scala 178:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_3; // @[Filter.scala 178:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_4; // @[Filter.scala 178:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_5; // @[Filter.scala 178:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_6; // @[Filter.scala 178:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_7; // @[Filter.scala 178:36]
  wire  KernelConvolution_io_valid_out; // @[Filter.scala 178:36]
  wire  KernelConvolution_1_clock; // @[Filter.scala 179:36]
  wire  KernelConvolution_1_reset; // @[Filter.scala 179:36]
  wire [4:0] KernelConvolution_1_io_kernelVal_in; // @[Filter.scala 179:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_0; // @[Filter.scala 179:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_1; // @[Filter.scala 179:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_2; // @[Filter.scala 179:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_3; // @[Filter.scala 179:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_4; // @[Filter.scala 179:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_5; // @[Filter.scala 179:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_6; // @[Filter.scala 179:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_7; // @[Filter.scala 179:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_0; // @[Filter.scala 179:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_1; // @[Filter.scala 179:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_2; // @[Filter.scala 179:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_3; // @[Filter.scala 179:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_4; // @[Filter.scala 179:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_5; // @[Filter.scala 179:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_6; // @[Filter.scala 179:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_7; // @[Filter.scala 179:36]
  wire  KernelConvolution_1_io_valid_out; // @[Filter.scala 179:36]
  wire  KernelConvolution_2_clock; // @[Filter.scala 180:36]
  wire  KernelConvolution_2_reset; // @[Filter.scala 180:36]
  wire [4:0] KernelConvolution_2_io_kernelVal_in; // @[Filter.scala 180:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_0; // @[Filter.scala 180:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_1; // @[Filter.scala 180:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_2; // @[Filter.scala 180:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_3; // @[Filter.scala 180:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_4; // @[Filter.scala 180:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_5; // @[Filter.scala 180:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_6; // @[Filter.scala 180:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_7; // @[Filter.scala 180:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_0; // @[Filter.scala 180:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_1; // @[Filter.scala 180:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_2; // @[Filter.scala 180:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_3; // @[Filter.scala 180:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_4; // @[Filter.scala 180:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_5; // @[Filter.scala 180:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_6; // @[Filter.scala 180:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_7; // @[Filter.scala 180:36]
  wire  KernelConvolution_2_io_valid_out; // @[Filter.scala 180:36]
  reg [3:0] kernelCounter; // @[Counter.scala 29:33]
  wire  kernelCountReset = kernelCounter == 4'h8; // @[Counter.scala 38:24]
  wire [3:0] _T_14 = kernelCounter + 4'h1; // @[Counter.scala 39:22]
  wire  _GEN_7259 = 3'h0 == io_SPI_filterIndex[2:0]; // @[Filter.scala 186:41]
  wire  _GEN_7260 = 4'h4 == kernelCounter; // @[Filter.scala 186:41]
  wire [4:0] _GEN_7 = _GEN_7259 & _GEN_7260 ? $signed(5'sh1) : $signed(5'sh0); // @[Filter.scala 186:41]
  wire  _GEN_7262 = 4'h5 == kernelCounter; // @[Filter.scala 186:41]
  wire [4:0] _GEN_8 = _GEN_7259 & _GEN_7262 ? $signed(5'sh0) : $signed(_GEN_7); // @[Filter.scala 186:41]
  wire  _GEN_7264 = 4'h6 == kernelCounter; // @[Filter.scala 186:41]
  wire [4:0] _GEN_9 = _GEN_7259 & _GEN_7264 ? $signed(5'sh0) : $signed(_GEN_8); // @[Filter.scala 186:41]
  wire  _GEN_7266 = 4'h7 == kernelCounter; // @[Filter.scala 186:41]
  wire [4:0] _GEN_10 = _GEN_7259 & _GEN_7266 ? $signed(5'sh0) : $signed(_GEN_9); // @[Filter.scala 186:41]
  wire  _GEN_7268 = 4'h8 == kernelCounter; // @[Filter.scala 186:41]
  wire [4:0] _GEN_11 = _GEN_7259 & _GEN_7268 ? $signed(5'sh0) : $signed(_GEN_10); // @[Filter.scala 186:41]
  wire  _GEN_7269 = 3'h1 == io_SPI_filterIndex[2:0]; // @[Filter.scala 186:41]
  wire  _GEN_7270 = 4'h0 == kernelCounter; // @[Filter.scala 186:41]
  wire [4:0] _GEN_12 = _GEN_7269 & _GEN_7270 ? $signed(5'sh1) : $signed(_GEN_11); // @[Filter.scala 186:41]
  wire  _GEN_7272 = 4'h1 == kernelCounter; // @[Filter.scala 186:41]
  wire [4:0] _GEN_13 = _GEN_7269 & _GEN_7272 ? $signed(5'sh1) : $signed(_GEN_12); // @[Filter.scala 186:41]
  wire  _GEN_7274 = 4'h2 == kernelCounter; // @[Filter.scala 186:41]
  wire [4:0] _GEN_14 = _GEN_7269 & _GEN_7274 ? $signed(5'sh1) : $signed(_GEN_13); // @[Filter.scala 186:41]
  wire  _GEN_7276 = 4'h3 == kernelCounter; // @[Filter.scala 186:41]
  wire [4:0] _GEN_15 = _GEN_7269 & _GEN_7276 ? $signed(5'sh1) : $signed(_GEN_14); // @[Filter.scala 186:41]
  wire [4:0] _GEN_16 = _GEN_7269 & _GEN_7260 ? $signed(5'sh1) : $signed(_GEN_15); // @[Filter.scala 186:41]
  wire [4:0] _GEN_17 = _GEN_7269 & _GEN_7262 ? $signed(5'sh1) : $signed(_GEN_16); // @[Filter.scala 186:41]
  wire [4:0] _GEN_18 = _GEN_7269 & _GEN_7264 ? $signed(5'sh1) : $signed(_GEN_17); // @[Filter.scala 186:41]
  wire [4:0] _GEN_19 = _GEN_7269 & _GEN_7266 ? $signed(5'sh1) : $signed(_GEN_18); // @[Filter.scala 186:41]
  wire [4:0] _GEN_20 = _GEN_7269 & _GEN_7268 ? $signed(5'sh1) : $signed(_GEN_19); // @[Filter.scala 186:41]
  wire  _GEN_7287 = 3'h2 == io_SPI_filterIndex[2:0]; // @[Filter.scala 186:41]
  wire [4:0] _GEN_21 = _GEN_7287 & _GEN_7270 ? $signed(5'sh1) : $signed(_GEN_20); // @[Filter.scala 186:41]
  wire [4:0] _GEN_22 = _GEN_7287 & _GEN_7272 ? $signed(5'sh2) : $signed(_GEN_21); // @[Filter.scala 186:41]
  wire [4:0] _GEN_23 = _GEN_7287 & _GEN_7274 ? $signed(5'sh1) : $signed(_GEN_22); // @[Filter.scala 186:41]
  wire [4:0] _GEN_24 = _GEN_7287 & _GEN_7276 ? $signed(5'sh2) : $signed(_GEN_23); // @[Filter.scala 186:41]
  wire [4:0] _GEN_25 = _GEN_7287 & _GEN_7260 ? $signed(5'sh4) : $signed(_GEN_24); // @[Filter.scala 186:41]
  wire [4:0] _GEN_26 = _GEN_7287 & _GEN_7262 ? $signed(5'sh2) : $signed(_GEN_25); // @[Filter.scala 186:41]
  wire [4:0] _GEN_27 = _GEN_7287 & _GEN_7264 ? $signed(5'sh1) : $signed(_GEN_26); // @[Filter.scala 186:41]
  wire [4:0] _GEN_28 = _GEN_7287 & _GEN_7266 ? $signed(5'sh2) : $signed(_GEN_27); // @[Filter.scala 186:41]
  wire [4:0] _GEN_29 = _GEN_7287 & _GEN_7268 ? $signed(5'sh1) : $signed(_GEN_28); // @[Filter.scala 186:41]
  wire  _GEN_7305 = 3'h3 == io_SPI_filterIndex[2:0]; // @[Filter.scala 186:41]
  wire [4:0] _GEN_30 = _GEN_7305 & _GEN_7270 ? $signed(5'sh0) : $signed(_GEN_29); // @[Filter.scala 186:41]
  wire [4:0] _GEN_31 = _GEN_7305 & _GEN_7272 ? $signed(-5'sh1) : $signed(_GEN_30); // @[Filter.scala 186:41]
  wire [4:0] _GEN_32 = _GEN_7305 & _GEN_7274 ? $signed(5'sh0) : $signed(_GEN_31); // @[Filter.scala 186:41]
  wire [4:0] _GEN_33 = _GEN_7305 & _GEN_7276 ? $signed(-5'sh1) : $signed(_GEN_32); // @[Filter.scala 186:41]
  wire [4:0] _GEN_34 = _GEN_7305 & _GEN_7260 ? $signed(5'sh4) : $signed(_GEN_33); // @[Filter.scala 186:41]
  wire [4:0] _GEN_35 = _GEN_7305 & _GEN_7262 ? $signed(-5'sh1) : $signed(_GEN_34); // @[Filter.scala 186:41]
  wire [4:0] _GEN_36 = _GEN_7305 & _GEN_7264 ? $signed(5'sh0) : $signed(_GEN_35); // @[Filter.scala 186:41]
  wire [4:0] _GEN_37 = _GEN_7305 & _GEN_7266 ? $signed(-5'sh1) : $signed(_GEN_36); // @[Filter.scala 186:41]
  wire [4:0] _GEN_38 = _GEN_7305 & _GEN_7268 ? $signed(5'sh0) : $signed(_GEN_37); // @[Filter.scala 186:41]
  wire  _GEN_7323 = 3'h4 == io_SPI_filterIndex[2:0]; // @[Filter.scala 186:41]
  wire [4:0] _GEN_39 = _GEN_7323 & _GEN_7270 ? $signed(-5'sh1) : $signed(_GEN_38); // @[Filter.scala 186:41]
  wire [4:0] _GEN_40 = _GEN_7323 & _GEN_7272 ? $signed(-5'sh1) : $signed(_GEN_39); // @[Filter.scala 186:41]
  wire [4:0] _GEN_41 = _GEN_7323 & _GEN_7274 ? $signed(-5'sh1) : $signed(_GEN_40); // @[Filter.scala 186:41]
  wire [4:0] _GEN_42 = _GEN_7323 & _GEN_7276 ? $signed(-5'sh1) : $signed(_GEN_41); // @[Filter.scala 186:41]
  wire [4:0] _GEN_43 = _GEN_7323 & _GEN_7260 ? $signed(5'sh8) : $signed(_GEN_42); // @[Filter.scala 186:41]
  wire [4:0] _GEN_44 = _GEN_7323 & _GEN_7262 ? $signed(-5'sh1) : $signed(_GEN_43); // @[Filter.scala 186:41]
  wire [4:0] _GEN_45 = _GEN_7323 & _GEN_7264 ? $signed(-5'sh1) : $signed(_GEN_44); // @[Filter.scala 186:41]
  wire [4:0] _GEN_46 = _GEN_7323 & _GEN_7266 ? $signed(-5'sh1) : $signed(_GEN_45); // @[Filter.scala 186:41]
  wire [4:0] _GEN_47 = _GEN_7323 & _GEN_7268 ? $signed(-5'sh1) : $signed(_GEN_46); // @[Filter.scala 186:41]
  wire  _GEN_7341 = 3'h5 == io_SPI_filterIndex[2:0]; // @[Filter.scala 186:41]
  wire [4:0] _GEN_48 = _GEN_7341 & _GEN_7270 ? $signed(5'sh0) : $signed(_GEN_47); // @[Filter.scala 186:41]
  wire [4:0] _GEN_49 = _GEN_7341 & _GEN_7272 ? $signed(-5'sh1) : $signed(_GEN_48); // @[Filter.scala 186:41]
  wire [4:0] _GEN_50 = _GEN_7341 & _GEN_7274 ? $signed(5'sh0) : $signed(_GEN_49); // @[Filter.scala 186:41]
  wire [4:0] _GEN_51 = _GEN_7341 & _GEN_7276 ? $signed(-5'sh1) : $signed(_GEN_50); // @[Filter.scala 186:41]
  wire [4:0] _GEN_52 = _GEN_7341 & _GEN_7260 ? $signed(5'sh5) : $signed(_GEN_51); // @[Filter.scala 186:41]
  wire [4:0] _GEN_53 = _GEN_7341 & _GEN_7262 ? $signed(-5'sh1) : $signed(_GEN_52); // @[Filter.scala 186:41]
  wire [4:0] _GEN_54 = _GEN_7341 & _GEN_7264 ? $signed(5'sh0) : $signed(_GEN_53); // @[Filter.scala 186:41]
  wire [4:0] _GEN_55 = _GEN_7341 & _GEN_7266 ? $signed(-5'sh1) : $signed(_GEN_54); // @[Filter.scala 186:41]
  reg [1:0] imageCounterX; // @[Counter.scala 29:33]
  wire  imageCounterXReset = imageCounterX == 2'h2; // @[Counter.scala 38:24]
  wire [1:0] _T_20 = imageCounterX + 2'h1; // @[Counter.scala 39:22]
  reg [1:0] imageCounterY; // @[Counter.scala 29:33]
  wire  _T_21 = imageCounterY == 2'h2; // @[Counter.scala 38:24]
  wire [1:0] _T_23 = imageCounterY + 2'h1; // @[Counter.scala 39:22]
  reg [31:0] pixelIndex; // @[Filter.scala 191:31]
  wire [32:0] _T_24 = {{1'd0}, pixelIndex}; // @[Filter.scala 194:31]
  wire [31:0] _GEN_0 = _T_24[31:0] % 32'h10; // @[Filter.scala 194:38]
  wire [4:0] _T_26 = _GEN_0[4:0]; // @[Filter.scala 194:38]
  wire [4:0] _GEN_7559 = {{3'd0}, imageCounterX}; // @[Filter.scala 194:53]
  wire [4:0] _T_28 = _T_26 + _GEN_7559; // @[Filter.scala 194:53]
  wire [4:0] _T_30 = _T_28 - 5'h1; // @[Filter.scala 194:69]
  wire [31:0] _T_33 = _T_24[31:0] / 32'h10; // @[Filter.scala 195:38]
  wire [31:0] _GEN_7560 = {{30'd0}, imageCounterY}; // @[Filter.scala 195:53]
  wire [31:0] _T_35 = _T_33 + _GEN_7560; // @[Filter.scala 195:53]
  wire [31:0] _T_37 = _T_35 - 32'h1; // @[Filter.scala 195:69]
  wire [36:0] _T_38 = _T_37 * 32'h10; // @[Filter.scala 196:42]
  wire [36:0] _GEN_7561 = {{32'd0}, _T_30}; // @[Filter.scala 196:57]
  wire [36:0] _T_40 = _T_38 + _GEN_7561; // @[Filter.scala 196:57]
  wire [3:0] _GEN_179 = 8'h8 == _T_40[7:0] ? 4'h0 : 4'hf; // @[Filter.scala 196:62]
  wire [3:0] _GEN_180 = 8'h9 == _T_40[7:0] ? 4'h0 : _GEN_179; // @[Filter.scala 196:62]
  wire [3:0] _GEN_181 = 8'ha == _T_40[7:0] ? 4'h0 : _GEN_180; // @[Filter.scala 196:62]
  wire [3:0] _GEN_182 = 8'hb == _T_40[7:0] ? 4'h0 : _GEN_181; // @[Filter.scala 196:62]
  wire [3:0] _GEN_183 = 8'hc == _T_40[7:0] ? 4'h0 : _GEN_182; // @[Filter.scala 196:62]
  wire [3:0] _GEN_184 = 8'hd == _T_40[7:0] ? 4'h0 : _GEN_183; // @[Filter.scala 196:62]
  wire [3:0] _GEN_185 = 8'he == _T_40[7:0] ? 4'h0 : _GEN_184; // @[Filter.scala 196:62]
  wire [3:0] _GEN_186 = 8'hf == _T_40[7:0] ? 4'h0 : _GEN_185; // @[Filter.scala 196:62]
  wire [3:0] _GEN_187 = 8'h10 == _T_40[7:0] ? 4'hf : _GEN_186; // @[Filter.scala 196:62]
  wire [3:0] _GEN_188 = 8'h11 == _T_40[7:0] ? 4'hf : _GEN_187; // @[Filter.scala 196:62]
  wire [3:0] _GEN_189 = 8'h12 == _T_40[7:0] ? 4'hf : _GEN_188; // @[Filter.scala 196:62]
  wire [3:0] _GEN_190 = 8'h13 == _T_40[7:0] ? 4'hf : _GEN_189; // @[Filter.scala 196:62]
  wire [3:0] _GEN_191 = 8'h14 == _T_40[7:0] ? 4'hf : _GEN_190; // @[Filter.scala 196:62]
  wire [3:0] _GEN_192 = 8'h15 == _T_40[7:0] ? 4'hf : _GEN_191; // @[Filter.scala 196:62]
  wire [3:0] _GEN_193 = 8'h16 == _T_40[7:0] ? 4'hf : _GEN_192; // @[Filter.scala 196:62]
  wire [3:0] _GEN_194 = 8'h17 == _T_40[7:0] ? 4'hf : _GEN_193; // @[Filter.scala 196:62]
  wire [3:0] _GEN_195 = 8'h18 == _T_40[7:0] ? 4'h0 : _GEN_194; // @[Filter.scala 196:62]
  wire [3:0] _GEN_196 = 8'h19 == _T_40[7:0] ? 4'h0 : _GEN_195; // @[Filter.scala 196:62]
  wire [3:0] _GEN_197 = 8'h1a == _T_40[7:0] ? 4'h0 : _GEN_196; // @[Filter.scala 196:62]
  wire [3:0] _GEN_198 = 8'h1b == _T_40[7:0] ? 4'h0 : _GEN_197; // @[Filter.scala 196:62]
  wire [3:0] _GEN_199 = 8'h1c == _T_40[7:0] ? 4'h0 : _GEN_198; // @[Filter.scala 196:62]
  wire [3:0] _GEN_200 = 8'h1d == _T_40[7:0] ? 4'h0 : _GEN_199; // @[Filter.scala 196:62]
  wire [3:0] _GEN_201 = 8'h1e == _T_40[7:0] ? 4'h0 : _GEN_200; // @[Filter.scala 196:62]
  wire [3:0] _GEN_202 = 8'h1f == _T_40[7:0] ? 4'h0 : _GEN_201; // @[Filter.scala 196:62]
  wire [3:0] _GEN_203 = 8'h20 == _T_40[7:0] ? 4'hf : _GEN_202; // @[Filter.scala 196:62]
  wire [3:0] _GEN_204 = 8'h21 == _T_40[7:0] ? 4'hf : _GEN_203; // @[Filter.scala 196:62]
  wire [3:0] _GEN_205 = 8'h22 == _T_40[7:0] ? 4'hf : _GEN_204; // @[Filter.scala 196:62]
  wire [3:0] _GEN_206 = 8'h23 == _T_40[7:0] ? 4'hf : _GEN_205; // @[Filter.scala 196:62]
  wire [3:0] _GEN_207 = 8'h24 == _T_40[7:0] ? 4'hf : _GEN_206; // @[Filter.scala 196:62]
  wire [3:0] _GEN_208 = 8'h25 == _T_40[7:0] ? 4'hf : _GEN_207; // @[Filter.scala 196:62]
  wire [3:0] _GEN_209 = 8'h26 == _T_40[7:0] ? 4'hf : _GEN_208; // @[Filter.scala 196:62]
  wire [3:0] _GEN_210 = 8'h27 == _T_40[7:0] ? 4'hf : _GEN_209; // @[Filter.scala 196:62]
  wire [3:0] _GEN_211 = 8'h28 == _T_40[7:0] ? 4'h0 : _GEN_210; // @[Filter.scala 196:62]
  wire [3:0] _GEN_212 = 8'h29 == _T_40[7:0] ? 4'h0 : _GEN_211; // @[Filter.scala 196:62]
  wire [3:0] _GEN_213 = 8'h2a == _T_40[7:0] ? 4'h0 : _GEN_212; // @[Filter.scala 196:62]
  wire [3:0] _GEN_214 = 8'h2b == _T_40[7:0] ? 4'h0 : _GEN_213; // @[Filter.scala 196:62]
  wire [3:0] _GEN_215 = 8'h2c == _T_40[7:0] ? 4'h0 : _GEN_214; // @[Filter.scala 196:62]
  wire [3:0] _GEN_216 = 8'h2d == _T_40[7:0] ? 4'h0 : _GEN_215; // @[Filter.scala 196:62]
  wire [3:0] _GEN_217 = 8'h2e == _T_40[7:0] ? 4'h0 : _GEN_216; // @[Filter.scala 196:62]
  wire [3:0] _GEN_218 = 8'h2f == _T_40[7:0] ? 4'h0 : _GEN_217; // @[Filter.scala 196:62]
  wire [3:0] _GEN_219 = 8'h30 == _T_40[7:0] ? 4'hf : _GEN_218; // @[Filter.scala 196:62]
  wire [3:0] _GEN_220 = 8'h31 == _T_40[7:0] ? 4'hf : _GEN_219; // @[Filter.scala 196:62]
  wire [3:0] _GEN_221 = 8'h32 == _T_40[7:0] ? 4'hf : _GEN_220; // @[Filter.scala 196:62]
  wire [3:0] _GEN_222 = 8'h33 == _T_40[7:0] ? 4'hf : _GEN_221; // @[Filter.scala 196:62]
  wire [3:0] _GEN_223 = 8'h34 == _T_40[7:0] ? 4'hf : _GEN_222; // @[Filter.scala 196:62]
  wire [3:0] _GEN_224 = 8'h35 == _T_40[7:0] ? 4'hf : _GEN_223; // @[Filter.scala 196:62]
  wire [3:0] _GEN_225 = 8'h36 == _T_40[7:0] ? 4'hf : _GEN_224; // @[Filter.scala 196:62]
  wire [3:0] _GEN_226 = 8'h37 == _T_40[7:0] ? 4'hf : _GEN_225; // @[Filter.scala 196:62]
  wire [3:0] _GEN_227 = 8'h38 == _T_40[7:0] ? 4'h0 : _GEN_226; // @[Filter.scala 196:62]
  wire [3:0] _GEN_228 = 8'h39 == _T_40[7:0] ? 4'h0 : _GEN_227; // @[Filter.scala 196:62]
  wire [3:0] _GEN_229 = 8'h3a == _T_40[7:0] ? 4'h0 : _GEN_228; // @[Filter.scala 196:62]
  wire [3:0] _GEN_230 = 8'h3b == _T_40[7:0] ? 4'h0 : _GEN_229; // @[Filter.scala 196:62]
  wire [3:0] _GEN_231 = 8'h3c == _T_40[7:0] ? 4'h0 : _GEN_230; // @[Filter.scala 196:62]
  wire [3:0] _GEN_232 = 8'h3d == _T_40[7:0] ? 4'h0 : _GEN_231; // @[Filter.scala 196:62]
  wire [3:0] _GEN_233 = 8'h3e == _T_40[7:0] ? 4'h0 : _GEN_232; // @[Filter.scala 196:62]
  wire [3:0] _GEN_234 = 8'h3f == _T_40[7:0] ? 4'h0 : _GEN_233; // @[Filter.scala 196:62]
  wire [3:0] _GEN_235 = 8'h40 == _T_40[7:0] ? 4'h0 : _GEN_234; // @[Filter.scala 196:62]
  wire [3:0] _GEN_236 = 8'h41 == _T_40[7:0] ? 4'h0 : _GEN_235; // @[Filter.scala 196:62]
  wire [3:0] _GEN_237 = 8'h42 == _T_40[7:0] ? 4'h0 : _GEN_236; // @[Filter.scala 196:62]
  wire [3:0] _GEN_238 = 8'h43 == _T_40[7:0] ? 4'h0 : _GEN_237; // @[Filter.scala 196:62]
  wire [3:0] _GEN_239 = 8'h44 == _T_40[7:0] ? 4'h0 : _GEN_238; // @[Filter.scala 196:62]
  wire [3:0] _GEN_240 = 8'h45 == _T_40[7:0] ? 4'h0 : _GEN_239; // @[Filter.scala 196:62]
  wire [3:0] _GEN_241 = 8'h46 == _T_40[7:0] ? 4'h0 : _GEN_240; // @[Filter.scala 196:62]
  wire [3:0] _GEN_242 = 8'h47 == _T_40[7:0] ? 4'h0 : _GEN_241; // @[Filter.scala 196:62]
  wire [3:0] _GEN_243 = 8'h48 == _T_40[7:0] ? 4'hf : _GEN_242; // @[Filter.scala 196:62]
  wire [3:0] _GEN_244 = 8'h49 == _T_40[7:0] ? 4'hf : _GEN_243; // @[Filter.scala 196:62]
  wire [3:0] _GEN_245 = 8'h4a == _T_40[7:0] ? 4'hf : _GEN_244; // @[Filter.scala 196:62]
  wire [3:0] _GEN_246 = 8'h4b == _T_40[7:0] ? 4'hf : _GEN_245; // @[Filter.scala 196:62]
  wire [3:0] _GEN_247 = 8'h4c == _T_40[7:0] ? 4'hf : _GEN_246; // @[Filter.scala 196:62]
  wire [3:0] _GEN_248 = 8'h4d == _T_40[7:0] ? 4'hf : _GEN_247; // @[Filter.scala 196:62]
  wire [3:0] _GEN_249 = 8'h4e == _T_40[7:0] ? 4'hf : _GEN_248; // @[Filter.scala 196:62]
  wire [3:0] _GEN_250 = 8'h4f == _T_40[7:0] ? 4'hf : _GEN_249; // @[Filter.scala 196:62]
  wire [3:0] _GEN_251 = 8'h50 == _T_40[7:0] ? 4'h0 : _GEN_250; // @[Filter.scala 196:62]
  wire [3:0] _GEN_252 = 8'h51 == _T_40[7:0] ? 4'h0 : _GEN_251; // @[Filter.scala 196:62]
  wire [3:0] _GEN_253 = 8'h52 == _T_40[7:0] ? 4'h0 : _GEN_252; // @[Filter.scala 196:62]
  wire [3:0] _GEN_254 = 8'h53 == _T_40[7:0] ? 4'h0 : _GEN_253; // @[Filter.scala 196:62]
  wire [3:0] _GEN_255 = 8'h54 == _T_40[7:0] ? 4'h0 : _GEN_254; // @[Filter.scala 196:62]
  wire [3:0] _GEN_256 = 8'h55 == _T_40[7:0] ? 4'h0 : _GEN_255; // @[Filter.scala 196:62]
  wire [3:0] _GEN_257 = 8'h56 == _T_40[7:0] ? 4'h0 : _GEN_256; // @[Filter.scala 196:62]
  wire [3:0] _GEN_258 = 8'h57 == _T_40[7:0] ? 4'h0 : _GEN_257; // @[Filter.scala 196:62]
  wire [3:0] _GEN_259 = 8'h58 == _T_40[7:0] ? 4'hf : _GEN_258; // @[Filter.scala 196:62]
  wire [3:0] _GEN_260 = 8'h59 == _T_40[7:0] ? 4'hf : _GEN_259; // @[Filter.scala 196:62]
  wire [3:0] _GEN_261 = 8'h5a == _T_40[7:0] ? 4'hf : _GEN_260; // @[Filter.scala 196:62]
  wire [3:0] _GEN_262 = 8'h5b == _T_40[7:0] ? 4'hf : _GEN_261; // @[Filter.scala 196:62]
  wire [3:0] _GEN_263 = 8'h5c == _T_40[7:0] ? 4'hf : _GEN_262; // @[Filter.scala 196:62]
  wire [3:0] _GEN_264 = 8'h5d == _T_40[7:0] ? 4'hf : _GEN_263; // @[Filter.scala 196:62]
  wire [3:0] _GEN_265 = 8'h5e == _T_40[7:0] ? 4'hf : _GEN_264; // @[Filter.scala 196:62]
  wire [3:0] _GEN_266 = 8'h5f == _T_40[7:0] ? 4'hf : _GEN_265; // @[Filter.scala 196:62]
  wire [3:0] _GEN_267 = 8'h60 == _T_40[7:0] ? 4'h0 : _GEN_266; // @[Filter.scala 196:62]
  wire [3:0] _GEN_268 = 8'h61 == _T_40[7:0] ? 4'h0 : _GEN_267; // @[Filter.scala 196:62]
  wire [3:0] _GEN_269 = 8'h62 == _T_40[7:0] ? 4'h0 : _GEN_268; // @[Filter.scala 196:62]
  wire [3:0] _GEN_270 = 8'h63 == _T_40[7:0] ? 4'h0 : _GEN_269; // @[Filter.scala 196:62]
  wire [3:0] _GEN_271 = 8'h64 == _T_40[7:0] ? 4'h0 : _GEN_270; // @[Filter.scala 196:62]
  wire [3:0] _GEN_272 = 8'h65 == _T_40[7:0] ? 4'h0 : _GEN_271; // @[Filter.scala 196:62]
  wire [3:0] _GEN_273 = 8'h66 == _T_40[7:0] ? 4'h0 : _GEN_272; // @[Filter.scala 196:62]
  wire [3:0] _GEN_274 = 8'h67 == _T_40[7:0] ? 4'h0 : _GEN_273; // @[Filter.scala 196:62]
  wire [3:0] _GEN_275 = 8'h68 == _T_40[7:0] ? 4'hf : _GEN_274; // @[Filter.scala 196:62]
  wire [3:0] _GEN_276 = 8'h69 == _T_40[7:0] ? 4'hf : _GEN_275; // @[Filter.scala 196:62]
  wire [3:0] _GEN_277 = 8'h6a == _T_40[7:0] ? 4'hf : _GEN_276; // @[Filter.scala 196:62]
  wire [3:0] _GEN_278 = 8'h6b == _T_40[7:0] ? 4'hf : _GEN_277; // @[Filter.scala 196:62]
  wire [3:0] _GEN_279 = 8'h6c == _T_40[7:0] ? 4'hf : _GEN_278; // @[Filter.scala 196:62]
  wire [3:0] _GEN_280 = 8'h6d == _T_40[7:0] ? 4'hf : _GEN_279; // @[Filter.scala 196:62]
  wire [3:0] _GEN_281 = 8'h6e == _T_40[7:0] ? 4'hf : _GEN_280; // @[Filter.scala 196:62]
  wire [3:0] _GEN_282 = 8'h6f == _T_40[7:0] ? 4'hf : _GEN_281; // @[Filter.scala 196:62]
  wire [3:0] _GEN_283 = 8'h70 == _T_40[7:0] ? 4'h0 : _GEN_282; // @[Filter.scala 196:62]
  wire [3:0] _GEN_284 = 8'h71 == _T_40[7:0] ? 4'h0 : _GEN_283; // @[Filter.scala 196:62]
  wire [3:0] _GEN_285 = 8'h72 == _T_40[7:0] ? 4'h0 : _GEN_284; // @[Filter.scala 196:62]
  wire [3:0] _GEN_286 = 8'h73 == _T_40[7:0] ? 4'h0 : _GEN_285; // @[Filter.scala 196:62]
  wire [3:0] _GEN_287 = 8'h74 == _T_40[7:0] ? 4'h0 : _GEN_286; // @[Filter.scala 196:62]
  wire [3:0] _GEN_288 = 8'h75 == _T_40[7:0] ? 4'h0 : _GEN_287; // @[Filter.scala 196:62]
  wire [3:0] _GEN_289 = 8'h76 == _T_40[7:0] ? 4'h0 : _GEN_288; // @[Filter.scala 196:62]
  wire [3:0] _GEN_290 = 8'h77 == _T_40[7:0] ? 4'h0 : _GEN_289; // @[Filter.scala 196:62]
  wire [3:0] _GEN_291 = 8'h78 == _T_40[7:0] ? 4'hf : _GEN_290; // @[Filter.scala 196:62]
  wire [3:0] _GEN_292 = 8'h79 == _T_40[7:0] ? 4'hf : _GEN_291; // @[Filter.scala 196:62]
  wire [3:0] _GEN_293 = 8'h7a == _T_40[7:0] ? 4'hf : _GEN_292; // @[Filter.scala 196:62]
  wire [3:0] _GEN_294 = 8'h7b == _T_40[7:0] ? 4'hf : _GEN_293; // @[Filter.scala 196:62]
  wire [3:0] _GEN_295 = 8'h7c == _T_40[7:0] ? 4'hf : _GEN_294; // @[Filter.scala 196:62]
  wire [3:0] _GEN_296 = 8'h7d == _T_40[7:0] ? 4'hf : _GEN_295; // @[Filter.scala 196:62]
  wire [3:0] _GEN_297 = 8'h7e == _T_40[7:0] ? 4'hf : _GEN_296; // @[Filter.scala 196:62]
  wire [3:0] _GEN_298 = 8'h7f == _T_40[7:0] ? 4'hf : _GEN_297; // @[Filter.scala 196:62]
  wire [3:0] _GEN_299 = 8'h80 == _T_40[7:0] ? 4'h0 : _GEN_298; // @[Filter.scala 196:62]
  wire [3:0] _GEN_300 = 8'h81 == _T_40[7:0] ? 4'h0 : _GEN_299; // @[Filter.scala 196:62]
  wire [3:0] _GEN_301 = 8'h82 == _T_40[7:0] ? 4'h0 : _GEN_300; // @[Filter.scala 196:62]
  wire [3:0] _GEN_302 = 8'h83 == _T_40[7:0] ? 4'h0 : _GEN_301; // @[Filter.scala 196:62]
  wire [3:0] _GEN_303 = 8'h84 == _T_40[7:0] ? 4'h0 : _GEN_302; // @[Filter.scala 196:62]
  wire [3:0] _GEN_304 = 8'h85 == _T_40[7:0] ? 4'h0 : _GEN_303; // @[Filter.scala 196:62]
  wire [3:0] _GEN_305 = 8'h86 == _T_40[7:0] ? 4'h0 : _GEN_304; // @[Filter.scala 196:62]
  wire [3:0] _GEN_306 = 8'h87 == _T_40[7:0] ? 4'h0 : _GEN_305; // @[Filter.scala 196:62]
  wire [3:0] _GEN_307 = 8'h88 == _T_40[7:0] ? 4'hf : _GEN_306; // @[Filter.scala 196:62]
  wire [3:0] _GEN_308 = 8'h89 == _T_40[7:0] ? 4'hf : _GEN_307; // @[Filter.scala 196:62]
  wire [3:0] _GEN_309 = 8'h8a == _T_40[7:0] ? 4'hf : _GEN_308; // @[Filter.scala 196:62]
  wire [3:0] _GEN_310 = 8'h8b == _T_40[7:0] ? 4'hf : _GEN_309; // @[Filter.scala 196:62]
  wire [3:0] _GEN_311 = 8'h8c == _T_40[7:0] ? 4'hf : _GEN_310; // @[Filter.scala 196:62]
  wire [3:0] _GEN_312 = 8'h8d == _T_40[7:0] ? 4'hf : _GEN_311; // @[Filter.scala 196:62]
  wire [3:0] _GEN_313 = 8'h8e == _T_40[7:0] ? 4'hf : _GEN_312; // @[Filter.scala 196:62]
  wire [3:0] _GEN_314 = 8'h8f == _T_40[7:0] ? 4'hf : _GEN_313; // @[Filter.scala 196:62]
  wire [4:0] _GEN_7562 = {{1'd0}, _GEN_314}; // @[Filter.scala 196:62]
  wire [8:0] _T_42 = _GEN_7562 * 5'h14; // @[Filter.scala 196:62]
  wire [3:0] _GEN_379 = 8'h40 == _T_40[7:0] ? 4'hf : 4'h0; // @[Filter.scala 196:102]
  wire [3:0] _GEN_380 = 8'h41 == _T_40[7:0] ? 4'hf : _GEN_379; // @[Filter.scala 196:102]
  wire [3:0] _GEN_381 = 8'h42 == _T_40[7:0] ? 4'hf : _GEN_380; // @[Filter.scala 196:102]
  wire [3:0] _GEN_382 = 8'h43 == _T_40[7:0] ? 4'hf : _GEN_381; // @[Filter.scala 196:102]
  wire [3:0] _GEN_383 = 8'h44 == _T_40[7:0] ? 4'hf : _GEN_382; // @[Filter.scala 196:102]
  wire [3:0] _GEN_384 = 8'h45 == _T_40[7:0] ? 4'hf : _GEN_383; // @[Filter.scala 196:102]
  wire [3:0] _GEN_385 = 8'h46 == _T_40[7:0] ? 4'hf : _GEN_384; // @[Filter.scala 196:102]
  wire [3:0] _GEN_386 = 8'h47 == _T_40[7:0] ? 4'hf : _GEN_385; // @[Filter.scala 196:102]
  wire [3:0] _GEN_387 = 8'h48 == _T_40[7:0] ? 4'hf : _GEN_386; // @[Filter.scala 196:102]
  wire [3:0] _GEN_388 = 8'h49 == _T_40[7:0] ? 4'hf : _GEN_387; // @[Filter.scala 196:102]
  wire [3:0] _GEN_389 = 8'h4a == _T_40[7:0] ? 4'hf : _GEN_388; // @[Filter.scala 196:102]
  wire [3:0] _GEN_390 = 8'h4b == _T_40[7:0] ? 4'hf : _GEN_389; // @[Filter.scala 196:102]
  wire [3:0] _GEN_391 = 8'h4c == _T_40[7:0] ? 4'hf : _GEN_390; // @[Filter.scala 196:102]
  wire [3:0] _GEN_392 = 8'h4d == _T_40[7:0] ? 4'hf : _GEN_391; // @[Filter.scala 196:102]
  wire [3:0] _GEN_393 = 8'h4e == _T_40[7:0] ? 4'hf : _GEN_392; // @[Filter.scala 196:102]
  wire [3:0] _GEN_394 = 8'h4f == _T_40[7:0] ? 4'hf : _GEN_393; // @[Filter.scala 196:102]
  wire [3:0] _GEN_395 = 8'h50 == _T_40[7:0] ? 4'hf : _GEN_394; // @[Filter.scala 196:102]
  wire [3:0] _GEN_396 = 8'h51 == _T_40[7:0] ? 4'hf : _GEN_395; // @[Filter.scala 196:102]
  wire [3:0] _GEN_397 = 8'h52 == _T_40[7:0] ? 4'hf : _GEN_396; // @[Filter.scala 196:102]
  wire [3:0] _GEN_398 = 8'h53 == _T_40[7:0] ? 4'hf : _GEN_397; // @[Filter.scala 196:102]
  wire [3:0] _GEN_399 = 8'h54 == _T_40[7:0] ? 4'hf : _GEN_398; // @[Filter.scala 196:102]
  wire [3:0] _GEN_400 = 8'h55 == _T_40[7:0] ? 4'hf : _GEN_399; // @[Filter.scala 196:102]
  wire [3:0] _GEN_401 = 8'h56 == _T_40[7:0] ? 4'hf : _GEN_400; // @[Filter.scala 196:102]
  wire [3:0] _GEN_402 = 8'h57 == _T_40[7:0] ? 4'hf : _GEN_401; // @[Filter.scala 196:102]
  wire [3:0] _GEN_403 = 8'h58 == _T_40[7:0] ? 4'hf : _GEN_402; // @[Filter.scala 196:102]
  wire [3:0] _GEN_404 = 8'h59 == _T_40[7:0] ? 4'hf : _GEN_403; // @[Filter.scala 196:102]
  wire [3:0] _GEN_405 = 8'h5a == _T_40[7:0] ? 4'hf : _GEN_404; // @[Filter.scala 196:102]
  wire [3:0] _GEN_406 = 8'h5b == _T_40[7:0] ? 4'hf : _GEN_405; // @[Filter.scala 196:102]
  wire [3:0] _GEN_407 = 8'h5c == _T_40[7:0] ? 4'hf : _GEN_406; // @[Filter.scala 196:102]
  wire [3:0] _GEN_408 = 8'h5d == _T_40[7:0] ? 4'hf : _GEN_407; // @[Filter.scala 196:102]
  wire [3:0] _GEN_409 = 8'h5e == _T_40[7:0] ? 4'hf : _GEN_408; // @[Filter.scala 196:102]
  wire [3:0] _GEN_410 = 8'h5f == _T_40[7:0] ? 4'hf : _GEN_409; // @[Filter.scala 196:102]
  wire [3:0] _GEN_411 = 8'h60 == _T_40[7:0] ? 4'hf : _GEN_410; // @[Filter.scala 196:102]
  wire [3:0] _GEN_412 = 8'h61 == _T_40[7:0] ? 4'hf : _GEN_411; // @[Filter.scala 196:102]
  wire [3:0] _GEN_413 = 8'h62 == _T_40[7:0] ? 4'hf : _GEN_412; // @[Filter.scala 196:102]
  wire [3:0] _GEN_414 = 8'h63 == _T_40[7:0] ? 4'hf : _GEN_413; // @[Filter.scala 196:102]
  wire [3:0] _GEN_415 = 8'h64 == _T_40[7:0] ? 4'hf : _GEN_414; // @[Filter.scala 196:102]
  wire [3:0] _GEN_416 = 8'h65 == _T_40[7:0] ? 4'hf : _GEN_415; // @[Filter.scala 196:102]
  wire [3:0] _GEN_417 = 8'h66 == _T_40[7:0] ? 4'hf : _GEN_416; // @[Filter.scala 196:102]
  wire [3:0] _GEN_418 = 8'h67 == _T_40[7:0] ? 4'hf : _GEN_417; // @[Filter.scala 196:102]
  wire [3:0] _GEN_419 = 8'h68 == _T_40[7:0] ? 4'hf : _GEN_418; // @[Filter.scala 196:102]
  wire [3:0] _GEN_420 = 8'h69 == _T_40[7:0] ? 4'hf : _GEN_419; // @[Filter.scala 196:102]
  wire [3:0] _GEN_421 = 8'h6a == _T_40[7:0] ? 4'hf : _GEN_420; // @[Filter.scala 196:102]
  wire [3:0] _GEN_422 = 8'h6b == _T_40[7:0] ? 4'hf : _GEN_421; // @[Filter.scala 196:102]
  wire [3:0] _GEN_423 = 8'h6c == _T_40[7:0] ? 4'hf : _GEN_422; // @[Filter.scala 196:102]
  wire [3:0] _GEN_424 = 8'h6d == _T_40[7:0] ? 4'hf : _GEN_423; // @[Filter.scala 196:102]
  wire [3:0] _GEN_425 = 8'h6e == _T_40[7:0] ? 4'hf : _GEN_424; // @[Filter.scala 196:102]
  wire [3:0] _GEN_426 = 8'h6f == _T_40[7:0] ? 4'hf : _GEN_425; // @[Filter.scala 196:102]
  wire [3:0] _GEN_427 = 8'h70 == _T_40[7:0] ? 4'hf : _GEN_426; // @[Filter.scala 196:102]
  wire [3:0] _GEN_428 = 8'h71 == _T_40[7:0] ? 4'hf : _GEN_427; // @[Filter.scala 196:102]
  wire [3:0] _GEN_429 = 8'h72 == _T_40[7:0] ? 4'hf : _GEN_428; // @[Filter.scala 196:102]
  wire [3:0] _GEN_430 = 8'h73 == _T_40[7:0] ? 4'hf : _GEN_429; // @[Filter.scala 196:102]
  wire [3:0] _GEN_431 = 8'h74 == _T_40[7:0] ? 4'hf : _GEN_430; // @[Filter.scala 196:102]
  wire [3:0] _GEN_432 = 8'h75 == _T_40[7:0] ? 4'hf : _GEN_431; // @[Filter.scala 196:102]
  wire [3:0] _GEN_433 = 8'h76 == _T_40[7:0] ? 4'hf : _GEN_432; // @[Filter.scala 196:102]
  wire [3:0] _GEN_434 = 8'h77 == _T_40[7:0] ? 4'hf : _GEN_433; // @[Filter.scala 196:102]
  wire [3:0] _GEN_435 = 8'h78 == _T_40[7:0] ? 4'hf : _GEN_434; // @[Filter.scala 196:102]
  wire [3:0] _GEN_436 = 8'h79 == _T_40[7:0] ? 4'hf : _GEN_435; // @[Filter.scala 196:102]
  wire [3:0] _GEN_437 = 8'h7a == _T_40[7:0] ? 4'hf : _GEN_436; // @[Filter.scala 196:102]
  wire [3:0] _GEN_438 = 8'h7b == _T_40[7:0] ? 4'hf : _GEN_437; // @[Filter.scala 196:102]
  wire [3:0] _GEN_439 = 8'h7c == _T_40[7:0] ? 4'hf : _GEN_438; // @[Filter.scala 196:102]
  wire [3:0] _GEN_440 = 8'h7d == _T_40[7:0] ? 4'hf : _GEN_439; // @[Filter.scala 196:102]
  wire [3:0] _GEN_441 = 8'h7e == _T_40[7:0] ? 4'hf : _GEN_440; // @[Filter.scala 196:102]
  wire [3:0] _GEN_442 = 8'h7f == _T_40[7:0] ? 4'hf : _GEN_441; // @[Filter.scala 196:102]
  wire [3:0] _GEN_443 = 8'h80 == _T_40[7:0] ? 4'hf : _GEN_442; // @[Filter.scala 196:102]
  wire [3:0] _GEN_444 = 8'h81 == _T_40[7:0] ? 4'hf : _GEN_443; // @[Filter.scala 196:102]
  wire [3:0] _GEN_445 = 8'h82 == _T_40[7:0] ? 4'hf : _GEN_444; // @[Filter.scala 196:102]
  wire [3:0] _GEN_446 = 8'h83 == _T_40[7:0] ? 4'hf : _GEN_445; // @[Filter.scala 196:102]
  wire [3:0] _GEN_447 = 8'h84 == _T_40[7:0] ? 4'hf : _GEN_446; // @[Filter.scala 196:102]
  wire [3:0] _GEN_448 = 8'h85 == _T_40[7:0] ? 4'hf : _GEN_447; // @[Filter.scala 196:102]
  wire [3:0] _GEN_449 = 8'h86 == _T_40[7:0] ? 4'hf : _GEN_448; // @[Filter.scala 196:102]
  wire [3:0] _GEN_450 = 8'h87 == _T_40[7:0] ? 4'hf : _GEN_449; // @[Filter.scala 196:102]
  wire [3:0] _GEN_451 = 8'h88 == _T_40[7:0] ? 4'hf : _GEN_450; // @[Filter.scala 196:102]
  wire [3:0] _GEN_452 = 8'h89 == _T_40[7:0] ? 4'hf : _GEN_451; // @[Filter.scala 196:102]
  wire [3:0] _GEN_453 = 8'h8a == _T_40[7:0] ? 4'hf : _GEN_452; // @[Filter.scala 196:102]
  wire [3:0] _GEN_454 = 8'h8b == _T_40[7:0] ? 4'hf : _GEN_453; // @[Filter.scala 196:102]
  wire [3:0] _GEN_455 = 8'h8c == _T_40[7:0] ? 4'hf : _GEN_454; // @[Filter.scala 196:102]
  wire [3:0] _GEN_456 = 8'h8d == _T_40[7:0] ? 4'hf : _GEN_455; // @[Filter.scala 196:102]
  wire [3:0] _GEN_457 = 8'h8e == _T_40[7:0] ? 4'hf : _GEN_456; // @[Filter.scala 196:102]
  wire [3:0] _GEN_458 = 8'h8f == _T_40[7:0] ? 4'hf : _GEN_457; // @[Filter.scala 196:102]
  wire [6:0] _GEN_7564 = {{3'd0}, _GEN_458}; // @[Filter.scala 196:102]
  wire [10:0] _T_47 = _GEN_7564 * 7'h46; // @[Filter.scala 196:102]
  wire [10:0] _GEN_7565 = {{2'd0}, _T_42}; // @[Filter.scala 196:69]
  wire [10:0] _T_49 = _GEN_7565 + _T_47; // @[Filter.scala 196:69]
  wire [3:0] _GEN_467 = 8'h8 == _T_40[7:0] ? 4'hf : 4'h0; // @[Filter.scala 196:142]
  wire [3:0] _GEN_468 = 8'h9 == _T_40[7:0] ? 4'hf : _GEN_467; // @[Filter.scala 196:142]
  wire [3:0] _GEN_469 = 8'ha == _T_40[7:0] ? 4'hf : _GEN_468; // @[Filter.scala 196:142]
  wire [3:0] _GEN_470 = 8'hb == _T_40[7:0] ? 4'hf : _GEN_469; // @[Filter.scala 196:142]
  wire [3:0] _GEN_471 = 8'hc == _T_40[7:0] ? 4'hf : _GEN_470; // @[Filter.scala 196:142]
  wire [3:0] _GEN_472 = 8'hd == _T_40[7:0] ? 4'hf : _GEN_471; // @[Filter.scala 196:142]
  wire [3:0] _GEN_473 = 8'he == _T_40[7:0] ? 4'hf : _GEN_472; // @[Filter.scala 196:142]
  wire [3:0] _GEN_474 = 8'hf == _T_40[7:0] ? 4'hf : _GEN_473; // @[Filter.scala 196:142]
  wire [3:0] _GEN_475 = 8'h10 == _T_40[7:0] ? 4'h0 : _GEN_474; // @[Filter.scala 196:142]
  wire [3:0] _GEN_476 = 8'h11 == _T_40[7:0] ? 4'h0 : _GEN_475; // @[Filter.scala 196:142]
  wire [3:0] _GEN_477 = 8'h12 == _T_40[7:0] ? 4'h0 : _GEN_476; // @[Filter.scala 196:142]
  wire [3:0] _GEN_478 = 8'h13 == _T_40[7:0] ? 4'h0 : _GEN_477; // @[Filter.scala 196:142]
  wire [3:0] _GEN_479 = 8'h14 == _T_40[7:0] ? 4'h0 : _GEN_478; // @[Filter.scala 196:142]
  wire [3:0] _GEN_480 = 8'h15 == _T_40[7:0] ? 4'h0 : _GEN_479; // @[Filter.scala 196:142]
  wire [3:0] _GEN_481 = 8'h16 == _T_40[7:0] ? 4'h0 : _GEN_480; // @[Filter.scala 196:142]
  wire [3:0] _GEN_482 = 8'h17 == _T_40[7:0] ? 4'h0 : _GEN_481; // @[Filter.scala 196:142]
  wire [3:0] _GEN_483 = 8'h18 == _T_40[7:0] ? 4'hf : _GEN_482; // @[Filter.scala 196:142]
  wire [3:0] _GEN_484 = 8'h19 == _T_40[7:0] ? 4'hf : _GEN_483; // @[Filter.scala 196:142]
  wire [3:0] _GEN_485 = 8'h1a == _T_40[7:0] ? 4'hf : _GEN_484; // @[Filter.scala 196:142]
  wire [3:0] _GEN_486 = 8'h1b == _T_40[7:0] ? 4'hf : _GEN_485; // @[Filter.scala 196:142]
  wire [3:0] _GEN_487 = 8'h1c == _T_40[7:0] ? 4'hf : _GEN_486; // @[Filter.scala 196:142]
  wire [3:0] _GEN_488 = 8'h1d == _T_40[7:0] ? 4'hf : _GEN_487; // @[Filter.scala 196:142]
  wire [3:0] _GEN_489 = 8'h1e == _T_40[7:0] ? 4'hf : _GEN_488; // @[Filter.scala 196:142]
  wire [3:0] _GEN_490 = 8'h1f == _T_40[7:0] ? 4'hf : _GEN_489; // @[Filter.scala 196:142]
  wire [3:0] _GEN_491 = 8'h20 == _T_40[7:0] ? 4'h0 : _GEN_490; // @[Filter.scala 196:142]
  wire [3:0] _GEN_492 = 8'h21 == _T_40[7:0] ? 4'h0 : _GEN_491; // @[Filter.scala 196:142]
  wire [3:0] _GEN_493 = 8'h22 == _T_40[7:0] ? 4'h0 : _GEN_492; // @[Filter.scala 196:142]
  wire [3:0] _GEN_494 = 8'h23 == _T_40[7:0] ? 4'h0 : _GEN_493; // @[Filter.scala 196:142]
  wire [3:0] _GEN_495 = 8'h24 == _T_40[7:0] ? 4'h0 : _GEN_494; // @[Filter.scala 196:142]
  wire [3:0] _GEN_496 = 8'h25 == _T_40[7:0] ? 4'h0 : _GEN_495; // @[Filter.scala 196:142]
  wire [3:0] _GEN_497 = 8'h26 == _T_40[7:0] ? 4'h0 : _GEN_496; // @[Filter.scala 196:142]
  wire [3:0] _GEN_498 = 8'h27 == _T_40[7:0] ? 4'h0 : _GEN_497; // @[Filter.scala 196:142]
  wire [3:0] _GEN_499 = 8'h28 == _T_40[7:0] ? 4'hf : _GEN_498; // @[Filter.scala 196:142]
  wire [3:0] _GEN_500 = 8'h29 == _T_40[7:0] ? 4'hf : _GEN_499; // @[Filter.scala 196:142]
  wire [3:0] _GEN_501 = 8'h2a == _T_40[7:0] ? 4'hf : _GEN_500; // @[Filter.scala 196:142]
  wire [3:0] _GEN_502 = 8'h2b == _T_40[7:0] ? 4'hf : _GEN_501; // @[Filter.scala 196:142]
  wire [3:0] _GEN_503 = 8'h2c == _T_40[7:0] ? 4'hf : _GEN_502; // @[Filter.scala 196:142]
  wire [3:0] _GEN_504 = 8'h2d == _T_40[7:0] ? 4'hf : _GEN_503; // @[Filter.scala 196:142]
  wire [3:0] _GEN_505 = 8'h2e == _T_40[7:0] ? 4'hf : _GEN_504; // @[Filter.scala 196:142]
  wire [3:0] _GEN_506 = 8'h2f == _T_40[7:0] ? 4'hf : _GEN_505; // @[Filter.scala 196:142]
  wire [3:0] _GEN_507 = 8'h30 == _T_40[7:0] ? 4'h0 : _GEN_506; // @[Filter.scala 196:142]
  wire [3:0] _GEN_508 = 8'h31 == _T_40[7:0] ? 4'h0 : _GEN_507; // @[Filter.scala 196:142]
  wire [3:0] _GEN_509 = 8'h32 == _T_40[7:0] ? 4'h0 : _GEN_508; // @[Filter.scala 196:142]
  wire [3:0] _GEN_510 = 8'h33 == _T_40[7:0] ? 4'h0 : _GEN_509; // @[Filter.scala 196:142]
  wire [3:0] _GEN_511 = 8'h34 == _T_40[7:0] ? 4'h0 : _GEN_510; // @[Filter.scala 196:142]
  wire [3:0] _GEN_512 = 8'h35 == _T_40[7:0] ? 4'h0 : _GEN_511; // @[Filter.scala 196:142]
  wire [3:0] _GEN_513 = 8'h36 == _T_40[7:0] ? 4'h0 : _GEN_512; // @[Filter.scala 196:142]
  wire [3:0] _GEN_514 = 8'h37 == _T_40[7:0] ? 4'h0 : _GEN_513; // @[Filter.scala 196:142]
  wire [3:0] _GEN_515 = 8'h38 == _T_40[7:0] ? 4'hf : _GEN_514; // @[Filter.scala 196:142]
  wire [3:0] _GEN_516 = 8'h39 == _T_40[7:0] ? 4'hf : _GEN_515; // @[Filter.scala 196:142]
  wire [3:0] _GEN_517 = 8'h3a == _T_40[7:0] ? 4'hf : _GEN_516; // @[Filter.scala 196:142]
  wire [3:0] _GEN_518 = 8'h3b == _T_40[7:0] ? 4'hf : _GEN_517; // @[Filter.scala 196:142]
  wire [3:0] _GEN_519 = 8'h3c == _T_40[7:0] ? 4'hf : _GEN_518; // @[Filter.scala 196:142]
  wire [3:0] _GEN_520 = 8'h3d == _T_40[7:0] ? 4'hf : _GEN_519; // @[Filter.scala 196:142]
  wire [3:0] _GEN_521 = 8'h3e == _T_40[7:0] ? 4'hf : _GEN_520; // @[Filter.scala 196:142]
  wire [3:0] _GEN_522 = 8'h3f == _T_40[7:0] ? 4'hf : _GEN_521; // @[Filter.scala 196:142]
  wire [3:0] _GEN_523 = 8'h40 == _T_40[7:0] ? 4'h0 : _GEN_522; // @[Filter.scala 196:142]
  wire [3:0] _GEN_524 = 8'h41 == _T_40[7:0] ? 4'h0 : _GEN_523; // @[Filter.scala 196:142]
  wire [3:0] _GEN_525 = 8'h42 == _T_40[7:0] ? 4'h0 : _GEN_524; // @[Filter.scala 196:142]
  wire [3:0] _GEN_526 = 8'h43 == _T_40[7:0] ? 4'h0 : _GEN_525; // @[Filter.scala 196:142]
  wire [3:0] _GEN_527 = 8'h44 == _T_40[7:0] ? 4'h0 : _GEN_526; // @[Filter.scala 196:142]
  wire [3:0] _GEN_528 = 8'h45 == _T_40[7:0] ? 4'h0 : _GEN_527; // @[Filter.scala 196:142]
  wire [3:0] _GEN_529 = 8'h46 == _T_40[7:0] ? 4'h0 : _GEN_528; // @[Filter.scala 196:142]
  wire [3:0] _GEN_530 = 8'h47 == _T_40[7:0] ? 4'h0 : _GEN_529; // @[Filter.scala 196:142]
  wire [3:0] _GEN_531 = 8'h48 == _T_40[7:0] ? 4'hf : _GEN_530; // @[Filter.scala 196:142]
  wire [3:0] _GEN_532 = 8'h49 == _T_40[7:0] ? 4'hf : _GEN_531; // @[Filter.scala 196:142]
  wire [3:0] _GEN_533 = 8'h4a == _T_40[7:0] ? 4'hf : _GEN_532; // @[Filter.scala 196:142]
  wire [3:0] _GEN_534 = 8'h4b == _T_40[7:0] ? 4'hf : _GEN_533; // @[Filter.scala 196:142]
  wire [3:0] _GEN_535 = 8'h4c == _T_40[7:0] ? 4'hf : _GEN_534; // @[Filter.scala 196:142]
  wire [3:0] _GEN_536 = 8'h4d == _T_40[7:0] ? 4'hf : _GEN_535; // @[Filter.scala 196:142]
  wire [3:0] _GEN_537 = 8'h4e == _T_40[7:0] ? 4'hf : _GEN_536; // @[Filter.scala 196:142]
  wire [3:0] _GEN_538 = 8'h4f == _T_40[7:0] ? 4'hf : _GEN_537; // @[Filter.scala 196:142]
  wire [3:0] _GEN_539 = 8'h50 == _T_40[7:0] ? 4'h0 : _GEN_538; // @[Filter.scala 196:142]
  wire [3:0] _GEN_540 = 8'h51 == _T_40[7:0] ? 4'h0 : _GEN_539; // @[Filter.scala 196:142]
  wire [3:0] _GEN_541 = 8'h52 == _T_40[7:0] ? 4'h0 : _GEN_540; // @[Filter.scala 196:142]
  wire [3:0] _GEN_542 = 8'h53 == _T_40[7:0] ? 4'h0 : _GEN_541; // @[Filter.scala 196:142]
  wire [3:0] _GEN_543 = 8'h54 == _T_40[7:0] ? 4'h0 : _GEN_542; // @[Filter.scala 196:142]
  wire [3:0] _GEN_544 = 8'h55 == _T_40[7:0] ? 4'h0 : _GEN_543; // @[Filter.scala 196:142]
  wire [3:0] _GEN_545 = 8'h56 == _T_40[7:0] ? 4'h0 : _GEN_544; // @[Filter.scala 196:142]
  wire [3:0] _GEN_546 = 8'h57 == _T_40[7:0] ? 4'h0 : _GEN_545; // @[Filter.scala 196:142]
  wire [3:0] _GEN_547 = 8'h58 == _T_40[7:0] ? 4'hf : _GEN_546; // @[Filter.scala 196:142]
  wire [3:0] _GEN_548 = 8'h59 == _T_40[7:0] ? 4'hf : _GEN_547; // @[Filter.scala 196:142]
  wire [3:0] _GEN_549 = 8'h5a == _T_40[7:0] ? 4'hf : _GEN_548; // @[Filter.scala 196:142]
  wire [3:0] _GEN_550 = 8'h5b == _T_40[7:0] ? 4'hf : _GEN_549; // @[Filter.scala 196:142]
  wire [3:0] _GEN_551 = 8'h5c == _T_40[7:0] ? 4'hf : _GEN_550; // @[Filter.scala 196:142]
  wire [3:0] _GEN_552 = 8'h5d == _T_40[7:0] ? 4'hf : _GEN_551; // @[Filter.scala 196:142]
  wire [3:0] _GEN_553 = 8'h5e == _T_40[7:0] ? 4'hf : _GEN_552; // @[Filter.scala 196:142]
  wire [3:0] _GEN_554 = 8'h5f == _T_40[7:0] ? 4'hf : _GEN_553; // @[Filter.scala 196:142]
  wire [3:0] _GEN_555 = 8'h60 == _T_40[7:0] ? 4'h0 : _GEN_554; // @[Filter.scala 196:142]
  wire [3:0] _GEN_556 = 8'h61 == _T_40[7:0] ? 4'h0 : _GEN_555; // @[Filter.scala 196:142]
  wire [3:0] _GEN_557 = 8'h62 == _T_40[7:0] ? 4'h0 : _GEN_556; // @[Filter.scala 196:142]
  wire [3:0] _GEN_558 = 8'h63 == _T_40[7:0] ? 4'h0 : _GEN_557; // @[Filter.scala 196:142]
  wire [3:0] _GEN_559 = 8'h64 == _T_40[7:0] ? 4'h0 : _GEN_558; // @[Filter.scala 196:142]
  wire [3:0] _GEN_560 = 8'h65 == _T_40[7:0] ? 4'h0 : _GEN_559; // @[Filter.scala 196:142]
  wire [3:0] _GEN_561 = 8'h66 == _T_40[7:0] ? 4'h0 : _GEN_560; // @[Filter.scala 196:142]
  wire [3:0] _GEN_562 = 8'h67 == _T_40[7:0] ? 4'h0 : _GEN_561; // @[Filter.scala 196:142]
  wire [3:0] _GEN_563 = 8'h68 == _T_40[7:0] ? 4'hf : _GEN_562; // @[Filter.scala 196:142]
  wire [3:0] _GEN_564 = 8'h69 == _T_40[7:0] ? 4'hf : _GEN_563; // @[Filter.scala 196:142]
  wire [3:0] _GEN_565 = 8'h6a == _T_40[7:0] ? 4'hf : _GEN_564; // @[Filter.scala 196:142]
  wire [3:0] _GEN_566 = 8'h6b == _T_40[7:0] ? 4'hf : _GEN_565; // @[Filter.scala 196:142]
  wire [3:0] _GEN_567 = 8'h6c == _T_40[7:0] ? 4'hf : _GEN_566; // @[Filter.scala 196:142]
  wire [3:0] _GEN_568 = 8'h6d == _T_40[7:0] ? 4'hf : _GEN_567; // @[Filter.scala 196:142]
  wire [3:0] _GEN_569 = 8'h6e == _T_40[7:0] ? 4'hf : _GEN_568; // @[Filter.scala 196:142]
  wire [3:0] _GEN_570 = 8'h6f == _T_40[7:0] ? 4'hf : _GEN_569; // @[Filter.scala 196:142]
  wire [3:0] _GEN_571 = 8'h70 == _T_40[7:0] ? 4'h0 : _GEN_570; // @[Filter.scala 196:142]
  wire [3:0] _GEN_572 = 8'h71 == _T_40[7:0] ? 4'h0 : _GEN_571; // @[Filter.scala 196:142]
  wire [3:0] _GEN_573 = 8'h72 == _T_40[7:0] ? 4'h0 : _GEN_572; // @[Filter.scala 196:142]
  wire [3:0] _GEN_574 = 8'h73 == _T_40[7:0] ? 4'h0 : _GEN_573; // @[Filter.scala 196:142]
  wire [3:0] _GEN_575 = 8'h74 == _T_40[7:0] ? 4'h0 : _GEN_574; // @[Filter.scala 196:142]
  wire [3:0] _GEN_576 = 8'h75 == _T_40[7:0] ? 4'h0 : _GEN_575; // @[Filter.scala 196:142]
  wire [3:0] _GEN_577 = 8'h76 == _T_40[7:0] ? 4'h0 : _GEN_576; // @[Filter.scala 196:142]
  wire [3:0] _GEN_578 = 8'h77 == _T_40[7:0] ? 4'h0 : _GEN_577; // @[Filter.scala 196:142]
  wire [3:0] _GEN_579 = 8'h78 == _T_40[7:0] ? 4'hf : _GEN_578; // @[Filter.scala 196:142]
  wire [3:0] _GEN_580 = 8'h79 == _T_40[7:0] ? 4'hf : _GEN_579; // @[Filter.scala 196:142]
  wire [3:0] _GEN_581 = 8'h7a == _T_40[7:0] ? 4'hf : _GEN_580; // @[Filter.scala 196:142]
  wire [3:0] _GEN_582 = 8'h7b == _T_40[7:0] ? 4'hf : _GEN_581; // @[Filter.scala 196:142]
  wire [3:0] _GEN_583 = 8'h7c == _T_40[7:0] ? 4'hf : _GEN_582; // @[Filter.scala 196:142]
  wire [3:0] _GEN_584 = 8'h7d == _T_40[7:0] ? 4'hf : _GEN_583; // @[Filter.scala 196:142]
  wire [3:0] _GEN_585 = 8'h7e == _T_40[7:0] ? 4'hf : _GEN_584; // @[Filter.scala 196:142]
  wire [3:0] _GEN_586 = 8'h7f == _T_40[7:0] ? 4'hf : _GEN_585; // @[Filter.scala 196:142]
  wire [3:0] _GEN_587 = 8'h80 == _T_40[7:0] ? 4'h0 : _GEN_586; // @[Filter.scala 196:142]
  wire [3:0] _GEN_588 = 8'h81 == _T_40[7:0] ? 4'h0 : _GEN_587; // @[Filter.scala 196:142]
  wire [3:0] _GEN_589 = 8'h82 == _T_40[7:0] ? 4'h0 : _GEN_588; // @[Filter.scala 196:142]
  wire [3:0] _GEN_590 = 8'h83 == _T_40[7:0] ? 4'h0 : _GEN_589; // @[Filter.scala 196:142]
  wire [3:0] _GEN_591 = 8'h84 == _T_40[7:0] ? 4'h0 : _GEN_590; // @[Filter.scala 196:142]
  wire [3:0] _GEN_592 = 8'h85 == _T_40[7:0] ? 4'h0 : _GEN_591; // @[Filter.scala 196:142]
  wire [3:0] _GEN_593 = 8'h86 == _T_40[7:0] ? 4'h0 : _GEN_592; // @[Filter.scala 196:142]
  wire [3:0] _GEN_594 = 8'h87 == _T_40[7:0] ? 4'h0 : _GEN_593; // @[Filter.scala 196:142]
  wire [3:0] _GEN_595 = 8'h88 == _T_40[7:0] ? 4'hf : _GEN_594; // @[Filter.scala 196:142]
  wire [3:0] _GEN_596 = 8'h89 == _T_40[7:0] ? 4'hf : _GEN_595; // @[Filter.scala 196:142]
  wire [3:0] _GEN_597 = 8'h8a == _T_40[7:0] ? 4'hf : _GEN_596; // @[Filter.scala 196:142]
  wire [3:0] _GEN_598 = 8'h8b == _T_40[7:0] ? 4'hf : _GEN_597; // @[Filter.scala 196:142]
  wire [3:0] _GEN_599 = 8'h8c == _T_40[7:0] ? 4'hf : _GEN_598; // @[Filter.scala 196:142]
  wire [3:0] _GEN_600 = 8'h8d == _T_40[7:0] ? 4'hf : _GEN_599; // @[Filter.scala 196:142]
  wire [3:0] _GEN_601 = 8'h8e == _T_40[7:0] ? 4'hf : _GEN_600; // @[Filter.scala 196:142]
  wire [3:0] _GEN_602 = 8'h8f == _T_40[7:0] ? 4'hf : _GEN_601; // @[Filter.scala 196:142]
  wire [7:0] _T_54 = _GEN_602 * 4'ha; // @[Filter.scala 196:142]
  wire [10:0] _GEN_7567 = {{3'd0}, _T_54}; // @[Filter.scala 196:109]
  wire [10:0] _T_56 = _T_49 + _GEN_7567; // @[Filter.scala 196:109]
  wire [10:0] _T_57 = _T_56 / 11'h64; // @[Filter.scala 196:150]
  wire  _T_59 = _T_30 >= 5'h10; // @[Filter.scala 199:31]
  wire  _T_63 = _T_37 >= 32'h9; // @[Filter.scala 199:63]
  wire  _T_64 = _T_59 | _T_63; // @[Filter.scala 199:58]
  wire [10:0] _GEN_747 = io_SPI_distort ? _T_57 : {{7'd0}, _GEN_314}; // @[Filter.scala 201:35]
  wire [10:0] _GEN_748 = _T_64 ? 11'h0 : _GEN_747; // @[Filter.scala 199:80]
  wire [10:0] _GEN_893 = io_SPI_distort ? _T_57 : {{7'd0}, _GEN_458}; // @[Filter.scala 201:35]
  wire [10:0] _GEN_894 = _T_64 ? 11'h0 : _GEN_893; // @[Filter.scala 199:80]
  wire [10:0] _GEN_1039 = io_SPI_distort ? _T_57 : {{7'd0}, _GEN_602}; // @[Filter.scala 201:35]
  wire [10:0] _GEN_1040 = _T_64 ? 11'h0 : _GEN_1039; // @[Filter.scala 199:80]
  wire [31:0] _T_92 = pixelIndex + 32'h1; // @[Filter.scala 194:31]
  wire [31:0] _GEN_1 = _T_92 % 32'h10; // @[Filter.scala 194:38]
  wire [4:0] _T_93 = _GEN_1[4:0]; // @[Filter.scala 194:38]
  wire [4:0] _T_95 = _T_93 + _GEN_7559; // @[Filter.scala 194:53]
  wire [4:0] _T_97 = _T_95 - 5'h1; // @[Filter.scala 194:69]
  wire [31:0] _T_100 = _T_92 / 32'h10; // @[Filter.scala 195:38]
  wire [31:0] _T_102 = _T_100 + _GEN_7560; // @[Filter.scala 195:53]
  wire [31:0] _T_104 = _T_102 - 32'h1; // @[Filter.scala 195:69]
  wire [36:0] _T_105 = _T_104 * 32'h10; // @[Filter.scala 196:42]
  wire [36:0] _GEN_7573 = {{32'd0}, _T_97}; // @[Filter.scala 196:57]
  wire [36:0] _T_107 = _T_105 + _GEN_7573; // @[Filter.scala 196:57]
  wire [3:0] _GEN_1049 = 8'h8 == _T_107[7:0] ? 4'h0 : 4'hf; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1050 = 8'h9 == _T_107[7:0] ? 4'h0 : _GEN_1049; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1051 = 8'ha == _T_107[7:0] ? 4'h0 : _GEN_1050; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1052 = 8'hb == _T_107[7:0] ? 4'h0 : _GEN_1051; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1053 = 8'hc == _T_107[7:0] ? 4'h0 : _GEN_1052; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1054 = 8'hd == _T_107[7:0] ? 4'h0 : _GEN_1053; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1055 = 8'he == _T_107[7:0] ? 4'h0 : _GEN_1054; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1056 = 8'hf == _T_107[7:0] ? 4'h0 : _GEN_1055; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1057 = 8'h10 == _T_107[7:0] ? 4'hf : _GEN_1056; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1058 = 8'h11 == _T_107[7:0] ? 4'hf : _GEN_1057; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1059 = 8'h12 == _T_107[7:0] ? 4'hf : _GEN_1058; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1060 = 8'h13 == _T_107[7:0] ? 4'hf : _GEN_1059; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1061 = 8'h14 == _T_107[7:0] ? 4'hf : _GEN_1060; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1062 = 8'h15 == _T_107[7:0] ? 4'hf : _GEN_1061; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1063 = 8'h16 == _T_107[7:0] ? 4'hf : _GEN_1062; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1064 = 8'h17 == _T_107[7:0] ? 4'hf : _GEN_1063; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1065 = 8'h18 == _T_107[7:0] ? 4'h0 : _GEN_1064; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1066 = 8'h19 == _T_107[7:0] ? 4'h0 : _GEN_1065; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1067 = 8'h1a == _T_107[7:0] ? 4'h0 : _GEN_1066; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1068 = 8'h1b == _T_107[7:0] ? 4'h0 : _GEN_1067; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1069 = 8'h1c == _T_107[7:0] ? 4'h0 : _GEN_1068; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1070 = 8'h1d == _T_107[7:0] ? 4'h0 : _GEN_1069; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1071 = 8'h1e == _T_107[7:0] ? 4'h0 : _GEN_1070; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1072 = 8'h1f == _T_107[7:0] ? 4'h0 : _GEN_1071; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1073 = 8'h20 == _T_107[7:0] ? 4'hf : _GEN_1072; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1074 = 8'h21 == _T_107[7:0] ? 4'hf : _GEN_1073; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1075 = 8'h22 == _T_107[7:0] ? 4'hf : _GEN_1074; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1076 = 8'h23 == _T_107[7:0] ? 4'hf : _GEN_1075; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1077 = 8'h24 == _T_107[7:0] ? 4'hf : _GEN_1076; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1078 = 8'h25 == _T_107[7:0] ? 4'hf : _GEN_1077; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1079 = 8'h26 == _T_107[7:0] ? 4'hf : _GEN_1078; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1080 = 8'h27 == _T_107[7:0] ? 4'hf : _GEN_1079; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1081 = 8'h28 == _T_107[7:0] ? 4'h0 : _GEN_1080; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1082 = 8'h29 == _T_107[7:0] ? 4'h0 : _GEN_1081; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1083 = 8'h2a == _T_107[7:0] ? 4'h0 : _GEN_1082; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1084 = 8'h2b == _T_107[7:0] ? 4'h0 : _GEN_1083; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1085 = 8'h2c == _T_107[7:0] ? 4'h0 : _GEN_1084; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1086 = 8'h2d == _T_107[7:0] ? 4'h0 : _GEN_1085; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1087 = 8'h2e == _T_107[7:0] ? 4'h0 : _GEN_1086; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1088 = 8'h2f == _T_107[7:0] ? 4'h0 : _GEN_1087; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1089 = 8'h30 == _T_107[7:0] ? 4'hf : _GEN_1088; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1090 = 8'h31 == _T_107[7:0] ? 4'hf : _GEN_1089; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1091 = 8'h32 == _T_107[7:0] ? 4'hf : _GEN_1090; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1092 = 8'h33 == _T_107[7:0] ? 4'hf : _GEN_1091; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1093 = 8'h34 == _T_107[7:0] ? 4'hf : _GEN_1092; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1094 = 8'h35 == _T_107[7:0] ? 4'hf : _GEN_1093; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1095 = 8'h36 == _T_107[7:0] ? 4'hf : _GEN_1094; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1096 = 8'h37 == _T_107[7:0] ? 4'hf : _GEN_1095; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1097 = 8'h38 == _T_107[7:0] ? 4'h0 : _GEN_1096; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1098 = 8'h39 == _T_107[7:0] ? 4'h0 : _GEN_1097; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1099 = 8'h3a == _T_107[7:0] ? 4'h0 : _GEN_1098; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1100 = 8'h3b == _T_107[7:0] ? 4'h0 : _GEN_1099; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1101 = 8'h3c == _T_107[7:0] ? 4'h0 : _GEN_1100; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1102 = 8'h3d == _T_107[7:0] ? 4'h0 : _GEN_1101; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1103 = 8'h3e == _T_107[7:0] ? 4'h0 : _GEN_1102; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1104 = 8'h3f == _T_107[7:0] ? 4'h0 : _GEN_1103; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1105 = 8'h40 == _T_107[7:0] ? 4'h0 : _GEN_1104; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1106 = 8'h41 == _T_107[7:0] ? 4'h0 : _GEN_1105; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1107 = 8'h42 == _T_107[7:0] ? 4'h0 : _GEN_1106; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1108 = 8'h43 == _T_107[7:0] ? 4'h0 : _GEN_1107; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1109 = 8'h44 == _T_107[7:0] ? 4'h0 : _GEN_1108; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1110 = 8'h45 == _T_107[7:0] ? 4'h0 : _GEN_1109; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1111 = 8'h46 == _T_107[7:0] ? 4'h0 : _GEN_1110; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1112 = 8'h47 == _T_107[7:0] ? 4'h0 : _GEN_1111; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1113 = 8'h48 == _T_107[7:0] ? 4'hf : _GEN_1112; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1114 = 8'h49 == _T_107[7:0] ? 4'hf : _GEN_1113; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1115 = 8'h4a == _T_107[7:0] ? 4'hf : _GEN_1114; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1116 = 8'h4b == _T_107[7:0] ? 4'hf : _GEN_1115; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1117 = 8'h4c == _T_107[7:0] ? 4'hf : _GEN_1116; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1118 = 8'h4d == _T_107[7:0] ? 4'hf : _GEN_1117; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1119 = 8'h4e == _T_107[7:0] ? 4'hf : _GEN_1118; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1120 = 8'h4f == _T_107[7:0] ? 4'hf : _GEN_1119; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1121 = 8'h50 == _T_107[7:0] ? 4'h0 : _GEN_1120; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1122 = 8'h51 == _T_107[7:0] ? 4'h0 : _GEN_1121; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1123 = 8'h52 == _T_107[7:0] ? 4'h0 : _GEN_1122; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1124 = 8'h53 == _T_107[7:0] ? 4'h0 : _GEN_1123; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1125 = 8'h54 == _T_107[7:0] ? 4'h0 : _GEN_1124; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1126 = 8'h55 == _T_107[7:0] ? 4'h0 : _GEN_1125; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1127 = 8'h56 == _T_107[7:0] ? 4'h0 : _GEN_1126; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1128 = 8'h57 == _T_107[7:0] ? 4'h0 : _GEN_1127; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1129 = 8'h58 == _T_107[7:0] ? 4'hf : _GEN_1128; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1130 = 8'h59 == _T_107[7:0] ? 4'hf : _GEN_1129; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1131 = 8'h5a == _T_107[7:0] ? 4'hf : _GEN_1130; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1132 = 8'h5b == _T_107[7:0] ? 4'hf : _GEN_1131; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1133 = 8'h5c == _T_107[7:0] ? 4'hf : _GEN_1132; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1134 = 8'h5d == _T_107[7:0] ? 4'hf : _GEN_1133; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1135 = 8'h5e == _T_107[7:0] ? 4'hf : _GEN_1134; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1136 = 8'h5f == _T_107[7:0] ? 4'hf : _GEN_1135; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1137 = 8'h60 == _T_107[7:0] ? 4'h0 : _GEN_1136; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1138 = 8'h61 == _T_107[7:0] ? 4'h0 : _GEN_1137; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1139 = 8'h62 == _T_107[7:0] ? 4'h0 : _GEN_1138; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1140 = 8'h63 == _T_107[7:0] ? 4'h0 : _GEN_1139; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1141 = 8'h64 == _T_107[7:0] ? 4'h0 : _GEN_1140; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1142 = 8'h65 == _T_107[7:0] ? 4'h0 : _GEN_1141; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1143 = 8'h66 == _T_107[7:0] ? 4'h0 : _GEN_1142; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1144 = 8'h67 == _T_107[7:0] ? 4'h0 : _GEN_1143; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1145 = 8'h68 == _T_107[7:0] ? 4'hf : _GEN_1144; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1146 = 8'h69 == _T_107[7:0] ? 4'hf : _GEN_1145; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1147 = 8'h6a == _T_107[7:0] ? 4'hf : _GEN_1146; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1148 = 8'h6b == _T_107[7:0] ? 4'hf : _GEN_1147; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1149 = 8'h6c == _T_107[7:0] ? 4'hf : _GEN_1148; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1150 = 8'h6d == _T_107[7:0] ? 4'hf : _GEN_1149; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1151 = 8'h6e == _T_107[7:0] ? 4'hf : _GEN_1150; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1152 = 8'h6f == _T_107[7:0] ? 4'hf : _GEN_1151; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1153 = 8'h70 == _T_107[7:0] ? 4'h0 : _GEN_1152; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1154 = 8'h71 == _T_107[7:0] ? 4'h0 : _GEN_1153; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1155 = 8'h72 == _T_107[7:0] ? 4'h0 : _GEN_1154; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1156 = 8'h73 == _T_107[7:0] ? 4'h0 : _GEN_1155; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1157 = 8'h74 == _T_107[7:0] ? 4'h0 : _GEN_1156; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1158 = 8'h75 == _T_107[7:0] ? 4'h0 : _GEN_1157; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1159 = 8'h76 == _T_107[7:0] ? 4'h0 : _GEN_1158; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1160 = 8'h77 == _T_107[7:0] ? 4'h0 : _GEN_1159; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1161 = 8'h78 == _T_107[7:0] ? 4'hf : _GEN_1160; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1162 = 8'h79 == _T_107[7:0] ? 4'hf : _GEN_1161; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1163 = 8'h7a == _T_107[7:0] ? 4'hf : _GEN_1162; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1164 = 8'h7b == _T_107[7:0] ? 4'hf : _GEN_1163; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1165 = 8'h7c == _T_107[7:0] ? 4'hf : _GEN_1164; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1166 = 8'h7d == _T_107[7:0] ? 4'hf : _GEN_1165; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1167 = 8'h7e == _T_107[7:0] ? 4'hf : _GEN_1166; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1168 = 8'h7f == _T_107[7:0] ? 4'hf : _GEN_1167; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1169 = 8'h80 == _T_107[7:0] ? 4'h0 : _GEN_1168; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1170 = 8'h81 == _T_107[7:0] ? 4'h0 : _GEN_1169; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1171 = 8'h82 == _T_107[7:0] ? 4'h0 : _GEN_1170; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1172 = 8'h83 == _T_107[7:0] ? 4'h0 : _GEN_1171; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1173 = 8'h84 == _T_107[7:0] ? 4'h0 : _GEN_1172; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1174 = 8'h85 == _T_107[7:0] ? 4'h0 : _GEN_1173; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1175 = 8'h86 == _T_107[7:0] ? 4'h0 : _GEN_1174; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1176 = 8'h87 == _T_107[7:0] ? 4'h0 : _GEN_1175; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1177 = 8'h88 == _T_107[7:0] ? 4'hf : _GEN_1176; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1178 = 8'h89 == _T_107[7:0] ? 4'hf : _GEN_1177; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1179 = 8'h8a == _T_107[7:0] ? 4'hf : _GEN_1178; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1180 = 8'h8b == _T_107[7:0] ? 4'hf : _GEN_1179; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1181 = 8'h8c == _T_107[7:0] ? 4'hf : _GEN_1180; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1182 = 8'h8d == _T_107[7:0] ? 4'hf : _GEN_1181; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1183 = 8'h8e == _T_107[7:0] ? 4'hf : _GEN_1182; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1184 = 8'h8f == _T_107[7:0] ? 4'hf : _GEN_1183; // @[Filter.scala 196:62]
  wire [4:0] _GEN_7574 = {{1'd0}, _GEN_1184}; // @[Filter.scala 196:62]
  wire [8:0] _T_109 = _GEN_7574 * 5'h14; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1249 = 8'h40 == _T_107[7:0] ? 4'hf : 4'h0; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1250 = 8'h41 == _T_107[7:0] ? 4'hf : _GEN_1249; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1251 = 8'h42 == _T_107[7:0] ? 4'hf : _GEN_1250; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1252 = 8'h43 == _T_107[7:0] ? 4'hf : _GEN_1251; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1253 = 8'h44 == _T_107[7:0] ? 4'hf : _GEN_1252; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1254 = 8'h45 == _T_107[7:0] ? 4'hf : _GEN_1253; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1255 = 8'h46 == _T_107[7:0] ? 4'hf : _GEN_1254; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1256 = 8'h47 == _T_107[7:0] ? 4'hf : _GEN_1255; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1257 = 8'h48 == _T_107[7:0] ? 4'hf : _GEN_1256; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1258 = 8'h49 == _T_107[7:0] ? 4'hf : _GEN_1257; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1259 = 8'h4a == _T_107[7:0] ? 4'hf : _GEN_1258; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1260 = 8'h4b == _T_107[7:0] ? 4'hf : _GEN_1259; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1261 = 8'h4c == _T_107[7:0] ? 4'hf : _GEN_1260; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1262 = 8'h4d == _T_107[7:0] ? 4'hf : _GEN_1261; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1263 = 8'h4e == _T_107[7:0] ? 4'hf : _GEN_1262; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1264 = 8'h4f == _T_107[7:0] ? 4'hf : _GEN_1263; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1265 = 8'h50 == _T_107[7:0] ? 4'hf : _GEN_1264; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1266 = 8'h51 == _T_107[7:0] ? 4'hf : _GEN_1265; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1267 = 8'h52 == _T_107[7:0] ? 4'hf : _GEN_1266; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1268 = 8'h53 == _T_107[7:0] ? 4'hf : _GEN_1267; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1269 = 8'h54 == _T_107[7:0] ? 4'hf : _GEN_1268; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1270 = 8'h55 == _T_107[7:0] ? 4'hf : _GEN_1269; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1271 = 8'h56 == _T_107[7:0] ? 4'hf : _GEN_1270; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1272 = 8'h57 == _T_107[7:0] ? 4'hf : _GEN_1271; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1273 = 8'h58 == _T_107[7:0] ? 4'hf : _GEN_1272; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1274 = 8'h59 == _T_107[7:0] ? 4'hf : _GEN_1273; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1275 = 8'h5a == _T_107[7:0] ? 4'hf : _GEN_1274; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1276 = 8'h5b == _T_107[7:0] ? 4'hf : _GEN_1275; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1277 = 8'h5c == _T_107[7:0] ? 4'hf : _GEN_1276; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1278 = 8'h5d == _T_107[7:0] ? 4'hf : _GEN_1277; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1279 = 8'h5e == _T_107[7:0] ? 4'hf : _GEN_1278; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1280 = 8'h5f == _T_107[7:0] ? 4'hf : _GEN_1279; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1281 = 8'h60 == _T_107[7:0] ? 4'hf : _GEN_1280; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1282 = 8'h61 == _T_107[7:0] ? 4'hf : _GEN_1281; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1283 = 8'h62 == _T_107[7:0] ? 4'hf : _GEN_1282; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1284 = 8'h63 == _T_107[7:0] ? 4'hf : _GEN_1283; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1285 = 8'h64 == _T_107[7:0] ? 4'hf : _GEN_1284; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1286 = 8'h65 == _T_107[7:0] ? 4'hf : _GEN_1285; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1287 = 8'h66 == _T_107[7:0] ? 4'hf : _GEN_1286; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1288 = 8'h67 == _T_107[7:0] ? 4'hf : _GEN_1287; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1289 = 8'h68 == _T_107[7:0] ? 4'hf : _GEN_1288; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1290 = 8'h69 == _T_107[7:0] ? 4'hf : _GEN_1289; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1291 = 8'h6a == _T_107[7:0] ? 4'hf : _GEN_1290; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1292 = 8'h6b == _T_107[7:0] ? 4'hf : _GEN_1291; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1293 = 8'h6c == _T_107[7:0] ? 4'hf : _GEN_1292; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1294 = 8'h6d == _T_107[7:0] ? 4'hf : _GEN_1293; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1295 = 8'h6e == _T_107[7:0] ? 4'hf : _GEN_1294; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1296 = 8'h6f == _T_107[7:0] ? 4'hf : _GEN_1295; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1297 = 8'h70 == _T_107[7:0] ? 4'hf : _GEN_1296; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1298 = 8'h71 == _T_107[7:0] ? 4'hf : _GEN_1297; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1299 = 8'h72 == _T_107[7:0] ? 4'hf : _GEN_1298; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1300 = 8'h73 == _T_107[7:0] ? 4'hf : _GEN_1299; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1301 = 8'h74 == _T_107[7:0] ? 4'hf : _GEN_1300; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1302 = 8'h75 == _T_107[7:0] ? 4'hf : _GEN_1301; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1303 = 8'h76 == _T_107[7:0] ? 4'hf : _GEN_1302; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1304 = 8'h77 == _T_107[7:0] ? 4'hf : _GEN_1303; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1305 = 8'h78 == _T_107[7:0] ? 4'hf : _GEN_1304; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1306 = 8'h79 == _T_107[7:0] ? 4'hf : _GEN_1305; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1307 = 8'h7a == _T_107[7:0] ? 4'hf : _GEN_1306; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1308 = 8'h7b == _T_107[7:0] ? 4'hf : _GEN_1307; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1309 = 8'h7c == _T_107[7:0] ? 4'hf : _GEN_1308; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1310 = 8'h7d == _T_107[7:0] ? 4'hf : _GEN_1309; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1311 = 8'h7e == _T_107[7:0] ? 4'hf : _GEN_1310; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1312 = 8'h7f == _T_107[7:0] ? 4'hf : _GEN_1311; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1313 = 8'h80 == _T_107[7:0] ? 4'hf : _GEN_1312; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1314 = 8'h81 == _T_107[7:0] ? 4'hf : _GEN_1313; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1315 = 8'h82 == _T_107[7:0] ? 4'hf : _GEN_1314; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1316 = 8'h83 == _T_107[7:0] ? 4'hf : _GEN_1315; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1317 = 8'h84 == _T_107[7:0] ? 4'hf : _GEN_1316; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1318 = 8'h85 == _T_107[7:0] ? 4'hf : _GEN_1317; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1319 = 8'h86 == _T_107[7:0] ? 4'hf : _GEN_1318; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1320 = 8'h87 == _T_107[7:0] ? 4'hf : _GEN_1319; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1321 = 8'h88 == _T_107[7:0] ? 4'hf : _GEN_1320; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1322 = 8'h89 == _T_107[7:0] ? 4'hf : _GEN_1321; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1323 = 8'h8a == _T_107[7:0] ? 4'hf : _GEN_1322; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1324 = 8'h8b == _T_107[7:0] ? 4'hf : _GEN_1323; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1325 = 8'h8c == _T_107[7:0] ? 4'hf : _GEN_1324; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1326 = 8'h8d == _T_107[7:0] ? 4'hf : _GEN_1325; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1327 = 8'h8e == _T_107[7:0] ? 4'hf : _GEN_1326; // @[Filter.scala 196:102]
  wire [3:0] _GEN_1328 = 8'h8f == _T_107[7:0] ? 4'hf : _GEN_1327; // @[Filter.scala 196:102]
  wire [6:0] _GEN_7576 = {{3'd0}, _GEN_1328}; // @[Filter.scala 196:102]
  wire [10:0] _T_114 = _GEN_7576 * 7'h46; // @[Filter.scala 196:102]
  wire [10:0] _GEN_7577 = {{2'd0}, _T_109}; // @[Filter.scala 196:69]
  wire [10:0] _T_116 = _GEN_7577 + _T_114; // @[Filter.scala 196:69]
  wire [3:0] _GEN_1337 = 8'h8 == _T_107[7:0] ? 4'hf : 4'h0; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1338 = 8'h9 == _T_107[7:0] ? 4'hf : _GEN_1337; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1339 = 8'ha == _T_107[7:0] ? 4'hf : _GEN_1338; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1340 = 8'hb == _T_107[7:0] ? 4'hf : _GEN_1339; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1341 = 8'hc == _T_107[7:0] ? 4'hf : _GEN_1340; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1342 = 8'hd == _T_107[7:0] ? 4'hf : _GEN_1341; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1343 = 8'he == _T_107[7:0] ? 4'hf : _GEN_1342; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1344 = 8'hf == _T_107[7:0] ? 4'hf : _GEN_1343; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1345 = 8'h10 == _T_107[7:0] ? 4'h0 : _GEN_1344; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1346 = 8'h11 == _T_107[7:0] ? 4'h0 : _GEN_1345; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1347 = 8'h12 == _T_107[7:0] ? 4'h0 : _GEN_1346; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1348 = 8'h13 == _T_107[7:0] ? 4'h0 : _GEN_1347; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1349 = 8'h14 == _T_107[7:0] ? 4'h0 : _GEN_1348; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1350 = 8'h15 == _T_107[7:0] ? 4'h0 : _GEN_1349; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1351 = 8'h16 == _T_107[7:0] ? 4'h0 : _GEN_1350; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1352 = 8'h17 == _T_107[7:0] ? 4'h0 : _GEN_1351; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1353 = 8'h18 == _T_107[7:0] ? 4'hf : _GEN_1352; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1354 = 8'h19 == _T_107[7:0] ? 4'hf : _GEN_1353; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1355 = 8'h1a == _T_107[7:0] ? 4'hf : _GEN_1354; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1356 = 8'h1b == _T_107[7:0] ? 4'hf : _GEN_1355; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1357 = 8'h1c == _T_107[7:0] ? 4'hf : _GEN_1356; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1358 = 8'h1d == _T_107[7:0] ? 4'hf : _GEN_1357; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1359 = 8'h1e == _T_107[7:0] ? 4'hf : _GEN_1358; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1360 = 8'h1f == _T_107[7:0] ? 4'hf : _GEN_1359; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1361 = 8'h20 == _T_107[7:0] ? 4'h0 : _GEN_1360; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1362 = 8'h21 == _T_107[7:0] ? 4'h0 : _GEN_1361; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1363 = 8'h22 == _T_107[7:0] ? 4'h0 : _GEN_1362; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1364 = 8'h23 == _T_107[7:0] ? 4'h0 : _GEN_1363; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1365 = 8'h24 == _T_107[7:0] ? 4'h0 : _GEN_1364; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1366 = 8'h25 == _T_107[7:0] ? 4'h0 : _GEN_1365; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1367 = 8'h26 == _T_107[7:0] ? 4'h0 : _GEN_1366; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1368 = 8'h27 == _T_107[7:0] ? 4'h0 : _GEN_1367; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1369 = 8'h28 == _T_107[7:0] ? 4'hf : _GEN_1368; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1370 = 8'h29 == _T_107[7:0] ? 4'hf : _GEN_1369; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1371 = 8'h2a == _T_107[7:0] ? 4'hf : _GEN_1370; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1372 = 8'h2b == _T_107[7:0] ? 4'hf : _GEN_1371; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1373 = 8'h2c == _T_107[7:0] ? 4'hf : _GEN_1372; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1374 = 8'h2d == _T_107[7:0] ? 4'hf : _GEN_1373; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1375 = 8'h2e == _T_107[7:0] ? 4'hf : _GEN_1374; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1376 = 8'h2f == _T_107[7:0] ? 4'hf : _GEN_1375; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1377 = 8'h30 == _T_107[7:0] ? 4'h0 : _GEN_1376; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1378 = 8'h31 == _T_107[7:0] ? 4'h0 : _GEN_1377; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1379 = 8'h32 == _T_107[7:0] ? 4'h0 : _GEN_1378; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1380 = 8'h33 == _T_107[7:0] ? 4'h0 : _GEN_1379; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1381 = 8'h34 == _T_107[7:0] ? 4'h0 : _GEN_1380; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1382 = 8'h35 == _T_107[7:0] ? 4'h0 : _GEN_1381; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1383 = 8'h36 == _T_107[7:0] ? 4'h0 : _GEN_1382; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1384 = 8'h37 == _T_107[7:0] ? 4'h0 : _GEN_1383; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1385 = 8'h38 == _T_107[7:0] ? 4'hf : _GEN_1384; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1386 = 8'h39 == _T_107[7:0] ? 4'hf : _GEN_1385; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1387 = 8'h3a == _T_107[7:0] ? 4'hf : _GEN_1386; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1388 = 8'h3b == _T_107[7:0] ? 4'hf : _GEN_1387; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1389 = 8'h3c == _T_107[7:0] ? 4'hf : _GEN_1388; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1390 = 8'h3d == _T_107[7:0] ? 4'hf : _GEN_1389; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1391 = 8'h3e == _T_107[7:0] ? 4'hf : _GEN_1390; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1392 = 8'h3f == _T_107[7:0] ? 4'hf : _GEN_1391; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1393 = 8'h40 == _T_107[7:0] ? 4'h0 : _GEN_1392; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1394 = 8'h41 == _T_107[7:0] ? 4'h0 : _GEN_1393; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1395 = 8'h42 == _T_107[7:0] ? 4'h0 : _GEN_1394; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1396 = 8'h43 == _T_107[7:0] ? 4'h0 : _GEN_1395; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1397 = 8'h44 == _T_107[7:0] ? 4'h0 : _GEN_1396; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1398 = 8'h45 == _T_107[7:0] ? 4'h0 : _GEN_1397; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1399 = 8'h46 == _T_107[7:0] ? 4'h0 : _GEN_1398; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1400 = 8'h47 == _T_107[7:0] ? 4'h0 : _GEN_1399; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1401 = 8'h48 == _T_107[7:0] ? 4'hf : _GEN_1400; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1402 = 8'h49 == _T_107[7:0] ? 4'hf : _GEN_1401; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1403 = 8'h4a == _T_107[7:0] ? 4'hf : _GEN_1402; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1404 = 8'h4b == _T_107[7:0] ? 4'hf : _GEN_1403; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1405 = 8'h4c == _T_107[7:0] ? 4'hf : _GEN_1404; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1406 = 8'h4d == _T_107[7:0] ? 4'hf : _GEN_1405; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1407 = 8'h4e == _T_107[7:0] ? 4'hf : _GEN_1406; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1408 = 8'h4f == _T_107[7:0] ? 4'hf : _GEN_1407; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1409 = 8'h50 == _T_107[7:0] ? 4'h0 : _GEN_1408; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1410 = 8'h51 == _T_107[7:0] ? 4'h0 : _GEN_1409; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1411 = 8'h52 == _T_107[7:0] ? 4'h0 : _GEN_1410; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1412 = 8'h53 == _T_107[7:0] ? 4'h0 : _GEN_1411; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1413 = 8'h54 == _T_107[7:0] ? 4'h0 : _GEN_1412; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1414 = 8'h55 == _T_107[7:0] ? 4'h0 : _GEN_1413; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1415 = 8'h56 == _T_107[7:0] ? 4'h0 : _GEN_1414; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1416 = 8'h57 == _T_107[7:0] ? 4'h0 : _GEN_1415; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1417 = 8'h58 == _T_107[7:0] ? 4'hf : _GEN_1416; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1418 = 8'h59 == _T_107[7:0] ? 4'hf : _GEN_1417; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1419 = 8'h5a == _T_107[7:0] ? 4'hf : _GEN_1418; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1420 = 8'h5b == _T_107[7:0] ? 4'hf : _GEN_1419; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1421 = 8'h5c == _T_107[7:0] ? 4'hf : _GEN_1420; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1422 = 8'h5d == _T_107[7:0] ? 4'hf : _GEN_1421; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1423 = 8'h5e == _T_107[7:0] ? 4'hf : _GEN_1422; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1424 = 8'h5f == _T_107[7:0] ? 4'hf : _GEN_1423; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1425 = 8'h60 == _T_107[7:0] ? 4'h0 : _GEN_1424; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1426 = 8'h61 == _T_107[7:0] ? 4'h0 : _GEN_1425; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1427 = 8'h62 == _T_107[7:0] ? 4'h0 : _GEN_1426; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1428 = 8'h63 == _T_107[7:0] ? 4'h0 : _GEN_1427; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1429 = 8'h64 == _T_107[7:0] ? 4'h0 : _GEN_1428; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1430 = 8'h65 == _T_107[7:0] ? 4'h0 : _GEN_1429; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1431 = 8'h66 == _T_107[7:0] ? 4'h0 : _GEN_1430; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1432 = 8'h67 == _T_107[7:0] ? 4'h0 : _GEN_1431; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1433 = 8'h68 == _T_107[7:0] ? 4'hf : _GEN_1432; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1434 = 8'h69 == _T_107[7:0] ? 4'hf : _GEN_1433; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1435 = 8'h6a == _T_107[7:0] ? 4'hf : _GEN_1434; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1436 = 8'h6b == _T_107[7:0] ? 4'hf : _GEN_1435; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1437 = 8'h6c == _T_107[7:0] ? 4'hf : _GEN_1436; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1438 = 8'h6d == _T_107[7:0] ? 4'hf : _GEN_1437; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1439 = 8'h6e == _T_107[7:0] ? 4'hf : _GEN_1438; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1440 = 8'h6f == _T_107[7:0] ? 4'hf : _GEN_1439; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1441 = 8'h70 == _T_107[7:0] ? 4'h0 : _GEN_1440; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1442 = 8'h71 == _T_107[7:0] ? 4'h0 : _GEN_1441; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1443 = 8'h72 == _T_107[7:0] ? 4'h0 : _GEN_1442; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1444 = 8'h73 == _T_107[7:0] ? 4'h0 : _GEN_1443; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1445 = 8'h74 == _T_107[7:0] ? 4'h0 : _GEN_1444; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1446 = 8'h75 == _T_107[7:0] ? 4'h0 : _GEN_1445; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1447 = 8'h76 == _T_107[7:0] ? 4'h0 : _GEN_1446; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1448 = 8'h77 == _T_107[7:0] ? 4'h0 : _GEN_1447; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1449 = 8'h78 == _T_107[7:0] ? 4'hf : _GEN_1448; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1450 = 8'h79 == _T_107[7:0] ? 4'hf : _GEN_1449; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1451 = 8'h7a == _T_107[7:0] ? 4'hf : _GEN_1450; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1452 = 8'h7b == _T_107[7:0] ? 4'hf : _GEN_1451; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1453 = 8'h7c == _T_107[7:0] ? 4'hf : _GEN_1452; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1454 = 8'h7d == _T_107[7:0] ? 4'hf : _GEN_1453; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1455 = 8'h7e == _T_107[7:0] ? 4'hf : _GEN_1454; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1456 = 8'h7f == _T_107[7:0] ? 4'hf : _GEN_1455; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1457 = 8'h80 == _T_107[7:0] ? 4'h0 : _GEN_1456; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1458 = 8'h81 == _T_107[7:0] ? 4'h0 : _GEN_1457; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1459 = 8'h82 == _T_107[7:0] ? 4'h0 : _GEN_1458; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1460 = 8'h83 == _T_107[7:0] ? 4'h0 : _GEN_1459; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1461 = 8'h84 == _T_107[7:0] ? 4'h0 : _GEN_1460; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1462 = 8'h85 == _T_107[7:0] ? 4'h0 : _GEN_1461; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1463 = 8'h86 == _T_107[7:0] ? 4'h0 : _GEN_1462; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1464 = 8'h87 == _T_107[7:0] ? 4'h0 : _GEN_1463; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1465 = 8'h88 == _T_107[7:0] ? 4'hf : _GEN_1464; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1466 = 8'h89 == _T_107[7:0] ? 4'hf : _GEN_1465; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1467 = 8'h8a == _T_107[7:0] ? 4'hf : _GEN_1466; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1468 = 8'h8b == _T_107[7:0] ? 4'hf : _GEN_1467; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1469 = 8'h8c == _T_107[7:0] ? 4'hf : _GEN_1468; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1470 = 8'h8d == _T_107[7:0] ? 4'hf : _GEN_1469; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1471 = 8'h8e == _T_107[7:0] ? 4'hf : _GEN_1470; // @[Filter.scala 196:142]
  wire [3:0] _GEN_1472 = 8'h8f == _T_107[7:0] ? 4'hf : _GEN_1471; // @[Filter.scala 196:142]
  wire [7:0] _T_121 = _GEN_1472 * 4'ha; // @[Filter.scala 196:142]
  wire [10:0] _GEN_7579 = {{3'd0}, _T_121}; // @[Filter.scala 196:109]
  wire [10:0] _T_123 = _T_116 + _GEN_7579; // @[Filter.scala 196:109]
  wire [10:0] _T_124 = _T_123 / 11'h64; // @[Filter.scala 196:150]
  wire  _T_126 = _T_97 >= 5'h10; // @[Filter.scala 199:31]
  wire  _T_130 = _T_104 >= 32'h9; // @[Filter.scala 199:63]
  wire  _T_131 = _T_126 | _T_130; // @[Filter.scala 199:58]
  wire [10:0] _GEN_1617 = io_SPI_distort ? _T_124 : {{7'd0}, _GEN_1184}; // @[Filter.scala 201:35]
  wire [10:0] _GEN_1618 = _T_131 ? 11'h0 : _GEN_1617; // @[Filter.scala 199:80]
  wire [10:0] _GEN_1763 = io_SPI_distort ? _T_124 : {{7'd0}, _GEN_1328}; // @[Filter.scala 201:35]
  wire [10:0] _GEN_1764 = _T_131 ? 11'h0 : _GEN_1763; // @[Filter.scala 199:80]
  wire [10:0] _GEN_1909 = io_SPI_distort ? _T_124 : {{7'd0}, _GEN_1472}; // @[Filter.scala 201:35]
  wire [10:0] _GEN_1910 = _T_131 ? 11'h0 : _GEN_1909; // @[Filter.scala 199:80]
  wire [31:0] _T_159 = pixelIndex + 32'h2; // @[Filter.scala 194:31]
  wire [31:0] _GEN_2 = _T_159 % 32'h10; // @[Filter.scala 194:38]
  wire [4:0] _T_160 = _GEN_2[4:0]; // @[Filter.scala 194:38]
  wire [4:0] _T_162 = _T_160 + _GEN_7559; // @[Filter.scala 194:53]
  wire [4:0] _T_164 = _T_162 - 5'h1; // @[Filter.scala 194:69]
  wire [31:0] _T_167 = _T_159 / 32'h10; // @[Filter.scala 195:38]
  wire [31:0] _T_169 = _T_167 + _GEN_7560; // @[Filter.scala 195:53]
  wire [31:0] _T_171 = _T_169 - 32'h1; // @[Filter.scala 195:69]
  wire [36:0] _T_172 = _T_171 * 32'h10; // @[Filter.scala 196:42]
  wire [36:0] _GEN_7585 = {{32'd0}, _T_164}; // @[Filter.scala 196:57]
  wire [36:0] _T_174 = _T_172 + _GEN_7585; // @[Filter.scala 196:57]
  wire [3:0] _GEN_1919 = 8'h8 == _T_174[7:0] ? 4'h0 : 4'hf; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1920 = 8'h9 == _T_174[7:0] ? 4'h0 : _GEN_1919; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1921 = 8'ha == _T_174[7:0] ? 4'h0 : _GEN_1920; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1922 = 8'hb == _T_174[7:0] ? 4'h0 : _GEN_1921; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1923 = 8'hc == _T_174[7:0] ? 4'h0 : _GEN_1922; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1924 = 8'hd == _T_174[7:0] ? 4'h0 : _GEN_1923; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1925 = 8'he == _T_174[7:0] ? 4'h0 : _GEN_1924; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1926 = 8'hf == _T_174[7:0] ? 4'h0 : _GEN_1925; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1927 = 8'h10 == _T_174[7:0] ? 4'hf : _GEN_1926; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1928 = 8'h11 == _T_174[7:0] ? 4'hf : _GEN_1927; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1929 = 8'h12 == _T_174[7:0] ? 4'hf : _GEN_1928; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1930 = 8'h13 == _T_174[7:0] ? 4'hf : _GEN_1929; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1931 = 8'h14 == _T_174[7:0] ? 4'hf : _GEN_1930; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1932 = 8'h15 == _T_174[7:0] ? 4'hf : _GEN_1931; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1933 = 8'h16 == _T_174[7:0] ? 4'hf : _GEN_1932; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1934 = 8'h17 == _T_174[7:0] ? 4'hf : _GEN_1933; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1935 = 8'h18 == _T_174[7:0] ? 4'h0 : _GEN_1934; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1936 = 8'h19 == _T_174[7:0] ? 4'h0 : _GEN_1935; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1937 = 8'h1a == _T_174[7:0] ? 4'h0 : _GEN_1936; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1938 = 8'h1b == _T_174[7:0] ? 4'h0 : _GEN_1937; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1939 = 8'h1c == _T_174[7:0] ? 4'h0 : _GEN_1938; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1940 = 8'h1d == _T_174[7:0] ? 4'h0 : _GEN_1939; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1941 = 8'h1e == _T_174[7:0] ? 4'h0 : _GEN_1940; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1942 = 8'h1f == _T_174[7:0] ? 4'h0 : _GEN_1941; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1943 = 8'h20 == _T_174[7:0] ? 4'hf : _GEN_1942; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1944 = 8'h21 == _T_174[7:0] ? 4'hf : _GEN_1943; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1945 = 8'h22 == _T_174[7:0] ? 4'hf : _GEN_1944; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1946 = 8'h23 == _T_174[7:0] ? 4'hf : _GEN_1945; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1947 = 8'h24 == _T_174[7:0] ? 4'hf : _GEN_1946; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1948 = 8'h25 == _T_174[7:0] ? 4'hf : _GEN_1947; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1949 = 8'h26 == _T_174[7:0] ? 4'hf : _GEN_1948; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1950 = 8'h27 == _T_174[7:0] ? 4'hf : _GEN_1949; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1951 = 8'h28 == _T_174[7:0] ? 4'h0 : _GEN_1950; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1952 = 8'h29 == _T_174[7:0] ? 4'h0 : _GEN_1951; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1953 = 8'h2a == _T_174[7:0] ? 4'h0 : _GEN_1952; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1954 = 8'h2b == _T_174[7:0] ? 4'h0 : _GEN_1953; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1955 = 8'h2c == _T_174[7:0] ? 4'h0 : _GEN_1954; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1956 = 8'h2d == _T_174[7:0] ? 4'h0 : _GEN_1955; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1957 = 8'h2e == _T_174[7:0] ? 4'h0 : _GEN_1956; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1958 = 8'h2f == _T_174[7:0] ? 4'h0 : _GEN_1957; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1959 = 8'h30 == _T_174[7:0] ? 4'hf : _GEN_1958; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1960 = 8'h31 == _T_174[7:0] ? 4'hf : _GEN_1959; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1961 = 8'h32 == _T_174[7:0] ? 4'hf : _GEN_1960; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1962 = 8'h33 == _T_174[7:0] ? 4'hf : _GEN_1961; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1963 = 8'h34 == _T_174[7:0] ? 4'hf : _GEN_1962; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1964 = 8'h35 == _T_174[7:0] ? 4'hf : _GEN_1963; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1965 = 8'h36 == _T_174[7:0] ? 4'hf : _GEN_1964; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1966 = 8'h37 == _T_174[7:0] ? 4'hf : _GEN_1965; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1967 = 8'h38 == _T_174[7:0] ? 4'h0 : _GEN_1966; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1968 = 8'h39 == _T_174[7:0] ? 4'h0 : _GEN_1967; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1969 = 8'h3a == _T_174[7:0] ? 4'h0 : _GEN_1968; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1970 = 8'h3b == _T_174[7:0] ? 4'h0 : _GEN_1969; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1971 = 8'h3c == _T_174[7:0] ? 4'h0 : _GEN_1970; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1972 = 8'h3d == _T_174[7:0] ? 4'h0 : _GEN_1971; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1973 = 8'h3e == _T_174[7:0] ? 4'h0 : _GEN_1972; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1974 = 8'h3f == _T_174[7:0] ? 4'h0 : _GEN_1973; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1975 = 8'h40 == _T_174[7:0] ? 4'h0 : _GEN_1974; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1976 = 8'h41 == _T_174[7:0] ? 4'h0 : _GEN_1975; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1977 = 8'h42 == _T_174[7:0] ? 4'h0 : _GEN_1976; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1978 = 8'h43 == _T_174[7:0] ? 4'h0 : _GEN_1977; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1979 = 8'h44 == _T_174[7:0] ? 4'h0 : _GEN_1978; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1980 = 8'h45 == _T_174[7:0] ? 4'h0 : _GEN_1979; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1981 = 8'h46 == _T_174[7:0] ? 4'h0 : _GEN_1980; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1982 = 8'h47 == _T_174[7:0] ? 4'h0 : _GEN_1981; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1983 = 8'h48 == _T_174[7:0] ? 4'hf : _GEN_1982; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1984 = 8'h49 == _T_174[7:0] ? 4'hf : _GEN_1983; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1985 = 8'h4a == _T_174[7:0] ? 4'hf : _GEN_1984; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1986 = 8'h4b == _T_174[7:0] ? 4'hf : _GEN_1985; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1987 = 8'h4c == _T_174[7:0] ? 4'hf : _GEN_1986; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1988 = 8'h4d == _T_174[7:0] ? 4'hf : _GEN_1987; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1989 = 8'h4e == _T_174[7:0] ? 4'hf : _GEN_1988; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1990 = 8'h4f == _T_174[7:0] ? 4'hf : _GEN_1989; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1991 = 8'h50 == _T_174[7:0] ? 4'h0 : _GEN_1990; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1992 = 8'h51 == _T_174[7:0] ? 4'h0 : _GEN_1991; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1993 = 8'h52 == _T_174[7:0] ? 4'h0 : _GEN_1992; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1994 = 8'h53 == _T_174[7:0] ? 4'h0 : _GEN_1993; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1995 = 8'h54 == _T_174[7:0] ? 4'h0 : _GEN_1994; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1996 = 8'h55 == _T_174[7:0] ? 4'h0 : _GEN_1995; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1997 = 8'h56 == _T_174[7:0] ? 4'h0 : _GEN_1996; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1998 = 8'h57 == _T_174[7:0] ? 4'h0 : _GEN_1997; // @[Filter.scala 196:62]
  wire [3:0] _GEN_1999 = 8'h58 == _T_174[7:0] ? 4'hf : _GEN_1998; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2000 = 8'h59 == _T_174[7:0] ? 4'hf : _GEN_1999; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2001 = 8'h5a == _T_174[7:0] ? 4'hf : _GEN_2000; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2002 = 8'h5b == _T_174[7:0] ? 4'hf : _GEN_2001; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2003 = 8'h5c == _T_174[7:0] ? 4'hf : _GEN_2002; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2004 = 8'h5d == _T_174[7:0] ? 4'hf : _GEN_2003; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2005 = 8'h5e == _T_174[7:0] ? 4'hf : _GEN_2004; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2006 = 8'h5f == _T_174[7:0] ? 4'hf : _GEN_2005; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2007 = 8'h60 == _T_174[7:0] ? 4'h0 : _GEN_2006; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2008 = 8'h61 == _T_174[7:0] ? 4'h0 : _GEN_2007; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2009 = 8'h62 == _T_174[7:0] ? 4'h0 : _GEN_2008; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2010 = 8'h63 == _T_174[7:0] ? 4'h0 : _GEN_2009; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2011 = 8'h64 == _T_174[7:0] ? 4'h0 : _GEN_2010; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2012 = 8'h65 == _T_174[7:0] ? 4'h0 : _GEN_2011; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2013 = 8'h66 == _T_174[7:0] ? 4'h0 : _GEN_2012; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2014 = 8'h67 == _T_174[7:0] ? 4'h0 : _GEN_2013; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2015 = 8'h68 == _T_174[7:0] ? 4'hf : _GEN_2014; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2016 = 8'h69 == _T_174[7:0] ? 4'hf : _GEN_2015; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2017 = 8'h6a == _T_174[7:0] ? 4'hf : _GEN_2016; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2018 = 8'h6b == _T_174[7:0] ? 4'hf : _GEN_2017; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2019 = 8'h6c == _T_174[7:0] ? 4'hf : _GEN_2018; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2020 = 8'h6d == _T_174[7:0] ? 4'hf : _GEN_2019; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2021 = 8'h6e == _T_174[7:0] ? 4'hf : _GEN_2020; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2022 = 8'h6f == _T_174[7:0] ? 4'hf : _GEN_2021; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2023 = 8'h70 == _T_174[7:0] ? 4'h0 : _GEN_2022; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2024 = 8'h71 == _T_174[7:0] ? 4'h0 : _GEN_2023; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2025 = 8'h72 == _T_174[7:0] ? 4'h0 : _GEN_2024; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2026 = 8'h73 == _T_174[7:0] ? 4'h0 : _GEN_2025; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2027 = 8'h74 == _T_174[7:0] ? 4'h0 : _GEN_2026; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2028 = 8'h75 == _T_174[7:0] ? 4'h0 : _GEN_2027; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2029 = 8'h76 == _T_174[7:0] ? 4'h0 : _GEN_2028; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2030 = 8'h77 == _T_174[7:0] ? 4'h0 : _GEN_2029; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2031 = 8'h78 == _T_174[7:0] ? 4'hf : _GEN_2030; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2032 = 8'h79 == _T_174[7:0] ? 4'hf : _GEN_2031; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2033 = 8'h7a == _T_174[7:0] ? 4'hf : _GEN_2032; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2034 = 8'h7b == _T_174[7:0] ? 4'hf : _GEN_2033; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2035 = 8'h7c == _T_174[7:0] ? 4'hf : _GEN_2034; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2036 = 8'h7d == _T_174[7:0] ? 4'hf : _GEN_2035; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2037 = 8'h7e == _T_174[7:0] ? 4'hf : _GEN_2036; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2038 = 8'h7f == _T_174[7:0] ? 4'hf : _GEN_2037; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2039 = 8'h80 == _T_174[7:0] ? 4'h0 : _GEN_2038; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2040 = 8'h81 == _T_174[7:0] ? 4'h0 : _GEN_2039; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2041 = 8'h82 == _T_174[7:0] ? 4'h0 : _GEN_2040; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2042 = 8'h83 == _T_174[7:0] ? 4'h0 : _GEN_2041; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2043 = 8'h84 == _T_174[7:0] ? 4'h0 : _GEN_2042; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2044 = 8'h85 == _T_174[7:0] ? 4'h0 : _GEN_2043; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2045 = 8'h86 == _T_174[7:0] ? 4'h0 : _GEN_2044; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2046 = 8'h87 == _T_174[7:0] ? 4'h0 : _GEN_2045; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2047 = 8'h88 == _T_174[7:0] ? 4'hf : _GEN_2046; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2048 = 8'h89 == _T_174[7:0] ? 4'hf : _GEN_2047; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2049 = 8'h8a == _T_174[7:0] ? 4'hf : _GEN_2048; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2050 = 8'h8b == _T_174[7:0] ? 4'hf : _GEN_2049; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2051 = 8'h8c == _T_174[7:0] ? 4'hf : _GEN_2050; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2052 = 8'h8d == _T_174[7:0] ? 4'hf : _GEN_2051; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2053 = 8'h8e == _T_174[7:0] ? 4'hf : _GEN_2052; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2054 = 8'h8f == _T_174[7:0] ? 4'hf : _GEN_2053; // @[Filter.scala 196:62]
  wire [4:0] _GEN_7586 = {{1'd0}, _GEN_2054}; // @[Filter.scala 196:62]
  wire [8:0] _T_176 = _GEN_7586 * 5'h14; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2119 = 8'h40 == _T_174[7:0] ? 4'hf : 4'h0; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2120 = 8'h41 == _T_174[7:0] ? 4'hf : _GEN_2119; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2121 = 8'h42 == _T_174[7:0] ? 4'hf : _GEN_2120; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2122 = 8'h43 == _T_174[7:0] ? 4'hf : _GEN_2121; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2123 = 8'h44 == _T_174[7:0] ? 4'hf : _GEN_2122; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2124 = 8'h45 == _T_174[7:0] ? 4'hf : _GEN_2123; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2125 = 8'h46 == _T_174[7:0] ? 4'hf : _GEN_2124; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2126 = 8'h47 == _T_174[7:0] ? 4'hf : _GEN_2125; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2127 = 8'h48 == _T_174[7:0] ? 4'hf : _GEN_2126; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2128 = 8'h49 == _T_174[7:0] ? 4'hf : _GEN_2127; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2129 = 8'h4a == _T_174[7:0] ? 4'hf : _GEN_2128; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2130 = 8'h4b == _T_174[7:0] ? 4'hf : _GEN_2129; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2131 = 8'h4c == _T_174[7:0] ? 4'hf : _GEN_2130; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2132 = 8'h4d == _T_174[7:0] ? 4'hf : _GEN_2131; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2133 = 8'h4e == _T_174[7:0] ? 4'hf : _GEN_2132; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2134 = 8'h4f == _T_174[7:0] ? 4'hf : _GEN_2133; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2135 = 8'h50 == _T_174[7:0] ? 4'hf : _GEN_2134; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2136 = 8'h51 == _T_174[7:0] ? 4'hf : _GEN_2135; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2137 = 8'h52 == _T_174[7:0] ? 4'hf : _GEN_2136; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2138 = 8'h53 == _T_174[7:0] ? 4'hf : _GEN_2137; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2139 = 8'h54 == _T_174[7:0] ? 4'hf : _GEN_2138; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2140 = 8'h55 == _T_174[7:0] ? 4'hf : _GEN_2139; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2141 = 8'h56 == _T_174[7:0] ? 4'hf : _GEN_2140; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2142 = 8'h57 == _T_174[7:0] ? 4'hf : _GEN_2141; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2143 = 8'h58 == _T_174[7:0] ? 4'hf : _GEN_2142; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2144 = 8'h59 == _T_174[7:0] ? 4'hf : _GEN_2143; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2145 = 8'h5a == _T_174[7:0] ? 4'hf : _GEN_2144; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2146 = 8'h5b == _T_174[7:0] ? 4'hf : _GEN_2145; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2147 = 8'h5c == _T_174[7:0] ? 4'hf : _GEN_2146; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2148 = 8'h5d == _T_174[7:0] ? 4'hf : _GEN_2147; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2149 = 8'h5e == _T_174[7:0] ? 4'hf : _GEN_2148; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2150 = 8'h5f == _T_174[7:0] ? 4'hf : _GEN_2149; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2151 = 8'h60 == _T_174[7:0] ? 4'hf : _GEN_2150; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2152 = 8'h61 == _T_174[7:0] ? 4'hf : _GEN_2151; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2153 = 8'h62 == _T_174[7:0] ? 4'hf : _GEN_2152; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2154 = 8'h63 == _T_174[7:0] ? 4'hf : _GEN_2153; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2155 = 8'h64 == _T_174[7:0] ? 4'hf : _GEN_2154; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2156 = 8'h65 == _T_174[7:0] ? 4'hf : _GEN_2155; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2157 = 8'h66 == _T_174[7:0] ? 4'hf : _GEN_2156; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2158 = 8'h67 == _T_174[7:0] ? 4'hf : _GEN_2157; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2159 = 8'h68 == _T_174[7:0] ? 4'hf : _GEN_2158; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2160 = 8'h69 == _T_174[7:0] ? 4'hf : _GEN_2159; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2161 = 8'h6a == _T_174[7:0] ? 4'hf : _GEN_2160; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2162 = 8'h6b == _T_174[7:0] ? 4'hf : _GEN_2161; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2163 = 8'h6c == _T_174[7:0] ? 4'hf : _GEN_2162; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2164 = 8'h6d == _T_174[7:0] ? 4'hf : _GEN_2163; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2165 = 8'h6e == _T_174[7:0] ? 4'hf : _GEN_2164; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2166 = 8'h6f == _T_174[7:0] ? 4'hf : _GEN_2165; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2167 = 8'h70 == _T_174[7:0] ? 4'hf : _GEN_2166; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2168 = 8'h71 == _T_174[7:0] ? 4'hf : _GEN_2167; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2169 = 8'h72 == _T_174[7:0] ? 4'hf : _GEN_2168; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2170 = 8'h73 == _T_174[7:0] ? 4'hf : _GEN_2169; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2171 = 8'h74 == _T_174[7:0] ? 4'hf : _GEN_2170; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2172 = 8'h75 == _T_174[7:0] ? 4'hf : _GEN_2171; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2173 = 8'h76 == _T_174[7:0] ? 4'hf : _GEN_2172; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2174 = 8'h77 == _T_174[7:0] ? 4'hf : _GEN_2173; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2175 = 8'h78 == _T_174[7:0] ? 4'hf : _GEN_2174; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2176 = 8'h79 == _T_174[7:0] ? 4'hf : _GEN_2175; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2177 = 8'h7a == _T_174[7:0] ? 4'hf : _GEN_2176; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2178 = 8'h7b == _T_174[7:0] ? 4'hf : _GEN_2177; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2179 = 8'h7c == _T_174[7:0] ? 4'hf : _GEN_2178; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2180 = 8'h7d == _T_174[7:0] ? 4'hf : _GEN_2179; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2181 = 8'h7e == _T_174[7:0] ? 4'hf : _GEN_2180; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2182 = 8'h7f == _T_174[7:0] ? 4'hf : _GEN_2181; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2183 = 8'h80 == _T_174[7:0] ? 4'hf : _GEN_2182; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2184 = 8'h81 == _T_174[7:0] ? 4'hf : _GEN_2183; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2185 = 8'h82 == _T_174[7:0] ? 4'hf : _GEN_2184; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2186 = 8'h83 == _T_174[7:0] ? 4'hf : _GEN_2185; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2187 = 8'h84 == _T_174[7:0] ? 4'hf : _GEN_2186; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2188 = 8'h85 == _T_174[7:0] ? 4'hf : _GEN_2187; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2189 = 8'h86 == _T_174[7:0] ? 4'hf : _GEN_2188; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2190 = 8'h87 == _T_174[7:0] ? 4'hf : _GEN_2189; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2191 = 8'h88 == _T_174[7:0] ? 4'hf : _GEN_2190; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2192 = 8'h89 == _T_174[7:0] ? 4'hf : _GEN_2191; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2193 = 8'h8a == _T_174[7:0] ? 4'hf : _GEN_2192; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2194 = 8'h8b == _T_174[7:0] ? 4'hf : _GEN_2193; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2195 = 8'h8c == _T_174[7:0] ? 4'hf : _GEN_2194; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2196 = 8'h8d == _T_174[7:0] ? 4'hf : _GEN_2195; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2197 = 8'h8e == _T_174[7:0] ? 4'hf : _GEN_2196; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2198 = 8'h8f == _T_174[7:0] ? 4'hf : _GEN_2197; // @[Filter.scala 196:102]
  wire [6:0] _GEN_7588 = {{3'd0}, _GEN_2198}; // @[Filter.scala 196:102]
  wire [10:0] _T_181 = _GEN_7588 * 7'h46; // @[Filter.scala 196:102]
  wire [10:0] _GEN_7589 = {{2'd0}, _T_176}; // @[Filter.scala 196:69]
  wire [10:0] _T_183 = _GEN_7589 + _T_181; // @[Filter.scala 196:69]
  wire [3:0] _GEN_2207 = 8'h8 == _T_174[7:0] ? 4'hf : 4'h0; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2208 = 8'h9 == _T_174[7:0] ? 4'hf : _GEN_2207; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2209 = 8'ha == _T_174[7:0] ? 4'hf : _GEN_2208; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2210 = 8'hb == _T_174[7:0] ? 4'hf : _GEN_2209; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2211 = 8'hc == _T_174[7:0] ? 4'hf : _GEN_2210; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2212 = 8'hd == _T_174[7:0] ? 4'hf : _GEN_2211; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2213 = 8'he == _T_174[7:0] ? 4'hf : _GEN_2212; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2214 = 8'hf == _T_174[7:0] ? 4'hf : _GEN_2213; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2215 = 8'h10 == _T_174[7:0] ? 4'h0 : _GEN_2214; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2216 = 8'h11 == _T_174[7:0] ? 4'h0 : _GEN_2215; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2217 = 8'h12 == _T_174[7:0] ? 4'h0 : _GEN_2216; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2218 = 8'h13 == _T_174[7:0] ? 4'h0 : _GEN_2217; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2219 = 8'h14 == _T_174[7:0] ? 4'h0 : _GEN_2218; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2220 = 8'h15 == _T_174[7:0] ? 4'h0 : _GEN_2219; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2221 = 8'h16 == _T_174[7:0] ? 4'h0 : _GEN_2220; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2222 = 8'h17 == _T_174[7:0] ? 4'h0 : _GEN_2221; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2223 = 8'h18 == _T_174[7:0] ? 4'hf : _GEN_2222; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2224 = 8'h19 == _T_174[7:0] ? 4'hf : _GEN_2223; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2225 = 8'h1a == _T_174[7:0] ? 4'hf : _GEN_2224; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2226 = 8'h1b == _T_174[7:0] ? 4'hf : _GEN_2225; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2227 = 8'h1c == _T_174[7:0] ? 4'hf : _GEN_2226; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2228 = 8'h1d == _T_174[7:0] ? 4'hf : _GEN_2227; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2229 = 8'h1e == _T_174[7:0] ? 4'hf : _GEN_2228; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2230 = 8'h1f == _T_174[7:0] ? 4'hf : _GEN_2229; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2231 = 8'h20 == _T_174[7:0] ? 4'h0 : _GEN_2230; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2232 = 8'h21 == _T_174[7:0] ? 4'h0 : _GEN_2231; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2233 = 8'h22 == _T_174[7:0] ? 4'h0 : _GEN_2232; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2234 = 8'h23 == _T_174[7:0] ? 4'h0 : _GEN_2233; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2235 = 8'h24 == _T_174[7:0] ? 4'h0 : _GEN_2234; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2236 = 8'h25 == _T_174[7:0] ? 4'h0 : _GEN_2235; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2237 = 8'h26 == _T_174[7:0] ? 4'h0 : _GEN_2236; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2238 = 8'h27 == _T_174[7:0] ? 4'h0 : _GEN_2237; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2239 = 8'h28 == _T_174[7:0] ? 4'hf : _GEN_2238; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2240 = 8'h29 == _T_174[7:0] ? 4'hf : _GEN_2239; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2241 = 8'h2a == _T_174[7:0] ? 4'hf : _GEN_2240; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2242 = 8'h2b == _T_174[7:0] ? 4'hf : _GEN_2241; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2243 = 8'h2c == _T_174[7:0] ? 4'hf : _GEN_2242; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2244 = 8'h2d == _T_174[7:0] ? 4'hf : _GEN_2243; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2245 = 8'h2e == _T_174[7:0] ? 4'hf : _GEN_2244; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2246 = 8'h2f == _T_174[7:0] ? 4'hf : _GEN_2245; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2247 = 8'h30 == _T_174[7:0] ? 4'h0 : _GEN_2246; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2248 = 8'h31 == _T_174[7:0] ? 4'h0 : _GEN_2247; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2249 = 8'h32 == _T_174[7:0] ? 4'h0 : _GEN_2248; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2250 = 8'h33 == _T_174[7:0] ? 4'h0 : _GEN_2249; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2251 = 8'h34 == _T_174[7:0] ? 4'h0 : _GEN_2250; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2252 = 8'h35 == _T_174[7:0] ? 4'h0 : _GEN_2251; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2253 = 8'h36 == _T_174[7:0] ? 4'h0 : _GEN_2252; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2254 = 8'h37 == _T_174[7:0] ? 4'h0 : _GEN_2253; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2255 = 8'h38 == _T_174[7:0] ? 4'hf : _GEN_2254; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2256 = 8'h39 == _T_174[7:0] ? 4'hf : _GEN_2255; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2257 = 8'h3a == _T_174[7:0] ? 4'hf : _GEN_2256; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2258 = 8'h3b == _T_174[7:0] ? 4'hf : _GEN_2257; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2259 = 8'h3c == _T_174[7:0] ? 4'hf : _GEN_2258; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2260 = 8'h3d == _T_174[7:0] ? 4'hf : _GEN_2259; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2261 = 8'h3e == _T_174[7:0] ? 4'hf : _GEN_2260; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2262 = 8'h3f == _T_174[7:0] ? 4'hf : _GEN_2261; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2263 = 8'h40 == _T_174[7:0] ? 4'h0 : _GEN_2262; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2264 = 8'h41 == _T_174[7:0] ? 4'h0 : _GEN_2263; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2265 = 8'h42 == _T_174[7:0] ? 4'h0 : _GEN_2264; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2266 = 8'h43 == _T_174[7:0] ? 4'h0 : _GEN_2265; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2267 = 8'h44 == _T_174[7:0] ? 4'h0 : _GEN_2266; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2268 = 8'h45 == _T_174[7:0] ? 4'h0 : _GEN_2267; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2269 = 8'h46 == _T_174[7:0] ? 4'h0 : _GEN_2268; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2270 = 8'h47 == _T_174[7:0] ? 4'h0 : _GEN_2269; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2271 = 8'h48 == _T_174[7:0] ? 4'hf : _GEN_2270; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2272 = 8'h49 == _T_174[7:0] ? 4'hf : _GEN_2271; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2273 = 8'h4a == _T_174[7:0] ? 4'hf : _GEN_2272; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2274 = 8'h4b == _T_174[7:0] ? 4'hf : _GEN_2273; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2275 = 8'h4c == _T_174[7:0] ? 4'hf : _GEN_2274; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2276 = 8'h4d == _T_174[7:0] ? 4'hf : _GEN_2275; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2277 = 8'h4e == _T_174[7:0] ? 4'hf : _GEN_2276; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2278 = 8'h4f == _T_174[7:0] ? 4'hf : _GEN_2277; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2279 = 8'h50 == _T_174[7:0] ? 4'h0 : _GEN_2278; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2280 = 8'h51 == _T_174[7:0] ? 4'h0 : _GEN_2279; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2281 = 8'h52 == _T_174[7:0] ? 4'h0 : _GEN_2280; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2282 = 8'h53 == _T_174[7:0] ? 4'h0 : _GEN_2281; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2283 = 8'h54 == _T_174[7:0] ? 4'h0 : _GEN_2282; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2284 = 8'h55 == _T_174[7:0] ? 4'h0 : _GEN_2283; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2285 = 8'h56 == _T_174[7:0] ? 4'h0 : _GEN_2284; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2286 = 8'h57 == _T_174[7:0] ? 4'h0 : _GEN_2285; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2287 = 8'h58 == _T_174[7:0] ? 4'hf : _GEN_2286; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2288 = 8'h59 == _T_174[7:0] ? 4'hf : _GEN_2287; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2289 = 8'h5a == _T_174[7:0] ? 4'hf : _GEN_2288; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2290 = 8'h5b == _T_174[7:0] ? 4'hf : _GEN_2289; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2291 = 8'h5c == _T_174[7:0] ? 4'hf : _GEN_2290; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2292 = 8'h5d == _T_174[7:0] ? 4'hf : _GEN_2291; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2293 = 8'h5e == _T_174[7:0] ? 4'hf : _GEN_2292; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2294 = 8'h5f == _T_174[7:0] ? 4'hf : _GEN_2293; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2295 = 8'h60 == _T_174[7:0] ? 4'h0 : _GEN_2294; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2296 = 8'h61 == _T_174[7:0] ? 4'h0 : _GEN_2295; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2297 = 8'h62 == _T_174[7:0] ? 4'h0 : _GEN_2296; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2298 = 8'h63 == _T_174[7:0] ? 4'h0 : _GEN_2297; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2299 = 8'h64 == _T_174[7:0] ? 4'h0 : _GEN_2298; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2300 = 8'h65 == _T_174[7:0] ? 4'h0 : _GEN_2299; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2301 = 8'h66 == _T_174[7:0] ? 4'h0 : _GEN_2300; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2302 = 8'h67 == _T_174[7:0] ? 4'h0 : _GEN_2301; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2303 = 8'h68 == _T_174[7:0] ? 4'hf : _GEN_2302; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2304 = 8'h69 == _T_174[7:0] ? 4'hf : _GEN_2303; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2305 = 8'h6a == _T_174[7:0] ? 4'hf : _GEN_2304; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2306 = 8'h6b == _T_174[7:0] ? 4'hf : _GEN_2305; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2307 = 8'h6c == _T_174[7:0] ? 4'hf : _GEN_2306; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2308 = 8'h6d == _T_174[7:0] ? 4'hf : _GEN_2307; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2309 = 8'h6e == _T_174[7:0] ? 4'hf : _GEN_2308; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2310 = 8'h6f == _T_174[7:0] ? 4'hf : _GEN_2309; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2311 = 8'h70 == _T_174[7:0] ? 4'h0 : _GEN_2310; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2312 = 8'h71 == _T_174[7:0] ? 4'h0 : _GEN_2311; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2313 = 8'h72 == _T_174[7:0] ? 4'h0 : _GEN_2312; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2314 = 8'h73 == _T_174[7:0] ? 4'h0 : _GEN_2313; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2315 = 8'h74 == _T_174[7:0] ? 4'h0 : _GEN_2314; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2316 = 8'h75 == _T_174[7:0] ? 4'h0 : _GEN_2315; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2317 = 8'h76 == _T_174[7:0] ? 4'h0 : _GEN_2316; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2318 = 8'h77 == _T_174[7:0] ? 4'h0 : _GEN_2317; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2319 = 8'h78 == _T_174[7:0] ? 4'hf : _GEN_2318; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2320 = 8'h79 == _T_174[7:0] ? 4'hf : _GEN_2319; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2321 = 8'h7a == _T_174[7:0] ? 4'hf : _GEN_2320; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2322 = 8'h7b == _T_174[7:0] ? 4'hf : _GEN_2321; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2323 = 8'h7c == _T_174[7:0] ? 4'hf : _GEN_2322; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2324 = 8'h7d == _T_174[7:0] ? 4'hf : _GEN_2323; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2325 = 8'h7e == _T_174[7:0] ? 4'hf : _GEN_2324; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2326 = 8'h7f == _T_174[7:0] ? 4'hf : _GEN_2325; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2327 = 8'h80 == _T_174[7:0] ? 4'h0 : _GEN_2326; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2328 = 8'h81 == _T_174[7:0] ? 4'h0 : _GEN_2327; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2329 = 8'h82 == _T_174[7:0] ? 4'h0 : _GEN_2328; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2330 = 8'h83 == _T_174[7:0] ? 4'h0 : _GEN_2329; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2331 = 8'h84 == _T_174[7:0] ? 4'h0 : _GEN_2330; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2332 = 8'h85 == _T_174[7:0] ? 4'h0 : _GEN_2331; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2333 = 8'h86 == _T_174[7:0] ? 4'h0 : _GEN_2332; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2334 = 8'h87 == _T_174[7:0] ? 4'h0 : _GEN_2333; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2335 = 8'h88 == _T_174[7:0] ? 4'hf : _GEN_2334; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2336 = 8'h89 == _T_174[7:0] ? 4'hf : _GEN_2335; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2337 = 8'h8a == _T_174[7:0] ? 4'hf : _GEN_2336; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2338 = 8'h8b == _T_174[7:0] ? 4'hf : _GEN_2337; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2339 = 8'h8c == _T_174[7:0] ? 4'hf : _GEN_2338; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2340 = 8'h8d == _T_174[7:0] ? 4'hf : _GEN_2339; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2341 = 8'h8e == _T_174[7:0] ? 4'hf : _GEN_2340; // @[Filter.scala 196:142]
  wire [3:0] _GEN_2342 = 8'h8f == _T_174[7:0] ? 4'hf : _GEN_2341; // @[Filter.scala 196:142]
  wire [7:0] _T_188 = _GEN_2342 * 4'ha; // @[Filter.scala 196:142]
  wire [10:0] _GEN_7591 = {{3'd0}, _T_188}; // @[Filter.scala 196:109]
  wire [10:0] _T_190 = _T_183 + _GEN_7591; // @[Filter.scala 196:109]
  wire [10:0] _T_191 = _T_190 / 11'h64; // @[Filter.scala 196:150]
  wire  _T_193 = _T_164 >= 5'h10; // @[Filter.scala 199:31]
  wire  _T_197 = _T_171 >= 32'h9; // @[Filter.scala 199:63]
  wire  _T_198 = _T_193 | _T_197; // @[Filter.scala 199:58]
  wire [10:0] _GEN_2487 = io_SPI_distort ? _T_191 : {{7'd0}, _GEN_2054}; // @[Filter.scala 201:35]
  wire [10:0] _GEN_2488 = _T_198 ? 11'h0 : _GEN_2487; // @[Filter.scala 199:80]
  wire [10:0] _GEN_2633 = io_SPI_distort ? _T_191 : {{7'd0}, _GEN_2198}; // @[Filter.scala 201:35]
  wire [10:0] _GEN_2634 = _T_198 ? 11'h0 : _GEN_2633; // @[Filter.scala 199:80]
  wire [10:0] _GEN_2779 = io_SPI_distort ? _T_191 : {{7'd0}, _GEN_2342}; // @[Filter.scala 201:35]
  wire [10:0] _GEN_2780 = _T_198 ? 11'h0 : _GEN_2779; // @[Filter.scala 199:80]
  wire [31:0] _T_226 = pixelIndex + 32'h3; // @[Filter.scala 194:31]
  wire [31:0] _GEN_3 = _T_226 % 32'h10; // @[Filter.scala 194:38]
  wire [4:0] _T_227 = _GEN_3[4:0]; // @[Filter.scala 194:38]
  wire [4:0] _T_229 = _T_227 + _GEN_7559; // @[Filter.scala 194:53]
  wire [4:0] _T_231 = _T_229 - 5'h1; // @[Filter.scala 194:69]
  wire [31:0] _T_234 = _T_226 / 32'h10; // @[Filter.scala 195:38]
  wire [31:0] _T_236 = _T_234 + _GEN_7560; // @[Filter.scala 195:53]
  wire [31:0] _T_238 = _T_236 - 32'h1; // @[Filter.scala 195:69]
  wire [36:0] _T_239 = _T_238 * 32'h10; // @[Filter.scala 196:42]
  wire [36:0] _GEN_7597 = {{32'd0}, _T_231}; // @[Filter.scala 196:57]
  wire [36:0] _T_241 = _T_239 + _GEN_7597; // @[Filter.scala 196:57]
  wire [3:0] _GEN_2789 = 8'h8 == _T_241[7:0] ? 4'h0 : 4'hf; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2790 = 8'h9 == _T_241[7:0] ? 4'h0 : _GEN_2789; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2791 = 8'ha == _T_241[7:0] ? 4'h0 : _GEN_2790; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2792 = 8'hb == _T_241[7:0] ? 4'h0 : _GEN_2791; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2793 = 8'hc == _T_241[7:0] ? 4'h0 : _GEN_2792; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2794 = 8'hd == _T_241[7:0] ? 4'h0 : _GEN_2793; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2795 = 8'he == _T_241[7:0] ? 4'h0 : _GEN_2794; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2796 = 8'hf == _T_241[7:0] ? 4'h0 : _GEN_2795; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2797 = 8'h10 == _T_241[7:0] ? 4'hf : _GEN_2796; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2798 = 8'h11 == _T_241[7:0] ? 4'hf : _GEN_2797; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2799 = 8'h12 == _T_241[7:0] ? 4'hf : _GEN_2798; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2800 = 8'h13 == _T_241[7:0] ? 4'hf : _GEN_2799; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2801 = 8'h14 == _T_241[7:0] ? 4'hf : _GEN_2800; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2802 = 8'h15 == _T_241[7:0] ? 4'hf : _GEN_2801; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2803 = 8'h16 == _T_241[7:0] ? 4'hf : _GEN_2802; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2804 = 8'h17 == _T_241[7:0] ? 4'hf : _GEN_2803; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2805 = 8'h18 == _T_241[7:0] ? 4'h0 : _GEN_2804; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2806 = 8'h19 == _T_241[7:0] ? 4'h0 : _GEN_2805; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2807 = 8'h1a == _T_241[7:0] ? 4'h0 : _GEN_2806; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2808 = 8'h1b == _T_241[7:0] ? 4'h0 : _GEN_2807; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2809 = 8'h1c == _T_241[7:0] ? 4'h0 : _GEN_2808; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2810 = 8'h1d == _T_241[7:0] ? 4'h0 : _GEN_2809; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2811 = 8'h1e == _T_241[7:0] ? 4'h0 : _GEN_2810; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2812 = 8'h1f == _T_241[7:0] ? 4'h0 : _GEN_2811; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2813 = 8'h20 == _T_241[7:0] ? 4'hf : _GEN_2812; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2814 = 8'h21 == _T_241[7:0] ? 4'hf : _GEN_2813; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2815 = 8'h22 == _T_241[7:0] ? 4'hf : _GEN_2814; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2816 = 8'h23 == _T_241[7:0] ? 4'hf : _GEN_2815; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2817 = 8'h24 == _T_241[7:0] ? 4'hf : _GEN_2816; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2818 = 8'h25 == _T_241[7:0] ? 4'hf : _GEN_2817; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2819 = 8'h26 == _T_241[7:0] ? 4'hf : _GEN_2818; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2820 = 8'h27 == _T_241[7:0] ? 4'hf : _GEN_2819; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2821 = 8'h28 == _T_241[7:0] ? 4'h0 : _GEN_2820; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2822 = 8'h29 == _T_241[7:0] ? 4'h0 : _GEN_2821; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2823 = 8'h2a == _T_241[7:0] ? 4'h0 : _GEN_2822; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2824 = 8'h2b == _T_241[7:0] ? 4'h0 : _GEN_2823; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2825 = 8'h2c == _T_241[7:0] ? 4'h0 : _GEN_2824; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2826 = 8'h2d == _T_241[7:0] ? 4'h0 : _GEN_2825; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2827 = 8'h2e == _T_241[7:0] ? 4'h0 : _GEN_2826; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2828 = 8'h2f == _T_241[7:0] ? 4'h0 : _GEN_2827; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2829 = 8'h30 == _T_241[7:0] ? 4'hf : _GEN_2828; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2830 = 8'h31 == _T_241[7:0] ? 4'hf : _GEN_2829; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2831 = 8'h32 == _T_241[7:0] ? 4'hf : _GEN_2830; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2832 = 8'h33 == _T_241[7:0] ? 4'hf : _GEN_2831; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2833 = 8'h34 == _T_241[7:0] ? 4'hf : _GEN_2832; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2834 = 8'h35 == _T_241[7:0] ? 4'hf : _GEN_2833; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2835 = 8'h36 == _T_241[7:0] ? 4'hf : _GEN_2834; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2836 = 8'h37 == _T_241[7:0] ? 4'hf : _GEN_2835; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2837 = 8'h38 == _T_241[7:0] ? 4'h0 : _GEN_2836; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2838 = 8'h39 == _T_241[7:0] ? 4'h0 : _GEN_2837; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2839 = 8'h3a == _T_241[7:0] ? 4'h0 : _GEN_2838; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2840 = 8'h3b == _T_241[7:0] ? 4'h0 : _GEN_2839; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2841 = 8'h3c == _T_241[7:0] ? 4'h0 : _GEN_2840; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2842 = 8'h3d == _T_241[7:0] ? 4'h0 : _GEN_2841; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2843 = 8'h3e == _T_241[7:0] ? 4'h0 : _GEN_2842; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2844 = 8'h3f == _T_241[7:0] ? 4'h0 : _GEN_2843; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2845 = 8'h40 == _T_241[7:0] ? 4'h0 : _GEN_2844; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2846 = 8'h41 == _T_241[7:0] ? 4'h0 : _GEN_2845; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2847 = 8'h42 == _T_241[7:0] ? 4'h0 : _GEN_2846; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2848 = 8'h43 == _T_241[7:0] ? 4'h0 : _GEN_2847; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2849 = 8'h44 == _T_241[7:0] ? 4'h0 : _GEN_2848; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2850 = 8'h45 == _T_241[7:0] ? 4'h0 : _GEN_2849; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2851 = 8'h46 == _T_241[7:0] ? 4'h0 : _GEN_2850; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2852 = 8'h47 == _T_241[7:0] ? 4'h0 : _GEN_2851; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2853 = 8'h48 == _T_241[7:0] ? 4'hf : _GEN_2852; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2854 = 8'h49 == _T_241[7:0] ? 4'hf : _GEN_2853; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2855 = 8'h4a == _T_241[7:0] ? 4'hf : _GEN_2854; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2856 = 8'h4b == _T_241[7:0] ? 4'hf : _GEN_2855; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2857 = 8'h4c == _T_241[7:0] ? 4'hf : _GEN_2856; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2858 = 8'h4d == _T_241[7:0] ? 4'hf : _GEN_2857; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2859 = 8'h4e == _T_241[7:0] ? 4'hf : _GEN_2858; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2860 = 8'h4f == _T_241[7:0] ? 4'hf : _GEN_2859; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2861 = 8'h50 == _T_241[7:0] ? 4'h0 : _GEN_2860; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2862 = 8'h51 == _T_241[7:0] ? 4'h0 : _GEN_2861; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2863 = 8'h52 == _T_241[7:0] ? 4'h0 : _GEN_2862; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2864 = 8'h53 == _T_241[7:0] ? 4'h0 : _GEN_2863; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2865 = 8'h54 == _T_241[7:0] ? 4'h0 : _GEN_2864; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2866 = 8'h55 == _T_241[7:0] ? 4'h0 : _GEN_2865; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2867 = 8'h56 == _T_241[7:0] ? 4'h0 : _GEN_2866; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2868 = 8'h57 == _T_241[7:0] ? 4'h0 : _GEN_2867; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2869 = 8'h58 == _T_241[7:0] ? 4'hf : _GEN_2868; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2870 = 8'h59 == _T_241[7:0] ? 4'hf : _GEN_2869; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2871 = 8'h5a == _T_241[7:0] ? 4'hf : _GEN_2870; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2872 = 8'h5b == _T_241[7:0] ? 4'hf : _GEN_2871; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2873 = 8'h5c == _T_241[7:0] ? 4'hf : _GEN_2872; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2874 = 8'h5d == _T_241[7:0] ? 4'hf : _GEN_2873; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2875 = 8'h5e == _T_241[7:0] ? 4'hf : _GEN_2874; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2876 = 8'h5f == _T_241[7:0] ? 4'hf : _GEN_2875; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2877 = 8'h60 == _T_241[7:0] ? 4'h0 : _GEN_2876; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2878 = 8'h61 == _T_241[7:0] ? 4'h0 : _GEN_2877; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2879 = 8'h62 == _T_241[7:0] ? 4'h0 : _GEN_2878; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2880 = 8'h63 == _T_241[7:0] ? 4'h0 : _GEN_2879; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2881 = 8'h64 == _T_241[7:0] ? 4'h0 : _GEN_2880; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2882 = 8'h65 == _T_241[7:0] ? 4'h0 : _GEN_2881; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2883 = 8'h66 == _T_241[7:0] ? 4'h0 : _GEN_2882; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2884 = 8'h67 == _T_241[7:0] ? 4'h0 : _GEN_2883; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2885 = 8'h68 == _T_241[7:0] ? 4'hf : _GEN_2884; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2886 = 8'h69 == _T_241[7:0] ? 4'hf : _GEN_2885; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2887 = 8'h6a == _T_241[7:0] ? 4'hf : _GEN_2886; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2888 = 8'h6b == _T_241[7:0] ? 4'hf : _GEN_2887; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2889 = 8'h6c == _T_241[7:0] ? 4'hf : _GEN_2888; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2890 = 8'h6d == _T_241[7:0] ? 4'hf : _GEN_2889; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2891 = 8'h6e == _T_241[7:0] ? 4'hf : _GEN_2890; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2892 = 8'h6f == _T_241[7:0] ? 4'hf : _GEN_2891; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2893 = 8'h70 == _T_241[7:0] ? 4'h0 : _GEN_2892; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2894 = 8'h71 == _T_241[7:0] ? 4'h0 : _GEN_2893; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2895 = 8'h72 == _T_241[7:0] ? 4'h0 : _GEN_2894; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2896 = 8'h73 == _T_241[7:0] ? 4'h0 : _GEN_2895; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2897 = 8'h74 == _T_241[7:0] ? 4'h0 : _GEN_2896; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2898 = 8'h75 == _T_241[7:0] ? 4'h0 : _GEN_2897; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2899 = 8'h76 == _T_241[7:0] ? 4'h0 : _GEN_2898; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2900 = 8'h77 == _T_241[7:0] ? 4'h0 : _GEN_2899; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2901 = 8'h78 == _T_241[7:0] ? 4'hf : _GEN_2900; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2902 = 8'h79 == _T_241[7:0] ? 4'hf : _GEN_2901; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2903 = 8'h7a == _T_241[7:0] ? 4'hf : _GEN_2902; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2904 = 8'h7b == _T_241[7:0] ? 4'hf : _GEN_2903; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2905 = 8'h7c == _T_241[7:0] ? 4'hf : _GEN_2904; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2906 = 8'h7d == _T_241[7:0] ? 4'hf : _GEN_2905; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2907 = 8'h7e == _T_241[7:0] ? 4'hf : _GEN_2906; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2908 = 8'h7f == _T_241[7:0] ? 4'hf : _GEN_2907; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2909 = 8'h80 == _T_241[7:0] ? 4'h0 : _GEN_2908; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2910 = 8'h81 == _T_241[7:0] ? 4'h0 : _GEN_2909; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2911 = 8'h82 == _T_241[7:0] ? 4'h0 : _GEN_2910; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2912 = 8'h83 == _T_241[7:0] ? 4'h0 : _GEN_2911; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2913 = 8'h84 == _T_241[7:0] ? 4'h0 : _GEN_2912; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2914 = 8'h85 == _T_241[7:0] ? 4'h0 : _GEN_2913; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2915 = 8'h86 == _T_241[7:0] ? 4'h0 : _GEN_2914; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2916 = 8'h87 == _T_241[7:0] ? 4'h0 : _GEN_2915; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2917 = 8'h88 == _T_241[7:0] ? 4'hf : _GEN_2916; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2918 = 8'h89 == _T_241[7:0] ? 4'hf : _GEN_2917; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2919 = 8'h8a == _T_241[7:0] ? 4'hf : _GEN_2918; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2920 = 8'h8b == _T_241[7:0] ? 4'hf : _GEN_2919; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2921 = 8'h8c == _T_241[7:0] ? 4'hf : _GEN_2920; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2922 = 8'h8d == _T_241[7:0] ? 4'hf : _GEN_2921; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2923 = 8'h8e == _T_241[7:0] ? 4'hf : _GEN_2922; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2924 = 8'h8f == _T_241[7:0] ? 4'hf : _GEN_2923; // @[Filter.scala 196:62]
  wire [4:0] _GEN_7598 = {{1'd0}, _GEN_2924}; // @[Filter.scala 196:62]
  wire [8:0] _T_243 = _GEN_7598 * 5'h14; // @[Filter.scala 196:62]
  wire [3:0] _GEN_2989 = 8'h40 == _T_241[7:0] ? 4'hf : 4'h0; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2990 = 8'h41 == _T_241[7:0] ? 4'hf : _GEN_2989; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2991 = 8'h42 == _T_241[7:0] ? 4'hf : _GEN_2990; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2992 = 8'h43 == _T_241[7:0] ? 4'hf : _GEN_2991; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2993 = 8'h44 == _T_241[7:0] ? 4'hf : _GEN_2992; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2994 = 8'h45 == _T_241[7:0] ? 4'hf : _GEN_2993; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2995 = 8'h46 == _T_241[7:0] ? 4'hf : _GEN_2994; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2996 = 8'h47 == _T_241[7:0] ? 4'hf : _GEN_2995; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2997 = 8'h48 == _T_241[7:0] ? 4'hf : _GEN_2996; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2998 = 8'h49 == _T_241[7:0] ? 4'hf : _GEN_2997; // @[Filter.scala 196:102]
  wire [3:0] _GEN_2999 = 8'h4a == _T_241[7:0] ? 4'hf : _GEN_2998; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3000 = 8'h4b == _T_241[7:0] ? 4'hf : _GEN_2999; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3001 = 8'h4c == _T_241[7:0] ? 4'hf : _GEN_3000; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3002 = 8'h4d == _T_241[7:0] ? 4'hf : _GEN_3001; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3003 = 8'h4e == _T_241[7:0] ? 4'hf : _GEN_3002; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3004 = 8'h4f == _T_241[7:0] ? 4'hf : _GEN_3003; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3005 = 8'h50 == _T_241[7:0] ? 4'hf : _GEN_3004; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3006 = 8'h51 == _T_241[7:0] ? 4'hf : _GEN_3005; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3007 = 8'h52 == _T_241[7:0] ? 4'hf : _GEN_3006; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3008 = 8'h53 == _T_241[7:0] ? 4'hf : _GEN_3007; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3009 = 8'h54 == _T_241[7:0] ? 4'hf : _GEN_3008; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3010 = 8'h55 == _T_241[7:0] ? 4'hf : _GEN_3009; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3011 = 8'h56 == _T_241[7:0] ? 4'hf : _GEN_3010; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3012 = 8'h57 == _T_241[7:0] ? 4'hf : _GEN_3011; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3013 = 8'h58 == _T_241[7:0] ? 4'hf : _GEN_3012; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3014 = 8'h59 == _T_241[7:0] ? 4'hf : _GEN_3013; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3015 = 8'h5a == _T_241[7:0] ? 4'hf : _GEN_3014; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3016 = 8'h5b == _T_241[7:0] ? 4'hf : _GEN_3015; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3017 = 8'h5c == _T_241[7:0] ? 4'hf : _GEN_3016; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3018 = 8'h5d == _T_241[7:0] ? 4'hf : _GEN_3017; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3019 = 8'h5e == _T_241[7:0] ? 4'hf : _GEN_3018; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3020 = 8'h5f == _T_241[7:0] ? 4'hf : _GEN_3019; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3021 = 8'h60 == _T_241[7:0] ? 4'hf : _GEN_3020; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3022 = 8'h61 == _T_241[7:0] ? 4'hf : _GEN_3021; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3023 = 8'h62 == _T_241[7:0] ? 4'hf : _GEN_3022; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3024 = 8'h63 == _T_241[7:0] ? 4'hf : _GEN_3023; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3025 = 8'h64 == _T_241[7:0] ? 4'hf : _GEN_3024; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3026 = 8'h65 == _T_241[7:0] ? 4'hf : _GEN_3025; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3027 = 8'h66 == _T_241[7:0] ? 4'hf : _GEN_3026; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3028 = 8'h67 == _T_241[7:0] ? 4'hf : _GEN_3027; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3029 = 8'h68 == _T_241[7:0] ? 4'hf : _GEN_3028; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3030 = 8'h69 == _T_241[7:0] ? 4'hf : _GEN_3029; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3031 = 8'h6a == _T_241[7:0] ? 4'hf : _GEN_3030; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3032 = 8'h6b == _T_241[7:0] ? 4'hf : _GEN_3031; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3033 = 8'h6c == _T_241[7:0] ? 4'hf : _GEN_3032; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3034 = 8'h6d == _T_241[7:0] ? 4'hf : _GEN_3033; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3035 = 8'h6e == _T_241[7:0] ? 4'hf : _GEN_3034; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3036 = 8'h6f == _T_241[7:0] ? 4'hf : _GEN_3035; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3037 = 8'h70 == _T_241[7:0] ? 4'hf : _GEN_3036; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3038 = 8'h71 == _T_241[7:0] ? 4'hf : _GEN_3037; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3039 = 8'h72 == _T_241[7:0] ? 4'hf : _GEN_3038; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3040 = 8'h73 == _T_241[7:0] ? 4'hf : _GEN_3039; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3041 = 8'h74 == _T_241[7:0] ? 4'hf : _GEN_3040; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3042 = 8'h75 == _T_241[7:0] ? 4'hf : _GEN_3041; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3043 = 8'h76 == _T_241[7:0] ? 4'hf : _GEN_3042; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3044 = 8'h77 == _T_241[7:0] ? 4'hf : _GEN_3043; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3045 = 8'h78 == _T_241[7:0] ? 4'hf : _GEN_3044; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3046 = 8'h79 == _T_241[7:0] ? 4'hf : _GEN_3045; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3047 = 8'h7a == _T_241[7:0] ? 4'hf : _GEN_3046; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3048 = 8'h7b == _T_241[7:0] ? 4'hf : _GEN_3047; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3049 = 8'h7c == _T_241[7:0] ? 4'hf : _GEN_3048; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3050 = 8'h7d == _T_241[7:0] ? 4'hf : _GEN_3049; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3051 = 8'h7e == _T_241[7:0] ? 4'hf : _GEN_3050; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3052 = 8'h7f == _T_241[7:0] ? 4'hf : _GEN_3051; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3053 = 8'h80 == _T_241[7:0] ? 4'hf : _GEN_3052; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3054 = 8'h81 == _T_241[7:0] ? 4'hf : _GEN_3053; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3055 = 8'h82 == _T_241[7:0] ? 4'hf : _GEN_3054; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3056 = 8'h83 == _T_241[7:0] ? 4'hf : _GEN_3055; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3057 = 8'h84 == _T_241[7:0] ? 4'hf : _GEN_3056; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3058 = 8'h85 == _T_241[7:0] ? 4'hf : _GEN_3057; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3059 = 8'h86 == _T_241[7:0] ? 4'hf : _GEN_3058; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3060 = 8'h87 == _T_241[7:0] ? 4'hf : _GEN_3059; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3061 = 8'h88 == _T_241[7:0] ? 4'hf : _GEN_3060; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3062 = 8'h89 == _T_241[7:0] ? 4'hf : _GEN_3061; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3063 = 8'h8a == _T_241[7:0] ? 4'hf : _GEN_3062; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3064 = 8'h8b == _T_241[7:0] ? 4'hf : _GEN_3063; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3065 = 8'h8c == _T_241[7:0] ? 4'hf : _GEN_3064; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3066 = 8'h8d == _T_241[7:0] ? 4'hf : _GEN_3065; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3067 = 8'h8e == _T_241[7:0] ? 4'hf : _GEN_3066; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3068 = 8'h8f == _T_241[7:0] ? 4'hf : _GEN_3067; // @[Filter.scala 196:102]
  wire [6:0] _GEN_7600 = {{3'd0}, _GEN_3068}; // @[Filter.scala 196:102]
  wire [10:0] _T_248 = _GEN_7600 * 7'h46; // @[Filter.scala 196:102]
  wire [10:0] _GEN_7601 = {{2'd0}, _T_243}; // @[Filter.scala 196:69]
  wire [10:0] _T_250 = _GEN_7601 + _T_248; // @[Filter.scala 196:69]
  wire [3:0] _GEN_3077 = 8'h8 == _T_241[7:0] ? 4'hf : 4'h0; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3078 = 8'h9 == _T_241[7:0] ? 4'hf : _GEN_3077; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3079 = 8'ha == _T_241[7:0] ? 4'hf : _GEN_3078; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3080 = 8'hb == _T_241[7:0] ? 4'hf : _GEN_3079; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3081 = 8'hc == _T_241[7:0] ? 4'hf : _GEN_3080; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3082 = 8'hd == _T_241[7:0] ? 4'hf : _GEN_3081; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3083 = 8'he == _T_241[7:0] ? 4'hf : _GEN_3082; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3084 = 8'hf == _T_241[7:0] ? 4'hf : _GEN_3083; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3085 = 8'h10 == _T_241[7:0] ? 4'h0 : _GEN_3084; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3086 = 8'h11 == _T_241[7:0] ? 4'h0 : _GEN_3085; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3087 = 8'h12 == _T_241[7:0] ? 4'h0 : _GEN_3086; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3088 = 8'h13 == _T_241[7:0] ? 4'h0 : _GEN_3087; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3089 = 8'h14 == _T_241[7:0] ? 4'h0 : _GEN_3088; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3090 = 8'h15 == _T_241[7:0] ? 4'h0 : _GEN_3089; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3091 = 8'h16 == _T_241[7:0] ? 4'h0 : _GEN_3090; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3092 = 8'h17 == _T_241[7:0] ? 4'h0 : _GEN_3091; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3093 = 8'h18 == _T_241[7:0] ? 4'hf : _GEN_3092; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3094 = 8'h19 == _T_241[7:0] ? 4'hf : _GEN_3093; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3095 = 8'h1a == _T_241[7:0] ? 4'hf : _GEN_3094; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3096 = 8'h1b == _T_241[7:0] ? 4'hf : _GEN_3095; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3097 = 8'h1c == _T_241[7:0] ? 4'hf : _GEN_3096; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3098 = 8'h1d == _T_241[7:0] ? 4'hf : _GEN_3097; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3099 = 8'h1e == _T_241[7:0] ? 4'hf : _GEN_3098; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3100 = 8'h1f == _T_241[7:0] ? 4'hf : _GEN_3099; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3101 = 8'h20 == _T_241[7:0] ? 4'h0 : _GEN_3100; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3102 = 8'h21 == _T_241[7:0] ? 4'h0 : _GEN_3101; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3103 = 8'h22 == _T_241[7:0] ? 4'h0 : _GEN_3102; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3104 = 8'h23 == _T_241[7:0] ? 4'h0 : _GEN_3103; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3105 = 8'h24 == _T_241[7:0] ? 4'h0 : _GEN_3104; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3106 = 8'h25 == _T_241[7:0] ? 4'h0 : _GEN_3105; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3107 = 8'h26 == _T_241[7:0] ? 4'h0 : _GEN_3106; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3108 = 8'h27 == _T_241[7:0] ? 4'h0 : _GEN_3107; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3109 = 8'h28 == _T_241[7:0] ? 4'hf : _GEN_3108; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3110 = 8'h29 == _T_241[7:0] ? 4'hf : _GEN_3109; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3111 = 8'h2a == _T_241[7:0] ? 4'hf : _GEN_3110; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3112 = 8'h2b == _T_241[7:0] ? 4'hf : _GEN_3111; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3113 = 8'h2c == _T_241[7:0] ? 4'hf : _GEN_3112; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3114 = 8'h2d == _T_241[7:0] ? 4'hf : _GEN_3113; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3115 = 8'h2e == _T_241[7:0] ? 4'hf : _GEN_3114; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3116 = 8'h2f == _T_241[7:0] ? 4'hf : _GEN_3115; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3117 = 8'h30 == _T_241[7:0] ? 4'h0 : _GEN_3116; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3118 = 8'h31 == _T_241[7:0] ? 4'h0 : _GEN_3117; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3119 = 8'h32 == _T_241[7:0] ? 4'h0 : _GEN_3118; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3120 = 8'h33 == _T_241[7:0] ? 4'h0 : _GEN_3119; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3121 = 8'h34 == _T_241[7:0] ? 4'h0 : _GEN_3120; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3122 = 8'h35 == _T_241[7:0] ? 4'h0 : _GEN_3121; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3123 = 8'h36 == _T_241[7:0] ? 4'h0 : _GEN_3122; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3124 = 8'h37 == _T_241[7:0] ? 4'h0 : _GEN_3123; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3125 = 8'h38 == _T_241[7:0] ? 4'hf : _GEN_3124; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3126 = 8'h39 == _T_241[7:0] ? 4'hf : _GEN_3125; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3127 = 8'h3a == _T_241[7:0] ? 4'hf : _GEN_3126; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3128 = 8'h3b == _T_241[7:0] ? 4'hf : _GEN_3127; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3129 = 8'h3c == _T_241[7:0] ? 4'hf : _GEN_3128; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3130 = 8'h3d == _T_241[7:0] ? 4'hf : _GEN_3129; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3131 = 8'h3e == _T_241[7:0] ? 4'hf : _GEN_3130; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3132 = 8'h3f == _T_241[7:0] ? 4'hf : _GEN_3131; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3133 = 8'h40 == _T_241[7:0] ? 4'h0 : _GEN_3132; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3134 = 8'h41 == _T_241[7:0] ? 4'h0 : _GEN_3133; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3135 = 8'h42 == _T_241[7:0] ? 4'h0 : _GEN_3134; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3136 = 8'h43 == _T_241[7:0] ? 4'h0 : _GEN_3135; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3137 = 8'h44 == _T_241[7:0] ? 4'h0 : _GEN_3136; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3138 = 8'h45 == _T_241[7:0] ? 4'h0 : _GEN_3137; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3139 = 8'h46 == _T_241[7:0] ? 4'h0 : _GEN_3138; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3140 = 8'h47 == _T_241[7:0] ? 4'h0 : _GEN_3139; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3141 = 8'h48 == _T_241[7:0] ? 4'hf : _GEN_3140; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3142 = 8'h49 == _T_241[7:0] ? 4'hf : _GEN_3141; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3143 = 8'h4a == _T_241[7:0] ? 4'hf : _GEN_3142; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3144 = 8'h4b == _T_241[7:0] ? 4'hf : _GEN_3143; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3145 = 8'h4c == _T_241[7:0] ? 4'hf : _GEN_3144; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3146 = 8'h4d == _T_241[7:0] ? 4'hf : _GEN_3145; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3147 = 8'h4e == _T_241[7:0] ? 4'hf : _GEN_3146; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3148 = 8'h4f == _T_241[7:0] ? 4'hf : _GEN_3147; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3149 = 8'h50 == _T_241[7:0] ? 4'h0 : _GEN_3148; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3150 = 8'h51 == _T_241[7:0] ? 4'h0 : _GEN_3149; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3151 = 8'h52 == _T_241[7:0] ? 4'h0 : _GEN_3150; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3152 = 8'h53 == _T_241[7:0] ? 4'h0 : _GEN_3151; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3153 = 8'h54 == _T_241[7:0] ? 4'h0 : _GEN_3152; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3154 = 8'h55 == _T_241[7:0] ? 4'h0 : _GEN_3153; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3155 = 8'h56 == _T_241[7:0] ? 4'h0 : _GEN_3154; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3156 = 8'h57 == _T_241[7:0] ? 4'h0 : _GEN_3155; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3157 = 8'h58 == _T_241[7:0] ? 4'hf : _GEN_3156; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3158 = 8'h59 == _T_241[7:0] ? 4'hf : _GEN_3157; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3159 = 8'h5a == _T_241[7:0] ? 4'hf : _GEN_3158; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3160 = 8'h5b == _T_241[7:0] ? 4'hf : _GEN_3159; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3161 = 8'h5c == _T_241[7:0] ? 4'hf : _GEN_3160; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3162 = 8'h5d == _T_241[7:0] ? 4'hf : _GEN_3161; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3163 = 8'h5e == _T_241[7:0] ? 4'hf : _GEN_3162; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3164 = 8'h5f == _T_241[7:0] ? 4'hf : _GEN_3163; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3165 = 8'h60 == _T_241[7:0] ? 4'h0 : _GEN_3164; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3166 = 8'h61 == _T_241[7:0] ? 4'h0 : _GEN_3165; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3167 = 8'h62 == _T_241[7:0] ? 4'h0 : _GEN_3166; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3168 = 8'h63 == _T_241[7:0] ? 4'h0 : _GEN_3167; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3169 = 8'h64 == _T_241[7:0] ? 4'h0 : _GEN_3168; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3170 = 8'h65 == _T_241[7:0] ? 4'h0 : _GEN_3169; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3171 = 8'h66 == _T_241[7:0] ? 4'h0 : _GEN_3170; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3172 = 8'h67 == _T_241[7:0] ? 4'h0 : _GEN_3171; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3173 = 8'h68 == _T_241[7:0] ? 4'hf : _GEN_3172; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3174 = 8'h69 == _T_241[7:0] ? 4'hf : _GEN_3173; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3175 = 8'h6a == _T_241[7:0] ? 4'hf : _GEN_3174; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3176 = 8'h6b == _T_241[7:0] ? 4'hf : _GEN_3175; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3177 = 8'h6c == _T_241[7:0] ? 4'hf : _GEN_3176; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3178 = 8'h6d == _T_241[7:0] ? 4'hf : _GEN_3177; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3179 = 8'h6e == _T_241[7:0] ? 4'hf : _GEN_3178; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3180 = 8'h6f == _T_241[7:0] ? 4'hf : _GEN_3179; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3181 = 8'h70 == _T_241[7:0] ? 4'h0 : _GEN_3180; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3182 = 8'h71 == _T_241[7:0] ? 4'h0 : _GEN_3181; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3183 = 8'h72 == _T_241[7:0] ? 4'h0 : _GEN_3182; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3184 = 8'h73 == _T_241[7:0] ? 4'h0 : _GEN_3183; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3185 = 8'h74 == _T_241[7:0] ? 4'h0 : _GEN_3184; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3186 = 8'h75 == _T_241[7:0] ? 4'h0 : _GEN_3185; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3187 = 8'h76 == _T_241[7:0] ? 4'h0 : _GEN_3186; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3188 = 8'h77 == _T_241[7:0] ? 4'h0 : _GEN_3187; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3189 = 8'h78 == _T_241[7:0] ? 4'hf : _GEN_3188; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3190 = 8'h79 == _T_241[7:0] ? 4'hf : _GEN_3189; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3191 = 8'h7a == _T_241[7:0] ? 4'hf : _GEN_3190; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3192 = 8'h7b == _T_241[7:0] ? 4'hf : _GEN_3191; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3193 = 8'h7c == _T_241[7:0] ? 4'hf : _GEN_3192; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3194 = 8'h7d == _T_241[7:0] ? 4'hf : _GEN_3193; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3195 = 8'h7e == _T_241[7:0] ? 4'hf : _GEN_3194; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3196 = 8'h7f == _T_241[7:0] ? 4'hf : _GEN_3195; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3197 = 8'h80 == _T_241[7:0] ? 4'h0 : _GEN_3196; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3198 = 8'h81 == _T_241[7:0] ? 4'h0 : _GEN_3197; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3199 = 8'h82 == _T_241[7:0] ? 4'h0 : _GEN_3198; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3200 = 8'h83 == _T_241[7:0] ? 4'h0 : _GEN_3199; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3201 = 8'h84 == _T_241[7:0] ? 4'h0 : _GEN_3200; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3202 = 8'h85 == _T_241[7:0] ? 4'h0 : _GEN_3201; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3203 = 8'h86 == _T_241[7:0] ? 4'h0 : _GEN_3202; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3204 = 8'h87 == _T_241[7:0] ? 4'h0 : _GEN_3203; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3205 = 8'h88 == _T_241[7:0] ? 4'hf : _GEN_3204; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3206 = 8'h89 == _T_241[7:0] ? 4'hf : _GEN_3205; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3207 = 8'h8a == _T_241[7:0] ? 4'hf : _GEN_3206; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3208 = 8'h8b == _T_241[7:0] ? 4'hf : _GEN_3207; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3209 = 8'h8c == _T_241[7:0] ? 4'hf : _GEN_3208; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3210 = 8'h8d == _T_241[7:0] ? 4'hf : _GEN_3209; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3211 = 8'h8e == _T_241[7:0] ? 4'hf : _GEN_3210; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3212 = 8'h8f == _T_241[7:0] ? 4'hf : _GEN_3211; // @[Filter.scala 196:142]
  wire [7:0] _T_255 = _GEN_3212 * 4'ha; // @[Filter.scala 196:142]
  wire [10:0] _GEN_7603 = {{3'd0}, _T_255}; // @[Filter.scala 196:109]
  wire [10:0] _T_257 = _T_250 + _GEN_7603; // @[Filter.scala 196:109]
  wire [10:0] _T_258 = _T_257 / 11'h64; // @[Filter.scala 196:150]
  wire  _T_260 = _T_231 >= 5'h10; // @[Filter.scala 199:31]
  wire  _T_264 = _T_238 >= 32'h9; // @[Filter.scala 199:63]
  wire  _T_265 = _T_260 | _T_264; // @[Filter.scala 199:58]
  wire [10:0] _GEN_3357 = io_SPI_distort ? _T_258 : {{7'd0}, _GEN_2924}; // @[Filter.scala 201:35]
  wire [10:0] _GEN_3358 = _T_265 ? 11'h0 : _GEN_3357; // @[Filter.scala 199:80]
  wire [10:0] _GEN_3503 = io_SPI_distort ? _T_258 : {{7'd0}, _GEN_3068}; // @[Filter.scala 201:35]
  wire [10:0] _GEN_3504 = _T_265 ? 11'h0 : _GEN_3503; // @[Filter.scala 199:80]
  wire [10:0] _GEN_3649 = io_SPI_distort ? _T_258 : {{7'd0}, _GEN_3212}; // @[Filter.scala 201:35]
  wire [10:0] _GEN_3650 = _T_265 ? 11'h0 : _GEN_3649; // @[Filter.scala 199:80]
  wire [31:0] _T_293 = pixelIndex + 32'h4; // @[Filter.scala 194:31]
  wire [31:0] _GEN_4 = _T_293 % 32'h10; // @[Filter.scala 194:38]
  wire [4:0] _T_294 = _GEN_4[4:0]; // @[Filter.scala 194:38]
  wire [4:0] _T_296 = _T_294 + _GEN_7559; // @[Filter.scala 194:53]
  wire [4:0] _T_298 = _T_296 - 5'h1; // @[Filter.scala 194:69]
  wire [31:0] _T_301 = _T_293 / 32'h10; // @[Filter.scala 195:38]
  wire [31:0] _T_303 = _T_301 + _GEN_7560; // @[Filter.scala 195:53]
  wire [31:0] _T_305 = _T_303 - 32'h1; // @[Filter.scala 195:69]
  wire [36:0] _T_306 = _T_305 * 32'h10; // @[Filter.scala 196:42]
  wire [36:0] _GEN_7609 = {{32'd0}, _T_298}; // @[Filter.scala 196:57]
  wire [36:0] _T_308 = _T_306 + _GEN_7609; // @[Filter.scala 196:57]
  wire [3:0] _GEN_3659 = 8'h8 == _T_308[7:0] ? 4'h0 : 4'hf; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3660 = 8'h9 == _T_308[7:0] ? 4'h0 : _GEN_3659; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3661 = 8'ha == _T_308[7:0] ? 4'h0 : _GEN_3660; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3662 = 8'hb == _T_308[7:0] ? 4'h0 : _GEN_3661; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3663 = 8'hc == _T_308[7:0] ? 4'h0 : _GEN_3662; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3664 = 8'hd == _T_308[7:0] ? 4'h0 : _GEN_3663; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3665 = 8'he == _T_308[7:0] ? 4'h0 : _GEN_3664; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3666 = 8'hf == _T_308[7:0] ? 4'h0 : _GEN_3665; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3667 = 8'h10 == _T_308[7:0] ? 4'hf : _GEN_3666; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3668 = 8'h11 == _T_308[7:0] ? 4'hf : _GEN_3667; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3669 = 8'h12 == _T_308[7:0] ? 4'hf : _GEN_3668; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3670 = 8'h13 == _T_308[7:0] ? 4'hf : _GEN_3669; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3671 = 8'h14 == _T_308[7:0] ? 4'hf : _GEN_3670; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3672 = 8'h15 == _T_308[7:0] ? 4'hf : _GEN_3671; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3673 = 8'h16 == _T_308[7:0] ? 4'hf : _GEN_3672; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3674 = 8'h17 == _T_308[7:0] ? 4'hf : _GEN_3673; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3675 = 8'h18 == _T_308[7:0] ? 4'h0 : _GEN_3674; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3676 = 8'h19 == _T_308[7:0] ? 4'h0 : _GEN_3675; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3677 = 8'h1a == _T_308[7:0] ? 4'h0 : _GEN_3676; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3678 = 8'h1b == _T_308[7:0] ? 4'h0 : _GEN_3677; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3679 = 8'h1c == _T_308[7:0] ? 4'h0 : _GEN_3678; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3680 = 8'h1d == _T_308[7:0] ? 4'h0 : _GEN_3679; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3681 = 8'h1e == _T_308[7:0] ? 4'h0 : _GEN_3680; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3682 = 8'h1f == _T_308[7:0] ? 4'h0 : _GEN_3681; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3683 = 8'h20 == _T_308[7:0] ? 4'hf : _GEN_3682; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3684 = 8'h21 == _T_308[7:0] ? 4'hf : _GEN_3683; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3685 = 8'h22 == _T_308[7:0] ? 4'hf : _GEN_3684; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3686 = 8'h23 == _T_308[7:0] ? 4'hf : _GEN_3685; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3687 = 8'h24 == _T_308[7:0] ? 4'hf : _GEN_3686; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3688 = 8'h25 == _T_308[7:0] ? 4'hf : _GEN_3687; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3689 = 8'h26 == _T_308[7:0] ? 4'hf : _GEN_3688; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3690 = 8'h27 == _T_308[7:0] ? 4'hf : _GEN_3689; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3691 = 8'h28 == _T_308[7:0] ? 4'h0 : _GEN_3690; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3692 = 8'h29 == _T_308[7:0] ? 4'h0 : _GEN_3691; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3693 = 8'h2a == _T_308[7:0] ? 4'h0 : _GEN_3692; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3694 = 8'h2b == _T_308[7:0] ? 4'h0 : _GEN_3693; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3695 = 8'h2c == _T_308[7:0] ? 4'h0 : _GEN_3694; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3696 = 8'h2d == _T_308[7:0] ? 4'h0 : _GEN_3695; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3697 = 8'h2e == _T_308[7:0] ? 4'h0 : _GEN_3696; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3698 = 8'h2f == _T_308[7:0] ? 4'h0 : _GEN_3697; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3699 = 8'h30 == _T_308[7:0] ? 4'hf : _GEN_3698; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3700 = 8'h31 == _T_308[7:0] ? 4'hf : _GEN_3699; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3701 = 8'h32 == _T_308[7:0] ? 4'hf : _GEN_3700; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3702 = 8'h33 == _T_308[7:0] ? 4'hf : _GEN_3701; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3703 = 8'h34 == _T_308[7:0] ? 4'hf : _GEN_3702; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3704 = 8'h35 == _T_308[7:0] ? 4'hf : _GEN_3703; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3705 = 8'h36 == _T_308[7:0] ? 4'hf : _GEN_3704; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3706 = 8'h37 == _T_308[7:0] ? 4'hf : _GEN_3705; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3707 = 8'h38 == _T_308[7:0] ? 4'h0 : _GEN_3706; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3708 = 8'h39 == _T_308[7:0] ? 4'h0 : _GEN_3707; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3709 = 8'h3a == _T_308[7:0] ? 4'h0 : _GEN_3708; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3710 = 8'h3b == _T_308[7:0] ? 4'h0 : _GEN_3709; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3711 = 8'h3c == _T_308[7:0] ? 4'h0 : _GEN_3710; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3712 = 8'h3d == _T_308[7:0] ? 4'h0 : _GEN_3711; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3713 = 8'h3e == _T_308[7:0] ? 4'h0 : _GEN_3712; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3714 = 8'h3f == _T_308[7:0] ? 4'h0 : _GEN_3713; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3715 = 8'h40 == _T_308[7:0] ? 4'h0 : _GEN_3714; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3716 = 8'h41 == _T_308[7:0] ? 4'h0 : _GEN_3715; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3717 = 8'h42 == _T_308[7:0] ? 4'h0 : _GEN_3716; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3718 = 8'h43 == _T_308[7:0] ? 4'h0 : _GEN_3717; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3719 = 8'h44 == _T_308[7:0] ? 4'h0 : _GEN_3718; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3720 = 8'h45 == _T_308[7:0] ? 4'h0 : _GEN_3719; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3721 = 8'h46 == _T_308[7:0] ? 4'h0 : _GEN_3720; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3722 = 8'h47 == _T_308[7:0] ? 4'h0 : _GEN_3721; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3723 = 8'h48 == _T_308[7:0] ? 4'hf : _GEN_3722; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3724 = 8'h49 == _T_308[7:0] ? 4'hf : _GEN_3723; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3725 = 8'h4a == _T_308[7:0] ? 4'hf : _GEN_3724; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3726 = 8'h4b == _T_308[7:0] ? 4'hf : _GEN_3725; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3727 = 8'h4c == _T_308[7:0] ? 4'hf : _GEN_3726; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3728 = 8'h4d == _T_308[7:0] ? 4'hf : _GEN_3727; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3729 = 8'h4e == _T_308[7:0] ? 4'hf : _GEN_3728; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3730 = 8'h4f == _T_308[7:0] ? 4'hf : _GEN_3729; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3731 = 8'h50 == _T_308[7:0] ? 4'h0 : _GEN_3730; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3732 = 8'h51 == _T_308[7:0] ? 4'h0 : _GEN_3731; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3733 = 8'h52 == _T_308[7:0] ? 4'h0 : _GEN_3732; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3734 = 8'h53 == _T_308[7:0] ? 4'h0 : _GEN_3733; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3735 = 8'h54 == _T_308[7:0] ? 4'h0 : _GEN_3734; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3736 = 8'h55 == _T_308[7:0] ? 4'h0 : _GEN_3735; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3737 = 8'h56 == _T_308[7:0] ? 4'h0 : _GEN_3736; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3738 = 8'h57 == _T_308[7:0] ? 4'h0 : _GEN_3737; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3739 = 8'h58 == _T_308[7:0] ? 4'hf : _GEN_3738; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3740 = 8'h59 == _T_308[7:0] ? 4'hf : _GEN_3739; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3741 = 8'h5a == _T_308[7:0] ? 4'hf : _GEN_3740; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3742 = 8'h5b == _T_308[7:0] ? 4'hf : _GEN_3741; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3743 = 8'h5c == _T_308[7:0] ? 4'hf : _GEN_3742; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3744 = 8'h5d == _T_308[7:0] ? 4'hf : _GEN_3743; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3745 = 8'h5e == _T_308[7:0] ? 4'hf : _GEN_3744; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3746 = 8'h5f == _T_308[7:0] ? 4'hf : _GEN_3745; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3747 = 8'h60 == _T_308[7:0] ? 4'h0 : _GEN_3746; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3748 = 8'h61 == _T_308[7:0] ? 4'h0 : _GEN_3747; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3749 = 8'h62 == _T_308[7:0] ? 4'h0 : _GEN_3748; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3750 = 8'h63 == _T_308[7:0] ? 4'h0 : _GEN_3749; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3751 = 8'h64 == _T_308[7:0] ? 4'h0 : _GEN_3750; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3752 = 8'h65 == _T_308[7:0] ? 4'h0 : _GEN_3751; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3753 = 8'h66 == _T_308[7:0] ? 4'h0 : _GEN_3752; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3754 = 8'h67 == _T_308[7:0] ? 4'h0 : _GEN_3753; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3755 = 8'h68 == _T_308[7:0] ? 4'hf : _GEN_3754; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3756 = 8'h69 == _T_308[7:0] ? 4'hf : _GEN_3755; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3757 = 8'h6a == _T_308[7:0] ? 4'hf : _GEN_3756; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3758 = 8'h6b == _T_308[7:0] ? 4'hf : _GEN_3757; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3759 = 8'h6c == _T_308[7:0] ? 4'hf : _GEN_3758; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3760 = 8'h6d == _T_308[7:0] ? 4'hf : _GEN_3759; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3761 = 8'h6e == _T_308[7:0] ? 4'hf : _GEN_3760; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3762 = 8'h6f == _T_308[7:0] ? 4'hf : _GEN_3761; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3763 = 8'h70 == _T_308[7:0] ? 4'h0 : _GEN_3762; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3764 = 8'h71 == _T_308[7:0] ? 4'h0 : _GEN_3763; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3765 = 8'h72 == _T_308[7:0] ? 4'h0 : _GEN_3764; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3766 = 8'h73 == _T_308[7:0] ? 4'h0 : _GEN_3765; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3767 = 8'h74 == _T_308[7:0] ? 4'h0 : _GEN_3766; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3768 = 8'h75 == _T_308[7:0] ? 4'h0 : _GEN_3767; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3769 = 8'h76 == _T_308[7:0] ? 4'h0 : _GEN_3768; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3770 = 8'h77 == _T_308[7:0] ? 4'h0 : _GEN_3769; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3771 = 8'h78 == _T_308[7:0] ? 4'hf : _GEN_3770; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3772 = 8'h79 == _T_308[7:0] ? 4'hf : _GEN_3771; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3773 = 8'h7a == _T_308[7:0] ? 4'hf : _GEN_3772; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3774 = 8'h7b == _T_308[7:0] ? 4'hf : _GEN_3773; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3775 = 8'h7c == _T_308[7:0] ? 4'hf : _GEN_3774; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3776 = 8'h7d == _T_308[7:0] ? 4'hf : _GEN_3775; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3777 = 8'h7e == _T_308[7:0] ? 4'hf : _GEN_3776; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3778 = 8'h7f == _T_308[7:0] ? 4'hf : _GEN_3777; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3779 = 8'h80 == _T_308[7:0] ? 4'h0 : _GEN_3778; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3780 = 8'h81 == _T_308[7:0] ? 4'h0 : _GEN_3779; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3781 = 8'h82 == _T_308[7:0] ? 4'h0 : _GEN_3780; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3782 = 8'h83 == _T_308[7:0] ? 4'h0 : _GEN_3781; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3783 = 8'h84 == _T_308[7:0] ? 4'h0 : _GEN_3782; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3784 = 8'h85 == _T_308[7:0] ? 4'h0 : _GEN_3783; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3785 = 8'h86 == _T_308[7:0] ? 4'h0 : _GEN_3784; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3786 = 8'h87 == _T_308[7:0] ? 4'h0 : _GEN_3785; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3787 = 8'h88 == _T_308[7:0] ? 4'hf : _GEN_3786; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3788 = 8'h89 == _T_308[7:0] ? 4'hf : _GEN_3787; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3789 = 8'h8a == _T_308[7:0] ? 4'hf : _GEN_3788; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3790 = 8'h8b == _T_308[7:0] ? 4'hf : _GEN_3789; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3791 = 8'h8c == _T_308[7:0] ? 4'hf : _GEN_3790; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3792 = 8'h8d == _T_308[7:0] ? 4'hf : _GEN_3791; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3793 = 8'h8e == _T_308[7:0] ? 4'hf : _GEN_3792; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3794 = 8'h8f == _T_308[7:0] ? 4'hf : _GEN_3793; // @[Filter.scala 196:62]
  wire [4:0] _GEN_7610 = {{1'd0}, _GEN_3794}; // @[Filter.scala 196:62]
  wire [8:0] _T_310 = _GEN_7610 * 5'h14; // @[Filter.scala 196:62]
  wire [3:0] _GEN_3859 = 8'h40 == _T_308[7:0] ? 4'hf : 4'h0; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3860 = 8'h41 == _T_308[7:0] ? 4'hf : _GEN_3859; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3861 = 8'h42 == _T_308[7:0] ? 4'hf : _GEN_3860; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3862 = 8'h43 == _T_308[7:0] ? 4'hf : _GEN_3861; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3863 = 8'h44 == _T_308[7:0] ? 4'hf : _GEN_3862; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3864 = 8'h45 == _T_308[7:0] ? 4'hf : _GEN_3863; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3865 = 8'h46 == _T_308[7:0] ? 4'hf : _GEN_3864; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3866 = 8'h47 == _T_308[7:0] ? 4'hf : _GEN_3865; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3867 = 8'h48 == _T_308[7:0] ? 4'hf : _GEN_3866; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3868 = 8'h49 == _T_308[7:0] ? 4'hf : _GEN_3867; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3869 = 8'h4a == _T_308[7:0] ? 4'hf : _GEN_3868; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3870 = 8'h4b == _T_308[7:0] ? 4'hf : _GEN_3869; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3871 = 8'h4c == _T_308[7:0] ? 4'hf : _GEN_3870; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3872 = 8'h4d == _T_308[7:0] ? 4'hf : _GEN_3871; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3873 = 8'h4e == _T_308[7:0] ? 4'hf : _GEN_3872; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3874 = 8'h4f == _T_308[7:0] ? 4'hf : _GEN_3873; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3875 = 8'h50 == _T_308[7:0] ? 4'hf : _GEN_3874; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3876 = 8'h51 == _T_308[7:0] ? 4'hf : _GEN_3875; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3877 = 8'h52 == _T_308[7:0] ? 4'hf : _GEN_3876; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3878 = 8'h53 == _T_308[7:0] ? 4'hf : _GEN_3877; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3879 = 8'h54 == _T_308[7:0] ? 4'hf : _GEN_3878; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3880 = 8'h55 == _T_308[7:0] ? 4'hf : _GEN_3879; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3881 = 8'h56 == _T_308[7:0] ? 4'hf : _GEN_3880; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3882 = 8'h57 == _T_308[7:0] ? 4'hf : _GEN_3881; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3883 = 8'h58 == _T_308[7:0] ? 4'hf : _GEN_3882; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3884 = 8'h59 == _T_308[7:0] ? 4'hf : _GEN_3883; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3885 = 8'h5a == _T_308[7:0] ? 4'hf : _GEN_3884; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3886 = 8'h5b == _T_308[7:0] ? 4'hf : _GEN_3885; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3887 = 8'h5c == _T_308[7:0] ? 4'hf : _GEN_3886; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3888 = 8'h5d == _T_308[7:0] ? 4'hf : _GEN_3887; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3889 = 8'h5e == _T_308[7:0] ? 4'hf : _GEN_3888; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3890 = 8'h5f == _T_308[7:0] ? 4'hf : _GEN_3889; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3891 = 8'h60 == _T_308[7:0] ? 4'hf : _GEN_3890; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3892 = 8'h61 == _T_308[7:0] ? 4'hf : _GEN_3891; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3893 = 8'h62 == _T_308[7:0] ? 4'hf : _GEN_3892; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3894 = 8'h63 == _T_308[7:0] ? 4'hf : _GEN_3893; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3895 = 8'h64 == _T_308[7:0] ? 4'hf : _GEN_3894; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3896 = 8'h65 == _T_308[7:0] ? 4'hf : _GEN_3895; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3897 = 8'h66 == _T_308[7:0] ? 4'hf : _GEN_3896; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3898 = 8'h67 == _T_308[7:0] ? 4'hf : _GEN_3897; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3899 = 8'h68 == _T_308[7:0] ? 4'hf : _GEN_3898; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3900 = 8'h69 == _T_308[7:0] ? 4'hf : _GEN_3899; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3901 = 8'h6a == _T_308[7:0] ? 4'hf : _GEN_3900; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3902 = 8'h6b == _T_308[7:0] ? 4'hf : _GEN_3901; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3903 = 8'h6c == _T_308[7:0] ? 4'hf : _GEN_3902; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3904 = 8'h6d == _T_308[7:0] ? 4'hf : _GEN_3903; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3905 = 8'h6e == _T_308[7:0] ? 4'hf : _GEN_3904; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3906 = 8'h6f == _T_308[7:0] ? 4'hf : _GEN_3905; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3907 = 8'h70 == _T_308[7:0] ? 4'hf : _GEN_3906; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3908 = 8'h71 == _T_308[7:0] ? 4'hf : _GEN_3907; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3909 = 8'h72 == _T_308[7:0] ? 4'hf : _GEN_3908; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3910 = 8'h73 == _T_308[7:0] ? 4'hf : _GEN_3909; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3911 = 8'h74 == _T_308[7:0] ? 4'hf : _GEN_3910; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3912 = 8'h75 == _T_308[7:0] ? 4'hf : _GEN_3911; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3913 = 8'h76 == _T_308[7:0] ? 4'hf : _GEN_3912; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3914 = 8'h77 == _T_308[7:0] ? 4'hf : _GEN_3913; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3915 = 8'h78 == _T_308[7:0] ? 4'hf : _GEN_3914; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3916 = 8'h79 == _T_308[7:0] ? 4'hf : _GEN_3915; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3917 = 8'h7a == _T_308[7:0] ? 4'hf : _GEN_3916; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3918 = 8'h7b == _T_308[7:0] ? 4'hf : _GEN_3917; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3919 = 8'h7c == _T_308[7:0] ? 4'hf : _GEN_3918; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3920 = 8'h7d == _T_308[7:0] ? 4'hf : _GEN_3919; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3921 = 8'h7e == _T_308[7:0] ? 4'hf : _GEN_3920; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3922 = 8'h7f == _T_308[7:0] ? 4'hf : _GEN_3921; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3923 = 8'h80 == _T_308[7:0] ? 4'hf : _GEN_3922; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3924 = 8'h81 == _T_308[7:0] ? 4'hf : _GEN_3923; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3925 = 8'h82 == _T_308[7:0] ? 4'hf : _GEN_3924; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3926 = 8'h83 == _T_308[7:0] ? 4'hf : _GEN_3925; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3927 = 8'h84 == _T_308[7:0] ? 4'hf : _GEN_3926; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3928 = 8'h85 == _T_308[7:0] ? 4'hf : _GEN_3927; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3929 = 8'h86 == _T_308[7:0] ? 4'hf : _GEN_3928; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3930 = 8'h87 == _T_308[7:0] ? 4'hf : _GEN_3929; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3931 = 8'h88 == _T_308[7:0] ? 4'hf : _GEN_3930; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3932 = 8'h89 == _T_308[7:0] ? 4'hf : _GEN_3931; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3933 = 8'h8a == _T_308[7:0] ? 4'hf : _GEN_3932; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3934 = 8'h8b == _T_308[7:0] ? 4'hf : _GEN_3933; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3935 = 8'h8c == _T_308[7:0] ? 4'hf : _GEN_3934; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3936 = 8'h8d == _T_308[7:0] ? 4'hf : _GEN_3935; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3937 = 8'h8e == _T_308[7:0] ? 4'hf : _GEN_3936; // @[Filter.scala 196:102]
  wire [3:0] _GEN_3938 = 8'h8f == _T_308[7:0] ? 4'hf : _GEN_3937; // @[Filter.scala 196:102]
  wire [6:0] _GEN_7612 = {{3'd0}, _GEN_3938}; // @[Filter.scala 196:102]
  wire [10:0] _T_315 = _GEN_7612 * 7'h46; // @[Filter.scala 196:102]
  wire [10:0] _GEN_7613 = {{2'd0}, _T_310}; // @[Filter.scala 196:69]
  wire [10:0] _T_317 = _GEN_7613 + _T_315; // @[Filter.scala 196:69]
  wire [3:0] _GEN_3947 = 8'h8 == _T_308[7:0] ? 4'hf : 4'h0; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3948 = 8'h9 == _T_308[7:0] ? 4'hf : _GEN_3947; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3949 = 8'ha == _T_308[7:0] ? 4'hf : _GEN_3948; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3950 = 8'hb == _T_308[7:0] ? 4'hf : _GEN_3949; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3951 = 8'hc == _T_308[7:0] ? 4'hf : _GEN_3950; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3952 = 8'hd == _T_308[7:0] ? 4'hf : _GEN_3951; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3953 = 8'he == _T_308[7:0] ? 4'hf : _GEN_3952; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3954 = 8'hf == _T_308[7:0] ? 4'hf : _GEN_3953; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3955 = 8'h10 == _T_308[7:0] ? 4'h0 : _GEN_3954; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3956 = 8'h11 == _T_308[7:0] ? 4'h0 : _GEN_3955; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3957 = 8'h12 == _T_308[7:0] ? 4'h0 : _GEN_3956; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3958 = 8'h13 == _T_308[7:0] ? 4'h0 : _GEN_3957; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3959 = 8'h14 == _T_308[7:0] ? 4'h0 : _GEN_3958; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3960 = 8'h15 == _T_308[7:0] ? 4'h0 : _GEN_3959; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3961 = 8'h16 == _T_308[7:0] ? 4'h0 : _GEN_3960; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3962 = 8'h17 == _T_308[7:0] ? 4'h0 : _GEN_3961; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3963 = 8'h18 == _T_308[7:0] ? 4'hf : _GEN_3962; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3964 = 8'h19 == _T_308[7:0] ? 4'hf : _GEN_3963; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3965 = 8'h1a == _T_308[7:0] ? 4'hf : _GEN_3964; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3966 = 8'h1b == _T_308[7:0] ? 4'hf : _GEN_3965; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3967 = 8'h1c == _T_308[7:0] ? 4'hf : _GEN_3966; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3968 = 8'h1d == _T_308[7:0] ? 4'hf : _GEN_3967; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3969 = 8'h1e == _T_308[7:0] ? 4'hf : _GEN_3968; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3970 = 8'h1f == _T_308[7:0] ? 4'hf : _GEN_3969; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3971 = 8'h20 == _T_308[7:0] ? 4'h0 : _GEN_3970; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3972 = 8'h21 == _T_308[7:0] ? 4'h0 : _GEN_3971; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3973 = 8'h22 == _T_308[7:0] ? 4'h0 : _GEN_3972; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3974 = 8'h23 == _T_308[7:0] ? 4'h0 : _GEN_3973; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3975 = 8'h24 == _T_308[7:0] ? 4'h0 : _GEN_3974; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3976 = 8'h25 == _T_308[7:0] ? 4'h0 : _GEN_3975; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3977 = 8'h26 == _T_308[7:0] ? 4'h0 : _GEN_3976; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3978 = 8'h27 == _T_308[7:0] ? 4'h0 : _GEN_3977; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3979 = 8'h28 == _T_308[7:0] ? 4'hf : _GEN_3978; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3980 = 8'h29 == _T_308[7:0] ? 4'hf : _GEN_3979; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3981 = 8'h2a == _T_308[7:0] ? 4'hf : _GEN_3980; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3982 = 8'h2b == _T_308[7:0] ? 4'hf : _GEN_3981; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3983 = 8'h2c == _T_308[7:0] ? 4'hf : _GEN_3982; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3984 = 8'h2d == _T_308[7:0] ? 4'hf : _GEN_3983; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3985 = 8'h2e == _T_308[7:0] ? 4'hf : _GEN_3984; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3986 = 8'h2f == _T_308[7:0] ? 4'hf : _GEN_3985; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3987 = 8'h30 == _T_308[7:0] ? 4'h0 : _GEN_3986; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3988 = 8'h31 == _T_308[7:0] ? 4'h0 : _GEN_3987; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3989 = 8'h32 == _T_308[7:0] ? 4'h0 : _GEN_3988; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3990 = 8'h33 == _T_308[7:0] ? 4'h0 : _GEN_3989; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3991 = 8'h34 == _T_308[7:0] ? 4'h0 : _GEN_3990; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3992 = 8'h35 == _T_308[7:0] ? 4'h0 : _GEN_3991; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3993 = 8'h36 == _T_308[7:0] ? 4'h0 : _GEN_3992; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3994 = 8'h37 == _T_308[7:0] ? 4'h0 : _GEN_3993; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3995 = 8'h38 == _T_308[7:0] ? 4'hf : _GEN_3994; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3996 = 8'h39 == _T_308[7:0] ? 4'hf : _GEN_3995; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3997 = 8'h3a == _T_308[7:0] ? 4'hf : _GEN_3996; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3998 = 8'h3b == _T_308[7:0] ? 4'hf : _GEN_3997; // @[Filter.scala 196:142]
  wire [3:0] _GEN_3999 = 8'h3c == _T_308[7:0] ? 4'hf : _GEN_3998; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4000 = 8'h3d == _T_308[7:0] ? 4'hf : _GEN_3999; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4001 = 8'h3e == _T_308[7:0] ? 4'hf : _GEN_4000; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4002 = 8'h3f == _T_308[7:0] ? 4'hf : _GEN_4001; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4003 = 8'h40 == _T_308[7:0] ? 4'h0 : _GEN_4002; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4004 = 8'h41 == _T_308[7:0] ? 4'h0 : _GEN_4003; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4005 = 8'h42 == _T_308[7:0] ? 4'h0 : _GEN_4004; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4006 = 8'h43 == _T_308[7:0] ? 4'h0 : _GEN_4005; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4007 = 8'h44 == _T_308[7:0] ? 4'h0 : _GEN_4006; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4008 = 8'h45 == _T_308[7:0] ? 4'h0 : _GEN_4007; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4009 = 8'h46 == _T_308[7:0] ? 4'h0 : _GEN_4008; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4010 = 8'h47 == _T_308[7:0] ? 4'h0 : _GEN_4009; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4011 = 8'h48 == _T_308[7:0] ? 4'hf : _GEN_4010; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4012 = 8'h49 == _T_308[7:0] ? 4'hf : _GEN_4011; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4013 = 8'h4a == _T_308[7:0] ? 4'hf : _GEN_4012; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4014 = 8'h4b == _T_308[7:0] ? 4'hf : _GEN_4013; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4015 = 8'h4c == _T_308[7:0] ? 4'hf : _GEN_4014; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4016 = 8'h4d == _T_308[7:0] ? 4'hf : _GEN_4015; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4017 = 8'h4e == _T_308[7:0] ? 4'hf : _GEN_4016; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4018 = 8'h4f == _T_308[7:0] ? 4'hf : _GEN_4017; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4019 = 8'h50 == _T_308[7:0] ? 4'h0 : _GEN_4018; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4020 = 8'h51 == _T_308[7:0] ? 4'h0 : _GEN_4019; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4021 = 8'h52 == _T_308[7:0] ? 4'h0 : _GEN_4020; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4022 = 8'h53 == _T_308[7:0] ? 4'h0 : _GEN_4021; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4023 = 8'h54 == _T_308[7:0] ? 4'h0 : _GEN_4022; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4024 = 8'h55 == _T_308[7:0] ? 4'h0 : _GEN_4023; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4025 = 8'h56 == _T_308[7:0] ? 4'h0 : _GEN_4024; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4026 = 8'h57 == _T_308[7:0] ? 4'h0 : _GEN_4025; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4027 = 8'h58 == _T_308[7:0] ? 4'hf : _GEN_4026; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4028 = 8'h59 == _T_308[7:0] ? 4'hf : _GEN_4027; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4029 = 8'h5a == _T_308[7:0] ? 4'hf : _GEN_4028; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4030 = 8'h5b == _T_308[7:0] ? 4'hf : _GEN_4029; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4031 = 8'h5c == _T_308[7:0] ? 4'hf : _GEN_4030; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4032 = 8'h5d == _T_308[7:0] ? 4'hf : _GEN_4031; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4033 = 8'h5e == _T_308[7:0] ? 4'hf : _GEN_4032; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4034 = 8'h5f == _T_308[7:0] ? 4'hf : _GEN_4033; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4035 = 8'h60 == _T_308[7:0] ? 4'h0 : _GEN_4034; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4036 = 8'h61 == _T_308[7:0] ? 4'h0 : _GEN_4035; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4037 = 8'h62 == _T_308[7:0] ? 4'h0 : _GEN_4036; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4038 = 8'h63 == _T_308[7:0] ? 4'h0 : _GEN_4037; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4039 = 8'h64 == _T_308[7:0] ? 4'h0 : _GEN_4038; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4040 = 8'h65 == _T_308[7:0] ? 4'h0 : _GEN_4039; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4041 = 8'h66 == _T_308[7:0] ? 4'h0 : _GEN_4040; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4042 = 8'h67 == _T_308[7:0] ? 4'h0 : _GEN_4041; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4043 = 8'h68 == _T_308[7:0] ? 4'hf : _GEN_4042; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4044 = 8'h69 == _T_308[7:0] ? 4'hf : _GEN_4043; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4045 = 8'h6a == _T_308[7:0] ? 4'hf : _GEN_4044; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4046 = 8'h6b == _T_308[7:0] ? 4'hf : _GEN_4045; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4047 = 8'h6c == _T_308[7:0] ? 4'hf : _GEN_4046; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4048 = 8'h6d == _T_308[7:0] ? 4'hf : _GEN_4047; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4049 = 8'h6e == _T_308[7:0] ? 4'hf : _GEN_4048; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4050 = 8'h6f == _T_308[7:0] ? 4'hf : _GEN_4049; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4051 = 8'h70 == _T_308[7:0] ? 4'h0 : _GEN_4050; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4052 = 8'h71 == _T_308[7:0] ? 4'h0 : _GEN_4051; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4053 = 8'h72 == _T_308[7:0] ? 4'h0 : _GEN_4052; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4054 = 8'h73 == _T_308[7:0] ? 4'h0 : _GEN_4053; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4055 = 8'h74 == _T_308[7:0] ? 4'h0 : _GEN_4054; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4056 = 8'h75 == _T_308[7:0] ? 4'h0 : _GEN_4055; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4057 = 8'h76 == _T_308[7:0] ? 4'h0 : _GEN_4056; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4058 = 8'h77 == _T_308[7:0] ? 4'h0 : _GEN_4057; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4059 = 8'h78 == _T_308[7:0] ? 4'hf : _GEN_4058; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4060 = 8'h79 == _T_308[7:0] ? 4'hf : _GEN_4059; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4061 = 8'h7a == _T_308[7:0] ? 4'hf : _GEN_4060; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4062 = 8'h7b == _T_308[7:0] ? 4'hf : _GEN_4061; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4063 = 8'h7c == _T_308[7:0] ? 4'hf : _GEN_4062; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4064 = 8'h7d == _T_308[7:0] ? 4'hf : _GEN_4063; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4065 = 8'h7e == _T_308[7:0] ? 4'hf : _GEN_4064; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4066 = 8'h7f == _T_308[7:0] ? 4'hf : _GEN_4065; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4067 = 8'h80 == _T_308[7:0] ? 4'h0 : _GEN_4066; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4068 = 8'h81 == _T_308[7:0] ? 4'h0 : _GEN_4067; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4069 = 8'h82 == _T_308[7:0] ? 4'h0 : _GEN_4068; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4070 = 8'h83 == _T_308[7:0] ? 4'h0 : _GEN_4069; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4071 = 8'h84 == _T_308[7:0] ? 4'h0 : _GEN_4070; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4072 = 8'h85 == _T_308[7:0] ? 4'h0 : _GEN_4071; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4073 = 8'h86 == _T_308[7:0] ? 4'h0 : _GEN_4072; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4074 = 8'h87 == _T_308[7:0] ? 4'h0 : _GEN_4073; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4075 = 8'h88 == _T_308[7:0] ? 4'hf : _GEN_4074; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4076 = 8'h89 == _T_308[7:0] ? 4'hf : _GEN_4075; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4077 = 8'h8a == _T_308[7:0] ? 4'hf : _GEN_4076; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4078 = 8'h8b == _T_308[7:0] ? 4'hf : _GEN_4077; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4079 = 8'h8c == _T_308[7:0] ? 4'hf : _GEN_4078; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4080 = 8'h8d == _T_308[7:0] ? 4'hf : _GEN_4079; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4081 = 8'h8e == _T_308[7:0] ? 4'hf : _GEN_4080; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4082 = 8'h8f == _T_308[7:0] ? 4'hf : _GEN_4081; // @[Filter.scala 196:142]
  wire [7:0] _T_322 = _GEN_4082 * 4'ha; // @[Filter.scala 196:142]
  wire [10:0] _GEN_7615 = {{3'd0}, _T_322}; // @[Filter.scala 196:109]
  wire [10:0] _T_324 = _T_317 + _GEN_7615; // @[Filter.scala 196:109]
  wire [10:0] _T_325 = _T_324 / 11'h64; // @[Filter.scala 196:150]
  wire  _T_327 = _T_298 >= 5'h10; // @[Filter.scala 199:31]
  wire  _T_331 = _T_305 >= 32'h9; // @[Filter.scala 199:63]
  wire  _T_332 = _T_327 | _T_331; // @[Filter.scala 199:58]
  wire [10:0] _GEN_4227 = io_SPI_distort ? _T_325 : {{7'd0}, _GEN_3794}; // @[Filter.scala 201:35]
  wire [10:0] _GEN_4228 = _T_332 ? 11'h0 : _GEN_4227; // @[Filter.scala 199:80]
  wire [10:0] _GEN_4373 = io_SPI_distort ? _T_325 : {{7'd0}, _GEN_3938}; // @[Filter.scala 201:35]
  wire [10:0] _GEN_4374 = _T_332 ? 11'h0 : _GEN_4373; // @[Filter.scala 199:80]
  wire [10:0] _GEN_4519 = io_SPI_distort ? _T_325 : {{7'd0}, _GEN_4082}; // @[Filter.scala 201:35]
  wire [10:0] _GEN_4520 = _T_332 ? 11'h0 : _GEN_4519; // @[Filter.scala 199:80]
  wire [31:0] _T_360 = pixelIndex + 32'h5; // @[Filter.scala 194:31]
  wire [31:0] _GEN_5 = _T_360 % 32'h10; // @[Filter.scala 194:38]
  wire [4:0] _T_361 = _GEN_5[4:0]; // @[Filter.scala 194:38]
  wire [4:0] _T_363 = _T_361 + _GEN_7559; // @[Filter.scala 194:53]
  wire [4:0] _T_365 = _T_363 - 5'h1; // @[Filter.scala 194:69]
  wire [31:0] _T_368 = _T_360 / 32'h10; // @[Filter.scala 195:38]
  wire [31:0] _T_370 = _T_368 + _GEN_7560; // @[Filter.scala 195:53]
  wire [31:0] _T_372 = _T_370 - 32'h1; // @[Filter.scala 195:69]
  wire [36:0] _T_373 = _T_372 * 32'h10; // @[Filter.scala 196:42]
  wire [36:0] _GEN_7621 = {{32'd0}, _T_365}; // @[Filter.scala 196:57]
  wire [36:0] _T_375 = _T_373 + _GEN_7621; // @[Filter.scala 196:57]
  wire [3:0] _GEN_4529 = 8'h8 == _T_375[7:0] ? 4'h0 : 4'hf; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4530 = 8'h9 == _T_375[7:0] ? 4'h0 : _GEN_4529; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4531 = 8'ha == _T_375[7:0] ? 4'h0 : _GEN_4530; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4532 = 8'hb == _T_375[7:0] ? 4'h0 : _GEN_4531; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4533 = 8'hc == _T_375[7:0] ? 4'h0 : _GEN_4532; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4534 = 8'hd == _T_375[7:0] ? 4'h0 : _GEN_4533; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4535 = 8'he == _T_375[7:0] ? 4'h0 : _GEN_4534; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4536 = 8'hf == _T_375[7:0] ? 4'h0 : _GEN_4535; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4537 = 8'h10 == _T_375[7:0] ? 4'hf : _GEN_4536; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4538 = 8'h11 == _T_375[7:0] ? 4'hf : _GEN_4537; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4539 = 8'h12 == _T_375[7:0] ? 4'hf : _GEN_4538; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4540 = 8'h13 == _T_375[7:0] ? 4'hf : _GEN_4539; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4541 = 8'h14 == _T_375[7:0] ? 4'hf : _GEN_4540; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4542 = 8'h15 == _T_375[7:0] ? 4'hf : _GEN_4541; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4543 = 8'h16 == _T_375[7:0] ? 4'hf : _GEN_4542; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4544 = 8'h17 == _T_375[7:0] ? 4'hf : _GEN_4543; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4545 = 8'h18 == _T_375[7:0] ? 4'h0 : _GEN_4544; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4546 = 8'h19 == _T_375[7:0] ? 4'h0 : _GEN_4545; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4547 = 8'h1a == _T_375[7:0] ? 4'h0 : _GEN_4546; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4548 = 8'h1b == _T_375[7:0] ? 4'h0 : _GEN_4547; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4549 = 8'h1c == _T_375[7:0] ? 4'h0 : _GEN_4548; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4550 = 8'h1d == _T_375[7:0] ? 4'h0 : _GEN_4549; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4551 = 8'h1e == _T_375[7:0] ? 4'h0 : _GEN_4550; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4552 = 8'h1f == _T_375[7:0] ? 4'h0 : _GEN_4551; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4553 = 8'h20 == _T_375[7:0] ? 4'hf : _GEN_4552; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4554 = 8'h21 == _T_375[7:0] ? 4'hf : _GEN_4553; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4555 = 8'h22 == _T_375[7:0] ? 4'hf : _GEN_4554; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4556 = 8'h23 == _T_375[7:0] ? 4'hf : _GEN_4555; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4557 = 8'h24 == _T_375[7:0] ? 4'hf : _GEN_4556; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4558 = 8'h25 == _T_375[7:0] ? 4'hf : _GEN_4557; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4559 = 8'h26 == _T_375[7:0] ? 4'hf : _GEN_4558; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4560 = 8'h27 == _T_375[7:0] ? 4'hf : _GEN_4559; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4561 = 8'h28 == _T_375[7:0] ? 4'h0 : _GEN_4560; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4562 = 8'h29 == _T_375[7:0] ? 4'h0 : _GEN_4561; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4563 = 8'h2a == _T_375[7:0] ? 4'h0 : _GEN_4562; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4564 = 8'h2b == _T_375[7:0] ? 4'h0 : _GEN_4563; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4565 = 8'h2c == _T_375[7:0] ? 4'h0 : _GEN_4564; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4566 = 8'h2d == _T_375[7:0] ? 4'h0 : _GEN_4565; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4567 = 8'h2e == _T_375[7:0] ? 4'h0 : _GEN_4566; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4568 = 8'h2f == _T_375[7:0] ? 4'h0 : _GEN_4567; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4569 = 8'h30 == _T_375[7:0] ? 4'hf : _GEN_4568; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4570 = 8'h31 == _T_375[7:0] ? 4'hf : _GEN_4569; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4571 = 8'h32 == _T_375[7:0] ? 4'hf : _GEN_4570; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4572 = 8'h33 == _T_375[7:0] ? 4'hf : _GEN_4571; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4573 = 8'h34 == _T_375[7:0] ? 4'hf : _GEN_4572; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4574 = 8'h35 == _T_375[7:0] ? 4'hf : _GEN_4573; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4575 = 8'h36 == _T_375[7:0] ? 4'hf : _GEN_4574; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4576 = 8'h37 == _T_375[7:0] ? 4'hf : _GEN_4575; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4577 = 8'h38 == _T_375[7:0] ? 4'h0 : _GEN_4576; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4578 = 8'h39 == _T_375[7:0] ? 4'h0 : _GEN_4577; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4579 = 8'h3a == _T_375[7:0] ? 4'h0 : _GEN_4578; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4580 = 8'h3b == _T_375[7:0] ? 4'h0 : _GEN_4579; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4581 = 8'h3c == _T_375[7:0] ? 4'h0 : _GEN_4580; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4582 = 8'h3d == _T_375[7:0] ? 4'h0 : _GEN_4581; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4583 = 8'h3e == _T_375[7:0] ? 4'h0 : _GEN_4582; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4584 = 8'h3f == _T_375[7:0] ? 4'h0 : _GEN_4583; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4585 = 8'h40 == _T_375[7:0] ? 4'h0 : _GEN_4584; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4586 = 8'h41 == _T_375[7:0] ? 4'h0 : _GEN_4585; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4587 = 8'h42 == _T_375[7:0] ? 4'h0 : _GEN_4586; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4588 = 8'h43 == _T_375[7:0] ? 4'h0 : _GEN_4587; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4589 = 8'h44 == _T_375[7:0] ? 4'h0 : _GEN_4588; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4590 = 8'h45 == _T_375[7:0] ? 4'h0 : _GEN_4589; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4591 = 8'h46 == _T_375[7:0] ? 4'h0 : _GEN_4590; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4592 = 8'h47 == _T_375[7:0] ? 4'h0 : _GEN_4591; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4593 = 8'h48 == _T_375[7:0] ? 4'hf : _GEN_4592; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4594 = 8'h49 == _T_375[7:0] ? 4'hf : _GEN_4593; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4595 = 8'h4a == _T_375[7:0] ? 4'hf : _GEN_4594; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4596 = 8'h4b == _T_375[7:0] ? 4'hf : _GEN_4595; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4597 = 8'h4c == _T_375[7:0] ? 4'hf : _GEN_4596; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4598 = 8'h4d == _T_375[7:0] ? 4'hf : _GEN_4597; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4599 = 8'h4e == _T_375[7:0] ? 4'hf : _GEN_4598; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4600 = 8'h4f == _T_375[7:0] ? 4'hf : _GEN_4599; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4601 = 8'h50 == _T_375[7:0] ? 4'h0 : _GEN_4600; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4602 = 8'h51 == _T_375[7:0] ? 4'h0 : _GEN_4601; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4603 = 8'h52 == _T_375[7:0] ? 4'h0 : _GEN_4602; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4604 = 8'h53 == _T_375[7:0] ? 4'h0 : _GEN_4603; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4605 = 8'h54 == _T_375[7:0] ? 4'h0 : _GEN_4604; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4606 = 8'h55 == _T_375[7:0] ? 4'h0 : _GEN_4605; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4607 = 8'h56 == _T_375[7:0] ? 4'h0 : _GEN_4606; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4608 = 8'h57 == _T_375[7:0] ? 4'h0 : _GEN_4607; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4609 = 8'h58 == _T_375[7:0] ? 4'hf : _GEN_4608; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4610 = 8'h59 == _T_375[7:0] ? 4'hf : _GEN_4609; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4611 = 8'h5a == _T_375[7:0] ? 4'hf : _GEN_4610; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4612 = 8'h5b == _T_375[7:0] ? 4'hf : _GEN_4611; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4613 = 8'h5c == _T_375[7:0] ? 4'hf : _GEN_4612; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4614 = 8'h5d == _T_375[7:0] ? 4'hf : _GEN_4613; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4615 = 8'h5e == _T_375[7:0] ? 4'hf : _GEN_4614; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4616 = 8'h5f == _T_375[7:0] ? 4'hf : _GEN_4615; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4617 = 8'h60 == _T_375[7:0] ? 4'h0 : _GEN_4616; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4618 = 8'h61 == _T_375[7:0] ? 4'h0 : _GEN_4617; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4619 = 8'h62 == _T_375[7:0] ? 4'h0 : _GEN_4618; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4620 = 8'h63 == _T_375[7:0] ? 4'h0 : _GEN_4619; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4621 = 8'h64 == _T_375[7:0] ? 4'h0 : _GEN_4620; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4622 = 8'h65 == _T_375[7:0] ? 4'h0 : _GEN_4621; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4623 = 8'h66 == _T_375[7:0] ? 4'h0 : _GEN_4622; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4624 = 8'h67 == _T_375[7:0] ? 4'h0 : _GEN_4623; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4625 = 8'h68 == _T_375[7:0] ? 4'hf : _GEN_4624; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4626 = 8'h69 == _T_375[7:0] ? 4'hf : _GEN_4625; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4627 = 8'h6a == _T_375[7:0] ? 4'hf : _GEN_4626; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4628 = 8'h6b == _T_375[7:0] ? 4'hf : _GEN_4627; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4629 = 8'h6c == _T_375[7:0] ? 4'hf : _GEN_4628; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4630 = 8'h6d == _T_375[7:0] ? 4'hf : _GEN_4629; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4631 = 8'h6e == _T_375[7:0] ? 4'hf : _GEN_4630; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4632 = 8'h6f == _T_375[7:0] ? 4'hf : _GEN_4631; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4633 = 8'h70 == _T_375[7:0] ? 4'h0 : _GEN_4632; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4634 = 8'h71 == _T_375[7:0] ? 4'h0 : _GEN_4633; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4635 = 8'h72 == _T_375[7:0] ? 4'h0 : _GEN_4634; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4636 = 8'h73 == _T_375[7:0] ? 4'h0 : _GEN_4635; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4637 = 8'h74 == _T_375[7:0] ? 4'h0 : _GEN_4636; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4638 = 8'h75 == _T_375[7:0] ? 4'h0 : _GEN_4637; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4639 = 8'h76 == _T_375[7:0] ? 4'h0 : _GEN_4638; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4640 = 8'h77 == _T_375[7:0] ? 4'h0 : _GEN_4639; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4641 = 8'h78 == _T_375[7:0] ? 4'hf : _GEN_4640; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4642 = 8'h79 == _T_375[7:0] ? 4'hf : _GEN_4641; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4643 = 8'h7a == _T_375[7:0] ? 4'hf : _GEN_4642; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4644 = 8'h7b == _T_375[7:0] ? 4'hf : _GEN_4643; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4645 = 8'h7c == _T_375[7:0] ? 4'hf : _GEN_4644; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4646 = 8'h7d == _T_375[7:0] ? 4'hf : _GEN_4645; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4647 = 8'h7e == _T_375[7:0] ? 4'hf : _GEN_4646; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4648 = 8'h7f == _T_375[7:0] ? 4'hf : _GEN_4647; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4649 = 8'h80 == _T_375[7:0] ? 4'h0 : _GEN_4648; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4650 = 8'h81 == _T_375[7:0] ? 4'h0 : _GEN_4649; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4651 = 8'h82 == _T_375[7:0] ? 4'h0 : _GEN_4650; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4652 = 8'h83 == _T_375[7:0] ? 4'h0 : _GEN_4651; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4653 = 8'h84 == _T_375[7:0] ? 4'h0 : _GEN_4652; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4654 = 8'h85 == _T_375[7:0] ? 4'h0 : _GEN_4653; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4655 = 8'h86 == _T_375[7:0] ? 4'h0 : _GEN_4654; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4656 = 8'h87 == _T_375[7:0] ? 4'h0 : _GEN_4655; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4657 = 8'h88 == _T_375[7:0] ? 4'hf : _GEN_4656; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4658 = 8'h89 == _T_375[7:0] ? 4'hf : _GEN_4657; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4659 = 8'h8a == _T_375[7:0] ? 4'hf : _GEN_4658; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4660 = 8'h8b == _T_375[7:0] ? 4'hf : _GEN_4659; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4661 = 8'h8c == _T_375[7:0] ? 4'hf : _GEN_4660; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4662 = 8'h8d == _T_375[7:0] ? 4'hf : _GEN_4661; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4663 = 8'h8e == _T_375[7:0] ? 4'hf : _GEN_4662; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4664 = 8'h8f == _T_375[7:0] ? 4'hf : _GEN_4663; // @[Filter.scala 196:62]
  wire [4:0] _GEN_7622 = {{1'd0}, _GEN_4664}; // @[Filter.scala 196:62]
  wire [8:0] _T_377 = _GEN_7622 * 5'h14; // @[Filter.scala 196:62]
  wire [3:0] _GEN_4729 = 8'h40 == _T_375[7:0] ? 4'hf : 4'h0; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4730 = 8'h41 == _T_375[7:0] ? 4'hf : _GEN_4729; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4731 = 8'h42 == _T_375[7:0] ? 4'hf : _GEN_4730; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4732 = 8'h43 == _T_375[7:0] ? 4'hf : _GEN_4731; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4733 = 8'h44 == _T_375[7:0] ? 4'hf : _GEN_4732; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4734 = 8'h45 == _T_375[7:0] ? 4'hf : _GEN_4733; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4735 = 8'h46 == _T_375[7:0] ? 4'hf : _GEN_4734; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4736 = 8'h47 == _T_375[7:0] ? 4'hf : _GEN_4735; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4737 = 8'h48 == _T_375[7:0] ? 4'hf : _GEN_4736; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4738 = 8'h49 == _T_375[7:0] ? 4'hf : _GEN_4737; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4739 = 8'h4a == _T_375[7:0] ? 4'hf : _GEN_4738; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4740 = 8'h4b == _T_375[7:0] ? 4'hf : _GEN_4739; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4741 = 8'h4c == _T_375[7:0] ? 4'hf : _GEN_4740; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4742 = 8'h4d == _T_375[7:0] ? 4'hf : _GEN_4741; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4743 = 8'h4e == _T_375[7:0] ? 4'hf : _GEN_4742; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4744 = 8'h4f == _T_375[7:0] ? 4'hf : _GEN_4743; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4745 = 8'h50 == _T_375[7:0] ? 4'hf : _GEN_4744; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4746 = 8'h51 == _T_375[7:0] ? 4'hf : _GEN_4745; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4747 = 8'h52 == _T_375[7:0] ? 4'hf : _GEN_4746; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4748 = 8'h53 == _T_375[7:0] ? 4'hf : _GEN_4747; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4749 = 8'h54 == _T_375[7:0] ? 4'hf : _GEN_4748; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4750 = 8'h55 == _T_375[7:0] ? 4'hf : _GEN_4749; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4751 = 8'h56 == _T_375[7:0] ? 4'hf : _GEN_4750; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4752 = 8'h57 == _T_375[7:0] ? 4'hf : _GEN_4751; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4753 = 8'h58 == _T_375[7:0] ? 4'hf : _GEN_4752; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4754 = 8'h59 == _T_375[7:0] ? 4'hf : _GEN_4753; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4755 = 8'h5a == _T_375[7:0] ? 4'hf : _GEN_4754; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4756 = 8'h5b == _T_375[7:0] ? 4'hf : _GEN_4755; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4757 = 8'h5c == _T_375[7:0] ? 4'hf : _GEN_4756; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4758 = 8'h5d == _T_375[7:0] ? 4'hf : _GEN_4757; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4759 = 8'h5e == _T_375[7:0] ? 4'hf : _GEN_4758; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4760 = 8'h5f == _T_375[7:0] ? 4'hf : _GEN_4759; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4761 = 8'h60 == _T_375[7:0] ? 4'hf : _GEN_4760; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4762 = 8'h61 == _T_375[7:0] ? 4'hf : _GEN_4761; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4763 = 8'h62 == _T_375[7:0] ? 4'hf : _GEN_4762; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4764 = 8'h63 == _T_375[7:0] ? 4'hf : _GEN_4763; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4765 = 8'h64 == _T_375[7:0] ? 4'hf : _GEN_4764; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4766 = 8'h65 == _T_375[7:0] ? 4'hf : _GEN_4765; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4767 = 8'h66 == _T_375[7:0] ? 4'hf : _GEN_4766; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4768 = 8'h67 == _T_375[7:0] ? 4'hf : _GEN_4767; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4769 = 8'h68 == _T_375[7:0] ? 4'hf : _GEN_4768; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4770 = 8'h69 == _T_375[7:0] ? 4'hf : _GEN_4769; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4771 = 8'h6a == _T_375[7:0] ? 4'hf : _GEN_4770; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4772 = 8'h6b == _T_375[7:0] ? 4'hf : _GEN_4771; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4773 = 8'h6c == _T_375[7:0] ? 4'hf : _GEN_4772; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4774 = 8'h6d == _T_375[7:0] ? 4'hf : _GEN_4773; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4775 = 8'h6e == _T_375[7:0] ? 4'hf : _GEN_4774; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4776 = 8'h6f == _T_375[7:0] ? 4'hf : _GEN_4775; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4777 = 8'h70 == _T_375[7:0] ? 4'hf : _GEN_4776; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4778 = 8'h71 == _T_375[7:0] ? 4'hf : _GEN_4777; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4779 = 8'h72 == _T_375[7:0] ? 4'hf : _GEN_4778; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4780 = 8'h73 == _T_375[7:0] ? 4'hf : _GEN_4779; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4781 = 8'h74 == _T_375[7:0] ? 4'hf : _GEN_4780; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4782 = 8'h75 == _T_375[7:0] ? 4'hf : _GEN_4781; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4783 = 8'h76 == _T_375[7:0] ? 4'hf : _GEN_4782; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4784 = 8'h77 == _T_375[7:0] ? 4'hf : _GEN_4783; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4785 = 8'h78 == _T_375[7:0] ? 4'hf : _GEN_4784; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4786 = 8'h79 == _T_375[7:0] ? 4'hf : _GEN_4785; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4787 = 8'h7a == _T_375[7:0] ? 4'hf : _GEN_4786; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4788 = 8'h7b == _T_375[7:0] ? 4'hf : _GEN_4787; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4789 = 8'h7c == _T_375[7:0] ? 4'hf : _GEN_4788; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4790 = 8'h7d == _T_375[7:0] ? 4'hf : _GEN_4789; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4791 = 8'h7e == _T_375[7:0] ? 4'hf : _GEN_4790; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4792 = 8'h7f == _T_375[7:0] ? 4'hf : _GEN_4791; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4793 = 8'h80 == _T_375[7:0] ? 4'hf : _GEN_4792; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4794 = 8'h81 == _T_375[7:0] ? 4'hf : _GEN_4793; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4795 = 8'h82 == _T_375[7:0] ? 4'hf : _GEN_4794; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4796 = 8'h83 == _T_375[7:0] ? 4'hf : _GEN_4795; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4797 = 8'h84 == _T_375[7:0] ? 4'hf : _GEN_4796; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4798 = 8'h85 == _T_375[7:0] ? 4'hf : _GEN_4797; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4799 = 8'h86 == _T_375[7:0] ? 4'hf : _GEN_4798; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4800 = 8'h87 == _T_375[7:0] ? 4'hf : _GEN_4799; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4801 = 8'h88 == _T_375[7:0] ? 4'hf : _GEN_4800; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4802 = 8'h89 == _T_375[7:0] ? 4'hf : _GEN_4801; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4803 = 8'h8a == _T_375[7:0] ? 4'hf : _GEN_4802; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4804 = 8'h8b == _T_375[7:0] ? 4'hf : _GEN_4803; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4805 = 8'h8c == _T_375[7:0] ? 4'hf : _GEN_4804; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4806 = 8'h8d == _T_375[7:0] ? 4'hf : _GEN_4805; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4807 = 8'h8e == _T_375[7:0] ? 4'hf : _GEN_4806; // @[Filter.scala 196:102]
  wire [3:0] _GEN_4808 = 8'h8f == _T_375[7:0] ? 4'hf : _GEN_4807; // @[Filter.scala 196:102]
  wire [6:0] _GEN_7624 = {{3'd0}, _GEN_4808}; // @[Filter.scala 196:102]
  wire [10:0] _T_382 = _GEN_7624 * 7'h46; // @[Filter.scala 196:102]
  wire [10:0] _GEN_7625 = {{2'd0}, _T_377}; // @[Filter.scala 196:69]
  wire [10:0] _T_384 = _GEN_7625 + _T_382; // @[Filter.scala 196:69]
  wire [3:0] _GEN_4817 = 8'h8 == _T_375[7:0] ? 4'hf : 4'h0; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4818 = 8'h9 == _T_375[7:0] ? 4'hf : _GEN_4817; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4819 = 8'ha == _T_375[7:0] ? 4'hf : _GEN_4818; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4820 = 8'hb == _T_375[7:0] ? 4'hf : _GEN_4819; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4821 = 8'hc == _T_375[7:0] ? 4'hf : _GEN_4820; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4822 = 8'hd == _T_375[7:0] ? 4'hf : _GEN_4821; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4823 = 8'he == _T_375[7:0] ? 4'hf : _GEN_4822; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4824 = 8'hf == _T_375[7:0] ? 4'hf : _GEN_4823; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4825 = 8'h10 == _T_375[7:0] ? 4'h0 : _GEN_4824; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4826 = 8'h11 == _T_375[7:0] ? 4'h0 : _GEN_4825; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4827 = 8'h12 == _T_375[7:0] ? 4'h0 : _GEN_4826; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4828 = 8'h13 == _T_375[7:0] ? 4'h0 : _GEN_4827; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4829 = 8'h14 == _T_375[7:0] ? 4'h0 : _GEN_4828; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4830 = 8'h15 == _T_375[7:0] ? 4'h0 : _GEN_4829; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4831 = 8'h16 == _T_375[7:0] ? 4'h0 : _GEN_4830; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4832 = 8'h17 == _T_375[7:0] ? 4'h0 : _GEN_4831; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4833 = 8'h18 == _T_375[7:0] ? 4'hf : _GEN_4832; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4834 = 8'h19 == _T_375[7:0] ? 4'hf : _GEN_4833; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4835 = 8'h1a == _T_375[7:0] ? 4'hf : _GEN_4834; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4836 = 8'h1b == _T_375[7:0] ? 4'hf : _GEN_4835; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4837 = 8'h1c == _T_375[7:0] ? 4'hf : _GEN_4836; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4838 = 8'h1d == _T_375[7:0] ? 4'hf : _GEN_4837; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4839 = 8'h1e == _T_375[7:0] ? 4'hf : _GEN_4838; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4840 = 8'h1f == _T_375[7:0] ? 4'hf : _GEN_4839; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4841 = 8'h20 == _T_375[7:0] ? 4'h0 : _GEN_4840; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4842 = 8'h21 == _T_375[7:0] ? 4'h0 : _GEN_4841; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4843 = 8'h22 == _T_375[7:0] ? 4'h0 : _GEN_4842; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4844 = 8'h23 == _T_375[7:0] ? 4'h0 : _GEN_4843; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4845 = 8'h24 == _T_375[7:0] ? 4'h0 : _GEN_4844; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4846 = 8'h25 == _T_375[7:0] ? 4'h0 : _GEN_4845; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4847 = 8'h26 == _T_375[7:0] ? 4'h0 : _GEN_4846; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4848 = 8'h27 == _T_375[7:0] ? 4'h0 : _GEN_4847; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4849 = 8'h28 == _T_375[7:0] ? 4'hf : _GEN_4848; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4850 = 8'h29 == _T_375[7:0] ? 4'hf : _GEN_4849; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4851 = 8'h2a == _T_375[7:0] ? 4'hf : _GEN_4850; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4852 = 8'h2b == _T_375[7:0] ? 4'hf : _GEN_4851; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4853 = 8'h2c == _T_375[7:0] ? 4'hf : _GEN_4852; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4854 = 8'h2d == _T_375[7:0] ? 4'hf : _GEN_4853; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4855 = 8'h2e == _T_375[7:0] ? 4'hf : _GEN_4854; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4856 = 8'h2f == _T_375[7:0] ? 4'hf : _GEN_4855; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4857 = 8'h30 == _T_375[7:0] ? 4'h0 : _GEN_4856; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4858 = 8'h31 == _T_375[7:0] ? 4'h0 : _GEN_4857; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4859 = 8'h32 == _T_375[7:0] ? 4'h0 : _GEN_4858; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4860 = 8'h33 == _T_375[7:0] ? 4'h0 : _GEN_4859; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4861 = 8'h34 == _T_375[7:0] ? 4'h0 : _GEN_4860; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4862 = 8'h35 == _T_375[7:0] ? 4'h0 : _GEN_4861; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4863 = 8'h36 == _T_375[7:0] ? 4'h0 : _GEN_4862; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4864 = 8'h37 == _T_375[7:0] ? 4'h0 : _GEN_4863; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4865 = 8'h38 == _T_375[7:0] ? 4'hf : _GEN_4864; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4866 = 8'h39 == _T_375[7:0] ? 4'hf : _GEN_4865; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4867 = 8'h3a == _T_375[7:0] ? 4'hf : _GEN_4866; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4868 = 8'h3b == _T_375[7:0] ? 4'hf : _GEN_4867; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4869 = 8'h3c == _T_375[7:0] ? 4'hf : _GEN_4868; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4870 = 8'h3d == _T_375[7:0] ? 4'hf : _GEN_4869; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4871 = 8'h3e == _T_375[7:0] ? 4'hf : _GEN_4870; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4872 = 8'h3f == _T_375[7:0] ? 4'hf : _GEN_4871; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4873 = 8'h40 == _T_375[7:0] ? 4'h0 : _GEN_4872; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4874 = 8'h41 == _T_375[7:0] ? 4'h0 : _GEN_4873; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4875 = 8'h42 == _T_375[7:0] ? 4'h0 : _GEN_4874; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4876 = 8'h43 == _T_375[7:0] ? 4'h0 : _GEN_4875; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4877 = 8'h44 == _T_375[7:0] ? 4'h0 : _GEN_4876; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4878 = 8'h45 == _T_375[7:0] ? 4'h0 : _GEN_4877; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4879 = 8'h46 == _T_375[7:0] ? 4'h0 : _GEN_4878; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4880 = 8'h47 == _T_375[7:0] ? 4'h0 : _GEN_4879; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4881 = 8'h48 == _T_375[7:0] ? 4'hf : _GEN_4880; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4882 = 8'h49 == _T_375[7:0] ? 4'hf : _GEN_4881; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4883 = 8'h4a == _T_375[7:0] ? 4'hf : _GEN_4882; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4884 = 8'h4b == _T_375[7:0] ? 4'hf : _GEN_4883; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4885 = 8'h4c == _T_375[7:0] ? 4'hf : _GEN_4884; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4886 = 8'h4d == _T_375[7:0] ? 4'hf : _GEN_4885; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4887 = 8'h4e == _T_375[7:0] ? 4'hf : _GEN_4886; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4888 = 8'h4f == _T_375[7:0] ? 4'hf : _GEN_4887; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4889 = 8'h50 == _T_375[7:0] ? 4'h0 : _GEN_4888; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4890 = 8'h51 == _T_375[7:0] ? 4'h0 : _GEN_4889; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4891 = 8'h52 == _T_375[7:0] ? 4'h0 : _GEN_4890; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4892 = 8'h53 == _T_375[7:0] ? 4'h0 : _GEN_4891; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4893 = 8'h54 == _T_375[7:0] ? 4'h0 : _GEN_4892; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4894 = 8'h55 == _T_375[7:0] ? 4'h0 : _GEN_4893; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4895 = 8'h56 == _T_375[7:0] ? 4'h0 : _GEN_4894; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4896 = 8'h57 == _T_375[7:0] ? 4'h0 : _GEN_4895; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4897 = 8'h58 == _T_375[7:0] ? 4'hf : _GEN_4896; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4898 = 8'h59 == _T_375[7:0] ? 4'hf : _GEN_4897; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4899 = 8'h5a == _T_375[7:0] ? 4'hf : _GEN_4898; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4900 = 8'h5b == _T_375[7:0] ? 4'hf : _GEN_4899; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4901 = 8'h5c == _T_375[7:0] ? 4'hf : _GEN_4900; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4902 = 8'h5d == _T_375[7:0] ? 4'hf : _GEN_4901; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4903 = 8'h5e == _T_375[7:0] ? 4'hf : _GEN_4902; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4904 = 8'h5f == _T_375[7:0] ? 4'hf : _GEN_4903; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4905 = 8'h60 == _T_375[7:0] ? 4'h0 : _GEN_4904; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4906 = 8'h61 == _T_375[7:0] ? 4'h0 : _GEN_4905; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4907 = 8'h62 == _T_375[7:0] ? 4'h0 : _GEN_4906; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4908 = 8'h63 == _T_375[7:0] ? 4'h0 : _GEN_4907; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4909 = 8'h64 == _T_375[7:0] ? 4'h0 : _GEN_4908; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4910 = 8'h65 == _T_375[7:0] ? 4'h0 : _GEN_4909; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4911 = 8'h66 == _T_375[7:0] ? 4'h0 : _GEN_4910; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4912 = 8'h67 == _T_375[7:0] ? 4'h0 : _GEN_4911; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4913 = 8'h68 == _T_375[7:0] ? 4'hf : _GEN_4912; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4914 = 8'h69 == _T_375[7:0] ? 4'hf : _GEN_4913; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4915 = 8'h6a == _T_375[7:0] ? 4'hf : _GEN_4914; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4916 = 8'h6b == _T_375[7:0] ? 4'hf : _GEN_4915; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4917 = 8'h6c == _T_375[7:0] ? 4'hf : _GEN_4916; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4918 = 8'h6d == _T_375[7:0] ? 4'hf : _GEN_4917; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4919 = 8'h6e == _T_375[7:0] ? 4'hf : _GEN_4918; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4920 = 8'h6f == _T_375[7:0] ? 4'hf : _GEN_4919; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4921 = 8'h70 == _T_375[7:0] ? 4'h0 : _GEN_4920; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4922 = 8'h71 == _T_375[7:0] ? 4'h0 : _GEN_4921; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4923 = 8'h72 == _T_375[7:0] ? 4'h0 : _GEN_4922; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4924 = 8'h73 == _T_375[7:0] ? 4'h0 : _GEN_4923; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4925 = 8'h74 == _T_375[7:0] ? 4'h0 : _GEN_4924; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4926 = 8'h75 == _T_375[7:0] ? 4'h0 : _GEN_4925; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4927 = 8'h76 == _T_375[7:0] ? 4'h0 : _GEN_4926; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4928 = 8'h77 == _T_375[7:0] ? 4'h0 : _GEN_4927; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4929 = 8'h78 == _T_375[7:0] ? 4'hf : _GEN_4928; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4930 = 8'h79 == _T_375[7:0] ? 4'hf : _GEN_4929; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4931 = 8'h7a == _T_375[7:0] ? 4'hf : _GEN_4930; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4932 = 8'h7b == _T_375[7:0] ? 4'hf : _GEN_4931; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4933 = 8'h7c == _T_375[7:0] ? 4'hf : _GEN_4932; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4934 = 8'h7d == _T_375[7:0] ? 4'hf : _GEN_4933; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4935 = 8'h7e == _T_375[7:0] ? 4'hf : _GEN_4934; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4936 = 8'h7f == _T_375[7:0] ? 4'hf : _GEN_4935; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4937 = 8'h80 == _T_375[7:0] ? 4'h0 : _GEN_4936; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4938 = 8'h81 == _T_375[7:0] ? 4'h0 : _GEN_4937; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4939 = 8'h82 == _T_375[7:0] ? 4'h0 : _GEN_4938; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4940 = 8'h83 == _T_375[7:0] ? 4'h0 : _GEN_4939; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4941 = 8'h84 == _T_375[7:0] ? 4'h0 : _GEN_4940; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4942 = 8'h85 == _T_375[7:0] ? 4'h0 : _GEN_4941; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4943 = 8'h86 == _T_375[7:0] ? 4'h0 : _GEN_4942; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4944 = 8'h87 == _T_375[7:0] ? 4'h0 : _GEN_4943; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4945 = 8'h88 == _T_375[7:0] ? 4'hf : _GEN_4944; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4946 = 8'h89 == _T_375[7:0] ? 4'hf : _GEN_4945; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4947 = 8'h8a == _T_375[7:0] ? 4'hf : _GEN_4946; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4948 = 8'h8b == _T_375[7:0] ? 4'hf : _GEN_4947; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4949 = 8'h8c == _T_375[7:0] ? 4'hf : _GEN_4948; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4950 = 8'h8d == _T_375[7:0] ? 4'hf : _GEN_4949; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4951 = 8'h8e == _T_375[7:0] ? 4'hf : _GEN_4950; // @[Filter.scala 196:142]
  wire [3:0] _GEN_4952 = 8'h8f == _T_375[7:0] ? 4'hf : _GEN_4951; // @[Filter.scala 196:142]
  wire [7:0] _T_389 = _GEN_4952 * 4'ha; // @[Filter.scala 196:142]
  wire [10:0] _GEN_7627 = {{3'd0}, _T_389}; // @[Filter.scala 196:109]
  wire [10:0] _T_391 = _T_384 + _GEN_7627; // @[Filter.scala 196:109]
  wire [10:0] _T_392 = _T_391 / 11'h64; // @[Filter.scala 196:150]
  wire  _T_394 = _T_365 >= 5'h10; // @[Filter.scala 199:31]
  wire  _T_398 = _T_372 >= 32'h9; // @[Filter.scala 199:63]
  wire  _T_399 = _T_394 | _T_398; // @[Filter.scala 199:58]
  wire [10:0] _GEN_5097 = io_SPI_distort ? _T_392 : {{7'd0}, _GEN_4664}; // @[Filter.scala 201:35]
  wire [10:0] _GEN_5098 = _T_399 ? 11'h0 : _GEN_5097; // @[Filter.scala 199:80]
  wire [10:0] _GEN_5243 = io_SPI_distort ? _T_392 : {{7'd0}, _GEN_4808}; // @[Filter.scala 201:35]
  wire [10:0] _GEN_5244 = _T_399 ? 11'h0 : _GEN_5243; // @[Filter.scala 199:80]
  wire [10:0] _GEN_5389 = io_SPI_distort ? _T_392 : {{7'd0}, _GEN_4952}; // @[Filter.scala 201:35]
  wire [10:0] _GEN_5390 = _T_399 ? 11'h0 : _GEN_5389; // @[Filter.scala 199:80]
  wire [31:0] _T_427 = pixelIndex + 32'h6; // @[Filter.scala 194:31]
  wire [31:0] _GEN_6 = _T_427 % 32'h10; // @[Filter.scala 194:38]
  wire [4:0] _T_428 = _GEN_6[4:0]; // @[Filter.scala 194:38]
  wire [4:0] _T_430 = _T_428 + _GEN_7559; // @[Filter.scala 194:53]
  wire [4:0] _T_432 = _T_430 - 5'h1; // @[Filter.scala 194:69]
  wire [31:0] _T_435 = _T_427 / 32'h10; // @[Filter.scala 195:38]
  wire [31:0] _T_437 = _T_435 + _GEN_7560; // @[Filter.scala 195:53]
  wire [31:0] _T_439 = _T_437 - 32'h1; // @[Filter.scala 195:69]
  wire [36:0] _T_440 = _T_439 * 32'h10; // @[Filter.scala 196:42]
  wire [36:0] _GEN_7633 = {{32'd0}, _T_432}; // @[Filter.scala 196:57]
  wire [36:0] _T_442 = _T_440 + _GEN_7633; // @[Filter.scala 196:57]
  wire [3:0] _GEN_5399 = 8'h8 == _T_442[7:0] ? 4'h0 : 4'hf; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5400 = 8'h9 == _T_442[7:0] ? 4'h0 : _GEN_5399; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5401 = 8'ha == _T_442[7:0] ? 4'h0 : _GEN_5400; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5402 = 8'hb == _T_442[7:0] ? 4'h0 : _GEN_5401; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5403 = 8'hc == _T_442[7:0] ? 4'h0 : _GEN_5402; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5404 = 8'hd == _T_442[7:0] ? 4'h0 : _GEN_5403; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5405 = 8'he == _T_442[7:0] ? 4'h0 : _GEN_5404; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5406 = 8'hf == _T_442[7:0] ? 4'h0 : _GEN_5405; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5407 = 8'h10 == _T_442[7:0] ? 4'hf : _GEN_5406; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5408 = 8'h11 == _T_442[7:0] ? 4'hf : _GEN_5407; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5409 = 8'h12 == _T_442[7:0] ? 4'hf : _GEN_5408; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5410 = 8'h13 == _T_442[7:0] ? 4'hf : _GEN_5409; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5411 = 8'h14 == _T_442[7:0] ? 4'hf : _GEN_5410; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5412 = 8'h15 == _T_442[7:0] ? 4'hf : _GEN_5411; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5413 = 8'h16 == _T_442[7:0] ? 4'hf : _GEN_5412; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5414 = 8'h17 == _T_442[7:0] ? 4'hf : _GEN_5413; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5415 = 8'h18 == _T_442[7:0] ? 4'h0 : _GEN_5414; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5416 = 8'h19 == _T_442[7:0] ? 4'h0 : _GEN_5415; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5417 = 8'h1a == _T_442[7:0] ? 4'h0 : _GEN_5416; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5418 = 8'h1b == _T_442[7:0] ? 4'h0 : _GEN_5417; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5419 = 8'h1c == _T_442[7:0] ? 4'h0 : _GEN_5418; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5420 = 8'h1d == _T_442[7:0] ? 4'h0 : _GEN_5419; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5421 = 8'h1e == _T_442[7:0] ? 4'h0 : _GEN_5420; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5422 = 8'h1f == _T_442[7:0] ? 4'h0 : _GEN_5421; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5423 = 8'h20 == _T_442[7:0] ? 4'hf : _GEN_5422; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5424 = 8'h21 == _T_442[7:0] ? 4'hf : _GEN_5423; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5425 = 8'h22 == _T_442[7:0] ? 4'hf : _GEN_5424; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5426 = 8'h23 == _T_442[7:0] ? 4'hf : _GEN_5425; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5427 = 8'h24 == _T_442[7:0] ? 4'hf : _GEN_5426; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5428 = 8'h25 == _T_442[7:0] ? 4'hf : _GEN_5427; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5429 = 8'h26 == _T_442[7:0] ? 4'hf : _GEN_5428; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5430 = 8'h27 == _T_442[7:0] ? 4'hf : _GEN_5429; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5431 = 8'h28 == _T_442[7:0] ? 4'h0 : _GEN_5430; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5432 = 8'h29 == _T_442[7:0] ? 4'h0 : _GEN_5431; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5433 = 8'h2a == _T_442[7:0] ? 4'h0 : _GEN_5432; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5434 = 8'h2b == _T_442[7:0] ? 4'h0 : _GEN_5433; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5435 = 8'h2c == _T_442[7:0] ? 4'h0 : _GEN_5434; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5436 = 8'h2d == _T_442[7:0] ? 4'h0 : _GEN_5435; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5437 = 8'h2e == _T_442[7:0] ? 4'h0 : _GEN_5436; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5438 = 8'h2f == _T_442[7:0] ? 4'h0 : _GEN_5437; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5439 = 8'h30 == _T_442[7:0] ? 4'hf : _GEN_5438; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5440 = 8'h31 == _T_442[7:0] ? 4'hf : _GEN_5439; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5441 = 8'h32 == _T_442[7:0] ? 4'hf : _GEN_5440; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5442 = 8'h33 == _T_442[7:0] ? 4'hf : _GEN_5441; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5443 = 8'h34 == _T_442[7:0] ? 4'hf : _GEN_5442; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5444 = 8'h35 == _T_442[7:0] ? 4'hf : _GEN_5443; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5445 = 8'h36 == _T_442[7:0] ? 4'hf : _GEN_5444; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5446 = 8'h37 == _T_442[7:0] ? 4'hf : _GEN_5445; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5447 = 8'h38 == _T_442[7:0] ? 4'h0 : _GEN_5446; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5448 = 8'h39 == _T_442[7:0] ? 4'h0 : _GEN_5447; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5449 = 8'h3a == _T_442[7:0] ? 4'h0 : _GEN_5448; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5450 = 8'h3b == _T_442[7:0] ? 4'h0 : _GEN_5449; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5451 = 8'h3c == _T_442[7:0] ? 4'h0 : _GEN_5450; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5452 = 8'h3d == _T_442[7:0] ? 4'h0 : _GEN_5451; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5453 = 8'h3e == _T_442[7:0] ? 4'h0 : _GEN_5452; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5454 = 8'h3f == _T_442[7:0] ? 4'h0 : _GEN_5453; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5455 = 8'h40 == _T_442[7:0] ? 4'h0 : _GEN_5454; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5456 = 8'h41 == _T_442[7:0] ? 4'h0 : _GEN_5455; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5457 = 8'h42 == _T_442[7:0] ? 4'h0 : _GEN_5456; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5458 = 8'h43 == _T_442[7:0] ? 4'h0 : _GEN_5457; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5459 = 8'h44 == _T_442[7:0] ? 4'h0 : _GEN_5458; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5460 = 8'h45 == _T_442[7:0] ? 4'h0 : _GEN_5459; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5461 = 8'h46 == _T_442[7:0] ? 4'h0 : _GEN_5460; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5462 = 8'h47 == _T_442[7:0] ? 4'h0 : _GEN_5461; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5463 = 8'h48 == _T_442[7:0] ? 4'hf : _GEN_5462; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5464 = 8'h49 == _T_442[7:0] ? 4'hf : _GEN_5463; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5465 = 8'h4a == _T_442[7:0] ? 4'hf : _GEN_5464; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5466 = 8'h4b == _T_442[7:0] ? 4'hf : _GEN_5465; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5467 = 8'h4c == _T_442[7:0] ? 4'hf : _GEN_5466; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5468 = 8'h4d == _T_442[7:0] ? 4'hf : _GEN_5467; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5469 = 8'h4e == _T_442[7:0] ? 4'hf : _GEN_5468; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5470 = 8'h4f == _T_442[7:0] ? 4'hf : _GEN_5469; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5471 = 8'h50 == _T_442[7:0] ? 4'h0 : _GEN_5470; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5472 = 8'h51 == _T_442[7:0] ? 4'h0 : _GEN_5471; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5473 = 8'h52 == _T_442[7:0] ? 4'h0 : _GEN_5472; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5474 = 8'h53 == _T_442[7:0] ? 4'h0 : _GEN_5473; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5475 = 8'h54 == _T_442[7:0] ? 4'h0 : _GEN_5474; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5476 = 8'h55 == _T_442[7:0] ? 4'h0 : _GEN_5475; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5477 = 8'h56 == _T_442[7:0] ? 4'h0 : _GEN_5476; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5478 = 8'h57 == _T_442[7:0] ? 4'h0 : _GEN_5477; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5479 = 8'h58 == _T_442[7:0] ? 4'hf : _GEN_5478; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5480 = 8'h59 == _T_442[7:0] ? 4'hf : _GEN_5479; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5481 = 8'h5a == _T_442[7:0] ? 4'hf : _GEN_5480; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5482 = 8'h5b == _T_442[7:0] ? 4'hf : _GEN_5481; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5483 = 8'h5c == _T_442[7:0] ? 4'hf : _GEN_5482; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5484 = 8'h5d == _T_442[7:0] ? 4'hf : _GEN_5483; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5485 = 8'h5e == _T_442[7:0] ? 4'hf : _GEN_5484; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5486 = 8'h5f == _T_442[7:0] ? 4'hf : _GEN_5485; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5487 = 8'h60 == _T_442[7:0] ? 4'h0 : _GEN_5486; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5488 = 8'h61 == _T_442[7:0] ? 4'h0 : _GEN_5487; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5489 = 8'h62 == _T_442[7:0] ? 4'h0 : _GEN_5488; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5490 = 8'h63 == _T_442[7:0] ? 4'h0 : _GEN_5489; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5491 = 8'h64 == _T_442[7:0] ? 4'h0 : _GEN_5490; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5492 = 8'h65 == _T_442[7:0] ? 4'h0 : _GEN_5491; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5493 = 8'h66 == _T_442[7:0] ? 4'h0 : _GEN_5492; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5494 = 8'h67 == _T_442[7:0] ? 4'h0 : _GEN_5493; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5495 = 8'h68 == _T_442[7:0] ? 4'hf : _GEN_5494; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5496 = 8'h69 == _T_442[7:0] ? 4'hf : _GEN_5495; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5497 = 8'h6a == _T_442[7:0] ? 4'hf : _GEN_5496; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5498 = 8'h6b == _T_442[7:0] ? 4'hf : _GEN_5497; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5499 = 8'h6c == _T_442[7:0] ? 4'hf : _GEN_5498; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5500 = 8'h6d == _T_442[7:0] ? 4'hf : _GEN_5499; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5501 = 8'h6e == _T_442[7:0] ? 4'hf : _GEN_5500; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5502 = 8'h6f == _T_442[7:0] ? 4'hf : _GEN_5501; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5503 = 8'h70 == _T_442[7:0] ? 4'h0 : _GEN_5502; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5504 = 8'h71 == _T_442[7:0] ? 4'h0 : _GEN_5503; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5505 = 8'h72 == _T_442[7:0] ? 4'h0 : _GEN_5504; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5506 = 8'h73 == _T_442[7:0] ? 4'h0 : _GEN_5505; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5507 = 8'h74 == _T_442[7:0] ? 4'h0 : _GEN_5506; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5508 = 8'h75 == _T_442[7:0] ? 4'h0 : _GEN_5507; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5509 = 8'h76 == _T_442[7:0] ? 4'h0 : _GEN_5508; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5510 = 8'h77 == _T_442[7:0] ? 4'h0 : _GEN_5509; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5511 = 8'h78 == _T_442[7:0] ? 4'hf : _GEN_5510; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5512 = 8'h79 == _T_442[7:0] ? 4'hf : _GEN_5511; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5513 = 8'h7a == _T_442[7:0] ? 4'hf : _GEN_5512; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5514 = 8'h7b == _T_442[7:0] ? 4'hf : _GEN_5513; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5515 = 8'h7c == _T_442[7:0] ? 4'hf : _GEN_5514; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5516 = 8'h7d == _T_442[7:0] ? 4'hf : _GEN_5515; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5517 = 8'h7e == _T_442[7:0] ? 4'hf : _GEN_5516; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5518 = 8'h7f == _T_442[7:0] ? 4'hf : _GEN_5517; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5519 = 8'h80 == _T_442[7:0] ? 4'h0 : _GEN_5518; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5520 = 8'h81 == _T_442[7:0] ? 4'h0 : _GEN_5519; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5521 = 8'h82 == _T_442[7:0] ? 4'h0 : _GEN_5520; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5522 = 8'h83 == _T_442[7:0] ? 4'h0 : _GEN_5521; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5523 = 8'h84 == _T_442[7:0] ? 4'h0 : _GEN_5522; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5524 = 8'h85 == _T_442[7:0] ? 4'h0 : _GEN_5523; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5525 = 8'h86 == _T_442[7:0] ? 4'h0 : _GEN_5524; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5526 = 8'h87 == _T_442[7:0] ? 4'h0 : _GEN_5525; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5527 = 8'h88 == _T_442[7:0] ? 4'hf : _GEN_5526; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5528 = 8'h89 == _T_442[7:0] ? 4'hf : _GEN_5527; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5529 = 8'h8a == _T_442[7:0] ? 4'hf : _GEN_5528; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5530 = 8'h8b == _T_442[7:0] ? 4'hf : _GEN_5529; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5531 = 8'h8c == _T_442[7:0] ? 4'hf : _GEN_5530; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5532 = 8'h8d == _T_442[7:0] ? 4'hf : _GEN_5531; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5533 = 8'h8e == _T_442[7:0] ? 4'hf : _GEN_5532; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5534 = 8'h8f == _T_442[7:0] ? 4'hf : _GEN_5533; // @[Filter.scala 196:62]
  wire [4:0] _GEN_7634 = {{1'd0}, _GEN_5534}; // @[Filter.scala 196:62]
  wire [8:0] _T_444 = _GEN_7634 * 5'h14; // @[Filter.scala 196:62]
  wire [3:0] _GEN_5599 = 8'h40 == _T_442[7:0] ? 4'hf : 4'h0; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5600 = 8'h41 == _T_442[7:0] ? 4'hf : _GEN_5599; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5601 = 8'h42 == _T_442[7:0] ? 4'hf : _GEN_5600; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5602 = 8'h43 == _T_442[7:0] ? 4'hf : _GEN_5601; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5603 = 8'h44 == _T_442[7:0] ? 4'hf : _GEN_5602; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5604 = 8'h45 == _T_442[7:0] ? 4'hf : _GEN_5603; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5605 = 8'h46 == _T_442[7:0] ? 4'hf : _GEN_5604; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5606 = 8'h47 == _T_442[7:0] ? 4'hf : _GEN_5605; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5607 = 8'h48 == _T_442[7:0] ? 4'hf : _GEN_5606; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5608 = 8'h49 == _T_442[7:0] ? 4'hf : _GEN_5607; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5609 = 8'h4a == _T_442[7:0] ? 4'hf : _GEN_5608; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5610 = 8'h4b == _T_442[7:0] ? 4'hf : _GEN_5609; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5611 = 8'h4c == _T_442[7:0] ? 4'hf : _GEN_5610; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5612 = 8'h4d == _T_442[7:0] ? 4'hf : _GEN_5611; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5613 = 8'h4e == _T_442[7:0] ? 4'hf : _GEN_5612; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5614 = 8'h4f == _T_442[7:0] ? 4'hf : _GEN_5613; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5615 = 8'h50 == _T_442[7:0] ? 4'hf : _GEN_5614; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5616 = 8'h51 == _T_442[7:0] ? 4'hf : _GEN_5615; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5617 = 8'h52 == _T_442[7:0] ? 4'hf : _GEN_5616; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5618 = 8'h53 == _T_442[7:0] ? 4'hf : _GEN_5617; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5619 = 8'h54 == _T_442[7:0] ? 4'hf : _GEN_5618; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5620 = 8'h55 == _T_442[7:0] ? 4'hf : _GEN_5619; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5621 = 8'h56 == _T_442[7:0] ? 4'hf : _GEN_5620; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5622 = 8'h57 == _T_442[7:0] ? 4'hf : _GEN_5621; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5623 = 8'h58 == _T_442[7:0] ? 4'hf : _GEN_5622; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5624 = 8'h59 == _T_442[7:0] ? 4'hf : _GEN_5623; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5625 = 8'h5a == _T_442[7:0] ? 4'hf : _GEN_5624; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5626 = 8'h5b == _T_442[7:0] ? 4'hf : _GEN_5625; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5627 = 8'h5c == _T_442[7:0] ? 4'hf : _GEN_5626; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5628 = 8'h5d == _T_442[7:0] ? 4'hf : _GEN_5627; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5629 = 8'h5e == _T_442[7:0] ? 4'hf : _GEN_5628; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5630 = 8'h5f == _T_442[7:0] ? 4'hf : _GEN_5629; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5631 = 8'h60 == _T_442[7:0] ? 4'hf : _GEN_5630; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5632 = 8'h61 == _T_442[7:0] ? 4'hf : _GEN_5631; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5633 = 8'h62 == _T_442[7:0] ? 4'hf : _GEN_5632; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5634 = 8'h63 == _T_442[7:0] ? 4'hf : _GEN_5633; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5635 = 8'h64 == _T_442[7:0] ? 4'hf : _GEN_5634; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5636 = 8'h65 == _T_442[7:0] ? 4'hf : _GEN_5635; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5637 = 8'h66 == _T_442[7:0] ? 4'hf : _GEN_5636; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5638 = 8'h67 == _T_442[7:0] ? 4'hf : _GEN_5637; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5639 = 8'h68 == _T_442[7:0] ? 4'hf : _GEN_5638; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5640 = 8'h69 == _T_442[7:0] ? 4'hf : _GEN_5639; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5641 = 8'h6a == _T_442[7:0] ? 4'hf : _GEN_5640; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5642 = 8'h6b == _T_442[7:0] ? 4'hf : _GEN_5641; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5643 = 8'h6c == _T_442[7:0] ? 4'hf : _GEN_5642; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5644 = 8'h6d == _T_442[7:0] ? 4'hf : _GEN_5643; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5645 = 8'h6e == _T_442[7:0] ? 4'hf : _GEN_5644; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5646 = 8'h6f == _T_442[7:0] ? 4'hf : _GEN_5645; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5647 = 8'h70 == _T_442[7:0] ? 4'hf : _GEN_5646; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5648 = 8'h71 == _T_442[7:0] ? 4'hf : _GEN_5647; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5649 = 8'h72 == _T_442[7:0] ? 4'hf : _GEN_5648; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5650 = 8'h73 == _T_442[7:0] ? 4'hf : _GEN_5649; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5651 = 8'h74 == _T_442[7:0] ? 4'hf : _GEN_5650; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5652 = 8'h75 == _T_442[7:0] ? 4'hf : _GEN_5651; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5653 = 8'h76 == _T_442[7:0] ? 4'hf : _GEN_5652; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5654 = 8'h77 == _T_442[7:0] ? 4'hf : _GEN_5653; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5655 = 8'h78 == _T_442[7:0] ? 4'hf : _GEN_5654; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5656 = 8'h79 == _T_442[7:0] ? 4'hf : _GEN_5655; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5657 = 8'h7a == _T_442[7:0] ? 4'hf : _GEN_5656; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5658 = 8'h7b == _T_442[7:0] ? 4'hf : _GEN_5657; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5659 = 8'h7c == _T_442[7:0] ? 4'hf : _GEN_5658; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5660 = 8'h7d == _T_442[7:0] ? 4'hf : _GEN_5659; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5661 = 8'h7e == _T_442[7:0] ? 4'hf : _GEN_5660; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5662 = 8'h7f == _T_442[7:0] ? 4'hf : _GEN_5661; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5663 = 8'h80 == _T_442[7:0] ? 4'hf : _GEN_5662; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5664 = 8'h81 == _T_442[7:0] ? 4'hf : _GEN_5663; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5665 = 8'h82 == _T_442[7:0] ? 4'hf : _GEN_5664; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5666 = 8'h83 == _T_442[7:0] ? 4'hf : _GEN_5665; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5667 = 8'h84 == _T_442[7:0] ? 4'hf : _GEN_5666; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5668 = 8'h85 == _T_442[7:0] ? 4'hf : _GEN_5667; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5669 = 8'h86 == _T_442[7:0] ? 4'hf : _GEN_5668; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5670 = 8'h87 == _T_442[7:0] ? 4'hf : _GEN_5669; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5671 = 8'h88 == _T_442[7:0] ? 4'hf : _GEN_5670; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5672 = 8'h89 == _T_442[7:0] ? 4'hf : _GEN_5671; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5673 = 8'h8a == _T_442[7:0] ? 4'hf : _GEN_5672; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5674 = 8'h8b == _T_442[7:0] ? 4'hf : _GEN_5673; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5675 = 8'h8c == _T_442[7:0] ? 4'hf : _GEN_5674; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5676 = 8'h8d == _T_442[7:0] ? 4'hf : _GEN_5675; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5677 = 8'h8e == _T_442[7:0] ? 4'hf : _GEN_5676; // @[Filter.scala 196:102]
  wire [3:0] _GEN_5678 = 8'h8f == _T_442[7:0] ? 4'hf : _GEN_5677; // @[Filter.scala 196:102]
  wire [6:0] _GEN_7636 = {{3'd0}, _GEN_5678}; // @[Filter.scala 196:102]
  wire [10:0] _T_449 = _GEN_7636 * 7'h46; // @[Filter.scala 196:102]
  wire [10:0] _GEN_7637 = {{2'd0}, _T_444}; // @[Filter.scala 196:69]
  wire [10:0] _T_451 = _GEN_7637 + _T_449; // @[Filter.scala 196:69]
  wire [3:0] _GEN_5687 = 8'h8 == _T_442[7:0] ? 4'hf : 4'h0; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5688 = 8'h9 == _T_442[7:0] ? 4'hf : _GEN_5687; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5689 = 8'ha == _T_442[7:0] ? 4'hf : _GEN_5688; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5690 = 8'hb == _T_442[7:0] ? 4'hf : _GEN_5689; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5691 = 8'hc == _T_442[7:0] ? 4'hf : _GEN_5690; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5692 = 8'hd == _T_442[7:0] ? 4'hf : _GEN_5691; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5693 = 8'he == _T_442[7:0] ? 4'hf : _GEN_5692; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5694 = 8'hf == _T_442[7:0] ? 4'hf : _GEN_5693; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5695 = 8'h10 == _T_442[7:0] ? 4'h0 : _GEN_5694; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5696 = 8'h11 == _T_442[7:0] ? 4'h0 : _GEN_5695; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5697 = 8'h12 == _T_442[7:0] ? 4'h0 : _GEN_5696; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5698 = 8'h13 == _T_442[7:0] ? 4'h0 : _GEN_5697; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5699 = 8'h14 == _T_442[7:0] ? 4'h0 : _GEN_5698; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5700 = 8'h15 == _T_442[7:0] ? 4'h0 : _GEN_5699; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5701 = 8'h16 == _T_442[7:0] ? 4'h0 : _GEN_5700; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5702 = 8'h17 == _T_442[7:0] ? 4'h0 : _GEN_5701; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5703 = 8'h18 == _T_442[7:0] ? 4'hf : _GEN_5702; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5704 = 8'h19 == _T_442[7:0] ? 4'hf : _GEN_5703; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5705 = 8'h1a == _T_442[7:0] ? 4'hf : _GEN_5704; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5706 = 8'h1b == _T_442[7:0] ? 4'hf : _GEN_5705; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5707 = 8'h1c == _T_442[7:0] ? 4'hf : _GEN_5706; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5708 = 8'h1d == _T_442[7:0] ? 4'hf : _GEN_5707; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5709 = 8'h1e == _T_442[7:0] ? 4'hf : _GEN_5708; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5710 = 8'h1f == _T_442[7:0] ? 4'hf : _GEN_5709; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5711 = 8'h20 == _T_442[7:0] ? 4'h0 : _GEN_5710; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5712 = 8'h21 == _T_442[7:0] ? 4'h0 : _GEN_5711; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5713 = 8'h22 == _T_442[7:0] ? 4'h0 : _GEN_5712; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5714 = 8'h23 == _T_442[7:0] ? 4'h0 : _GEN_5713; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5715 = 8'h24 == _T_442[7:0] ? 4'h0 : _GEN_5714; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5716 = 8'h25 == _T_442[7:0] ? 4'h0 : _GEN_5715; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5717 = 8'h26 == _T_442[7:0] ? 4'h0 : _GEN_5716; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5718 = 8'h27 == _T_442[7:0] ? 4'h0 : _GEN_5717; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5719 = 8'h28 == _T_442[7:0] ? 4'hf : _GEN_5718; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5720 = 8'h29 == _T_442[7:0] ? 4'hf : _GEN_5719; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5721 = 8'h2a == _T_442[7:0] ? 4'hf : _GEN_5720; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5722 = 8'h2b == _T_442[7:0] ? 4'hf : _GEN_5721; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5723 = 8'h2c == _T_442[7:0] ? 4'hf : _GEN_5722; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5724 = 8'h2d == _T_442[7:0] ? 4'hf : _GEN_5723; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5725 = 8'h2e == _T_442[7:0] ? 4'hf : _GEN_5724; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5726 = 8'h2f == _T_442[7:0] ? 4'hf : _GEN_5725; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5727 = 8'h30 == _T_442[7:0] ? 4'h0 : _GEN_5726; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5728 = 8'h31 == _T_442[7:0] ? 4'h0 : _GEN_5727; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5729 = 8'h32 == _T_442[7:0] ? 4'h0 : _GEN_5728; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5730 = 8'h33 == _T_442[7:0] ? 4'h0 : _GEN_5729; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5731 = 8'h34 == _T_442[7:0] ? 4'h0 : _GEN_5730; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5732 = 8'h35 == _T_442[7:0] ? 4'h0 : _GEN_5731; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5733 = 8'h36 == _T_442[7:0] ? 4'h0 : _GEN_5732; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5734 = 8'h37 == _T_442[7:0] ? 4'h0 : _GEN_5733; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5735 = 8'h38 == _T_442[7:0] ? 4'hf : _GEN_5734; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5736 = 8'h39 == _T_442[7:0] ? 4'hf : _GEN_5735; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5737 = 8'h3a == _T_442[7:0] ? 4'hf : _GEN_5736; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5738 = 8'h3b == _T_442[7:0] ? 4'hf : _GEN_5737; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5739 = 8'h3c == _T_442[7:0] ? 4'hf : _GEN_5738; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5740 = 8'h3d == _T_442[7:0] ? 4'hf : _GEN_5739; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5741 = 8'h3e == _T_442[7:0] ? 4'hf : _GEN_5740; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5742 = 8'h3f == _T_442[7:0] ? 4'hf : _GEN_5741; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5743 = 8'h40 == _T_442[7:0] ? 4'h0 : _GEN_5742; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5744 = 8'h41 == _T_442[7:0] ? 4'h0 : _GEN_5743; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5745 = 8'h42 == _T_442[7:0] ? 4'h0 : _GEN_5744; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5746 = 8'h43 == _T_442[7:0] ? 4'h0 : _GEN_5745; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5747 = 8'h44 == _T_442[7:0] ? 4'h0 : _GEN_5746; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5748 = 8'h45 == _T_442[7:0] ? 4'h0 : _GEN_5747; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5749 = 8'h46 == _T_442[7:0] ? 4'h0 : _GEN_5748; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5750 = 8'h47 == _T_442[7:0] ? 4'h0 : _GEN_5749; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5751 = 8'h48 == _T_442[7:0] ? 4'hf : _GEN_5750; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5752 = 8'h49 == _T_442[7:0] ? 4'hf : _GEN_5751; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5753 = 8'h4a == _T_442[7:0] ? 4'hf : _GEN_5752; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5754 = 8'h4b == _T_442[7:0] ? 4'hf : _GEN_5753; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5755 = 8'h4c == _T_442[7:0] ? 4'hf : _GEN_5754; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5756 = 8'h4d == _T_442[7:0] ? 4'hf : _GEN_5755; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5757 = 8'h4e == _T_442[7:0] ? 4'hf : _GEN_5756; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5758 = 8'h4f == _T_442[7:0] ? 4'hf : _GEN_5757; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5759 = 8'h50 == _T_442[7:0] ? 4'h0 : _GEN_5758; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5760 = 8'h51 == _T_442[7:0] ? 4'h0 : _GEN_5759; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5761 = 8'h52 == _T_442[7:0] ? 4'h0 : _GEN_5760; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5762 = 8'h53 == _T_442[7:0] ? 4'h0 : _GEN_5761; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5763 = 8'h54 == _T_442[7:0] ? 4'h0 : _GEN_5762; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5764 = 8'h55 == _T_442[7:0] ? 4'h0 : _GEN_5763; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5765 = 8'h56 == _T_442[7:0] ? 4'h0 : _GEN_5764; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5766 = 8'h57 == _T_442[7:0] ? 4'h0 : _GEN_5765; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5767 = 8'h58 == _T_442[7:0] ? 4'hf : _GEN_5766; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5768 = 8'h59 == _T_442[7:0] ? 4'hf : _GEN_5767; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5769 = 8'h5a == _T_442[7:0] ? 4'hf : _GEN_5768; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5770 = 8'h5b == _T_442[7:0] ? 4'hf : _GEN_5769; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5771 = 8'h5c == _T_442[7:0] ? 4'hf : _GEN_5770; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5772 = 8'h5d == _T_442[7:0] ? 4'hf : _GEN_5771; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5773 = 8'h5e == _T_442[7:0] ? 4'hf : _GEN_5772; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5774 = 8'h5f == _T_442[7:0] ? 4'hf : _GEN_5773; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5775 = 8'h60 == _T_442[7:0] ? 4'h0 : _GEN_5774; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5776 = 8'h61 == _T_442[7:0] ? 4'h0 : _GEN_5775; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5777 = 8'h62 == _T_442[7:0] ? 4'h0 : _GEN_5776; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5778 = 8'h63 == _T_442[7:0] ? 4'h0 : _GEN_5777; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5779 = 8'h64 == _T_442[7:0] ? 4'h0 : _GEN_5778; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5780 = 8'h65 == _T_442[7:0] ? 4'h0 : _GEN_5779; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5781 = 8'h66 == _T_442[7:0] ? 4'h0 : _GEN_5780; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5782 = 8'h67 == _T_442[7:0] ? 4'h0 : _GEN_5781; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5783 = 8'h68 == _T_442[7:0] ? 4'hf : _GEN_5782; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5784 = 8'h69 == _T_442[7:0] ? 4'hf : _GEN_5783; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5785 = 8'h6a == _T_442[7:0] ? 4'hf : _GEN_5784; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5786 = 8'h6b == _T_442[7:0] ? 4'hf : _GEN_5785; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5787 = 8'h6c == _T_442[7:0] ? 4'hf : _GEN_5786; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5788 = 8'h6d == _T_442[7:0] ? 4'hf : _GEN_5787; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5789 = 8'h6e == _T_442[7:0] ? 4'hf : _GEN_5788; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5790 = 8'h6f == _T_442[7:0] ? 4'hf : _GEN_5789; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5791 = 8'h70 == _T_442[7:0] ? 4'h0 : _GEN_5790; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5792 = 8'h71 == _T_442[7:0] ? 4'h0 : _GEN_5791; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5793 = 8'h72 == _T_442[7:0] ? 4'h0 : _GEN_5792; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5794 = 8'h73 == _T_442[7:0] ? 4'h0 : _GEN_5793; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5795 = 8'h74 == _T_442[7:0] ? 4'h0 : _GEN_5794; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5796 = 8'h75 == _T_442[7:0] ? 4'h0 : _GEN_5795; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5797 = 8'h76 == _T_442[7:0] ? 4'h0 : _GEN_5796; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5798 = 8'h77 == _T_442[7:0] ? 4'h0 : _GEN_5797; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5799 = 8'h78 == _T_442[7:0] ? 4'hf : _GEN_5798; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5800 = 8'h79 == _T_442[7:0] ? 4'hf : _GEN_5799; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5801 = 8'h7a == _T_442[7:0] ? 4'hf : _GEN_5800; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5802 = 8'h7b == _T_442[7:0] ? 4'hf : _GEN_5801; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5803 = 8'h7c == _T_442[7:0] ? 4'hf : _GEN_5802; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5804 = 8'h7d == _T_442[7:0] ? 4'hf : _GEN_5803; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5805 = 8'h7e == _T_442[7:0] ? 4'hf : _GEN_5804; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5806 = 8'h7f == _T_442[7:0] ? 4'hf : _GEN_5805; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5807 = 8'h80 == _T_442[7:0] ? 4'h0 : _GEN_5806; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5808 = 8'h81 == _T_442[7:0] ? 4'h0 : _GEN_5807; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5809 = 8'h82 == _T_442[7:0] ? 4'h0 : _GEN_5808; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5810 = 8'h83 == _T_442[7:0] ? 4'h0 : _GEN_5809; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5811 = 8'h84 == _T_442[7:0] ? 4'h0 : _GEN_5810; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5812 = 8'h85 == _T_442[7:0] ? 4'h0 : _GEN_5811; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5813 = 8'h86 == _T_442[7:0] ? 4'h0 : _GEN_5812; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5814 = 8'h87 == _T_442[7:0] ? 4'h0 : _GEN_5813; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5815 = 8'h88 == _T_442[7:0] ? 4'hf : _GEN_5814; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5816 = 8'h89 == _T_442[7:0] ? 4'hf : _GEN_5815; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5817 = 8'h8a == _T_442[7:0] ? 4'hf : _GEN_5816; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5818 = 8'h8b == _T_442[7:0] ? 4'hf : _GEN_5817; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5819 = 8'h8c == _T_442[7:0] ? 4'hf : _GEN_5818; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5820 = 8'h8d == _T_442[7:0] ? 4'hf : _GEN_5819; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5821 = 8'h8e == _T_442[7:0] ? 4'hf : _GEN_5820; // @[Filter.scala 196:142]
  wire [3:0] _GEN_5822 = 8'h8f == _T_442[7:0] ? 4'hf : _GEN_5821; // @[Filter.scala 196:142]
  wire [7:0] _T_456 = _GEN_5822 * 4'ha; // @[Filter.scala 196:142]
  wire [10:0] _GEN_7639 = {{3'd0}, _T_456}; // @[Filter.scala 196:109]
  wire [10:0] _T_458 = _T_451 + _GEN_7639; // @[Filter.scala 196:109]
  wire [10:0] _T_459 = _T_458 / 11'h64; // @[Filter.scala 196:150]
  wire  _T_461 = _T_432 >= 5'h10; // @[Filter.scala 199:31]
  wire  _T_465 = _T_439 >= 32'h9; // @[Filter.scala 199:63]
  wire  _T_466 = _T_461 | _T_465; // @[Filter.scala 199:58]
  wire [10:0] _GEN_5967 = io_SPI_distort ? _T_459 : {{7'd0}, _GEN_5534}; // @[Filter.scala 201:35]
  wire [10:0] _GEN_5968 = _T_466 ? 11'h0 : _GEN_5967; // @[Filter.scala 199:80]
  wire [10:0] _GEN_6113 = io_SPI_distort ? _T_459 : {{7'd0}, _GEN_5678}; // @[Filter.scala 201:35]
  wire [10:0] _GEN_6114 = _T_466 ? 11'h0 : _GEN_6113; // @[Filter.scala 199:80]
  wire [10:0] _GEN_6259 = io_SPI_distort ? _T_459 : {{7'd0}, _GEN_5822}; // @[Filter.scala 201:35]
  wire [10:0] _GEN_6260 = _T_466 ? 11'h0 : _GEN_6259; // @[Filter.scala 199:80]
  wire [31:0] _T_494 = pixelIndex + 32'h7; // @[Filter.scala 194:31]
  wire [31:0] _GEN_56 = _T_494 % 32'h10; // @[Filter.scala 194:38]
  wire [4:0] _T_495 = _GEN_56[4:0]; // @[Filter.scala 194:38]
  wire [4:0] _T_497 = _T_495 + _GEN_7559; // @[Filter.scala 194:53]
  wire [4:0] _T_499 = _T_497 - 5'h1; // @[Filter.scala 194:69]
  wire [31:0] _T_502 = _T_494 / 32'h10; // @[Filter.scala 195:38]
  wire [31:0] _T_504 = _T_502 + _GEN_7560; // @[Filter.scala 195:53]
  wire [31:0] _T_506 = _T_504 - 32'h1; // @[Filter.scala 195:69]
  wire [36:0] _T_507 = _T_506 * 32'h10; // @[Filter.scala 196:42]
  wire [36:0] _GEN_7645 = {{32'd0}, _T_499}; // @[Filter.scala 196:57]
  wire [36:0] _T_509 = _T_507 + _GEN_7645; // @[Filter.scala 196:57]
  wire [3:0] _GEN_6269 = 8'h8 == _T_509[7:0] ? 4'h0 : 4'hf; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6270 = 8'h9 == _T_509[7:0] ? 4'h0 : _GEN_6269; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6271 = 8'ha == _T_509[7:0] ? 4'h0 : _GEN_6270; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6272 = 8'hb == _T_509[7:0] ? 4'h0 : _GEN_6271; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6273 = 8'hc == _T_509[7:0] ? 4'h0 : _GEN_6272; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6274 = 8'hd == _T_509[7:0] ? 4'h0 : _GEN_6273; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6275 = 8'he == _T_509[7:0] ? 4'h0 : _GEN_6274; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6276 = 8'hf == _T_509[7:0] ? 4'h0 : _GEN_6275; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6277 = 8'h10 == _T_509[7:0] ? 4'hf : _GEN_6276; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6278 = 8'h11 == _T_509[7:0] ? 4'hf : _GEN_6277; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6279 = 8'h12 == _T_509[7:0] ? 4'hf : _GEN_6278; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6280 = 8'h13 == _T_509[7:0] ? 4'hf : _GEN_6279; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6281 = 8'h14 == _T_509[7:0] ? 4'hf : _GEN_6280; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6282 = 8'h15 == _T_509[7:0] ? 4'hf : _GEN_6281; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6283 = 8'h16 == _T_509[7:0] ? 4'hf : _GEN_6282; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6284 = 8'h17 == _T_509[7:0] ? 4'hf : _GEN_6283; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6285 = 8'h18 == _T_509[7:0] ? 4'h0 : _GEN_6284; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6286 = 8'h19 == _T_509[7:0] ? 4'h0 : _GEN_6285; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6287 = 8'h1a == _T_509[7:0] ? 4'h0 : _GEN_6286; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6288 = 8'h1b == _T_509[7:0] ? 4'h0 : _GEN_6287; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6289 = 8'h1c == _T_509[7:0] ? 4'h0 : _GEN_6288; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6290 = 8'h1d == _T_509[7:0] ? 4'h0 : _GEN_6289; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6291 = 8'h1e == _T_509[7:0] ? 4'h0 : _GEN_6290; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6292 = 8'h1f == _T_509[7:0] ? 4'h0 : _GEN_6291; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6293 = 8'h20 == _T_509[7:0] ? 4'hf : _GEN_6292; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6294 = 8'h21 == _T_509[7:0] ? 4'hf : _GEN_6293; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6295 = 8'h22 == _T_509[7:0] ? 4'hf : _GEN_6294; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6296 = 8'h23 == _T_509[7:0] ? 4'hf : _GEN_6295; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6297 = 8'h24 == _T_509[7:0] ? 4'hf : _GEN_6296; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6298 = 8'h25 == _T_509[7:0] ? 4'hf : _GEN_6297; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6299 = 8'h26 == _T_509[7:0] ? 4'hf : _GEN_6298; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6300 = 8'h27 == _T_509[7:0] ? 4'hf : _GEN_6299; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6301 = 8'h28 == _T_509[7:0] ? 4'h0 : _GEN_6300; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6302 = 8'h29 == _T_509[7:0] ? 4'h0 : _GEN_6301; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6303 = 8'h2a == _T_509[7:0] ? 4'h0 : _GEN_6302; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6304 = 8'h2b == _T_509[7:0] ? 4'h0 : _GEN_6303; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6305 = 8'h2c == _T_509[7:0] ? 4'h0 : _GEN_6304; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6306 = 8'h2d == _T_509[7:0] ? 4'h0 : _GEN_6305; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6307 = 8'h2e == _T_509[7:0] ? 4'h0 : _GEN_6306; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6308 = 8'h2f == _T_509[7:0] ? 4'h0 : _GEN_6307; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6309 = 8'h30 == _T_509[7:0] ? 4'hf : _GEN_6308; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6310 = 8'h31 == _T_509[7:0] ? 4'hf : _GEN_6309; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6311 = 8'h32 == _T_509[7:0] ? 4'hf : _GEN_6310; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6312 = 8'h33 == _T_509[7:0] ? 4'hf : _GEN_6311; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6313 = 8'h34 == _T_509[7:0] ? 4'hf : _GEN_6312; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6314 = 8'h35 == _T_509[7:0] ? 4'hf : _GEN_6313; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6315 = 8'h36 == _T_509[7:0] ? 4'hf : _GEN_6314; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6316 = 8'h37 == _T_509[7:0] ? 4'hf : _GEN_6315; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6317 = 8'h38 == _T_509[7:0] ? 4'h0 : _GEN_6316; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6318 = 8'h39 == _T_509[7:0] ? 4'h0 : _GEN_6317; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6319 = 8'h3a == _T_509[7:0] ? 4'h0 : _GEN_6318; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6320 = 8'h3b == _T_509[7:0] ? 4'h0 : _GEN_6319; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6321 = 8'h3c == _T_509[7:0] ? 4'h0 : _GEN_6320; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6322 = 8'h3d == _T_509[7:0] ? 4'h0 : _GEN_6321; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6323 = 8'h3e == _T_509[7:0] ? 4'h0 : _GEN_6322; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6324 = 8'h3f == _T_509[7:0] ? 4'h0 : _GEN_6323; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6325 = 8'h40 == _T_509[7:0] ? 4'h0 : _GEN_6324; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6326 = 8'h41 == _T_509[7:0] ? 4'h0 : _GEN_6325; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6327 = 8'h42 == _T_509[7:0] ? 4'h0 : _GEN_6326; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6328 = 8'h43 == _T_509[7:0] ? 4'h0 : _GEN_6327; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6329 = 8'h44 == _T_509[7:0] ? 4'h0 : _GEN_6328; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6330 = 8'h45 == _T_509[7:0] ? 4'h0 : _GEN_6329; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6331 = 8'h46 == _T_509[7:0] ? 4'h0 : _GEN_6330; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6332 = 8'h47 == _T_509[7:0] ? 4'h0 : _GEN_6331; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6333 = 8'h48 == _T_509[7:0] ? 4'hf : _GEN_6332; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6334 = 8'h49 == _T_509[7:0] ? 4'hf : _GEN_6333; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6335 = 8'h4a == _T_509[7:0] ? 4'hf : _GEN_6334; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6336 = 8'h4b == _T_509[7:0] ? 4'hf : _GEN_6335; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6337 = 8'h4c == _T_509[7:0] ? 4'hf : _GEN_6336; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6338 = 8'h4d == _T_509[7:0] ? 4'hf : _GEN_6337; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6339 = 8'h4e == _T_509[7:0] ? 4'hf : _GEN_6338; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6340 = 8'h4f == _T_509[7:0] ? 4'hf : _GEN_6339; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6341 = 8'h50 == _T_509[7:0] ? 4'h0 : _GEN_6340; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6342 = 8'h51 == _T_509[7:0] ? 4'h0 : _GEN_6341; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6343 = 8'h52 == _T_509[7:0] ? 4'h0 : _GEN_6342; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6344 = 8'h53 == _T_509[7:0] ? 4'h0 : _GEN_6343; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6345 = 8'h54 == _T_509[7:0] ? 4'h0 : _GEN_6344; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6346 = 8'h55 == _T_509[7:0] ? 4'h0 : _GEN_6345; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6347 = 8'h56 == _T_509[7:0] ? 4'h0 : _GEN_6346; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6348 = 8'h57 == _T_509[7:0] ? 4'h0 : _GEN_6347; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6349 = 8'h58 == _T_509[7:0] ? 4'hf : _GEN_6348; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6350 = 8'h59 == _T_509[7:0] ? 4'hf : _GEN_6349; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6351 = 8'h5a == _T_509[7:0] ? 4'hf : _GEN_6350; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6352 = 8'h5b == _T_509[7:0] ? 4'hf : _GEN_6351; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6353 = 8'h5c == _T_509[7:0] ? 4'hf : _GEN_6352; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6354 = 8'h5d == _T_509[7:0] ? 4'hf : _GEN_6353; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6355 = 8'h5e == _T_509[7:0] ? 4'hf : _GEN_6354; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6356 = 8'h5f == _T_509[7:0] ? 4'hf : _GEN_6355; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6357 = 8'h60 == _T_509[7:0] ? 4'h0 : _GEN_6356; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6358 = 8'h61 == _T_509[7:0] ? 4'h0 : _GEN_6357; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6359 = 8'h62 == _T_509[7:0] ? 4'h0 : _GEN_6358; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6360 = 8'h63 == _T_509[7:0] ? 4'h0 : _GEN_6359; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6361 = 8'h64 == _T_509[7:0] ? 4'h0 : _GEN_6360; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6362 = 8'h65 == _T_509[7:0] ? 4'h0 : _GEN_6361; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6363 = 8'h66 == _T_509[7:0] ? 4'h0 : _GEN_6362; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6364 = 8'h67 == _T_509[7:0] ? 4'h0 : _GEN_6363; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6365 = 8'h68 == _T_509[7:0] ? 4'hf : _GEN_6364; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6366 = 8'h69 == _T_509[7:0] ? 4'hf : _GEN_6365; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6367 = 8'h6a == _T_509[7:0] ? 4'hf : _GEN_6366; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6368 = 8'h6b == _T_509[7:0] ? 4'hf : _GEN_6367; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6369 = 8'h6c == _T_509[7:0] ? 4'hf : _GEN_6368; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6370 = 8'h6d == _T_509[7:0] ? 4'hf : _GEN_6369; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6371 = 8'h6e == _T_509[7:0] ? 4'hf : _GEN_6370; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6372 = 8'h6f == _T_509[7:0] ? 4'hf : _GEN_6371; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6373 = 8'h70 == _T_509[7:0] ? 4'h0 : _GEN_6372; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6374 = 8'h71 == _T_509[7:0] ? 4'h0 : _GEN_6373; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6375 = 8'h72 == _T_509[7:0] ? 4'h0 : _GEN_6374; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6376 = 8'h73 == _T_509[7:0] ? 4'h0 : _GEN_6375; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6377 = 8'h74 == _T_509[7:0] ? 4'h0 : _GEN_6376; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6378 = 8'h75 == _T_509[7:0] ? 4'h0 : _GEN_6377; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6379 = 8'h76 == _T_509[7:0] ? 4'h0 : _GEN_6378; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6380 = 8'h77 == _T_509[7:0] ? 4'h0 : _GEN_6379; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6381 = 8'h78 == _T_509[7:0] ? 4'hf : _GEN_6380; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6382 = 8'h79 == _T_509[7:0] ? 4'hf : _GEN_6381; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6383 = 8'h7a == _T_509[7:0] ? 4'hf : _GEN_6382; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6384 = 8'h7b == _T_509[7:0] ? 4'hf : _GEN_6383; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6385 = 8'h7c == _T_509[7:0] ? 4'hf : _GEN_6384; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6386 = 8'h7d == _T_509[7:0] ? 4'hf : _GEN_6385; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6387 = 8'h7e == _T_509[7:0] ? 4'hf : _GEN_6386; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6388 = 8'h7f == _T_509[7:0] ? 4'hf : _GEN_6387; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6389 = 8'h80 == _T_509[7:0] ? 4'h0 : _GEN_6388; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6390 = 8'h81 == _T_509[7:0] ? 4'h0 : _GEN_6389; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6391 = 8'h82 == _T_509[7:0] ? 4'h0 : _GEN_6390; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6392 = 8'h83 == _T_509[7:0] ? 4'h0 : _GEN_6391; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6393 = 8'h84 == _T_509[7:0] ? 4'h0 : _GEN_6392; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6394 = 8'h85 == _T_509[7:0] ? 4'h0 : _GEN_6393; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6395 = 8'h86 == _T_509[7:0] ? 4'h0 : _GEN_6394; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6396 = 8'h87 == _T_509[7:0] ? 4'h0 : _GEN_6395; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6397 = 8'h88 == _T_509[7:0] ? 4'hf : _GEN_6396; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6398 = 8'h89 == _T_509[7:0] ? 4'hf : _GEN_6397; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6399 = 8'h8a == _T_509[7:0] ? 4'hf : _GEN_6398; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6400 = 8'h8b == _T_509[7:0] ? 4'hf : _GEN_6399; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6401 = 8'h8c == _T_509[7:0] ? 4'hf : _GEN_6400; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6402 = 8'h8d == _T_509[7:0] ? 4'hf : _GEN_6401; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6403 = 8'h8e == _T_509[7:0] ? 4'hf : _GEN_6402; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6404 = 8'h8f == _T_509[7:0] ? 4'hf : _GEN_6403; // @[Filter.scala 196:62]
  wire [4:0] _GEN_7646 = {{1'd0}, _GEN_6404}; // @[Filter.scala 196:62]
  wire [8:0] _T_511 = _GEN_7646 * 5'h14; // @[Filter.scala 196:62]
  wire [3:0] _GEN_6469 = 8'h40 == _T_509[7:0] ? 4'hf : 4'h0; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6470 = 8'h41 == _T_509[7:0] ? 4'hf : _GEN_6469; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6471 = 8'h42 == _T_509[7:0] ? 4'hf : _GEN_6470; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6472 = 8'h43 == _T_509[7:0] ? 4'hf : _GEN_6471; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6473 = 8'h44 == _T_509[7:0] ? 4'hf : _GEN_6472; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6474 = 8'h45 == _T_509[7:0] ? 4'hf : _GEN_6473; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6475 = 8'h46 == _T_509[7:0] ? 4'hf : _GEN_6474; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6476 = 8'h47 == _T_509[7:0] ? 4'hf : _GEN_6475; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6477 = 8'h48 == _T_509[7:0] ? 4'hf : _GEN_6476; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6478 = 8'h49 == _T_509[7:0] ? 4'hf : _GEN_6477; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6479 = 8'h4a == _T_509[7:0] ? 4'hf : _GEN_6478; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6480 = 8'h4b == _T_509[7:0] ? 4'hf : _GEN_6479; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6481 = 8'h4c == _T_509[7:0] ? 4'hf : _GEN_6480; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6482 = 8'h4d == _T_509[7:0] ? 4'hf : _GEN_6481; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6483 = 8'h4e == _T_509[7:0] ? 4'hf : _GEN_6482; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6484 = 8'h4f == _T_509[7:0] ? 4'hf : _GEN_6483; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6485 = 8'h50 == _T_509[7:0] ? 4'hf : _GEN_6484; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6486 = 8'h51 == _T_509[7:0] ? 4'hf : _GEN_6485; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6487 = 8'h52 == _T_509[7:0] ? 4'hf : _GEN_6486; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6488 = 8'h53 == _T_509[7:0] ? 4'hf : _GEN_6487; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6489 = 8'h54 == _T_509[7:0] ? 4'hf : _GEN_6488; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6490 = 8'h55 == _T_509[7:0] ? 4'hf : _GEN_6489; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6491 = 8'h56 == _T_509[7:0] ? 4'hf : _GEN_6490; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6492 = 8'h57 == _T_509[7:0] ? 4'hf : _GEN_6491; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6493 = 8'h58 == _T_509[7:0] ? 4'hf : _GEN_6492; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6494 = 8'h59 == _T_509[7:0] ? 4'hf : _GEN_6493; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6495 = 8'h5a == _T_509[7:0] ? 4'hf : _GEN_6494; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6496 = 8'h5b == _T_509[7:0] ? 4'hf : _GEN_6495; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6497 = 8'h5c == _T_509[7:0] ? 4'hf : _GEN_6496; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6498 = 8'h5d == _T_509[7:0] ? 4'hf : _GEN_6497; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6499 = 8'h5e == _T_509[7:0] ? 4'hf : _GEN_6498; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6500 = 8'h5f == _T_509[7:0] ? 4'hf : _GEN_6499; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6501 = 8'h60 == _T_509[7:0] ? 4'hf : _GEN_6500; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6502 = 8'h61 == _T_509[7:0] ? 4'hf : _GEN_6501; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6503 = 8'h62 == _T_509[7:0] ? 4'hf : _GEN_6502; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6504 = 8'h63 == _T_509[7:0] ? 4'hf : _GEN_6503; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6505 = 8'h64 == _T_509[7:0] ? 4'hf : _GEN_6504; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6506 = 8'h65 == _T_509[7:0] ? 4'hf : _GEN_6505; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6507 = 8'h66 == _T_509[7:0] ? 4'hf : _GEN_6506; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6508 = 8'h67 == _T_509[7:0] ? 4'hf : _GEN_6507; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6509 = 8'h68 == _T_509[7:0] ? 4'hf : _GEN_6508; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6510 = 8'h69 == _T_509[7:0] ? 4'hf : _GEN_6509; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6511 = 8'h6a == _T_509[7:0] ? 4'hf : _GEN_6510; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6512 = 8'h6b == _T_509[7:0] ? 4'hf : _GEN_6511; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6513 = 8'h6c == _T_509[7:0] ? 4'hf : _GEN_6512; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6514 = 8'h6d == _T_509[7:0] ? 4'hf : _GEN_6513; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6515 = 8'h6e == _T_509[7:0] ? 4'hf : _GEN_6514; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6516 = 8'h6f == _T_509[7:0] ? 4'hf : _GEN_6515; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6517 = 8'h70 == _T_509[7:0] ? 4'hf : _GEN_6516; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6518 = 8'h71 == _T_509[7:0] ? 4'hf : _GEN_6517; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6519 = 8'h72 == _T_509[7:0] ? 4'hf : _GEN_6518; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6520 = 8'h73 == _T_509[7:0] ? 4'hf : _GEN_6519; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6521 = 8'h74 == _T_509[7:0] ? 4'hf : _GEN_6520; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6522 = 8'h75 == _T_509[7:0] ? 4'hf : _GEN_6521; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6523 = 8'h76 == _T_509[7:0] ? 4'hf : _GEN_6522; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6524 = 8'h77 == _T_509[7:0] ? 4'hf : _GEN_6523; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6525 = 8'h78 == _T_509[7:0] ? 4'hf : _GEN_6524; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6526 = 8'h79 == _T_509[7:0] ? 4'hf : _GEN_6525; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6527 = 8'h7a == _T_509[7:0] ? 4'hf : _GEN_6526; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6528 = 8'h7b == _T_509[7:0] ? 4'hf : _GEN_6527; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6529 = 8'h7c == _T_509[7:0] ? 4'hf : _GEN_6528; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6530 = 8'h7d == _T_509[7:0] ? 4'hf : _GEN_6529; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6531 = 8'h7e == _T_509[7:0] ? 4'hf : _GEN_6530; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6532 = 8'h7f == _T_509[7:0] ? 4'hf : _GEN_6531; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6533 = 8'h80 == _T_509[7:0] ? 4'hf : _GEN_6532; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6534 = 8'h81 == _T_509[7:0] ? 4'hf : _GEN_6533; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6535 = 8'h82 == _T_509[7:0] ? 4'hf : _GEN_6534; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6536 = 8'h83 == _T_509[7:0] ? 4'hf : _GEN_6535; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6537 = 8'h84 == _T_509[7:0] ? 4'hf : _GEN_6536; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6538 = 8'h85 == _T_509[7:0] ? 4'hf : _GEN_6537; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6539 = 8'h86 == _T_509[7:0] ? 4'hf : _GEN_6538; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6540 = 8'h87 == _T_509[7:0] ? 4'hf : _GEN_6539; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6541 = 8'h88 == _T_509[7:0] ? 4'hf : _GEN_6540; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6542 = 8'h89 == _T_509[7:0] ? 4'hf : _GEN_6541; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6543 = 8'h8a == _T_509[7:0] ? 4'hf : _GEN_6542; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6544 = 8'h8b == _T_509[7:0] ? 4'hf : _GEN_6543; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6545 = 8'h8c == _T_509[7:0] ? 4'hf : _GEN_6544; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6546 = 8'h8d == _T_509[7:0] ? 4'hf : _GEN_6545; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6547 = 8'h8e == _T_509[7:0] ? 4'hf : _GEN_6546; // @[Filter.scala 196:102]
  wire [3:0] _GEN_6548 = 8'h8f == _T_509[7:0] ? 4'hf : _GEN_6547; // @[Filter.scala 196:102]
  wire [6:0] _GEN_7648 = {{3'd0}, _GEN_6548}; // @[Filter.scala 196:102]
  wire [10:0] _T_516 = _GEN_7648 * 7'h46; // @[Filter.scala 196:102]
  wire [10:0] _GEN_7649 = {{2'd0}, _T_511}; // @[Filter.scala 196:69]
  wire [10:0] _T_518 = _GEN_7649 + _T_516; // @[Filter.scala 196:69]
  wire [3:0] _GEN_6557 = 8'h8 == _T_509[7:0] ? 4'hf : 4'h0; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6558 = 8'h9 == _T_509[7:0] ? 4'hf : _GEN_6557; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6559 = 8'ha == _T_509[7:0] ? 4'hf : _GEN_6558; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6560 = 8'hb == _T_509[7:0] ? 4'hf : _GEN_6559; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6561 = 8'hc == _T_509[7:0] ? 4'hf : _GEN_6560; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6562 = 8'hd == _T_509[7:0] ? 4'hf : _GEN_6561; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6563 = 8'he == _T_509[7:0] ? 4'hf : _GEN_6562; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6564 = 8'hf == _T_509[7:0] ? 4'hf : _GEN_6563; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6565 = 8'h10 == _T_509[7:0] ? 4'h0 : _GEN_6564; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6566 = 8'h11 == _T_509[7:0] ? 4'h0 : _GEN_6565; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6567 = 8'h12 == _T_509[7:0] ? 4'h0 : _GEN_6566; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6568 = 8'h13 == _T_509[7:0] ? 4'h0 : _GEN_6567; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6569 = 8'h14 == _T_509[7:0] ? 4'h0 : _GEN_6568; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6570 = 8'h15 == _T_509[7:0] ? 4'h0 : _GEN_6569; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6571 = 8'h16 == _T_509[7:0] ? 4'h0 : _GEN_6570; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6572 = 8'h17 == _T_509[7:0] ? 4'h0 : _GEN_6571; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6573 = 8'h18 == _T_509[7:0] ? 4'hf : _GEN_6572; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6574 = 8'h19 == _T_509[7:0] ? 4'hf : _GEN_6573; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6575 = 8'h1a == _T_509[7:0] ? 4'hf : _GEN_6574; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6576 = 8'h1b == _T_509[7:0] ? 4'hf : _GEN_6575; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6577 = 8'h1c == _T_509[7:0] ? 4'hf : _GEN_6576; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6578 = 8'h1d == _T_509[7:0] ? 4'hf : _GEN_6577; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6579 = 8'h1e == _T_509[7:0] ? 4'hf : _GEN_6578; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6580 = 8'h1f == _T_509[7:0] ? 4'hf : _GEN_6579; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6581 = 8'h20 == _T_509[7:0] ? 4'h0 : _GEN_6580; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6582 = 8'h21 == _T_509[7:0] ? 4'h0 : _GEN_6581; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6583 = 8'h22 == _T_509[7:0] ? 4'h0 : _GEN_6582; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6584 = 8'h23 == _T_509[7:0] ? 4'h0 : _GEN_6583; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6585 = 8'h24 == _T_509[7:0] ? 4'h0 : _GEN_6584; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6586 = 8'h25 == _T_509[7:0] ? 4'h0 : _GEN_6585; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6587 = 8'h26 == _T_509[7:0] ? 4'h0 : _GEN_6586; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6588 = 8'h27 == _T_509[7:0] ? 4'h0 : _GEN_6587; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6589 = 8'h28 == _T_509[7:0] ? 4'hf : _GEN_6588; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6590 = 8'h29 == _T_509[7:0] ? 4'hf : _GEN_6589; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6591 = 8'h2a == _T_509[7:0] ? 4'hf : _GEN_6590; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6592 = 8'h2b == _T_509[7:0] ? 4'hf : _GEN_6591; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6593 = 8'h2c == _T_509[7:0] ? 4'hf : _GEN_6592; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6594 = 8'h2d == _T_509[7:0] ? 4'hf : _GEN_6593; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6595 = 8'h2e == _T_509[7:0] ? 4'hf : _GEN_6594; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6596 = 8'h2f == _T_509[7:0] ? 4'hf : _GEN_6595; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6597 = 8'h30 == _T_509[7:0] ? 4'h0 : _GEN_6596; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6598 = 8'h31 == _T_509[7:0] ? 4'h0 : _GEN_6597; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6599 = 8'h32 == _T_509[7:0] ? 4'h0 : _GEN_6598; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6600 = 8'h33 == _T_509[7:0] ? 4'h0 : _GEN_6599; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6601 = 8'h34 == _T_509[7:0] ? 4'h0 : _GEN_6600; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6602 = 8'h35 == _T_509[7:0] ? 4'h0 : _GEN_6601; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6603 = 8'h36 == _T_509[7:0] ? 4'h0 : _GEN_6602; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6604 = 8'h37 == _T_509[7:0] ? 4'h0 : _GEN_6603; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6605 = 8'h38 == _T_509[7:0] ? 4'hf : _GEN_6604; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6606 = 8'h39 == _T_509[7:0] ? 4'hf : _GEN_6605; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6607 = 8'h3a == _T_509[7:0] ? 4'hf : _GEN_6606; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6608 = 8'h3b == _T_509[7:0] ? 4'hf : _GEN_6607; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6609 = 8'h3c == _T_509[7:0] ? 4'hf : _GEN_6608; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6610 = 8'h3d == _T_509[7:0] ? 4'hf : _GEN_6609; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6611 = 8'h3e == _T_509[7:0] ? 4'hf : _GEN_6610; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6612 = 8'h3f == _T_509[7:0] ? 4'hf : _GEN_6611; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6613 = 8'h40 == _T_509[7:0] ? 4'h0 : _GEN_6612; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6614 = 8'h41 == _T_509[7:0] ? 4'h0 : _GEN_6613; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6615 = 8'h42 == _T_509[7:0] ? 4'h0 : _GEN_6614; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6616 = 8'h43 == _T_509[7:0] ? 4'h0 : _GEN_6615; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6617 = 8'h44 == _T_509[7:0] ? 4'h0 : _GEN_6616; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6618 = 8'h45 == _T_509[7:0] ? 4'h0 : _GEN_6617; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6619 = 8'h46 == _T_509[7:0] ? 4'h0 : _GEN_6618; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6620 = 8'h47 == _T_509[7:0] ? 4'h0 : _GEN_6619; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6621 = 8'h48 == _T_509[7:0] ? 4'hf : _GEN_6620; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6622 = 8'h49 == _T_509[7:0] ? 4'hf : _GEN_6621; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6623 = 8'h4a == _T_509[7:0] ? 4'hf : _GEN_6622; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6624 = 8'h4b == _T_509[7:0] ? 4'hf : _GEN_6623; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6625 = 8'h4c == _T_509[7:0] ? 4'hf : _GEN_6624; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6626 = 8'h4d == _T_509[7:0] ? 4'hf : _GEN_6625; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6627 = 8'h4e == _T_509[7:0] ? 4'hf : _GEN_6626; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6628 = 8'h4f == _T_509[7:0] ? 4'hf : _GEN_6627; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6629 = 8'h50 == _T_509[7:0] ? 4'h0 : _GEN_6628; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6630 = 8'h51 == _T_509[7:0] ? 4'h0 : _GEN_6629; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6631 = 8'h52 == _T_509[7:0] ? 4'h0 : _GEN_6630; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6632 = 8'h53 == _T_509[7:0] ? 4'h0 : _GEN_6631; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6633 = 8'h54 == _T_509[7:0] ? 4'h0 : _GEN_6632; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6634 = 8'h55 == _T_509[7:0] ? 4'h0 : _GEN_6633; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6635 = 8'h56 == _T_509[7:0] ? 4'h0 : _GEN_6634; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6636 = 8'h57 == _T_509[7:0] ? 4'h0 : _GEN_6635; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6637 = 8'h58 == _T_509[7:0] ? 4'hf : _GEN_6636; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6638 = 8'h59 == _T_509[7:0] ? 4'hf : _GEN_6637; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6639 = 8'h5a == _T_509[7:0] ? 4'hf : _GEN_6638; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6640 = 8'h5b == _T_509[7:0] ? 4'hf : _GEN_6639; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6641 = 8'h5c == _T_509[7:0] ? 4'hf : _GEN_6640; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6642 = 8'h5d == _T_509[7:0] ? 4'hf : _GEN_6641; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6643 = 8'h5e == _T_509[7:0] ? 4'hf : _GEN_6642; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6644 = 8'h5f == _T_509[7:0] ? 4'hf : _GEN_6643; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6645 = 8'h60 == _T_509[7:0] ? 4'h0 : _GEN_6644; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6646 = 8'h61 == _T_509[7:0] ? 4'h0 : _GEN_6645; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6647 = 8'h62 == _T_509[7:0] ? 4'h0 : _GEN_6646; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6648 = 8'h63 == _T_509[7:0] ? 4'h0 : _GEN_6647; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6649 = 8'h64 == _T_509[7:0] ? 4'h0 : _GEN_6648; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6650 = 8'h65 == _T_509[7:0] ? 4'h0 : _GEN_6649; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6651 = 8'h66 == _T_509[7:0] ? 4'h0 : _GEN_6650; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6652 = 8'h67 == _T_509[7:0] ? 4'h0 : _GEN_6651; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6653 = 8'h68 == _T_509[7:0] ? 4'hf : _GEN_6652; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6654 = 8'h69 == _T_509[7:0] ? 4'hf : _GEN_6653; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6655 = 8'h6a == _T_509[7:0] ? 4'hf : _GEN_6654; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6656 = 8'h6b == _T_509[7:0] ? 4'hf : _GEN_6655; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6657 = 8'h6c == _T_509[7:0] ? 4'hf : _GEN_6656; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6658 = 8'h6d == _T_509[7:0] ? 4'hf : _GEN_6657; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6659 = 8'h6e == _T_509[7:0] ? 4'hf : _GEN_6658; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6660 = 8'h6f == _T_509[7:0] ? 4'hf : _GEN_6659; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6661 = 8'h70 == _T_509[7:0] ? 4'h0 : _GEN_6660; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6662 = 8'h71 == _T_509[7:0] ? 4'h0 : _GEN_6661; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6663 = 8'h72 == _T_509[7:0] ? 4'h0 : _GEN_6662; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6664 = 8'h73 == _T_509[7:0] ? 4'h0 : _GEN_6663; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6665 = 8'h74 == _T_509[7:0] ? 4'h0 : _GEN_6664; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6666 = 8'h75 == _T_509[7:0] ? 4'h0 : _GEN_6665; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6667 = 8'h76 == _T_509[7:0] ? 4'h0 : _GEN_6666; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6668 = 8'h77 == _T_509[7:0] ? 4'h0 : _GEN_6667; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6669 = 8'h78 == _T_509[7:0] ? 4'hf : _GEN_6668; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6670 = 8'h79 == _T_509[7:0] ? 4'hf : _GEN_6669; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6671 = 8'h7a == _T_509[7:0] ? 4'hf : _GEN_6670; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6672 = 8'h7b == _T_509[7:0] ? 4'hf : _GEN_6671; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6673 = 8'h7c == _T_509[7:0] ? 4'hf : _GEN_6672; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6674 = 8'h7d == _T_509[7:0] ? 4'hf : _GEN_6673; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6675 = 8'h7e == _T_509[7:0] ? 4'hf : _GEN_6674; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6676 = 8'h7f == _T_509[7:0] ? 4'hf : _GEN_6675; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6677 = 8'h80 == _T_509[7:0] ? 4'h0 : _GEN_6676; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6678 = 8'h81 == _T_509[7:0] ? 4'h0 : _GEN_6677; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6679 = 8'h82 == _T_509[7:0] ? 4'h0 : _GEN_6678; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6680 = 8'h83 == _T_509[7:0] ? 4'h0 : _GEN_6679; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6681 = 8'h84 == _T_509[7:0] ? 4'h0 : _GEN_6680; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6682 = 8'h85 == _T_509[7:0] ? 4'h0 : _GEN_6681; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6683 = 8'h86 == _T_509[7:0] ? 4'h0 : _GEN_6682; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6684 = 8'h87 == _T_509[7:0] ? 4'h0 : _GEN_6683; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6685 = 8'h88 == _T_509[7:0] ? 4'hf : _GEN_6684; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6686 = 8'h89 == _T_509[7:0] ? 4'hf : _GEN_6685; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6687 = 8'h8a == _T_509[7:0] ? 4'hf : _GEN_6686; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6688 = 8'h8b == _T_509[7:0] ? 4'hf : _GEN_6687; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6689 = 8'h8c == _T_509[7:0] ? 4'hf : _GEN_6688; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6690 = 8'h8d == _T_509[7:0] ? 4'hf : _GEN_6689; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6691 = 8'h8e == _T_509[7:0] ? 4'hf : _GEN_6690; // @[Filter.scala 196:142]
  wire [3:0] _GEN_6692 = 8'h8f == _T_509[7:0] ? 4'hf : _GEN_6691; // @[Filter.scala 196:142]
  wire [7:0] _T_523 = _GEN_6692 * 4'ha; // @[Filter.scala 196:142]
  wire [10:0] _GEN_7651 = {{3'd0}, _T_523}; // @[Filter.scala 196:109]
  wire [10:0] _T_525 = _T_518 + _GEN_7651; // @[Filter.scala 196:109]
  wire [10:0] _T_526 = _T_525 / 11'h64; // @[Filter.scala 196:150]
  wire  _T_528 = _T_499 >= 5'h10; // @[Filter.scala 199:31]
  wire  _T_532 = _T_506 >= 32'h9; // @[Filter.scala 199:63]
  wire  _T_533 = _T_528 | _T_532; // @[Filter.scala 199:58]
  wire [10:0] _GEN_6837 = io_SPI_distort ? _T_526 : {{7'd0}, _GEN_6404}; // @[Filter.scala 201:35]
  wire [10:0] _GEN_6838 = _T_533 ? 11'h0 : _GEN_6837; // @[Filter.scala 199:80]
  wire [10:0] _GEN_6983 = io_SPI_distort ? _T_526 : {{7'd0}, _GEN_6548}; // @[Filter.scala 201:35]
  wire [10:0] _GEN_6984 = _T_533 ? 11'h0 : _GEN_6983; // @[Filter.scala 199:80]
  wire [10:0] _GEN_7129 = io_SPI_distort ? _T_526 : {{7'd0}, _GEN_6692}; // @[Filter.scala 201:35]
  wire [10:0] _GEN_7130 = _T_533 ? 11'h0 : _GEN_7129; // @[Filter.scala 199:80]
  reg [8:0] pixOut_0_0; // @[Filter.scala 210:32]
  reg [8:0] pixOut_0_1; // @[Filter.scala 210:32]
  reg [8:0] pixOut_0_2; // @[Filter.scala 210:32]
  reg [8:0] pixOut_0_3; // @[Filter.scala 210:32]
  reg [8:0] pixOut_0_4; // @[Filter.scala 210:32]
  reg [8:0] pixOut_0_5; // @[Filter.scala 210:32]
  reg [8:0] pixOut_0_6; // @[Filter.scala 210:32]
  reg [8:0] pixOut_0_7; // @[Filter.scala 210:32]
  reg [8:0] pixOut_1_0; // @[Filter.scala 210:87]
  reg [8:0] pixOut_1_1; // @[Filter.scala 210:87]
  reg [8:0] pixOut_1_2; // @[Filter.scala 210:87]
  reg [8:0] pixOut_1_3; // @[Filter.scala 210:87]
  reg [8:0] pixOut_1_4; // @[Filter.scala 210:87]
  reg [8:0] pixOut_1_5; // @[Filter.scala 210:87]
  reg [8:0] pixOut_1_6; // @[Filter.scala 210:87]
  reg [8:0] pixOut_1_7; // @[Filter.scala 210:87]
  reg [8:0] pixOut_2_0; // @[Filter.scala 210:142]
  reg [8:0] pixOut_2_1; // @[Filter.scala 210:142]
  reg [8:0] pixOut_2_2; // @[Filter.scala 210:142]
  reg [8:0] pixOut_2_3; // @[Filter.scala 210:142]
  reg [8:0] pixOut_2_4; // @[Filter.scala 210:142]
  reg [8:0] pixOut_2_5; // @[Filter.scala 210:142]
  reg [8:0] pixOut_2_6; // @[Filter.scala 210:142]
  reg [8:0] pixOut_2_7; // @[Filter.scala 210:142]
  reg  validOut; // @[Filter.scala 211:29]
  wire [7:0] _GEN_7132 = 3'h1 == io_SPI_filterIndex[2:0] ? $signed(8'sh9) : $signed(8'sh1); // @[Filter.scala 215:64]
  wire [7:0] _GEN_7133 = 3'h2 == io_SPI_filterIndex[2:0] ? $signed(8'sh10) : $signed(_GEN_7132); // @[Filter.scala 215:64]
  wire [7:0] _GEN_7134 = 3'h3 == io_SPI_filterIndex[2:0] ? $signed(8'sh1) : $signed(_GEN_7133); // @[Filter.scala 215:64]
  wire [7:0] _GEN_7135 = 3'h4 == io_SPI_filterIndex[2:0] ? $signed(8'sh1) : $signed(_GEN_7134); // @[Filter.scala 215:64]
  wire [7:0] _GEN_7136 = 3'h5 == io_SPI_filterIndex[2:0] ? $signed(8'sh1) : $signed(_GEN_7135); // @[Filter.scala 215:64]
  wire [8:0] _GEN_7655 = {{1{_GEN_7136[7]}},_GEN_7136}; // @[Filter.scala 215:64]
  wire [9:0] _T_564 = $signed(KernelConvolution_io_pixelVal_out_0) / $signed(_GEN_7655); // @[Filter.scala 215:64]
  wire  _T_565 = $signed(pixOut_0_0) < 9'sh0; // @[Filter.scala 217:30]
  wire  _T_568 = $signed(pixOut_0_0) > 9'shf; // @[Filter.scala 222:36]
  wire [8:0] _GEN_7138 = _T_568 ? 9'hf : pixOut_0_0; // @[Filter.scala 224:44]
  wire [8:0] _GEN_7140 = _T_565 ? 9'h0 : _GEN_7138; // @[Filter.scala 219:43]
  wire [9:0] _T_575 = $signed(KernelConvolution_io_pixelVal_out_1) / $signed(_GEN_7655); // @[Filter.scala 215:64]
  wire  _T_576 = $signed(pixOut_0_1) < 9'sh0; // @[Filter.scala 217:30]
  wire  _T_579 = $signed(pixOut_0_1) > 9'shf; // @[Filter.scala 222:36]
  wire [8:0] _GEN_7143 = _T_579 ? 9'hf : pixOut_0_1; // @[Filter.scala 224:44]
  wire [8:0] _GEN_7145 = _T_576 ? 9'h0 : _GEN_7143; // @[Filter.scala 219:43]
  wire [9:0] _T_586 = $signed(KernelConvolution_io_pixelVal_out_2) / $signed(_GEN_7655); // @[Filter.scala 215:64]
  wire  _T_587 = $signed(pixOut_0_2) < 9'sh0; // @[Filter.scala 217:30]
  wire  _T_590 = $signed(pixOut_0_2) > 9'shf; // @[Filter.scala 222:36]
  wire [8:0] _GEN_7148 = _T_590 ? 9'hf : pixOut_0_2; // @[Filter.scala 224:44]
  wire [8:0] _GEN_7150 = _T_587 ? 9'h0 : _GEN_7148; // @[Filter.scala 219:43]
  wire [9:0] _T_597 = $signed(KernelConvolution_io_pixelVal_out_3) / $signed(_GEN_7655); // @[Filter.scala 215:64]
  wire  _T_598 = $signed(pixOut_0_3) < 9'sh0; // @[Filter.scala 217:30]
  wire  _T_601 = $signed(pixOut_0_3) > 9'shf; // @[Filter.scala 222:36]
  wire [8:0] _GEN_7153 = _T_601 ? 9'hf : pixOut_0_3; // @[Filter.scala 224:44]
  wire [8:0] _GEN_7155 = _T_598 ? 9'h0 : _GEN_7153; // @[Filter.scala 219:43]
  wire [9:0] _T_608 = $signed(KernelConvolution_io_pixelVal_out_4) / $signed(_GEN_7655); // @[Filter.scala 215:64]
  wire  _T_609 = $signed(pixOut_0_4) < 9'sh0; // @[Filter.scala 217:30]
  wire  _T_612 = $signed(pixOut_0_4) > 9'shf; // @[Filter.scala 222:36]
  wire [8:0] _GEN_7158 = _T_612 ? 9'hf : pixOut_0_4; // @[Filter.scala 224:44]
  wire [8:0] _GEN_7160 = _T_609 ? 9'h0 : _GEN_7158; // @[Filter.scala 219:43]
  wire [9:0] _T_619 = $signed(KernelConvolution_io_pixelVal_out_5) / $signed(_GEN_7655); // @[Filter.scala 215:64]
  wire  _T_620 = $signed(pixOut_0_5) < 9'sh0; // @[Filter.scala 217:30]
  wire  _T_623 = $signed(pixOut_0_5) > 9'shf; // @[Filter.scala 222:36]
  wire [8:0] _GEN_7163 = _T_623 ? 9'hf : pixOut_0_5; // @[Filter.scala 224:44]
  wire [8:0] _GEN_7165 = _T_620 ? 9'h0 : _GEN_7163; // @[Filter.scala 219:43]
  wire [9:0] _T_630 = $signed(KernelConvolution_io_pixelVal_out_6) / $signed(_GEN_7655); // @[Filter.scala 215:64]
  wire  _T_631 = $signed(pixOut_0_6) < 9'sh0; // @[Filter.scala 217:30]
  wire  _T_634 = $signed(pixOut_0_6) > 9'shf; // @[Filter.scala 222:36]
  wire [8:0] _GEN_7168 = _T_634 ? 9'hf : pixOut_0_6; // @[Filter.scala 224:44]
  wire [8:0] _GEN_7170 = _T_631 ? 9'h0 : _GEN_7168; // @[Filter.scala 219:43]
  wire [9:0] _T_641 = $signed(KernelConvolution_io_pixelVal_out_7) / $signed(_GEN_7655); // @[Filter.scala 215:64]
  wire  _T_642 = $signed(pixOut_0_7) < 9'sh0; // @[Filter.scala 217:30]
  wire  _T_645 = $signed(pixOut_0_7) > 9'shf; // @[Filter.scala 222:36]
  wire [8:0] _GEN_7173 = _T_645 ? 9'hf : pixOut_0_7; // @[Filter.scala 224:44]
  wire [8:0] _GEN_7175 = _T_642 ? 9'h0 : _GEN_7173; // @[Filter.scala 219:43]
  wire [9:0] _T_652 = $signed(KernelConvolution_1_io_pixelVal_out_0) / $signed(_GEN_7655); // @[Filter.scala 215:64]
  wire  _T_653 = $signed(pixOut_1_0) < 9'sh0; // @[Filter.scala 217:30]
  wire  _T_656 = $signed(pixOut_1_0) > 9'shf; // @[Filter.scala 222:36]
  wire [8:0] _GEN_7178 = _T_656 ? 9'hf : pixOut_1_0; // @[Filter.scala 224:44]
  wire [8:0] _GEN_7180 = _T_653 ? 9'h0 : _GEN_7178; // @[Filter.scala 219:43]
  wire [9:0] _T_663 = $signed(KernelConvolution_1_io_pixelVal_out_1) / $signed(_GEN_7655); // @[Filter.scala 215:64]
  wire  _T_664 = $signed(pixOut_1_1) < 9'sh0; // @[Filter.scala 217:30]
  wire  _T_667 = $signed(pixOut_1_1) > 9'shf; // @[Filter.scala 222:36]
  wire [8:0] _GEN_7183 = _T_667 ? 9'hf : pixOut_1_1; // @[Filter.scala 224:44]
  wire [8:0] _GEN_7185 = _T_664 ? 9'h0 : _GEN_7183; // @[Filter.scala 219:43]
  wire [9:0] _T_674 = $signed(KernelConvolution_1_io_pixelVal_out_2) / $signed(_GEN_7655); // @[Filter.scala 215:64]
  wire  _T_675 = $signed(pixOut_1_2) < 9'sh0; // @[Filter.scala 217:30]
  wire  _T_678 = $signed(pixOut_1_2) > 9'shf; // @[Filter.scala 222:36]
  wire [8:0] _GEN_7188 = _T_678 ? 9'hf : pixOut_1_2; // @[Filter.scala 224:44]
  wire [8:0] _GEN_7190 = _T_675 ? 9'h0 : _GEN_7188; // @[Filter.scala 219:43]
  wire [9:0] _T_685 = $signed(KernelConvolution_1_io_pixelVal_out_3) / $signed(_GEN_7655); // @[Filter.scala 215:64]
  wire  _T_686 = $signed(pixOut_1_3) < 9'sh0; // @[Filter.scala 217:30]
  wire  _T_689 = $signed(pixOut_1_3) > 9'shf; // @[Filter.scala 222:36]
  wire [8:0] _GEN_7193 = _T_689 ? 9'hf : pixOut_1_3; // @[Filter.scala 224:44]
  wire [8:0] _GEN_7195 = _T_686 ? 9'h0 : _GEN_7193; // @[Filter.scala 219:43]
  wire [9:0] _T_696 = $signed(KernelConvolution_1_io_pixelVal_out_4) / $signed(_GEN_7655); // @[Filter.scala 215:64]
  wire  _T_697 = $signed(pixOut_1_4) < 9'sh0; // @[Filter.scala 217:30]
  wire  _T_700 = $signed(pixOut_1_4) > 9'shf; // @[Filter.scala 222:36]
  wire [8:0] _GEN_7198 = _T_700 ? 9'hf : pixOut_1_4; // @[Filter.scala 224:44]
  wire [8:0] _GEN_7200 = _T_697 ? 9'h0 : _GEN_7198; // @[Filter.scala 219:43]
  wire [9:0] _T_707 = $signed(KernelConvolution_1_io_pixelVal_out_5) / $signed(_GEN_7655); // @[Filter.scala 215:64]
  wire  _T_708 = $signed(pixOut_1_5) < 9'sh0; // @[Filter.scala 217:30]
  wire  _T_711 = $signed(pixOut_1_5) > 9'shf; // @[Filter.scala 222:36]
  wire [8:0] _GEN_7203 = _T_711 ? 9'hf : pixOut_1_5; // @[Filter.scala 224:44]
  wire [8:0] _GEN_7205 = _T_708 ? 9'h0 : _GEN_7203; // @[Filter.scala 219:43]
  wire [9:0] _T_718 = $signed(KernelConvolution_1_io_pixelVal_out_6) / $signed(_GEN_7655); // @[Filter.scala 215:64]
  wire  _T_719 = $signed(pixOut_1_6) < 9'sh0; // @[Filter.scala 217:30]
  wire  _T_722 = $signed(pixOut_1_6) > 9'shf; // @[Filter.scala 222:36]
  wire [8:0] _GEN_7208 = _T_722 ? 9'hf : pixOut_1_6; // @[Filter.scala 224:44]
  wire [8:0] _GEN_7210 = _T_719 ? 9'h0 : _GEN_7208; // @[Filter.scala 219:43]
  wire [9:0] _T_729 = $signed(KernelConvolution_1_io_pixelVal_out_7) / $signed(_GEN_7655); // @[Filter.scala 215:64]
  wire  _T_730 = $signed(pixOut_1_7) < 9'sh0; // @[Filter.scala 217:30]
  wire  _T_733 = $signed(pixOut_1_7) > 9'shf; // @[Filter.scala 222:36]
  wire [8:0] _GEN_7213 = _T_733 ? 9'hf : pixOut_1_7; // @[Filter.scala 224:44]
  wire [8:0] _GEN_7215 = _T_730 ? 9'h0 : _GEN_7213; // @[Filter.scala 219:43]
  wire [9:0] _T_740 = $signed(KernelConvolution_2_io_pixelVal_out_0) / $signed(_GEN_7655); // @[Filter.scala 215:64]
  wire  _T_741 = $signed(pixOut_2_0) < 9'sh0; // @[Filter.scala 217:30]
  wire  _T_744 = $signed(pixOut_2_0) > 9'shf; // @[Filter.scala 222:36]
  wire [8:0] _GEN_7218 = _T_744 ? 9'hf : pixOut_2_0; // @[Filter.scala 224:44]
  wire [8:0] _GEN_7220 = _T_741 ? 9'h0 : _GEN_7218; // @[Filter.scala 219:43]
  wire [9:0] _T_751 = $signed(KernelConvolution_2_io_pixelVal_out_1) / $signed(_GEN_7655); // @[Filter.scala 215:64]
  wire  _T_752 = $signed(pixOut_2_1) < 9'sh0; // @[Filter.scala 217:30]
  wire  _T_755 = $signed(pixOut_2_1) > 9'shf; // @[Filter.scala 222:36]
  wire [8:0] _GEN_7223 = _T_755 ? 9'hf : pixOut_2_1; // @[Filter.scala 224:44]
  wire [8:0] _GEN_7225 = _T_752 ? 9'h0 : _GEN_7223; // @[Filter.scala 219:43]
  wire [9:0] _T_762 = $signed(KernelConvolution_2_io_pixelVal_out_2) / $signed(_GEN_7655); // @[Filter.scala 215:64]
  wire  _T_763 = $signed(pixOut_2_2) < 9'sh0; // @[Filter.scala 217:30]
  wire  _T_766 = $signed(pixOut_2_2) > 9'shf; // @[Filter.scala 222:36]
  wire [8:0] _GEN_7228 = _T_766 ? 9'hf : pixOut_2_2; // @[Filter.scala 224:44]
  wire [8:0] _GEN_7230 = _T_763 ? 9'h0 : _GEN_7228; // @[Filter.scala 219:43]
  wire [9:0] _T_773 = $signed(KernelConvolution_2_io_pixelVal_out_3) / $signed(_GEN_7655); // @[Filter.scala 215:64]
  wire  _T_774 = $signed(pixOut_2_3) < 9'sh0; // @[Filter.scala 217:30]
  wire  _T_777 = $signed(pixOut_2_3) > 9'shf; // @[Filter.scala 222:36]
  wire [8:0] _GEN_7233 = _T_777 ? 9'hf : pixOut_2_3; // @[Filter.scala 224:44]
  wire [8:0] _GEN_7235 = _T_774 ? 9'h0 : _GEN_7233; // @[Filter.scala 219:43]
  wire [9:0] _T_784 = $signed(KernelConvolution_2_io_pixelVal_out_4) / $signed(_GEN_7655); // @[Filter.scala 215:64]
  wire  _T_785 = $signed(pixOut_2_4) < 9'sh0; // @[Filter.scala 217:30]
  wire  _T_788 = $signed(pixOut_2_4) > 9'shf; // @[Filter.scala 222:36]
  wire [8:0] _GEN_7238 = _T_788 ? 9'hf : pixOut_2_4; // @[Filter.scala 224:44]
  wire [8:0] _GEN_7240 = _T_785 ? 9'h0 : _GEN_7238; // @[Filter.scala 219:43]
  wire [9:0] _T_795 = $signed(KernelConvolution_2_io_pixelVal_out_5) / $signed(_GEN_7655); // @[Filter.scala 215:64]
  wire  _T_796 = $signed(pixOut_2_5) < 9'sh0; // @[Filter.scala 217:30]
  wire  _T_799 = $signed(pixOut_2_5) > 9'shf; // @[Filter.scala 222:36]
  wire [8:0] _GEN_7243 = _T_799 ? 9'hf : pixOut_2_5; // @[Filter.scala 224:44]
  wire [8:0] _GEN_7245 = _T_796 ? 9'h0 : _GEN_7243; // @[Filter.scala 219:43]
  wire [9:0] _T_806 = $signed(KernelConvolution_2_io_pixelVal_out_6) / $signed(_GEN_7655); // @[Filter.scala 215:64]
  wire  _T_807 = $signed(pixOut_2_6) < 9'sh0; // @[Filter.scala 217:30]
  wire  _T_810 = $signed(pixOut_2_6) > 9'shf; // @[Filter.scala 222:36]
  wire [8:0] _GEN_7248 = _T_810 ? 9'hf : pixOut_2_6; // @[Filter.scala 224:44]
  wire [8:0] _GEN_7250 = _T_807 ? 9'h0 : _GEN_7248; // @[Filter.scala 219:43]
  wire [9:0] _T_817 = $signed(KernelConvolution_2_io_pixelVal_out_7) / $signed(_GEN_7655); // @[Filter.scala 215:64]
  wire  _T_818 = $signed(pixOut_2_7) < 9'sh0; // @[Filter.scala 217:30]
  wire  _T_821 = $signed(pixOut_2_7) > 9'shf; // @[Filter.scala 222:36]
  wire [8:0] _GEN_7253 = _T_821 ? 9'hf : pixOut_2_7; // @[Filter.scala 224:44]
  wire [8:0] _GEN_7255 = _T_818 ? 9'h0 : _GEN_7253; // @[Filter.scala 219:43]
  wire [31:0] _T_829 = pixelIndex + 32'h8; // @[Filter.scala 239:34]
  wire [8:0] _T_830 = 5'h10 * 5'h9; // @[Filter.scala 240:42]
  wire [31:0] _GEN_7679 = {{23'd0}, _T_830}; // @[Filter.scala 240:25]
  wire  _T_831 = pixelIndex == _GEN_7679; // @[Filter.scala 240:25]
  KernelConvolution KernelConvolution ( // @[Filter.scala 178:36]
    .clock(KernelConvolution_clock),
    .reset(KernelConvolution_reset),
    .io_kernelVal_in(KernelConvolution_io_kernelVal_in),
    .io_pixelVal_in_0(KernelConvolution_io_pixelVal_in_0),
    .io_pixelVal_in_1(KernelConvolution_io_pixelVal_in_1),
    .io_pixelVal_in_2(KernelConvolution_io_pixelVal_in_2),
    .io_pixelVal_in_3(KernelConvolution_io_pixelVal_in_3),
    .io_pixelVal_in_4(KernelConvolution_io_pixelVal_in_4),
    .io_pixelVal_in_5(KernelConvolution_io_pixelVal_in_5),
    .io_pixelVal_in_6(KernelConvolution_io_pixelVal_in_6),
    .io_pixelVal_in_7(KernelConvolution_io_pixelVal_in_7),
    .io_pixelVal_out_0(KernelConvolution_io_pixelVal_out_0),
    .io_pixelVal_out_1(KernelConvolution_io_pixelVal_out_1),
    .io_pixelVal_out_2(KernelConvolution_io_pixelVal_out_2),
    .io_pixelVal_out_3(KernelConvolution_io_pixelVal_out_3),
    .io_pixelVal_out_4(KernelConvolution_io_pixelVal_out_4),
    .io_pixelVal_out_5(KernelConvolution_io_pixelVal_out_5),
    .io_pixelVal_out_6(KernelConvolution_io_pixelVal_out_6),
    .io_pixelVal_out_7(KernelConvolution_io_pixelVal_out_7),
    .io_valid_out(KernelConvolution_io_valid_out)
  );
  KernelConvolution KernelConvolution_1 ( // @[Filter.scala 179:36]
    .clock(KernelConvolution_1_clock),
    .reset(KernelConvolution_1_reset),
    .io_kernelVal_in(KernelConvolution_1_io_kernelVal_in),
    .io_pixelVal_in_0(KernelConvolution_1_io_pixelVal_in_0),
    .io_pixelVal_in_1(KernelConvolution_1_io_pixelVal_in_1),
    .io_pixelVal_in_2(KernelConvolution_1_io_pixelVal_in_2),
    .io_pixelVal_in_3(KernelConvolution_1_io_pixelVal_in_3),
    .io_pixelVal_in_4(KernelConvolution_1_io_pixelVal_in_4),
    .io_pixelVal_in_5(KernelConvolution_1_io_pixelVal_in_5),
    .io_pixelVal_in_6(KernelConvolution_1_io_pixelVal_in_6),
    .io_pixelVal_in_7(KernelConvolution_1_io_pixelVal_in_7),
    .io_pixelVal_out_0(KernelConvolution_1_io_pixelVal_out_0),
    .io_pixelVal_out_1(KernelConvolution_1_io_pixelVal_out_1),
    .io_pixelVal_out_2(KernelConvolution_1_io_pixelVal_out_2),
    .io_pixelVal_out_3(KernelConvolution_1_io_pixelVal_out_3),
    .io_pixelVal_out_4(KernelConvolution_1_io_pixelVal_out_4),
    .io_pixelVal_out_5(KernelConvolution_1_io_pixelVal_out_5),
    .io_pixelVal_out_6(KernelConvolution_1_io_pixelVal_out_6),
    .io_pixelVal_out_7(KernelConvolution_1_io_pixelVal_out_7),
    .io_valid_out(KernelConvolution_1_io_valid_out)
  );
  KernelConvolution KernelConvolution_2 ( // @[Filter.scala 180:36]
    .clock(KernelConvolution_2_clock),
    .reset(KernelConvolution_2_reset),
    .io_kernelVal_in(KernelConvolution_2_io_kernelVal_in),
    .io_pixelVal_in_0(KernelConvolution_2_io_pixelVal_in_0),
    .io_pixelVal_in_1(KernelConvolution_2_io_pixelVal_in_1),
    .io_pixelVal_in_2(KernelConvolution_2_io_pixelVal_in_2),
    .io_pixelVal_in_3(KernelConvolution_2_io_pixelVal_in_3),
    .io_pixelVal_in_4(KernelConvolution_2_io_pixelVal_in_4),
    .io_pixelVal_in_5(KernelConvolution_2_io_pixelVal_in_5),
    .io_pixelVal_in_6(KernelConvolution_2_io_pixelVal_in_6),
    .io_pixelVal_in_7(KernelConvolution_2_io_pixelVal_in_7),
    .io_pixelVal_out_0(KernelConvolution_2_io_pixelVal_out_0),
    .io_pixelVal_out_1(KernelConvolution_2_io_pixelVal_out_1),
    .io_pixelVal_out_2(KernelConvolution_2_io_pixelVal_out_2),
    .io_pixelVal_out_3(KernelConvolution_2_io_pixelVal_out_3),
    .io_pixelVal_out_4(KernelConvolution_2_io_pixelVal_out_4),
    .io_pixelVal_out_5(KernelConvolution_2_io_pixelVal_out_5),
    .io_pixelVal_out_6(KernelConvolution_2_io_pixelVal_out_6),
    .io_pixelVal_out_7(KernelConvolution_2_io_pixelVal_out_7),
    .io_valid_out(KernelConvolution_2_io_valid_out)
  );
  assign io_pixelVal_out_0_0 = _GEN_7140[3:0]; // @[Filter.scala 218:35 Filter.scala 220:37 Filter.scala 223:35 Filter.scala 225:35 Filter.scala 227:35 Filter.scala 229:35]
  assign io_pixelVal_out_0_1 = _GEN_7145[3:0]; // @[Filter.scala 218:35 Filter.scala 220:37 Filter.scala 223:35 Filter.scala 225:35 Filter.scala 227:35 Filter.scala 229:35]
  assign io_pixelVal_out_0_2 = _GEN_7150[3:0]; // @[Filter.scala 218:35 Filter.scala 220:37 Filter.scala 223:35 Filter.scala 225:35 Filter.scala 227:35 Filter.scala 229:35]
  assign io_pixelVal_out_0_3 = _GEN_7155[3:0]; // @[Filter.scala 218:35 Filter.scala 220:37 Filter.scala 223:35 Filter.scala 225:35 Filter.scala 227:35 Filter.scala 229:35]
  assign io_pixelVal_out_0_4 = _GEN_7160[3:0]; // @[Filter.scala 218:35 Filter.scala 220:37 Filter.scala 223:35 Filter.scala 225:35 Filter.scala 227:35 Filter.scala 229:35]
  assign io_pixelVal_out_0_5 = _GEN_7165[3:0]; // @[Filter.scala 218:35 Filter.scala 220:37 Filter.scala 223:35 Filter.scala 225:35 Filter.scala 227:35 Filter.scala 229:35]
  assign io_pixelVal_out_0_6 = _GEN_7170[3:0]; // @[Filter.scala 218:35 Filter.scala 220:37 Filter.scala 223:35 Filter.scala 225:35 Filter.scala 227:35 Filter.scala 229:35]
  assign io_pixelVal_out_0_7 = _GEN_7175[3:0]; // @[Filter.scala 218:35 Filter.scala 220:37 Filter.scala 223:35 Filter.scala 225:35 Filter.scala 227:35 Filter.scala 229:35]
  assign io_pixelVal_out_1_0 = _GEN_7180[3:0]; // @[Filter.scala 218:35 Filter.scala 220:37 Filter.scala 223:35 Filter.scala 225:35 Filter.scala 227:35 Filter.scala 229:35]
  assign io_pixelVal_out_1_1 = _GEN_7185[3:0]; // @[Filter.scala 218:35 Filter.scala 220:37 Filter.scala 223:35 Filter.scala 225:35 Filter.scala 227:35 Filter.scala 229:35]
  assign io_pixelVal_out_1_2 = _GEN_7190[3:0]; // @[Filter.scala 218:35 Filter.scala 220:37 Filter.scala 223:35 Filter.scala 225:35 Filter.scala 227:35 Filter.scala 229:35]
  assign io_pixelVal_out_1_3 = _GEN_7195[3:0]; // @[Filter.scala 218:35 Filter.scala 220:37 Filter.scala 223:35 Filter.scala 225:35 Filter.scala 227:35 Filter.scala 229:35]
  assign io_pixelVal_out_1_4 = _GEN_7200[3:0]; // @[Filter.scala 218:35 Filter.scala 220:37 Filter.scala 223:35 Filter.scala 225:35 Filter.scala 227:35 Filter.scala 229:35]
  assign io_pixelVal_out_1_5 = _GEN_7205[3:0]; // @[Filter.scala 218:35 Filter.scala 220:37 Filter.scala 223:35 Filter.scala 225:35 Filter.scala 227:35 Filter.scala 229:35]
  assign io_pixelVal_out_1_6 = _GEN_7210[3:0]; // @[Filter.scala 218:35 Filter.scala 220:37 Filter.scala 223:35 Filter.scala 225:35 Filter.scala 227:35 Filter.scala 229:35]
  assign io_pixelVal_out_1_7 = _GEN_7215[3:0]; // @[Filter.scala 218:35 Filter.scala 220:37 Filter.scala 223:35 Filter.scala 225:35 Filter.scala 227:35 Filter.scala 229:35]
  assign io_pixelVal_out_2_0 = _GEN_7220[3:0]; // @[Filter.scala 218:35 Filter.scala 220:37 Filter.scala 223:35 Filter.scala 225:35 Filter.scala 227:35 Filter.scala 229:35]
  assign io_pixelVal_out_2_1 = _GEN_7225[3:0]; // @[Filter.scala 218:35 Filter.scala 220:37 Filter.scala 223:35 Filter.scala 225:35 Filter.scala 227:35 Filter.scala 229:35]
  assign io_pixelVal_out_2_2 = _GEN_7230[3:0]; // @[Filter.scala 218:35 Filter.scala 220:37 Filter.scala 223:35 Filter.scala 225:35 Filter.scala 227:35 Filter.scala 229:35]
  assign io_pixelVal_out_2_3 = _GEN_7235[3:0]; // @[Filter.scala 218:35 Filter.scala 220:37 Filter.scala 223:35 Filter.scala 225:35 Filter.scala 227:35 Filter.scala 229:35]
  assign io_pixelVal_out_2_4 = _GEN_7240[3:0]; // @[Filter.scala 218:35 Filter.scala 220:37 Filter.scala 223:35 Filter.scala 225:35 Filter.scala 227:35 Filter.scala 229:35]
  assign io_pixelVal_out_2_5 = _GEN_7245[3:0]; // @[Filter.scala 218:35 Filter.scala 220:37 Filter.scala 223:35 Filter.scala 225:35 Filter.scala 227:35 Filter.scala 229:35]
  assign io_pixelVal_out_2_6 = _GEN_7250[3:0]; // @[Filter.scala 218:35 Filter.scala 220:37 Filter.scala 223:35 Filter.scala 225:35 Filter.scala 227:35 Filter.scala 229:35]
  assign io_pixelVal_out_2_7 = _GEN_7255[3:0]; // @[Filter.scala 218:35 Filter.scala 220:37 Filter.scala 223:35 Filter.scala 225:35 Filter.scala 227:35 Filter.scala 229:35]
  assign io_valid_out = validOut; // @[Filter.scala 236:18]
  assign KernelConvolution_clock = clock;
  assign KernelConvolution_reset = reset;
  assign KernelConvolution_io_kernelVal_in = _GEN_7341 & _GEN_7268 ? $signed(5'sh0) : $signed(_GEN_55); // @[Filter.scala 186:41]
  assign KernelConvolution_io_pixelVal_in_0 = _GEN_748[3:0]; // @[Filter.scala 200:53 Filter.scala 202:51 Filter.scala 204:51]
  assign KernelConvolution_io_pixelVal_in_1 = _GEN_1618[3:0]; // @[Filter.scala 200:53 Filter.scala 202:51 Filter.scala 204:51]
  assign KernelConvolution_io_pixelVal_in_2 = _GEN_2488[3:0]; // @[Filter.scala 200:53 Filter.scala 202:51 Filter.scala 204:51]
  assign KernelConvolution_io_pixelVal_in_3 = _GEN_3358[3:0]; // @[Filter.scala 200:53 Filter.scala 202:51 Filter.scala 204:51]
  assign KernelConvolution_io_pixelVal_in_4 = _GEN_4228[3:0]; // @[Filter.scala 200:53 Filter.scala 202:51 Filter.scala 204:51]
  assign KernelConvolution_io_pixelVal_in_5 = _GEN_5098[3:0]; // @[Filter.scala 200:53 Filter.scala 202:51 Filter.scala 204:51]
  assign KernelConvolution_io_pixelVal_in_6 = _GEN_5968[3:0]; // @[Filter.scala 200:53 Filter.scala 202:51 Filter.scala 204:51]
  assign KernelConvolution_io_pixelVal_in_7 = _GEN_6838[3:0]; // @[Filter.scala 200:53 Filter.scala 202:51 Filter.scala 204:51]
  assign KernelConvolution_1_clock = clock;
  assign KernelConvolution_1_reset = reset;
  assign KernelConvolution_1_io_kernelVal_in = _GEN_7341 & _GEN_7268 ? $signed(5'sh0) : $signed(_GEN_55); // @[Filter.scala 186:41]
  assign KernelConvolution_1_io_pixelVal_in_0 = _GEN_894[3:0]; // @[Filter.scala 200:53 Filter.scala 202:51 Filter.scala 204:51]
  assign KernelConvolution_1_io_pixelVal_in_1 = _GEN_1764[3:0]; // @[Filter.scala 200:53 Filter.scala 202:51 Filter.scala 204:51]
  assign KernelConvolution_1_io_pixelVal_in_2 = _GEN_2634[3:0]; // @[Filter.scala 200:53 Filter.scala 202:51 Filter.scala 204:51]
  assign KernelConvolution_1_io_pixelVal_in_3 = _GEN_3504[3:0]; // @[Filter.scala 200:53 Filter.scala 202:51 Filter.scala 204:51]
  assign KernelConvolution_1_io_pixelVal_in_4 = _GEN_4374[3:0]; // @[Filter.scala 200:53 Filter.scala 202:51 Filter.scala 204:51]
  assign KernelConvolution_1_io_pixelVal_in_5 = _GEN_5244[3:0]; // @[Filter.scala 200:53 Filter.scala 202:51 Filter.scala 204:51]
  assign KernelConvolution_1_io_pixelVal_in_6 = _GEN_6114[3:0]; // @[Filter.scala 200:53 Filter.scala 202:51 Filter.scala 204:51]
  assign KernelConvolution_1_io_pixelVal_in_7 = _GEN_6984[3:0]; // @[Filter.scala 200:53 Filter.scala 202:51 Filter.scala 204:51]
  assign KernelConvolution_2_clock = clock;
  assign KernelConvolution_2_reset = reset;
  assign KernelConvolution_2_io_kernelVal_in = _GEN_7341 & _GEN_7268 ? $signed(5'sh0) : $signed(_GEN_55); // @[Filter.scala 186:41]
  assign KernelConvolution_2_io_pixelVal_in_0 = _GEN_1040[3:0]; // @[Filter.scala 200:53 Filter.scala 202:51 Filter.scala 204:51]
  assign KernelConvolution_2_io_pixelVal_in_1 = _GEN_1910[3:0]; // @[Filter.scala 200:53 Filter.scala 202:51 Filter.scala 204:51]
  assign KernelConvolution_2_io_pixelVal_in_2 = _GEN_2780[3:0]; // @[Filter.scala 200:53 Filter.scala 202:51 Filter.scala 204:51]
  assign KernelConvolution_2_io_pixelVal_in_3 = _GEN_3650[3:0]; // @[Filter.scala 200:53 Filter.scala 202:51 Filter.scala 204:51]
  assign KernelConvolution_2_io_pixelVal_in_4 = _GEN_4520[3:0]; // @[Filter.scala 200:53 Filter.scala 202:51 Filter.scala 204:51]
  assign KernelConvolution_2_io_pixelVal_in_5 = _GEN_5390[3:0]; // @[Filter.scala 200:53 Filter.scala 202:51 Filter.scala 204:51]
  assign KernelConvolution_2_io_pixelVal_in_6 = _GEN_6260[3:0]; // @[Filter.scala 200:53 Filter.scala 202:51 Filter.scala 204:51]
  assign KernelConvolution_2_io_pixelVal_in_7 = _GEN_7130[3:0]; // @[Filter.scala 200:53 Filter.scala 202:51 Filter.scala 204:51]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  kernelCounter = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  imageCounterX = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  imageCounterY = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  pixelIndex = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  pixOut_0_0 = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  pixOut_0_1 = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  pixOut_0_2 = _RAND_6[8:0];
  _RAND_7 = {1{`RANDOM}};
  pixOut_0_3 = _RAND_7[8:0];
  _RAND_8 = {1{`RANDOM}};
  pixOut_0_4 = _RAND_8[8:0];
  _RAND_9 = {1{`RANDOM}};
  pixOut_0_5 = _RAND_9[8:0];
  _RAND_10 = {1{`RANDOM}};
  pixOut_0_6 = _RAND_10[8:0];
  _RAND_11 = {1{`RANDOM}};
  pixOut_0_7 = _RAND_11[8:0];
  _RAND_12 = {1{`RANDOM}};
  pixOut_1_0 = _RAND_12[8:0];
  _RAND_13 = {1{`RANDOM}};
  pixOut_1_1 = _RAND_13[8:0];
  _RAND_14 = {1{`RANDOM}};
  pixOut_1_2 = _RAND_14[8:0];
  _RAND_15 = {1{`RANDOM}};
  pixOut_1_3 = _RAND_15[8:0];
  _RAND_16 = {1{`RANDOM}};
  pixOut_1_4 = _RAND_16[8:0];
  _RAND_17 = {1{`RANDOM}};
  pixOut_1_5 = _RAND_17[8:0];
  _RAND_18 = {1{`RANDOM}};
  pixOut_1_6 = _RAND_18[8:0];
  _RAND_19 = {1{`RANDOM}};
  pixOut_1_7 = _RAND_19[8:0];
  _RAND_20 = {1{`RANDOM}};
  pixOut_2_0 = _RAND_20[8:0];
  _RAND_21 = {1{`RANDOM}};
  pixOut_2_1 = _RAND_21[8:0];
  _RAND_22 = {1{`RANDOM}};
  pixOut_2_2 = _RAND_22[8:0];
  _RAND_23 = {1{`RANDOM}};
  pixOut_2_3 = _RAND_23[8:0];
  _RAND_24 = {1{`RANDOM}};
  pixOut_2_4 = _RAND_24[8:0];
  _RAND_25 = {1{`RANDOM}};
  pixOut_2_5 = _RAND_25[8:0];
  _RAND_26 = {1{`RANDOM}};
  pixOut_2_6 = _RAND_26[8:0];
  _RAND_27 = {1{`RANDOM}};
  pixOut_2_7 = _RAND_27[8:0];
  _RAND_28 = {1{`RANDOM}};
  validOut = _RAND_28[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      kernelCounter <= 4'h0;
    end else if (kernelCountReset) begin
      kernelCounter <= 4'h0;
    end else begin
      kernelCounter <= _T_14;
    end
    if (reset) begin
      imageCounterX <= 2'h0;
    end else if (imageCounterXReset) begin
      imageCounterX <= 2'h0;
    end else begin
      imageCounterX <= _T_20;
    end
    if (reset) begin
      imageCounterY <= 2'h0;
    end else if (imageCounterXReset) begin
      if (_T_21) begin
        imageCounterY <= 2'h0;
      end else begin
        imageCounterY <= _T_23;
      end
    end
    if (reset) begin
      pixelIndex <= 32'h0;
    end else if (kernelCountReset) begin
      if (_T_831) begin
        pixelIndex <= 32'h0;
      end else begin
        pixelIndex <= _T_829;
      end
    end
    if (reset) begin
      pixOut_0_0 <= 9'sh0;
    end else begin
      pixOut_0_0 <= _T_564[8:0];
    end
    if (reset) begin
      pixOut_0_1 <= 9'sh0;
    end else begin
      pixOut_0_1 <= _T_575[8:0];
    end
    if (reset) begin
      pixOut_0_2 <= 9'sh0;
    end else begin
      pixOut_0_2 <= _T_586[8:0];
    end
    if (reset) begin
      pixOut_0_3 <= 9'sh0;
    end else begin
      pixOut_0_3 <= _T_597[8:0];
    end
    if (reset) begin
      pixOut_0_4 <= 9'sh0;
    end else begin
      pixOut_0_4 <= _T_608[8:0];
    end
    if (reset) begin
      pixOut_0_5 <= 9'sh0;
    end else begin
      pixOut_0_5 <= _T_619[8:0];
    end
    if (reset) begin
      pixOut_0_6 <= 9'sh0;
    end else begin
      pixOut_0_6 <= _T_630[8:0];
    end
    if (reset) begin
      pixOut_0_7 <= 9'sh0;
    end else begin
      pixOut_0_7 <= _T_641[8:0];
    end
    if (reset) begin
      pixOut_1_0 <= 9'sh0;
    end else begin
      pixOut_1_0 <= _T_652[8:0];
    end
    if (reset) begin
      pixOut_1_1 <= 9'sh0;
    end else begin
      pixOut_1_1 <= _T_663[8:0];
    end
    if (reset) begin
      pixOut_1_2 <= 9'sh0;
    end else begin
      pixOut_1_2 <= _T_674[8:0];
    end
    if (reset) begin
      pixOut_1_3 <= 9'sh0;
    end else begin
      pixOut_1_3 <= _T_685[8:0];
    end
    if (reset) begin
      pixOut_1_4 <= 9'sh0;
    end else begin
      pixOut_1_4 <= _T_696[8:0];
    end
    if (reset) begin
      pixOut_1_5 <= 9'sh0;
    end else begin
      pixOut_1_5 <= _T_707[8:0];
    end
    if (reset) begin
      pixOut_1_6 <= 9'sh0;
    end else begin
      pixOut_1_6 <= _T_718[8:0];
    end
    if (reset) begin
      pixOut_1_7 <= 9'sh0;
    end else begin
      pixOut_1_7 <= _T_729[8:0];
    end
    if (reset) begin
      pixOut_2_0 <= 9'sh0;
    end else begin
      pixOut_2_0 <= _T_740[8:0];
    end
    if (reset) begin
      pixOut_2_1 <= 9'sh0;
    end else begin
      pixOut_2_1 <= _T_751[8:0];
    end
    if (reset) begin
      pixOut_2_2 <= 9'sh0;
    end else begin
      pixOut_2_2 <= _T_762[8:0];
    end
    if (reset) begin
      pixOut_2_3 <= 9'sh0;
    end else begin
      pixOut_2_3 <= _T_773[8:0];
    end
    if (reset) begin
      pixOut_2_4 <= 9'sh0;
    end else begin
      pixOut_2_4 <= _T_784[8:0];
    end
    if (reset) begin
      pixOut_2_5 <= 9'sh0;
    end else begin
      pixOut_2_5 <= _T_795[8:0];
    end
    if (reset) begin
      pixOut_2_6 <= 9'sh0;
    end else begin
      pixOut_2_6 <= _T_806[8:0];
    end
    if (reset) begin
      pixOut_2_7 <= 9'sh0;
    end else begin
      pixOut_2_7 <= _T_817[8:0];
    end
    if (reset) begin
      validOut <= 1'h0;
    end else begin
      validOut <= KernelConvolution_io_valid_out;
    end
  end
endmodule
module VideoBuffer(
  input         clock,
  input         reset,
  input  [3:0]  io_pixelVal_in_0_0,
  input  [3:0]  io_pixelVal_in_0_1,
  input  [3:0]  io_pixelVal_in_0_2,
  input  [3:0]  io_pixelVal_in_0_3,
  input  [3:0]  io_pixelVal_in_0_4,
  input  [3:0]  io_pixelVal_in_0_5,
  input  [3:0]  io_pixelVal_in_0_6,
  input  [3:0]  io_pixelVal_in_0_7,
  input  [3:0]  io_pixelVal_in_1_0,
  input  [3:0]  io_pixelVal_in_1_1,
  input  [3:0]  io_pixelVal_in_1_2,
  input  [3:0]  io_pixelVal_in_1_3,
  input  [3:0]  io_pixelVal_in_1_4,
  input  [3:0]  io_pixelVal_in_1_5,
  input  [3:0]  io_pixelVal_in_1_6,
  input  [3:0]  io_pixelVal_in_1_7,
  input  [3:0]  io_pixelVal_in_2_0,
  input  [3:0]  io_pixelVal_in_2_1,
  input  [3:0]  io_pixelVal_in_2_2,
  input  [3:0]  io_pixelVal_in_2_3,
  input  [3:0]  io_pixelVal_in_2_4,
  input  [3:0]  io_pixelVal_in_2_5,
  input  [3:0]  io_pixelVal_in_2_6,
  input  [3:0]  io_pixelVal_in_2_7,
  input         io_valid_in,
  input  [10:0] io_rowIndex,
  input  [10:0] io_colIndex,
  output [3:0]  io_pixelVal_out_0,
  output [3:0]  io_pixelVal_out_1,
  output [3:0]  io_pixelVal_out_2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] image_0_0; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_1; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_2; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_3; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_4; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_5; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_6; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_7; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_8; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_9; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_10; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_11; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_12; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_13; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_14; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_15; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_16; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_17; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_18; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_19; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_20; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_21; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_22; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_23; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_24; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_25; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_26; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_27; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_28; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_29; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_30; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_31; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_32; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_33; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_34; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_35; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_36; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_37; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_38; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_39; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_40; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_41; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_42; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_43; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_44; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_45; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_46; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_47; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_48; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_49; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_50; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_51; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_52; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_53; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_54; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_55; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_56; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_57; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_58; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_59; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_60; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_61; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_62; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_63; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_64; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_65; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_66; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_67; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_68; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_69; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_70; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_71; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_72; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_73; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_74; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_75; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_76; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_77; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_78; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_79; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_80; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_81; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_82; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_83; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_84; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_85; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_86; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_87; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_88; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_89; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_90; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_91; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_92; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_93; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_94; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_95; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_96; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_97; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_98; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_99; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_100; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_101; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_102; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_103; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_104; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_105; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_106; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_107; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_108; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_109; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_110; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_111; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_112; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_113; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_114; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_115; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_116; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_117; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_118; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_119; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_120; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_121; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_122; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_123; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_124; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_125; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_126; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_127; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_128; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_129; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_130; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_131; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_132; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_133; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_134; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_135; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_136; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_137; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_138; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_139; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_140; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_141; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_142; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_143; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_1_0; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_1; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_2; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_3; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_4; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_5; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_6; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_7; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_8; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_9; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_10; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_11; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_12; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_13; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_14; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_15; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_16; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_17; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_18; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_19; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_20; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_21; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_22; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_23; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_24; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_25; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_26; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_27; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_28; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_29; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_30; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_31; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_32; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_33; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_34; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_35; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_36; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_37; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_38; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_39; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_40; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_41; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_42; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_43; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_44; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_45; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_46; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_47; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_48; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_49; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_50; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_51; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_52; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_53; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_54; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_55; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_56; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_57; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_58; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_59; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_60; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_61; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_62; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_63; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_64; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_65; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_66; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_67; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_68; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_69; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_70; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_71; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_72; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_73; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_74; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_75; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_76; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_77; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_78; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_79; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_80; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_81; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_82; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_83; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_84; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_85; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_86; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_87; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_88; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_89; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_90; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_91; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_92; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_93; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_94; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_95; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_96; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_97; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_98; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_99; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_100; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_101; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_102; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_103; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_104; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_105; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_106; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_107; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_108; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_109; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_110; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_111; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_112; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_113; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_114; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_115; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_116; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_117; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_118; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_119; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_120; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_121; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_122; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_123; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_124; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_125; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_126; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_127; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_128; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_129; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_130; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_131; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_132; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_133; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_134; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_135; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_136; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_137; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_138; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_139; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_140; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_141; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_142; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_143; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_2_0; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_1; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_2; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_3; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_4; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_5; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_6; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_7; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_8; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_9; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_10; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_11; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_12; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_13; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_14; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_15; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_16; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_17; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_18; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_19; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_20; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_21; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_22; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_23; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_24; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_25; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_26; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_27; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_28; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_29; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_30; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_31; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_32; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_33; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_34; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_35; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_36; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_37; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_38; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_39; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_40; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_41; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_42; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_43; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_44; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_45; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_46; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_47; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_48; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_49; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_50; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_51; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_52; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_53; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_54; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_55; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_56; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_57; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_58; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_59; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_60; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_61; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_62; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_63; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_64; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_65; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_66; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_67; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_68; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_69; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_70; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_71; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_72; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_73; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_74; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_75; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_76; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_77; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_78; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_79; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_80; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_81; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_82; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_83; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_84; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_85; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_86; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_87; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_88; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_89; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_90; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_91; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_92; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_93; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_94; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_95; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_96; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_97; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_98; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_99; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_100; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_101; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_102; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_103; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_104; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_105; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_106; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_107; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_108; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_109; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_110; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_111; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_112; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_113; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_114; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_115; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_116; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_117; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_118; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_119; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_120; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_121; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_122; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_123; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_124; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_125; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_126; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_127; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_128; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_129; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_130; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_131; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_132; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_133; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_134; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_135; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_136; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_137; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_138; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_139; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_140; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_141; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_142; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_143; // @[VideoBuffer.scala 21:25]
  reg [31:0] pixelIndex; // @[VideoBuffer.scala 24:33]
  wire [15:0] _T_3 = io_rowIndex * 11'h10; // @[VideoBuffer.scala 27:54]
  wire [15:0] _GEN_4322 = {{5'd0}, io_colIndex}; // @[VideoBuffer.scala 27:69]
  wire [15:0] _T_5 = _T_3 + _GEN_4322; // @[VideoBuffer.scala 27:69]
  wire [3:0] _GEN_1 = 8'h1 == _T_5[7:0] ? image_0_1 : image_0_0; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2 = 8'h2 == _T_5[7:0] ? image_0_2 : _GEN_1; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3 = 8'h3 == _T_5[7:0] ? image_0_3 : _GEN_2; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4 = 8'h4 == _T_5[7:0] ? image_0_4 : _GEN_3; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_5 = 8'h5 == _T_5[7:0] ? image_0_5 : _GEN_4; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_6 = 8'h6 == _T_5[7:0] ? image_0_6 : _GEN_5; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_7 = 8'h7 == _T_5[7:0] ? image_0_7 : _GEN_6; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_8 = 8'h8 == _T_5[7:0] ? image_0_8 : _GEN_7; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_9 = 8'h9 == _T_5[7:0] ? image_0_9 : _GEN_8; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_10 = 8'ha == _T_5[7:0] ? image_0_10 : _GEN_9; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_11 = 8'hb == _T_5[7:0] ? image_0_11 : _GEN_10; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_12 = 8'hc == _T_5[7:0] ? image_0_12 : _GEN_11; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_13 = 8'hd == _T_5[7:0] ? image_0_13 : _GEN_12; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_14 = 8'he == _T_5[7:0] ? image_0_14 : _GEN_13; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_15 = 8'hf == _T_5[7:0] ? image_0_15 : _GEN_14; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_16 = 8'h10 == _T_5[7:0] ? image_0_16 : _GEN_15; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_17 = 8'h11 == _T_5[7:0] ? image_0_17 : _GEN_16; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_18 = 8'h12 == _T_5[7:0] ? image_0_18 : _GEN_17; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_19 = 8'h13 == _T_5[7:0] ? image_0_19 : _GEN_18; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_20 = 8'h14 == _T_5[7:0] ? image_0_20 : _GEN_19; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_21 = 8'h15 == _T_5[7:0] ? image_0_21 : _GEN_20; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_22 = 8'h16 == _T_5[7:0] ? image_0_22 : _GEN_21; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_23 = 8'h17 == _T_5[7:0] ? image_0_23 : _GEN_22; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_24 = 8'h18 == _T_5[7:0] ? image_0_24 : _GEN_23; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_25 = 8'h19 == _T_5[7:0] ? image_0_25 : _GEN_24; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_26 = 8'h1a == _T_5[7:0] ? image_0_26 : _GEN_25; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_27 = 8'h1b == _T_5[7:0] ? image_0_27 : _GEN_26; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_28 = 8'h1c == _T_5[7:0] ? image_0_28 : _GEN_27; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_29 = 8'h1d == _T_5[7:0] ? image_0_29 : _GEN_28; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_30 = 8'h1e == _T_5[7:0] ? image_0_30 : _GEN_29; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_31 = 8'h1f == _T_5[7:0] ? image_0_31 : _GEN_30; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_32 = 8'h20 == _T_5[7:0] ? image_0_32 : _GEN_31; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_33 = 8'h21 == _T_5[7:0] ? image_0_33 : _GEN_32; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_34 = 8'h22 == _T_5[7:0] ? image_0_34 : _GEN_33; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_35 = 8'h23 == _T_5[7:0] ? image_0_35 : _GEN_34; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_36 = 8'h24 == _T_5[7:0] ? image_0_36 : _GEN_35; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_37 = 8'h25 == _T_5[7:0] ? image_0_37 : _GEN_36; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_38 = 8'h26 == _T_5[7:0] ? image_0_38 : _GEN_37; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_39 = 8'h27 == _T_5[7:0] ? image_0_39 : _GEN_38; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_40 = 8'h28 == _T_5[7:0] ? image_0_40 : _GEN_39; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_41 = 8'h29 == _T_5[7:0] ? image_0_41 : _GEN_40; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_42 = 8'h2a == _T_5[7:0] ? image_0_42 : _GEN_41; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_43 = 8'h2b == _T_5[7:0] ? image_0_43 : _GEN_42; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_44 = 8'h2c == _T_5[7:0] ? image_0_44 : _GEN_43; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_45 = 8'h2d == _T_5[7:0] ? image_0_45 : _GEN_44; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_46 = 8'h2e == _T_5[7:0] ? image_0_46 : _GEN_45; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_47 = 8'h2f == _T_5[7:0] ? image_0_47 : _GEN_46; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_48 = 8'h30 == _T_5[7:0] ? image_0_48 : _GEN_47; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_49 = 8'h31 == _T_5[7:0] ? image_0_49 : _GEN_48; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_50 = 8'h32 == _T_5[7:0] ? image_0_50 : _GEN_49; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_51 = 8'h33 == _T_5[7:0] ? image_0_51 : _GEN_50; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_52 = 8'h34 == _T_5[7:0] ? image_0_52 : _GEN_51; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_53 = 8'h35 == _T_5[7:0] ? image_0_53 : _GEN_52; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_54 = 8'h36 == _T_5[7:0] ? image_0_54 : _GEN_53; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_55 = 8'h37 == _T_5[7:0] ? image_0_55 : _GEN_54; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_56 = 8'h38 == _T_5[7:0] ? image_0_56 : _GEN_55; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_57 = 8'h39 == _T_5[7:0] ? image_0_57 : _GEN_56; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_58 = 8'h3a == _T_5[7:0] ? image_0_58 : _GEN_57; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_59 = 8'h3b == _T_5[7:0] ? image_0_59 : _GEN_58; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_60 = 8'h3c == _T_5[7:0] ? image_0_60 : _GEN_59; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_61 = 8'h3d == _T_5[7:0] ? image_0_61 : _GEN_60; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_62 = 8'h3e == _T_5[7:0] ? image_0_62 : _GEN_61; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_63 = 8'h3f == _T_5[7:0] ? image_0_63 : _GEN_62; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_64 = 8'h40 == _T_5[7:0] ? image_0_64 : _GEN_63; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_65 = 8'h41 == _T_5[7:0] ? image_0_65 : _GEN_64; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_66 = 8'h42 == _T_5[7:0] ? image_0_66 : _GEN_65; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_67 = 8'h43 == _T_5[7:0] ? image_0_67 : _GEN_66; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_68 = 8'h44 == _T_5[7:0] ? image_0_68 : _GEN_67; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_69 = 8'h45 == _T_5[7:0] ? image_0_69 : _GEN_68; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_70 = 8'h46 == _T_5[7:0] ? image_0_70 : _GEN_69; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_71 = 8'h47 == _T_5[7:0] ? image_0_71 : _GEN_70; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_72 = 8'h48 == _T_5[7:0] ? image_0_72 : _GEN_71; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_73 = 8'h49 == _T_5[7:0] ? image_0_73 : _GEN_72; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_74 = 8'h4a == _T_5[7:0] ? image_0_74 : _GEN_73; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_75 = 8'h4b == _T_5[7:0] ? image_0_75 : _GEN_74; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_76 = 8'h4c == _T_5[7:0] ? image_0_76 : _GEN_75; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_77 = 8'h4d == _T_5[7:0] ? image_0_77 : _GEN_76; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_78 = 8'h4e == _T_5[7:0] ? image_0_78 : _GEN_77; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_79 = 8'h4f == _T_5[7:0] ? image_0_79 : _GEN_78; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_80 = 8'h50 == _T_5[7:0] ? image_0_80 : _GEN_79; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_81 = 8'h51 == _T_5[7:0] ? image_0_81 : _GEN_80; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_82 = 8'h52 == _T_5[7:0] ? image_0_82 : _GEN_81; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_83 = 8'h53 == _T_5[7:0] ? image_0_83 : _GEN_82; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_84 = 8'h54 == _T_5[7:0] ? image_0_84 : _GEN_83; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_85 = 8'h55 == _T_5[7:0] ? image_0_85 : _GEN_84; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_86 = 8'h56 == _T_5[7:0] ? image_0_86 : _GEN_85; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_87 = 8'h57 == _T_5[7:0] ? image_0_87 : _GEN_86; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_88 = 8'h58 == _T_5[7:0] ? image_0_88 : _GEN_87; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_89 = 8'h59 == _T_5[7:0] ? image_0_89 : _GEN_88; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_90 = 8'h5a == _T_5[7:0] ? image_0_90 : _GEN_89; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_91 = 8'h5b == _T_5[7:0] ? image_0_91 : _GEN_90; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_92 = 8'h5c == _T_5[7:0] ? image_0_92 : _GEN_91; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_93 = 8'h5d == _T_5[7:0] ? image_0_93 : _GEN_92; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_94 = 8'h5e == _T_5[7:0] ? image_0_94 : _GEN_93; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_95 = 8'h5f == _T_5[7:0] ? image_0_95 : _GEN_94; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_96 = 8'h60 == _T_5[7:0] ? image_0_96 : _GEN_95; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_97 = 8'h61 == _T_5[7:0] ? image_0_97 : _GEN_96; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_98 = 8'h62 == _T_5[7:0] ? image_0_98 : _GEN_97; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_99 = 8'h63 == _T_5[7:0] ? image_0_99 : _GEN_98; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_100 = 8'h64 == _T_5[7:0] ? image_0_100 : _GEN_99; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_101 = 8'h65 == _T_5[7:0] ? image_0_101 : _GEN_100; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_102 = 8'h66 == _T_5[7:0] ? image_0_102 : _GEN_101; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_103 = 8'h67 == _T_5[7:0] ? image_0_103 : _GEN_102; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_104 = 8'h68 == _T_5[7:0] ? image_0_104 : _GEN_103; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_105 = 8'h69 == _T_5[7:0] ? image_0_105 : _GEN_104; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_106 = 8'h6a == _T_5[7:0] ? image_0_106 : _GEN_105; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_107 = 8'h6b == _T_5[7:0] ? image_0_107 : _GEN_106; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_108 = 8'h6c == _T_5[7:0] ? image_0_108 : _GEN_107; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_109 = 8'h6d == _T_5[7:0] ? image_0_109 : _GEN_108; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_110 = 8'h6e == _T_5[7:0] ? image_0_110 : _GEN_109; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_111 = 8'h6f == _T_5[7:0] ? image_0_111 : _GEN_110; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_112 = 8'h70 == _T_5[7:0] ? image_0_112 : _GEN_111; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_113 = 8'h71 == _T_5[7:0] ? image_0_113 : _GEN_112; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_114 = 8'h72 == _T_5[7:0] ? image_0_114 : _GEN_113; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_115 = 8'h73 == _T_5[7:0] ? image_0_115 : _GEN_114; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_116 = 8'h74 == _T_5[7:0] ? image_0_116 : _GEN_115; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_117 = 8'h75 == _T_5[7:0] ? image_0_117 : _GEN_116; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_118 = 8'h76 == _T_5[7:0] ? image_0_118 : _GEN_117; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_119 = 8'h77 == _T_5[7:0] ? image_0_119 : _GEN_118; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_120 = 8'h78 == _T_5[7:0] ? image_0_120 : _GEN_119; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_121 = 8'h79 == _T_5[7:0] ? image_0_121 : _GEN_120; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_122 = 8'h7a == _T_5[7:0] ? image_0_122 : _GEN_121; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_123 = 8'h7b == _T_5[7:0] ? image_0_123 : _GEN_122; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_124 = 8'h7c == _T_5[7:0] ? image_0_124 : _GEN_123; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_125 = 8'h7d == _T_5[7:0] ? image_0_125 : _GEN_124; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_126 = 8'h7e == _T_5[7:0] ? image_0_126 : _GEN_125; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_127 = 8'h7f == _T_5[7:0] ? image_0_127 : _GEN_126; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_128 = 8'h80 == _T_5[7:0] ? image_0_128 : _GEN_127; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_129 = 8'h81 == _T_5[7:0] ? image_0_129 : _GEN_128; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_130 = 8'h82 == _T_5[7:0] ? image_0_130 : _GEN_129; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_131 = 8'h83 == _T_5[7:0] ? image_0_131 : _GEN_130; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_132 = 8'h84 == _T_5[7:0] ? image_0_132 : _GEN_131; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_133 = 8'h85 == _T_5[7:0] ? image_0_133 : _GEN_132; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_134 = 8'h86 == _T_5[7:0] ? image_0_134 : _GEN_133; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_135 = 8'h87 == _T_5[7:0] ? image_0_135 : _GEN_134; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_136 = 8'h88 == _T_5[7:0] ? image_0_136 : _GEN_135; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_137 = 8'h89 == _T_5[7:0] ? image_0_137 : _GEN_136; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_138 = 8'h8a == _T_5[7:0] ? image_0_138 : _GEN_137; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_139 = 8'h8b == _T_5[7:0] ? image_0_139 : _GEN_138; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_140 = 8'h8c == _T_5[7:0] ? image_0_140 : _GEN_139; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_141 = 8'h8d == _T_5[7:0] ? image_0_141 : _GEN_140; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_142 = 8'h8e == _T_5[7:0] ? image_0_142 : _GEN_141; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_145 = 8'h1 == _T_5[7:0] ? image_1_1 : image_1_0; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_146 = 8'h2 == _T_5[7:0] ? image_1_2 : _GEN_145; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_147 = 8'h3 == _T_5[7:0] ? image_1_3 : _GEN_146; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_148 = 8'h4 == _T_5[7:0] ? image_1_4 : _GEN_147; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_149 = 8'h5 == _T_5[7:0] ? image_1_5 : _GEN_148; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_150 = 8'h6 == _T_5[7:0] ? image_1_6 : _GEN_149; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_151 = 8'h7 == _T_5[7:0] ? image_1_7 : _GEN_150; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_152 = 8'h8 == _T_5[7:0] ? image_1_8 : _GEN_151; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_153 = 8'h9 == _T_5[7:0] ? image_1_9 : _GEN_152; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_154 = 8'ha == _T_5[7:0] ? image_1_10 : _GEN_153; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_155 = 8'hb == _T_5[7:0] ? image_1_11 : _GEN_154; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_156 = 8'hc == _T_5[7:0] ? image_1_12 : _GEN_155; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_157 = 8'hd == _T_5[7:0] ? image_1_13 : _GEN_156; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_158 = 8'he == _T_5[7:0] ? image_1_14 : _GEN_157; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_159 = 8'hf == _T_5[7:0] ? image_1_15 : _GEN_158; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_160 = 8'h10 == _T_5[7:0] ? image_1_16 : _GEN_159; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_161 = 8'h11 == _T_5[7:0] ? image_1_17 : _GEN_160; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_162 = 8'h12 == _T_5[7:0] ? image_1_18 : _GEN_161; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_163 = 8'h13 == _T_5[7:0] ? image_1_19 : _GEN_162; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_164 = 8'h14 == _T_5[7:0] ? image_1_20 : _GEN_163; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_165 = 8'h15 == _T_5[7:0] ? image_1_21 : _GEN_164; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_166 = 8'h16 == _T_5[7:0] ? image_1_22 : _GEN_165; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_167 = 8'h17 == _T_5[7:0] ? image_1_23 : _GEN_166; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_168 = 8'h18 == _T_5[7:0] ? image_1_24 : _GEN_167; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_169 = 8'h19 == _T_5[7:0] ? image_1_25 : _GEN_168; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_170 = 8'h1a == _T_5[7:0] ? image_1_26 : _GEN_169; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_171 = 8'h1b == _T_5[7:0] ? image_1_27 : _GEN_170; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_172 = 8'h1c == _T_5[7:0] ? image_1_28 : _GEN_171; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_173 = 8'h1d == _T_5[7:0] ? image_1_29 : _GEN_172; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_174 = 8'h1e == _T_5[7:0] ? image_1_30 : _GEN_173; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_175 = 8'h1f == _T_5[7:0] ? image_1_31 : _GEN_174; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_176 = 8'h20 == _T_5[7:0] ? image_1_32 : _GEN_175; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_177 = 8'h21 == _T_5[7:0] ? image_1_33 : _GEN_176; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_178 = 8'h22 == _T_5[7:0] ? image_1_34 : _GEN_177; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_179 = 8'h23 == _T_5[7:0] ? image_1_35 : _GEN_178; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_180 = 8'h24 == _T_5[7:0] ? image_1_36 : _GEN_179; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_181 = 8'h25 == _T_5[7:0] ? image_1_37 : _GEN_180; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_182 = 8'h26 == _T_5[7:0] ? image_1_38 : _GEN_181; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_183 = 8'h27 == _T_5[7:0] ? image_1_39 : _GEN_182; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_184 = 8'h28 == _T_5[7:0] ? image_1_40 : _GEN_183; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_185 = 8'h29 == _T_5[7:0] ? image_1_41 : _GEN_184; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_186 = 8'h2a == _T_5[7:0] ? image_1_42 : _GEN_185; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_187 = 8'h2b == _T_5[7:0] ? image_1_43 : _GEN_186; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_188 = 8'h2c == _T_5[7:0] ? image_1_44 : _GEN_187; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_189 = 8'h2d == _T_5[7:0] ? image_1_45 : _GEN_188; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_190 = 8'h2e == _T_5[7:0] ? image_1_46 : _GEN_189; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_191 = 8'h2f == _T_5[7:0] ? image_1_47 : _GEN_190; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_192 = 8'h30 == _T_5[7:0] ? image_1_48 : _GEN_191; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_193 = 8'h31 == _T_5[7:0] ? image_1_49 : _GEN_192; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_194 = 8'h32 == _T_5[7:0] ? image_1_50 : _GEN_193; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_195 = 8'h33 == _T_5[7:0] ? image_1_51 : _GEN_194; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_196 = 8'h34 == _T_5[7:0] ? image_1_52 : _GEN_195; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_197 = 8'h35 == _T_5[7:0] ? image_1_53 : _GEN_196; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_198 = 8'h36 == _T_5[7:0] ? image_1_54 : _GEN_197; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_199 = 8'h37 == _T_5[7:0] ? image_1_55 : _GEN_198; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_200 = 8'h38 == _T_5[7:0] ? image_1_56 : _GEN_199; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_201 = 8'h39 == _T_5[7:0] ? image_1_57 : _GEN_200; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_202 = 8'h3a == _T_5[7:0] ? image_1_58 : _GEN_201; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_203 = 8'h3b == _T_5[7:0] ? image_1_59 : _GEN_202; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_204 = 8'h3c == _T_5[7:0] ? image_1_60 : _GEN_203; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_205 = 8'h3d == _T_5[7:0] ? image_1_61 : _GEN_204; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_206 = 8'h3e == _T_5[7:0] ? image_1_62 : _GEN_205; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_207 = 8'h3f == _T_5[7:0] ? image_1_63 : _GEN_206; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_208 = 8'h40 == _T_5[7:0] ? image_1_64 : _GEN_207; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_209 = 8'h41 == _T_5[7:0] ? image_1_65 : _GEN_208; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_210 = 8'h42 == _T_5[7:0] ? image_1_66 : _GEN_209; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_211 = 8'h43 == _T_5[7:0] ? image_1_67 : _GEN_210; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_212 = 8'h44 == _T_5[7:0] ? image_1_68 : _GEN_211; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_213 = 8'h45 == _T_5[7:0] ? image_1_69 : _GEN_212; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_214 = 8'h46 == _T_5[7:0] ? image_1_70 : _GEN_213; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_215 = 8'h47 == _T_5[7:0] ? image_1_71 : _GEN_214; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_216 = 8'h48 == _T_5[7:0] ? image_1_72 : _GEN_215; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_217 = 8'h49 == _T_5[7:0] ? image_1_73 : _GEN_216; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_218 = 8'h4a == _T_5[7:0] ? image_1_74 : _GEN_217; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_219 = 8'h4b == _T_5[7:0] ? image_1_75 : _GEN_218; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_220 = 8'h4c == _T_5[7:0] ? image_1_76 : _GEN_219; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_221 = 8'h4d == _T_5[7:0] ? image_1_77 : _GEN_220; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_222 = 8'h4e == _T_5[7:0] ? image_1_78 : _GEN_221; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_223 = 8'h4f == _T_5[7:0] ? image_1_79 : _GEN_222; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_224 = 8'h50 == _T_5[7:0] ? image_1_80 : _GEN_223; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_225 = 8'h51 == _T_5[7:0] ? image_1_81 : _GEN_224; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_226 = 8'h52 == _T_5[7:0] ? image_1_82 : _GEN_225; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_227 = 8'h53 == _T_5[7:0] ? image_1_83 : _GEN_226; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_228 = 8'h54 == _T_5[7:0] ? image_1_84 : _GEN_227; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_229 = 8'h55 == _T_5[7:0] ? image_1_85 : _GEN_228; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_230 = 8'h56 == _T_5[7:0] ? image_1_86 : _GEN_229; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_231 = 8'h57 == _T_5[7:0] ? image_1_87 : _GEN_230; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_232 = 8'h58 == _T_5[7:0] ? image_1_88 : _GEN_231; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_233 = 8'h59 == _T_5[7:0] ? image_1_89 : _GEN_232; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_234 = 8'h5a == _T_5[7:0] ? image_1_90 : _GEN_233; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_235 = 8'h5b == _T_5[7:0] ? image_1_91 : _GEN_234; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_236 = 8'h5c == _T_5[7:0] ? image_1_92 : _GEN_235; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_237 = 8'h5d == _T_5[7:0] ? image_1_93 : _GEN_236; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_238 = 8'h5e == _T_5[7:0] ? image_1_94 : _GEN_237; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_239 = 8'h5f == _T_5[7:0] ? image_1_95 : _GEN_238; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_240 = 8'h60 == _T_5[7:0] ? image_1_96 : _GEN_239; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_241 = 8'h61 == _T_5[7:0] ? image_1_97 : _GEN_240; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_242 = 8'h62 == _T_5[7:0] ? image_1_98 : _GEN_241; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_243 = 8'h63 == _T_5[7:0] ? image_1_99 : _GEN_242; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_244 = 8'h64 == _T_5[7:0] ? image_1_100 : _GEN_243; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_245 = 8'h65 == _T_5[7:0] ? image_1_101 : _GEN_244; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_246 = 8'h66 == _T_5[7:0] ? image_1_102 : _GEN_245; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_247 = 8'h67 == _T_5[7:0] ? image_1_103 : _GEN_246; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_248 = 8'h68 == _T_5[7:0] ? image_1_104 : _GEN_247; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_249 = 8'h69 == _T_5[7:0] ? image_1_105 : _GEN_248; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_250 = 8'h6a == _T_5[7:0] ? image_1_106 : _GEN_249; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_251 = 8'h6b == _T_5[7:0] ? image_1_107 : _GEN_250; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_252 = 8'h6c == _T_5[7:0] ? image_1_108 : _GEN_251; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_253 = 8'h6d == _T_5[7:0] ? image_1_109 : _GEN_252; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_254 = 8'h6e == _T_5[7:0] ? image_1_110 : _GEN_253; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_255 = 8'h6f == _T_5[7:0] ? image_1_111 : _GEN_254; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_256 = 8'h70 == _T_5[7:0] ? image_1_112 : _GEN_255; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_257 = 8'h71 == _T_5[7:0] ? image_1_113 : _GEN_256; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_258 = 8'h72 == _T_5[7:0] ? image_1_114 : _GEN_257; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_259 = 8'h73 == _T_5[7:0] ? image_1_115 : _GEN_258; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_260 = 8'h74 == _T_5[7:0] ? image_1_116 : _GEN_259; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_261 = 8'h75 == _T_5[7:0] ? image_1_117 : _GEN_260; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_262 = 8'h76 == _T_5[7:0] ? image_1_118 : _GEN_261; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_263 = 8'h77 == _T_5[7:0] ? image_1_119 : _GEN_262; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_264 = 8'h78 == _T_5[7:0] ? image_1_120 : _GEN_263; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_265 = 8'h79 == _T_5[7:0] ? image_1_121 : _GEN_264; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_266 = 8'h7a == _T_5[7:0] ? image_1_122 : _GEN_265; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_267 = 8'h7b == _T_5[7:0] ? image_1_123 : _GEN_266; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_268 = 8'h7c == _T_5[7:0] ? image_1_124 : _GEN_267; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_269 = 8'h7d == _T_5[7:0] ? image_1_125 : _GEN_268; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_270 = 8'h7e == _T_5[7:0] ? image_1_126 : _GEN_269; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_271 = 8'h7f == _T_5[7:0] ? image_1_127 : _GEN_270; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_272 = 8'h80 == _T_5[7:0] ? image_1_128 : _GEN_271; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_273 = 8'h81 == _T_5[7:0] ? image_1_129 : _GEN_272; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_274 = 8'h82 == _T_5[7:0] ? image_1_130 : _GEN_273; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_275 = 8'h83 == _T_5[7:0] ? image_1_131 : _GEN_274; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_276 = 8'h84 == _T_5[7:0] ? image_1_132 : _GEN_275; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_277 = 8'h85 == _T_5[7:0] ? image_1_133 : _GEN_276; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_278 = 8'h86 == _T_5[7:0] ? image_1_134 : _GEN_277; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_279 = 8'h87 == _T_5[7:0] ? image_1_135 : _GEN_278; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_280 = 8'h88 == _T_5[7:0] ? image_1_136 : _GEN_279; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_281 = 8'h89 == _T_5[7:0] ? image_1_137 : _GEN_280; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_282 = 8'h8a == _T_5[7:0] ? image_1_138 : _GEN_281; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_283 = 8'h8b == _T_5[7:0] ? image_1_139 : _GEN_282; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_284 = 8'h8c == _T_5[7:0] ? image_1_140 : _GEN_283; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_285 = 8'h8d == _T_5[7:0] ? image_1_141 : _GEN_284; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_286 = 8'h8e == _T_5[7:0] ? image_1_142 : _GEN_285; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_289 = 8'h1 == _T_5[7:0] ? image_2_1 : image_2_0; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_290 = 8'h2 == _T_5[7:0] ? image_2_2 : _GEN_289; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_291 = 8'h3 == _T_5[7:0] ? image_2_3 : _GEN_290; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_292 = 8'h4 == _T_5[7:0] ? image_2_4 : _GEN_291; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_293 = 8'h5 == _T_5[7:0] ? image_2_5 : _GEN_292; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_294 = 8'h6 == _T_5[7:0] ? image_2_6 : _GEN_293; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_295 = 8'h7 == _T_5[7:0] ? image_2_7 : _GEN_294; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_296 = 8'h8 == _T_5[7:0] ? image_2_8 : _GEN_295; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_297 = 8'h9 == _T_5[7:0] ? image_2_9 : _GEN_296; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_298 = 8'ha == _T_5[7:0] ? image_2_10 : _GEN_297; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_299 = 8'hb == _T_5[7:0] ? image_2_11 : _GEN_298; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_300 = 8'hc == _T_5[7:0] ? image_2_12 : _GEN_299; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_301 = 8'hd == _T_5[7:0] ? image_2_13 : _GEN_300; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_302 = 8'he == _T_5[7:0] ? image_2_14 : _GEN_301; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_303 = 8'hf == _T_5[7:0] ? image_2_15 : _GEN_302; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_304 = 8'h10 == _T_5[7:0] ? image_2_16 : _GEN_303; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_305 = 8'h11 == _T_5[7:0] ? image_2_17 : _GEN_304; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_306 = 8'h12 == _T_5[7:0] ? image_2_18 : _GEN_305; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_307 = 8'h13 == _T_5[7:0] ? image_2_19 : _GEN_306; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_308 = 8'h14 == _T_5[7:0] ? image_2_20 : _GEN_307; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_309 = 8'h15 == _T_5[7:0] ? image_2_21 : _GEN_308; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_310 = 8'h16 == _T_5[7:0] ? image_2_22 : _GEN_309; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_311 = 8'h17 == _T_5[7:0] ? image_2_23 : _GEN_310; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_312 = 8'h18 == _T_5[7:0] ? image_2_24 : _GEN_311; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_313 = 8'h19 == _T_5[7:0] ? image_2_25 : _GEN_312; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_314 = 8'h1a == _T_5[7:0] ? image_2_26 : _GEN_313; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_315 = 8'h1b == _T_5[7:0] ? image_2_27 : _GEN_314; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_316 = 8'h1c == _T_5[7:0] ? image_2_28 : _GEN_315; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_317 = 8'h1d == _T_5[7:0] ? image_2_29 : _GEN_316; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_318 = 8'h1e == _T_5[7:0] ? image_2_30 : _GEN_317; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_319 = 8'h1f == _T_5[7:0] ? image_2_31 : _GEN_318; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_320 = 8'h20 == _T_5[7:0] ? image_2_32 : _GEN_319; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_321 = 8'h21 == _T_5[7:0] ? image_2_33 : _GEN_320; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_322 = 8'h22 == _T_5[7:0] ? image_2_34 : _GEN_321; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_323 = 8'h23 == _T_5[7:0] ? image_2_35 : _GEN_322; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_324 = 8'h24 == _T_5[7:0] ? image_2_36 : _GEN_323; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_325 = 8'h25 == _T_5[7:0] ? image_2_37 : _GEN_324; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_326 = 8'h26 == _T_5[7:0] ? image_2_38 : _GEN_325; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_327 = 8'h27 == _T_5[7:0] ? image_2_39 : _GEN_326; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_328 = 8'h28 == _T_5[7:0] ? image_2_40 : _GEN_327; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_329 = 8'h29 == _T_5[7:0] ? image_2_41 : _GEN_328; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_330 = 8'h2a == _T_5[7:0] ? image_2_42 : _GEN_329; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_331 = 8'h2b == _T_5[7:0] ? image_2_43 : _GEN_330; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_332 = 8'h2c == _T_5[7:0] ? image_2_44 : _GEN_331; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_333 = 8'h2d == _T_5[7:0] ? image_2_45 : _GEN_332; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_334 = 8'h2e == _T_5[7:0] ? image_2_46 : _GEN_333; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_335 = 8'h2f == _T_5[7:0] ? image_2_47 : _GEN_334; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_336 = 8'h30 == _T_5[7:0] ? image_2_48 : _GEN_335; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_337 = 8'h31 == _T_5[7:0] ? image_2_49 : _GEN_336; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_338 = 8'h32 == _T_5[7:0] ? image_2_50 : _GEN_337; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_339 = 8'h33 == _T_5[7:0] ? image_2_51 : _GEN_338; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_340 = 8'h34 == _T_5[7:0] ? image_2_52 : _GEN_339; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_341 = 8'h35 == _T_5[7:0] ? image_2_53 : _GEN_340; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_342 = 8'h36 == _T_5[7:0] ? image_2_54 : _GEN_341; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_343 = 8'h37 == _T_5[7:0] ? image_2_55 : _GEN_342; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_344 = 8'h38 == _T_5[7:0] ? image_2_56 : _GEN_343; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_345 = 8'h39 == _T_5[7:0] ? image_2_57 : _GEN_344; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_346 = 8'h3a == _T_5[7:0] ? image_2_58 : _GEN_345; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_347 = 8'h3b == _T_5[7:0] ? image_2_59 : _GEN_346; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_348 = 8'h3c == _T_5[7:0] ? image_2_60 : _GEN_347; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_349 = 8'h3d == _T_5[7:0] ? image_2_61 : _GEN_348; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_350 = 8'h3e == _T_5[7:0] ? image_2_62 : _GEN_349; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_351 = 8'h3f == _T_5[7:0] ? image_2_63 : _GEN_350; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_352 = 8'h40 == _T_5[7:0] ? image_2_64 : _GEN_351; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_353 = 8'h41 == _T_5[7:0] ? image_2_65 : _GEN_352; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_354 = 8'h42 == _T_5[7:0] ? image_2_66 : _GEN_353; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_355 = 8'h43 == _T_5[7:0] ? image_2_67 : _GEN_354; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_356 = 8'h44 == _T_5[7:0] ? image_2_68 : _GEN_355; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_357 = 8'h45 == _T_5[7:0] ? image_2_69 : _GEN_356; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_358 = 8'h46 == _T_5[7:0] ? image_2_70 : _GEN_357; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_359 = 8'h47 == _T_5[7:0] ? image_2_71 : _GEN_358; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_360 = 8'h48 == _T_5[7:0] ? image_2_72 : _GEN_359; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_361 = 8'h49 == _T_5[7:0] ? image_2_73 : _GEN_360; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_362 = 8'h4a == _T_5[7:0] ? image_2_74 : _GEN_361; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_363 = 8'h4b == _T_5[7:0] ? image_2_75 : _GEN_362; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_364 = 8'h4c == _T_5[7:0] ? image_2_76 : _GEN_363; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_365 = 8'h4d == _T_5[7:0] ? image_2_77 : _GEN_364; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_366 = 8'h4e == _T_5[7:0] ? image_2_78 : _GEN_365; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_367 = 8'h4f == _T_5[7:0] ? image_2_79 : _GEN_366; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_368 = 8'h50 == _T_5[7:0] ? image_2_80 : _GEN_367; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_369 = 8'h51 == _T_5[7:0] ? image_2_81 : _GEN_368; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_370 = 8'h52 == _T_5[7:0] ? image_2_82 : _GEN_369; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_371 = 8'h53 == _T_5[7:0] ? image_2_83 : _GEN_370; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_372 = 8'h54 == _T_5[7:0] ? image_2_84 : _GEN_371; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_373 = 8'h55 == _T_5[7:0] ? image_2_85 : _GEN_372; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_374 = 8'h56 == _T_5[7:0] ? image_2_86 : _GEN_373; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_375 = 8'h57 == _T_5[7:0] ? image_2_87 : _GEN_374; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_376 = 8'h58 == _T_5[7:0] ? image_2_88 : _GEN_375; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_377 = 8'h59 == _T_5[7:0] ? image_2_89 : _GEN_376; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_378 = 8'h5a == _T_5[7:0] ? image_2_90 : _GEN_377; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_379 = 8'h5b == _T_5[7:0] ? image_2_91 : _GEN_378; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_380 = 8'h5c == _T_5[7:0] ? image_2_92 : _GEN_379; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_381 = 8'h5d == _T_5[7:0] ? image_2_93 : _GEN_380; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_382 = 8'h5e == _T_5[7:0] ? image_2_94 : _GEN_381; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_383 = 8'h5f == _T_5[7:0] ? image_2_95 : _GEN_382; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_384 = 8'h60 == _T_5[7:0] ? image_2_96 : _GEN_383; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_385 = 8'h61 == _T_5[7:0] ? image_2_97 : _GEN_384; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_386 = 8'h62 == _T_5[7:0] ? image_2_98 : _GEN_385; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_387 = 8'h63 == _T_5[7:0] ? image_2_99 : _GEN_386; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_388 = 8'h64 == _T_5[7:0] ? image_2_100 : _GEN_387; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_389 = 8'h65 == _T_5[7:0] ? image_2_101 : _GEN_388; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_390 = 8'h66 == _T_5[7:0] ? image_2_102 : _GEN_389; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_391 = 8'h67 == _T_5[7:0] ? image_2_103 : _GEN_390; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_392 = 8'h68 == _T_5[7:0] ? image_2_104 : _GEN_391; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_393 = 8'h69 == _T_5[7:0] ? image_2_105 : _GEN_392; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_394 = 8'h6a == _T_5[7:0] ? image_2_106 : _GEN_393; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_395 = 8'h6b == _T_5[7:0] ? image_2_107 : _GEN_394; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_396 = 8'h6c == _T_5[7:0] ? image_2_108 : _GEN_395; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_397 = 8'h6d == _T_5[7:0] ? image_2_109 : _GEN_396; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_398 = 8'h6e == _T_5[7:0] ? image_2_110 : _GEN_397; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_399 = 8'h6f == _T_5[7:0] ? image_2_111 : _GEN_398; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_400 = 8'h70 == _T_5[7:0] ? image_2_112 : _GEN_399; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_401 = 8'h71 == _T_5[7:0] ? image_2_113 : _GEN_400; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_402 = 8'h72 == _T_5[7:0] ? image_2_114 : _GEN_401; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_403 = 8'h73 == _T_5[7:0] ? image_2_115 : _GEN_402; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_404 = 8'h74 == _T_5[7:0] ? image_2_116 : _GEN_403; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_405 = 8'h75 == _T_5[7:0] ? image_2_117 : _GEN_404; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_406 = 8'h76 == _T_5[7:0] ? image_2_118 : _GEN_405; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_407 = 8'h77 == _T_5[7:0] ? image_2_119 : _GEN_406; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_408 = 8'h78 == _T_5[7:0] ? image_2_120 : _GEN_407; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_409 = 8'h79 == _T_5[7:0] ? image_2_121 : _GEN_408; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_410 = 8'h7a == _T_5[7:0] ? image_2_122 : _GEN_409; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_411 = 8'h7b == _T_5[7:0] ? image_2_123 : _GEN_410; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_412 = 8'h7c == _T_5[7:0] ? image_2_124 : _GEN_411; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_413 = 8'h7d == _T_5[7:0] ? image_2_125 : _GEN_412; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_414 = 8'h7e == _T_5[7:0] ? image_2_126 : _GEN_413; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_415 = 8'h7f == _T_5[7:0] ? image_2_127 : _GEN_414; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_416 = 8'h80 == _T_5[7:0] ? image_2_128 : _GEN_415; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_417 = 8'h81 == _T_5[7:0] ? image_2_129 : _GEN_416; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_418 = 8'h82 == _T_5[7:0] ? image_2_130 : _GEN_417; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_419 = 8'h83 == _T_5[7:0] ? image_2_131 : _GEN_418; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_420 = 8'h84 == _T_5[7:0] ? image_2_132 : _GEN_419; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_421 = 8'h85 == _T_5[7:0] ? image_2_133 : _GEN_420; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_422 = 8'h86 == _T_5[7:0] ? image_2_134 : _GEN_421; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_423 = 8'h87 == _T_5[7:0] ? image_2_135 : _GEN_422; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_424 = 8'h88 == _T_5[7:0] ? image_2_136 : _GEN_423; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_425 = 8'h89 == _T_5[7:0] ? image_2_137 : _GEN_424; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_426 = 8'h8a == _T_5[7:0] ? image_2_138 : _GEN_425; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_427 = 8'h8b == _T_5[7:0] ? image_2_139 : _GEN_426; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_428 = 8'h8c == _T_5[7:0] ? image_2_140 : _GEN_427; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_429 = 8'h8d == _T_5[7:0] ? image_2_141 : _GEN_428; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_430 = 8'h8e == _T_5[7:0] ? image_2_142 : _GEN_429; // @[VideoBuffer.scala 27:30]
  wire [32:0] _T_15 = {{1'd0}, pixelIndex}; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_19 = pixelIndex + 32'h1; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_22 = pixelIndex + 32'h2; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_25 = pixelIndex + 32'h3; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_28 = pixelIndex + 32'h4; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_31 = pixelIndex + 32'h5; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_34 = pixelIndex + 32'h6; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_37 = pixelIndex + 32'h7; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_88 = pixelIndex + 32'h8; // @[VideoBuffer.scala 36:34]
  wire [8:0] _T_89 = 5'h10 * 5'h9; // @[VideoBuffer.scala 37:42]
  wire [31:0] _GEN_4325 = {{23'd0}, _T_89}; // @[VideoBuffer.scala 37:25]
  wire  _T_90 = pixelIndex == _GEN_4325; // @[VideoBuffer.scala 37:25]
  assign io_pixelVal_out_0 = 8'h8f == _T_5[7:0] ? image_0_143 : _GEN_142; // @[VideoBuffer.scala 27:30]
  assign io_pixelVal_out_1 = 8'h8f == _T_5[7:0] ? image_1_143 : _GEN_286; // @[VideoBuffer.scala 27:30]
  assign io_pixelVal_out_2 = 8'h8f == _T_5[7:0] ? image_2_143 : _GEN_430; // @[VideoBuffer.scala 27:30]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  image_0_0 = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  image_0_1 = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  image_0_2 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  image_0_3 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  image_0_4 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  image_0_5 = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  image_0_6 = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  image_0_7 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  image_0_8 = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  image_0_9 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  image_0_10 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  image_0_11 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  image_0_12 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  image_0_13 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  image_0_14 = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  image_0_15 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  image_0_16 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  image_0_17 = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  image_0_18 = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  image_0_19 = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  image_0_20 = _RAND_20[3:0];
  _RAND_21 = {1{`RANDOM}};
  image_0_21 = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  image_0_22 = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  image_0_23 = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  image_0_24 = _RAND_24[3:0];
  _RAND_25 = {1{`RANDOM}};
  image_0_25 = _RAND_25[3:0];
  _RAND_26 = {1{`RANDOM}};
  image_0_26 = _RAND_26[3:0];
  _RAND_27 = {1{`RANDOM}};
  image_0_27 = _RAND_27[3:0];
  _RAND_28 = {1{`RANDOM}};
  image_0_28 = _RAND_28[3:0];
  _RAND_29 = {1{`RANDOM}};
  image_0_29 = _RAND_29[3:0];
  _RAND_30 = {1{`RANDOM}};
  image_0_30 = _RAND_30[3:0];
  _RAND_31 = {1{`RANDOM}};
  image_0_31 = _RAND_31[3:0];
  _RAND_32 = {1{`RANDOM}};
  image_0_32 = _RAND_32[3:0];
  _RAND_33 = {1{`RANDOM}};
  image_0_33 = _RAND_33[3:0];
  _RAND_34 = {1{`RANDOM}};
  image_0_34 = _RAND_34[3:0];
  _RAND_35 = {1{`RANDOM}};
  image_0_35 = _RAND_35[3:0];
  _RAND_36 = {1{`RANDOM}};
  image_0_36 = _RAND_36[3:0];
  _RAND_37 = {1{`RANDOM}};
  image_0_37 = _RAND_37[3:0];
  _RAND_38 = {1{`RANDOM}};
  image_0_38 = _RAND_38[3:0];
  _RAND_39 = {1{`RANDOM}};
  image_0_39 = _RAND_39[3:0];
  _RAND_40 = {1{`RANDOM}};
  image_0_40 = _RAND_40[3:0];
  _RAND_41 = {1{`RANDOM}};
  image_0_41 = _RAND_41[3:0];
  _RAND_42 = {1{`RANDOM}};
  image_0_42 = _RAND_42[3:0];
  _RAND_43 = {1{`RANDOM}};
  image_0_43 = _RAND_43[3:0];
  _RAND_44 = {1{`RANDOM}};
  image_0_44 = _RAND_44[3:0];
  _RAND_45 = {1{`RANDOM}};
  image_0_45 = _RAND_45[3:0];
  _RAND_46 = {1{`RANDOM}};
  image_0_46 = _RAND_46[3:0];
  _RAND_47 = {1{`RANDOM}};
  image_0_47 = _RAND_47[3:0];
  _RAND_48 = {1{`RANDOM}};
  image_0_48 = _RAND_48[3:0];
  _RAND_49 = {1{`RANDOM}};
  image_0_49 = _RAND_49[3:0];
  _RAND_50 = {1{`RANDOM}};
  image_0_50 = _RAND_50[3:0];
  _RAND_51 = {1{`RANDOM}};
  image_0_51 = _RAND_51[3:0];
  _RAND_52 = {1{`RANDOM}};
  image_0_52 = _RAND_52[3:0];
  _RAND_53 = {1{`RANDOM}};
  image_0_53 = _RAND_53[3:0];
  _RAND_54 = {1{`RANDOM}};
  image_0_54 = _RAND_54[3:0];
  _RAND_55 = {1{`RANDOM}};
  image_0_55 = _RAND_55[3:0];
  _RAND_56 = {1{`RANDOM}};
  image_0_56 = _RAND_56[3:0];
  _RAND_57 = {1{`RANDOM}};
  image_0_57 = _RAND_57[3:0];
  _RAND_58 = {1{`RANDOM}};
  image_0_58 = _RAND_58[3:0];
  _RAND_59 = {1{`RANDOM}};
  image_0_59 = _RAND_59[3:0];
  _RAND_60 = {1{`RANDOM}};
  image_0_60 = _RAND_60[3:0];
  _RAND_61 = {1{`RANDOM}};
  image_0_61 = _RAND_61[3:0];
  _RAND_62 = {1{`RANDOM}};
  image_0_62 = _RAND_62[3:0];
  _RAND_63 = {1{`RANDOM}};
  image_0_63 = _RAND_63[3:0];
  _RAND_64 = {1{`RANDOM}};
  image_0_64 = _RAND_64[3:0];
  _RAND_65 = {1{`RANDOM}};
  image_0_65 = _RAND_65[3:0];
  _RAND_66 = {1{`RANDOM}};
  image_0_66 = _RAND_66[3:0];
  _RAND_67 = {1{`RANDOM}};
  image_0_67 = _RAND_67[3:0];
  _RAND_68 = {1{`RANDOM}};
  image_0_68 = _RAND_68[3:0];
  _RAND_69 = {1{`RANDOM}};
  image_0_69 = _RAND_69[3:0];
  _RAND_70 = {1{`RANDOM}};
  image_0_70 = _RAND_70[3:0];
  _RAND_71 = {1{`RANDOM}};
  image_0_71 = _RAND_71[3:0];
  _RAND_72 = {1{`RANDOM}};
  image_0_72 = _RAND_72[3:0];
  _RAND_73 = {1{`RANDOM}};
  image_0_73 = _RAND_73[3:0];
  _RAND_74 = {1{`RANDOM}};
  image_0_74 = _RAND_74[3:0];
  _RAND_75 = {1{`RANDOM}};
  image_0_75 = _RAND_75[3:0];
  _RAND_76 = {1{`RANDOM}};
  image_0_76 = _RAND_76[3:0];
  _RAND_77 = {1{`RANDOM}};
  image_0_77 = _RAND_77[3:0];
  _RAND_78 = {1{`RANDOM}};
  image_0_78 = _RAND_78[3:0];
  _RAND_79 = {1{`RANDOM}};
  image_0_79 = _RAND_79[3:0];
  _RAND_80 = {1{`RANDOM}};
  image_0_80 = _RAND_80[3:0];
  _RAND_81 = {1{`RANDOM}};
  image_0_81 = _RAND_81[3:0];
  _RAND_82 = {1{`RANDOM}};
  image_0_82 = _RAND_82[3:0];
  _RAND_83 = {1{`RANDOM}};
  image_0_83 = _RAND_83[3:0];
  _RAND_84 = {1{`RANDOM}};
  image_0_84 = _RAND_84[3:0];
  _RAND_85 = {1{`RANDOM}};
  image_0_85 = _RAND_85[3:0];
  _RAND_86 = {1{`RANDOM}};
  image_0_86 = _RAND_86[3:0];
  _RAND_87 = {1{`RANDOM}};
  image_0_87 = _RAND_87[3:0];
  _RAND_88 = {1{`RANDOM}};
  image_0_88 = _RAND_88[3:0];
  _RAND_89 = {1{`RANDOM}};
  image_0_89 = _RAND_89[3:0];
  _RAND_90 = {1{`RANDOM}};
  image_0_90 = _RAND_90[3:0];
  _RAND_91 = {1{`RANDOM}};
  image_0_91 = _RAND_91[3:0];
  _RAND_92 = {1{`RANDOM}};
  image_0_92 = _RAND_92[3:0];
  _RAND_93 = {1{`RANDOM}};
  image_0_93 = _RAND_93[3:0];
  _RAND_94 = {1{`RANDOM}};
  image_0_94 = _RAND_94[3:0];
  _RAND_95 = {1{`RANDOM}};
  image_0_95 = _RAND_95[3:0];
  _RAND_96 = {1{`RANDOM}};
  image_0_96 = _RAND_96[3:0];
  _RAND_97 = {1{`RANDOM}};
  image_0_97 = _RAND_97[3:0];
  _RAND_98 = {1{`RANDOM}};
  image_0_98 = _RAND_98[3:0];
  _RAND_99 = {1{`RANDOM}};
  image_0_99 = _RAND_99[3:0];
  _RAND_100 = {1{`RANDOM}};
  image_0_100 = _RAND_100[3:0];
  _RAND_101 = {1{`RANDOM}};
  image_0_101 = _RAND_101[3:0];
  _RAND_102 = {1{`RANDOM}};
  image_0_102 = _RAND_102[3:0];
  _RAND_103 = {1{`RANDOM}};
  image_0_103 = _RAND_103[3:0];
  _RAND_104 = {1{`RANDOM}};
  image_0_104 = _RAND_104[3:0];
  _RAND_105 = {1{`RANDOM}};
  image_0_105 = _RAND_105[3:0];
  _RAND_106 = {1{`RANDOM}};
  image_0_106 = _RAND_106[3:0];
  _RAND_107 = {1{`RANDOM}};
  image_0_107 = _RAND_107[3:0];
  _RAND_108 = {1{`RANDOM}};
  image_0_108 = _RAND_108[3:0];
  _RAND_109 = {1{`RANDOM}};
  image_0_109 = _RAND_109[3:0];
  _RAND_110 = {1{`RANDOM}};
  image_0_110 = _RAND_110[3:0];
  _RAND_111 = {1{`RANDOM}};
  image_0_111 = _RAND_111[3:0];
  _RAND_112 = {1{`RANDOM}};
  image_0_112 = _RAND_112[3:0];
  _RAND_113 = {1{`RANDOM}};
  image_0_113 = _RAND_113[3:0];
  _RAND_114 = {1{`RANDOM}};
  image_0_114 = _RAND_114[3:0];
  _RAND_115 = {1{`RANDOM}};
  image_0_115 = _RAND_115[3:0];
  _RAND_116 = {1{`RANDOM}};
  image_0_116 = _RAND_116[3:0];
  _RAND_117 = {1{`RANDOM}};
  image_0_117 = _RAND_117[3:0];
  _RAND_118 = {1{`RANDOM}};
  image_0_118 = _RAND_118[3:0];
  _RAND_119 = {1{`RANDOM}};
  image_0_119 = _RAND_119[3:0];
  _RAND_120 = {1{`RANDOM}};
  image_0_120 = _RAND_120[3:0];
  _RAND_121 = {1{`RANDOM}};
  image_0_121 = _RAND_121[3:0];
  _RAND_122 = {1{`RANDOM}};
  image_0_122 = _RAND_122[3:0];
  _RAND_123 = {1{`RANDOM}};
  image_0_123 = _RAND_123[3:0];
  _RAND_124 = {1{`RANDOM}};
  image_0_124 = _RAND_124[3:0];
  _RAND_125 = {1{`RANDOM}};
  image_0_125 = _RAND_125[3:0];
  _RAND_126 = {1{`RANDOM}};
  image_0_126 = _RAND_126[3:0];
  _RAND_127 = {1{`RANDOM}};
  image_0_127 = _RAND_127[3:0];
  _RAND_128 = {1{`RANDOM}};
  image_0_128 = _RAND_128[3:0];
  _RAND_129 = {1{`RANDOM}};
  image_0_129 = _RAND_129[3:0];
  _RAND_130 = {1{`RANDOM}};
  image_0_130 = _RAND_130[3:0];
  _RAND_131 = {1{`RANDOM}};
  image_0_131 = _RAND_131[3:0];
  _RAND_132 = {1{`RANDOM}};
  image_0_132 = _RAND_132[3:0];
  _RAND_133 = {1{`RANDOM}};
  image_0_133 = _RAND_133[3:0];
  _RAND_134 = {1{`RANDOM}};
  image_0_134 = _RAND_134[3:0];
  _RAND_135 = {1{`RANDOM}};
  image_0_135 = _RAND_135[3:0];
  _RAND_136 = {1{`RANDOM}};
  image_0_136 = _RAND_136[3:0];
  _RAND_137 = {1{`RANDOM}};
  image_0_137 = _RAND_137[3:0];
  _RAND_138 = {1{`RANDOM}};
  image_0_138 = _RAND_138[3:0];
  _RAND_139 = {1{`RANDOM}};
  image_0_139 = _RAND_139[3:0];
  _RAND_140 = {1{`RANDOM}};
  image_0_140 = _RAND_140[3:0];
  _RAND_141 = {1{`RANDOM}};
  image_0_141 = _RAND_141[3:0];
  _RAND_142 = {1{`RANDOM}};
  image_0_142 = _RAND_142[3:0];
  _RAND_143 = {1{`RANDOM}};
  image_0_143 = _RAND_143[3:0];
  _RAND_144 = {1{`RANDOM}};
  image_1_0 = _RAND_144[3:0];
  _RAND_145 = {1{`RANDOM}};
  image_1_1 = _RAND_145[3:0];
  _RAND_146 = {1{`RANDOM}};
  image_1_2 = _RAND_146[3:0];
  _RAND_147 = {1{`RANDOM}};
  image_1_3 = _RAND_147[3:0];
  _RAND_148 = {1{`RANDOM}};
  image_1_4 = _RAND_148[3:0];
  _RAND_149 = {1{`RANDOM}};
  image_1_5 = _RAND_149[3:0];
  _RAND_150 = {1{`RANDOM}};
  image_1_6 = _RAND_150[3:0];
  _RAND_151 = {1{`RANDOM}};
  image_1_7 = _RAND_151[3:0];
  _RAND_152 = {1{`RANDOM}};
  image_1_8 = _RAND_152[3:0];
  _RAND_153 = {1{`RANDOM}};
  image_1_9 = _RAND_153[3:0];
  _RAND_154 = {1{`RANDOM}};
  image_1_10 = _RAND_154[3:0];
  _RAND_155 = {1{`RANDOM}};
  image_1_11 = _RAND_155[3:0];
  _RAND_156 = {1{`RANDOM}};
  image_1_12 = _RAND_156[3:0];
  _RAND_157 = {1{`RANDOM}};
  image_1_13 = _RAND_157[3:0];
  _RAND_158 = {1{`RANDOM}};
  image_1_14 = _RAND_158[3:0];
  _RAND_159 = {1{`RANDOM}};
  image_1_15 = _RAND_159[3:0];
  _RAND_160 = {1{`RANDOM}};
  image_1_16 = _RAND_160[3:0];
  _RAND_161 = {1{`RANDOM}};
  image_1_17 = _RAND_161[3:0];
  _RAND_162 = {1{`RANDOM}};
  image_1_18 = _RAND_162[3:0];
  _RAND_163 = {1{`RANDOM}};
  image_1_19 = _RAND_163[3:0];
  _RAND_164 = {1{`RANDOM}};
  image_1_20 = _RAND_164[3:0];
  _RAND_165 = {1{`RANDOM}};
  image_1_21 = _RAND_165[3:0];
  _RAND_166 = {1{`RANDOM}};
  image_1_22 = _RAND_166[3:0];
  _RAND_167 = {1{`RANDOM}};
  image_1_23 = _RAND_167[3:0];
  _RAND_168 = {1{`RANDOM}};
  image_1_24 = _RAND_168[3:0];
  _RAND_169 = {1{`RANDOM}};
  image_1_25 = _RAND_169[3:0];
  _RAND_170 = {1{`RANDOM}};
  image_1_26 = _RAND_170[3:0];
  _RAND_171 = {1{`RANDOM}};
  image_1_27 = _RAND_171[3:0];
  _RAND_172 = {1{`RANDOM}};
  image_1_28 = _RAND_172[3:0];
  _RAND_173 = {1{`RANDOM}};
  image_1_29 = _RAND_173[3:0];
  _RAND_174 = {1{`RANDOM}};
  image_1_30 = _RAND_174[3:0];
  _RAND_175 = {1{`RANDOM}};
  image_1_31 = _RAND_175[3:0];
  _RAND_176 = {1{`RANDOM}};
  image_1_32 = _RAND_176[3:0];
  _RAND_177 = {1{`RANDOM}};
  image_1_33 = _RAND_177[3:0];
  _RAND_178 = {1{`RANDOM}};
  image_1_34 = _RAND_178[3:0];
  _RAND_179 = {1{`RANDOM}};
  image_1_35 = _RAND_179[3:0];
  _RAND_180 = {1{`RANDOM}};
  image_1_36 = _RAND_180[3:0];
  _RAND_181 = {1{`RANDOM}};
  image_1_37 = _RAND_181[3:0];
  _RAND_182 = {1{`RANDOM}};
  image_1_38 = _RAND_182[3:0];
  _RAND_183 = {1{`RANDOM}};
  image_1_39 = _RAND_183[3:0];
  _RAND_184 = {1{`RANDOM}};
  image_1_40 = _RAND_184[3:0];
  _RAND_185 = {1{`RANDOM}};
  image_1_41 = _RAND_185[3:0];
  _RAND_186 = {1{`RANDOM}};
  image_1_42 = _RAND_186[3:0];
  _RAND_187 = {1{`RANDOM}};
  image_1_43 = _RAND_187[3:0];
  _RAND_188 = {1{`RANDOM}};
  image_1_44 = _RAND_188[3:0];
  _RAND_189 = {1{`RANDOM}};
  image_1_45 = _RAND_189[3:0];
  _RAND_190 = {1{`RANDOM}};
  image_1_46 = _RAND_190[3:0];
  _RAND_191 = {1{`RANDOM}};
  image_1_47 = _RAND_191[3:0];
  _RAND_192 = {1{`RANDOM}};
  image_1_48 = _RAND_192[3:0];
  _RAND_193 = {1{`RANDOM}};
  image_1_49 = _RAND_193[3:0];
  _RAND_194 = {1{`RANDOM}};
  image_1_50 = _RAND_194[3:0];
  _RAND_195 = {1{`RANDOM}};
  image_1_51 = _RAND_195[3:0];
  _RAND_196 = {1{`RANDOM}};
  image_1_52 = _RAND_196[3:0];
  _RAND_197 = {1{`RANDOM}};
  image_1_53 = _RAND_197[3:0];
  _RAND_198 = {1{`RANDOM}};
  image_1_54 = _RAND_198[3:0];
  _RAND_199 = {1{`RANDOM}};
  image_1_55 = _RAND_199[3:0];
  _RAND_200 = {1{`RANDOM}};
  image_1_56 = _RAND_200[3:0];
  _RAND_201 = {1{`RANDOM}};
  image_1_57 = _RAND_201[3:0];
  _RAND_202 = {1{`RANDOM}};
  image_1_58 = _RAND_202[3:0];
  _RAND_203 = {1{`RANDOM}};
  image_1_59 = _RAND_203[3:0];
  _RAND_204 = {1{`RANDOM}};
  image_1_60 = _RAND_204[3:0];
  _RAND_205 = {1{`RANDOM}};
  image_1_61 = _RAND_205[3:0];
  _RAND_206 = {1{`RANDOM}};
  image_1_62 = _RAND_206[3:0];
  _RAND_207 = {1{`RANDOM}};
  image_1_63 = _RAND_207[3:0];
  _RAND_208 = {1{`RANDOM}};
  image_1_64 = _RAND_208[3:0];
  _RAND_209 = {1{`RANDOM}};
  image_1_65 = _RAND_209[3:0];
  _RAND_210 = {1{`RANDOM}};
  image_1_66 = _RAND_210[3:0];
  _RAND_211 = {1{`RANDOM}};
  image_1_67 = _RAND_211[3:0];
  _RAND_212 = {1{`RANDOM}};
  image_1_68 = _RAND_212[3:0];
  _RAND_213 = {1{`RANDOM}};
  image_1_69 = _RAND_213[3:0];
  _RAND_214 = {1{`RANDOM}};
  image_1_70 = _RAND_214[3:0];
  _RAND_215 = {1{`RANDOM}};
  image_1_71 = _RAND_215[3:0];
  _RAND_216 = {1{`RANDOM}};
  image_1_72 = _RAND_216[3:0];
  _RAND_217 = {1{`RANDOM}};
  image_1_73 = _RAND_217[3:0];
  _RAND_218 = {1{`RANDOM}};
  image_1_74 = _RAND_218[3:0];
  _RAND_219 = {1{`RANDOM}};
  image_1_75 = _RAND_219[3:0];
  _RAND_220 = {1{`RANDOM}};
  image_1_76 = _RAND_220[3:0];
  _RAND_221 = {1{`RANDOM}};
  image_1_77 = _RAND_221[3:0];
  _RAND_222 = {1{`RANDOM}};
  image_1_78 = _RAND_222[3:0];
  _RAND_223 = {1{`RANDOM}};
  image_1_79 = _RAND_223[3:0];
  _RAND_224 = {1{`RANDOM}};
  image_1_80 = _RAND_224[3:0];
  _RAND_225 = {1{`RANDOM}};
  image_1_81 = _RAND_225[3:0];
  _RAND_226 = {1{`RANDOM}};
  image_1_82 = _RAND_226[3:0];
  _RAND_227 = {1{`RANDOM}};
  image_1_83 = _RAND_227[3:0];
  _RAND_228 = {1{`RANDOM}};
  image_1_84 = _RAND_228[3:0];
  _RAND_229 = {1{`RANDOM}};
  image_1_85 = _RAND_229[3:0];
  _RAND_230 = {1{`RANDOM}};
  image_1_86 = _RAND_230[3:0];
  _RAND_231 = {1{`RANDOM}};
  image_1_87 = _RAND_231[3:0];
  _RAND_232 = {1{`RANDOM}};
  image_1_88 = _RAND_232[3:0];
  _RAND_233 = {1{`RANDOM}};
  image_1_89 = _RAND_233[3:0];
  _RAND_234 = {1{`RANDOM}};
  image_1_90 = _RAND_234[3:0];
  _RAND_235 = {1{`RANDOM}};
  image_1_91 = _RAND_235[3:0];
  _RAND_236 = {1{`RANDOM}};
  image_1_92 = _RAND_236[3:0];
  _RAND_237 = {1{`RANDOM}};
  image_1_93 = _RAND_237[3:0];
  _RAND_238 = {1{`RANDOM}};
  image_1_94 = _RAND_238[3:0];
  _RAND_239 = {1{`RANDOM}};
  image_1_95 = _RAND_239[3:0];
  _RAND_240 = {1{`RANDOM}};
  image_1_96 = _RAND_240[3:0];
  _RAND_241 = {1{`RANDOM}};
  image_1_97 = _RAND_241[3:0];
  _RAND_242 = {1{`RANDOM}};
  image_1_98 = _RAND_242[3:0];
  _RAND_243 = {1{`RANDOM}};
  image_1_99 = _RAND_243[3:0];
  _RAND_244 = {1{`RANDOM}};
  image_1_100 = _RAND_244[3:0];
  _RAND_245 = {1{`RANDOM}};
  image_1_101 = _RAND_245[3:0];
  _RAND_246 = {1{`RANDOM}};
  image_1_102 = _RAND_246[3:0];
  _RAND_247 = {1{`RANDOM}};
  image_1_103 = _RAND_247[3:0];
  _RAND_248 = {1{`RANDOM}};
  image_1_104 = _RAND_248[3:0];
  _RAND_249 = {1{`RANDOM}};
  image_1_105 = _RAND_249[3:0];
  _RAND_250 = {1{`RANDOM}};
  image_1_106 = _RAND_250[3:0];
  _RAND_251 = {1{`RANDOM}};
  image_1_107 = _RAND_251[3:0];
  _RAND_252 = {1{`RANDOM}};
  image_1_108 = _RAND_252[3:0];
  _RAND_253 = {1{`RANDOM}};
  image_1_109 = _RAND_253[3:0];
  _RAND_254 = {1{`RANDOM}};
  image_1_110 = _RAND_254[3:0];
  _RAND_255 = {1{`RANDOM}};
  image_1_111 = _RAND_255[3:0];
  _RAND_256 = {1{`RANDOM}};
  image_1_112 = _RAND_256[3:0];
  _RAND_257 = {1{`RANDOM}};
  image_1_113 = _RAND_257[3:0];
  _RAND_258 = {1{`RANDOM}};
  image_1_114 = _RAND_258[3:0];
  _RAND_259 = {1{`RANDOM}};
  image_1_115 = _RAND_259[3:0];
  _RAND_260 = {1{`RANDOM}};
  image_1_116 = _RAND_260[3:0];
  _RAND_261 = {1{`RANDOM}};
  image_1_117 = _RAND_261[3:0];
  _RAND_262 = {1{`RANDOM}};
  image_1_118 = _RAND_262[3:0];
  _RAND_263 = {1{`RANDOM}};
  image_1_119 = _RAND_263[3:0];
  _RAND_264 = {1{`RANDOM}};
  image_1_120 = _RAND_264[3:0];
  _RAND_265 = {1{`RANDOM}};
  image_1_121 = _RAND_265[3:0];
  _RAND_266 = {1{`RANDOM}};
  image_1_122 = _RAND_266[3:0];
  _RAND_267 = {1{`RANDOM}};
  image_1_123 = _RAND_267[3:0];
  _RAND_268 = {1{`RANDOM}};
  image_1_124 = _RAND_268[3:0];
  _RAND_269 = {1{`RANDOM}};
  image_1_125 = _RAND_269[3:0];
  _RAND_270 = {1{`RANDOM}};
  image_1_126 = _RAND_270[3:0];
  _RAND_271 = {1{`RANDOM}};
  image_1_127 = _RAND_271[3:0];
  _RAND_272 = {1{`RANDOM}};
  image_1_128 = _RAND_272[3:0];
  _RAND_273 = {1{`RANDOM}};
  image_1_129 = _RAND_273[3:0];
  _RAND_274 = {1{`RANDOM}};
  image_1_130 = _RAND_274[3:0];
  _RAND_275 = {1{`RANDOM}};
  image_1_131 = _RAND_275[3:0];
  _RAND_276 = {1{`RANDOM}};
  image_1_132 = _RAND_276[3:0];
  _RAND_277 = {1{`RANDOM}};
  image_1_133 = _RAND_277[3:0];
  _RAND_278 = {1{`RANDOM}};
  image_1_134 = _RAND_278[3:0];
  _RAND_279 = {1{`RANDOM}};
  image_1_135 = _RAND_279[3:0];
  _RAND_280 = {1{`RANDOM}};
  image_1_136 = _RAND_280[3:0];
  _RAND_281 = {1{`RANDOM}};
  image_1_137 = _RAND_281[3:0];
  _RAND_282 = {1{`RANDOM}};
  image_1_138 = _RAND_282[3:0];
  _RAND_283 = {1{`RANDOM}};
  image_1_139 = _RAND_283[3:0];
  _RAND_284 = {1{`RANDOM}};
  image_1_140 = _RAND_284[3:0];
  _RAND_285 = {1{`RANDOM}};
  image_1_141 = _RAND_285[3:0];
  _RAND_286 = {1{`RANDOM}};
  image_1_142 = _RAND_286[3:0];
  _RAND_287 = {1{`RANDOM}};
  image_1_143 = _RAND_287[3:0];
  _RAND_288 = {1{`RANDOM}};
  image_2_0 = _RAND_288[3:0];
  _RAND_289 = {1{`RANDOM}};
  image_2_1 = _RAND_289[3:0];
  _RAND_290 = {1{`RANDOM}};
  image_2_2 = _RAND_290[3:0];
  _RAND_291 = {1{`RANDOM}};
  image_2_3 = _RAND_291[3:0];
  _RAND_292 = {1{`RANDOM}};
  image_2_4 = _RAND_292[3:0];
  _RAND_293 = {1{`RANDOM}};
  image_2_5 = _RAND_293[3:0];
  _RAND_294 = {1{`RANDOM}};
  image_2_6 = _RAND_294[3:0];
  _RAND_295 = {1{`RANDOM}};
  image_2_7 = _RAND_295[3:0];
  _RAND_296 = {1{`RANDOM}};
  image_2_8 = _RAND_296[3:0];
  _RAND_297 = {1{`RANDOM}};
  image_2_9 = _RAND_297[3:0];
  _RAND_298 = {1{`RANDOM}};
  image_2_10 = _RAND_298[3:0];
  _RAND_299 = {1{`RANDOM}};
  image_2_11 = _RAND_299[3:0];
  _RAND_300 = {1{`RANDOM}};
  image_2_12 = _RAND_300[3:0];
  _RAND_301 = {1{`RANDOM}};
  image_2_13 = _RAND_301[3:0];
  _RAND_302 = {1{`RANDOM}};
  image_2_14 = _RAND_302[3:0];
  _RAND_303 = {1{`RANDOM}};
  image_2_15 = _RAND_303[3:0];
  _RAND_304 = {1{`RANDOM}};
  image_2_16 = _RAND_304[3:0];
  _RAND_305 = {1{`RANDOM}};
  image_2_17 = _RAND_305[3:0];
  _RAND_306 = {1{`RANDOM}};
  image_2_18 = _RAND_306[3:0];
  _RAND_307 = {1{`RANDOM}};
  image_2_19 = _RAND_307[3:0];
  _RAND_308 = {1{`RANDOM}};
  image_2_20 = _RAND_308[3:0];
  _RAND_309 = {1{`RANDOM}};
  image_2_21 = _RAND_309[3:0];
  _RAND_310 = {1{`RANDOM}};
  image_2_22 = _RAND_310[3:0];
  _RAND_311 = {1{`RANDOM}};
  image_2_23 = _RAND_311[3:0];
  _RAND_312 = {1{`RANDOM}};
  image_2_24 = _RAND_312[3:0];
  _RAND_313 = {1{`RANDOM}};
  image_2_25 = _RAND_313[3:0];
  _RAND_314 = {1{`RANDOM}};
  image_2_26 = _RAND_314[3:0];
  _RAND_315 = {1{`RANDOM}};
  image_2_27 = _RAND_315[3:0];
  _RAND_316 = {1{`RANDOM}};
  image_2_28 = _RAND_316[3:0];
  _RAND_317 = {1{`RANDOM}};
  image_2_29 = _RAND_317[3:0];
  _RAND_318 = {1{`RANDOM}};
  image_2_30 = _RAND_318[3:0];
  _RAND_319 = {1{`RANDOM}};
  image_2_31 = _RAND_319[3:0];
  _RAND_320 = {1{`RANDOM}};
  image_2_32 = _RAND_320[3:0];
  _RAND_321 = {1{`RANDOM}};
  image_2_33 = _RAND_321[3:0];
  _RAND_322 = {1{`RANDOM}};
  image_2_34 = _RAND_322[3:0];
  _RAND_323 = {1{`RANDOM}};
  image_2_35 = _RAND_323[3:0];
  _RAND_324 = {1{`RANDOM}};
  image_2_36 = _RAND_324[3:0];
  _RAND_325 = {1{`RANDOM}};
  image_2_37 = _RAND_325[3:0];
  _RAND_326 = {1{`RANDOM}};
  image_2_38 = _RAND_326[3:0];
  _RAND_327 = {1{`RANDOM}};
  image_2_39 = _RAND_327[3:0];
  _RAND_328 = {1{`RANDOM}};
  image_2_40 = _RAND_328[3:0];
  _RAND_329 = {1{`RANDOM}};
  image_2_41 = _RAND_329[3:0];
  _RAND_330 = {1{`RANDOM}};
  image_2_42 = _RAND_330[3:0];
  _RAND_331 = {1{`RANDOM}};
  image_2_43 = _RAND_331[3:0];
  _RAND_332 = {1{`RANDOM}};
  image_2_44 = _RAND_332[3:0];
  _RAND_333 = {1{`RANDOM}};
  image_2_45 = _RAND_333[3:0];
  _RAND_334 = {1{`RANDOM}};
  image_2_46 = _RAND_334[3:0];
  _RAND_335 = {1{`RANDOM}};
  image_2_47 = _RAND_335[3:0];
  _RAND_336 = {1{`RANDOM}};
  image_2_48 = _RAND_336[3:0];
  _RAND_337 = {1{`RANDOM}};
  image_2_49 = _RAND_337[3:0];
  _RAND_338 = {1{`RANDOM}};
  image_2_50 = _RAND_338[3:0];
  _RAND_339 = {1{`RANDOM}};
  image_2_51 = _RAND_339[3:0];
  _RAND_340 = {1{`RANDOM}};
  image_2_52 = _RAND_340[3:0];
  _RAND_341 = {1{`RANDOM}};
  image_2_53 = _RAND_341[3:0];
  _RAND_342 = {1{`RANDOM}};
  image_2_54 = _RAND_342[3:0];
  _RAND_343 = {1{`RANDOM}};
  image_2_55 = _RAND_343[3:0];
  _RAND_344 = {1{`RANDOM}};
  image_2_56 = _RAND_344[3:0];
  _RAND_345 = {1{`RANDOM}};
  image_2_57 = _RAND_345[3:0];
  _RAND_346 = {1{`RANDOM}};
  image_2_58 = _RAND_346[3:0];
  _RAND_347 = {1{`RANDOM}};
  image_2_59 = _RAND_347[3:0];
  _RAND_348 = {1{`RANDOM}};
  image_2_60 = _RAND_348[3:0];
  _RAND_349 = {1{`RANDOM}};
  image_2_61 = _RAND_349[3:0];
  _RAND_350 = {1{`RANDOM}};
  image_2_62 = _RAND_350[3:0];
  _RAND_351 = {1{`RANDOM}};
  image_2_63 = _RAND_351[3:0];
  _RAND_352 = {1{`RANDOM}};
  image_2_64 = _RAND_352[3:0];
  _RAND_353 = {1{`RANDOM}};
  image_2_65 = _RAND_353[3:0];
  _RAND_354 = {1{`RANDOM}};
  image_2_66 = _RAND_354[3:0];
  _RAND_355 = {1{`RANDOM}};
  image_2_67 = _RAND_355[3:0];
  _RAND_356 = {1{`RANDOM}};
  image_2_68 = _RAND_356[3:0];
  _RAND_357 = {1{`RANDOM}};
  image_2_69 = _RAND_357[3:0];
  _RAND_358 = {1{`RANDOM}};
  image_2_70 = _RAND_358[3:0];
  _RAND_359 = {1{`RANDOM}};
  image_2_71 = _RAND_359[3:0];
  _RAND_360 = {1{`RANDOM}};
  image_2_72 = _RAND_360[3:0];
  _RAND_361 = {1{`RANDOM}};
  image_2_73 = _RAND_361[3:0];
  _RAND_362 = {1{`RANDOM}};
  image_2_74 = _RAND_362[3:0];
  _RAND_363 = {1{`RANDOM}};
  image_2_75 = _RAND_363[3:0];
  _RAND_364 = {1{`RANDOM}};
  image_2_76 = _RAND_364[3:0];
  _RAND_365 = {1{`RANDOM}};
  image_2_77 = _RAND_365[3:0];
  _RAND_366 = {1{`RANDOM}};
  image_2_78 = _RAND_366[3:0];
  _RAND_367 = {1{`RANDOM}};
  image_2_79 = _RAND_367[3:0];
  _RAND_368 = {1{`RANDOM}};
  image_2_80 = _RAND_368[3:0];
  _RAND_369 = {1{`RANDOM}};
  image_2_81 = _RAND_369[3:0];
  _RAND_370 = {1{`RANDOM}};
  image_2_82 = _RAND_370[3:0];
  _RAND_371 = {1{`RANDOM}};
  image_2_83 = _RAND_371[3:0];
  _RAND_372 = {1{`RANDOM}};
  image_2_84 = _RAND_372[3:0];
  _RAND_373 = {1{`RANDOM}};
  image_2_85 = _RAND_373[3:0];
  _RAND_374 = {1{`RANDOM}};
  image_2_86 = _RAND_374[3:0];
  _RAND_375 = {1{`RANDOM}};
  image_2_87 = _RAND_375[3:0];
  _RAND_376 = {1{`RANDOM}};
  image_2_88 = _RAND_376[3:0];
  _RAND_377 = {1{`RANDOM}};
  image_2_89 = _RAND_377[3:0];
  _RAND_378 = {1{`RANDOM}};
  image_2_90 = _RAND_378[3:0];
  _RAND_379 = {1{`RANDOM}};
  image_2_91 = _RAND_379[3:0];
  _RAND_380 = {1{`RANDOM}};
  image_2_92 = _RAND_380[3:0];
  _RAND_381 = {1{`RANDOM}};
  image_2_93 = _RAND_381[3:0];
  _RAND_382 = {1{`RANDOM}};
  image_2_94 = _RAND_382[3:0];
  _RAND_383 = {1{`RANDOM}};
  image_2_95 = _RAND_383[3:0];
  _RAND_384 = {1{`RANDOM}};
  image_2_96 = _RAND_384[3:0];
  _RAND_385 = {1{`RANDOM}};
  image_2_97 = _RAND_385[3:0];
  _RAND_386 = {1{`RANDOM}};
  image_2_98 = _RAND_386[3:0];
  _RAND_387 = {1{`RANDOM}};
  image_2_99 = _RAND_387[3:0];
  _RAND_388 = {1{`RANDOM}};
  image_2_100 = _RAND_388[3:0];
  _RAND_389 = {1{`RANDOM}};
  image_2_101 = _RAND_389[3:0];
  _RAND_390 = {1{`RANDOM}};
  image_2_102 = _RAND_390[3:0];
  _RAND_391 = {1{`RANDOM}};
  image_2_103 = _RAND_391[3:0];
  _RAND_392 = {1{`RANDOM}};
  image_2_104 = _RAND_392[3:0];
  _RAND_393 = {1{`RANDOM}};
  image_2_105 = _RAND_393[3:0];
  _RAND_394 = {1{`RANDOM}};
  image_2_106 = _RAND_394[3:0];
  _RAND_395 = {1{`RANDOM}};
  image_2_107 = _RAND_395[3:0];
  _RAND_396 = {1{`RANDOM}};
  image_2_108 = _RAND_396[3:0];
  _RAND_397 = {1{`RANDOM}};
  image_2_109 = _RAND_397[3:0];
  _RAND_398 = {1{`RANDOM}};
  image_2_110 = _RAND_398[3:0];
  _RAND_399 = {1{`RANDOM}};
  image_2_111 = _RAND_399[3:0];
  _RAND_400 = {1{`RANDOM}};
  image_2_112 = _RAND_400[3:0];
  _RAND_401 = {1{`RANDOM}};
  image_2_113 = _RAND_401[3:0];
  _RAND_402 = {1{`RANDOM}};
  image_2_114 = _RAND_402[3:0];
  _RAND_403 = {1{`RANDOM}};
  image_2_115 = _RAND_403[3:0];
  _RAND_404 = {1{`RANDOM}};
  image_2_116 = _RAND_404[3:0];
  _RAND_405 = {1{`RANDOM}};
  image_2_117 = _RAND_405[3:0];
  _RAND_406 = {1{`RANDOM}};
  image_2_118 = _RAND_406[3:0];
  _RAND_407 = {1{`RANDOM}};
  image_2_119 = _RAND_407[3:0];
  _RAND_408 = {1{`RANDOM}};
  image_2_120 = _RAND_408[3:0];
  _RAND_409 = {1{`RANDOM}};
  image_2_121 = _RAND_409[3:0];
  _RAND_410 = {1{`RANDOM}};
  image_2_122 = _RAND_410[3:0];
  _RAND_411 = {1{`RANDOM}};
  image_2_123 = _RAND_411[3:0];
  _RAND_412 = {1{`RANDOM}};
  image_2_124 = _RAND_412[3:0];
  _RAND_413 = {1{`RANDOM}};
  image_2_125 = _RAND_413[3:0];
  _RAND_414 = {1{`RANDOM}};
  image_2_126 = _RAND_414[3:0];
  _RAND_415 = {1{`RANDOM}};
  image_2_127 = _RAND_415[3:0];
  _RAND_416 = {1{`RANDOM}};
  image_2_128 = _RAND_416[3:0];
  _RAND_417 = {1{`RANDOM}};
  image_2_129 = _RAND_417[3:0];
  _RAND_418 = {1{`RANDOM}};
  image_2_130 = _RAND_418[3:0];
  _RAND_419 = {1{`RANDOM}};
  image_2_131 = _RAND_419[3:0];
  _RAND_420 = {1{`RANDOM}};
  image_2_132 = _RAND_420[3:0];
  _RAND_421 = {1{`RANDOM}};
  image_2_133 = _RAND_421[3:0];
  _RAND_422 = {1{`RANDOM}};
  image_2_134 = _RAND_422[3:0];
  _RAND_423 = {1{`RANDOM}};
  image_2_135 = _RAND_423[3:0];
  _RAND_424 = {1{`RANDOM}};
  image_2_136 = _RAND_424[3:0];
  _RAND_425 = {1{`RANDOM}};
  image_2_137 = _RAND_425[3:0];
  _RAND_426 = {1{`RANDOM}};
  image_2_138 = _RAND_426[3:0];
  _RAND_427 = {1{`RANDOM}};
  image_2_139 = _RAND_427[3:0];
  _RAND_428 = {1{`RANDOM}};
  image_2_140 = _RAND_428[3:0];
  _RAND_429 = {1{`RANDOM}};
  image_2_141 = _RAND_429[3:0];
  _RAND_430 = {1{`RANDOM}};
  image_2_142 = _RAND_430[3:0];
  _RAND_431 = {1{`RANDOM}};
  image_2_143 = _RAND_431[3:0];
  _RAND_432 = {1{`RANDOM}};
  pixelIndex = _RAND_432[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      image_0_0 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h0 == _T_37[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_7;
      end else if (8'h0 == _T_34[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_6;
      end else if (8'h0 == _T_31[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_5;
      end else if (8'h0 == _T_28[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_4;
      end else if (8'h0 == _T_25[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_3;
      end else if (8'h0 == _T_22[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_2;
      end else if (8'h0 == _T_19[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_1;
      end else if (8'h0 == _T_15[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_1 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1 == _T_37[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_7;
      end else if (8'h1 == _T_34[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_6;
      end else if (8'h1 == _T_31[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_5;
      end else if (8'h1 == _T_28[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_4;
      end else if (8'h1 == _T_25[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_3;
      end else if (8'h1 == _T_22[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_2;
      end else if (8'h1 == _T_19[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_1;
      end else if (8'h1 == _T_15[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_2 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2 == _T_37[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_7;
      end else if (8'h2 == _T_34[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_6;
      end else if (8'h2 == _T_31[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_5;
      end else if (8'h2 == _T_28[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_4;
      end else if (8'h2 == _T_25[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_3;
      end else if (8'h2 == _T_22[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_2;
      end else if (8'h2 == _T_19[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_1;
      end else if (8'h2 == _T_15[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_3 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3 == _T_37[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_7;
      end else if (8'h3 == _T_34[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_6;
      end else if (8'h3 == _T_31[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_5;
      end else if (8'h3 == _T_28[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_4;
      end else if (8'h3 == _T_25[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_3;
      end else if (8'h3 == _T_22[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_2;
      end else if (8'h3 == _T_19[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_1;
      end else if (8'h3 == _T_15[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_4 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4 == _T_37[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_7;
      end else if (8'h4 == _T_34[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_6;
      end else if (8'h4 == _T_31[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_5;
      end else if (8'h4 == _T_28[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_4;
      end else if (8'h4 == _T_25[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_3;
      end else if (8'h4 == _T_22[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_2;
      end else if (8'h4 == _T_19[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_1;
      end else if (8'h4 == _T_15[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_5 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5 == _T_37[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_7;
      end else if (8'h5 == _T_34[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_6;
      end else if (8'h5 == _T_31[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_5;
      end else if (8'h5 == _T_28[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_4;
      end else if (8'h5 == _T_25[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_3;
      end else if (8'h5 == _T_22[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_2;
      end else if (8'h5 == _T_19[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_1;
      end else if (8'h5 == _T_15[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_6 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6 == _T_37[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_7;
      end else if (8'h6 == _T_34[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_6;
      end else if (8'h6 == _T_31[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_5;
      end else if (8'h6 == _T_28[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_4;
      end else if (8'h6 == _T_25[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_3;
      end else if (8'h6 == _T_22[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_2;
      end else if (8'h6 == _T_19[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_1;
      end else if (8'h6 == _T_15[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_7 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7 == _T_37[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_7;
      end else if (8'h7 == _T_34[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_6;
      end else if (8'h7 == _T_31[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_5;
      end else if (8'h7 == _T_28[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_4;
      end else if (8'h7 == _T_25[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_3;
      end else if (8'h7 == _T_22[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_2;
      end else if (8'h7 == _T_19[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_1;
      end else if (8'h7 == _T_15[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_8 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8 == _T_37[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_7;
      end else if (8'h8 == _T_34[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_6;
      end else if (8'h8 == _T_31[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_5;
      end else if (8'h8 == _T_28[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_4;
      end else if (8'h8 == _T_25[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_3;
      end else if (8'h8 == _T_22[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_2;
      end else if (8'h8 == _T_19[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_1;
      end else if (8'h8 == _T_15[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_9 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h9 == _T_37[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_7;
      end else if (8'h9 == _T_34[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_6;
      end else if (8'h9 == _T_31[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_5;
      end else if (8'h9 == _T_28[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_4;
      end else if (8'h9 == _T_25[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_3;
      end else if (8'h9 == _T_22[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_2;
      end else if (8'h9 == _T_19[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_1;
      end else if (8'h9 == _T_15[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_10 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha == _T_37[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_7;
      end else if (8'ha == _T_34[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_6;
      end else if (8'ha == _T_31[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_5;
      end else if (8'ha == _T_28[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_4;
      end else if (8'ha == _T_25[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_3;
      end else if (8'ha == _T_22[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_2;
      end else if (8'ha == _T_19[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_1;
      end else if (8'ha == _T_15[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_11 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb == _T_37[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_7;
      end else if (8'hb == _T_34[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_6;
      end else if (8'hb == _T_31[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_5;
      end else if (8'hb == _T_28[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_4;
      end else if (8'hb == _T_25[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_3;
      end else if (8'hb == _T_22[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_2;
      end else if (8'hb == _T_19[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_1;
      end else if (8'hb == _T_15[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_12 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hc == _T_37[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_7;
      end else if (8'hc == _T_34[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_6;
      end else if (8'hc == _T_31[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_5;
      end else if (8'hc == _T_28[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_4;
      end else if (8'hc == _T_25[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_3;
      end else if (8'hc == _T_22[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_2;
      end else if (8'hc == _T_19[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_1;
      end else if (8'hc == _T_15[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_13 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hd == _T_37[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_7;
      end else if (8'hd == _T_34[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_6;
      end else if (8'hd == _T_31[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_5;
      end else if (8'hd == _T_28[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_4;
      end else if (8'hd == _T_25[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_3;
      end else if (8'hd == _T_22[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_2;
      end else if (8'hd == _T_19[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_1;
      end else if (8'hd == _T_15[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_14 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'he == _T_37[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_7;
      end else if (8'he == _T_34[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_6;
      end else if (8'he == _T_31[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_5;
      end else if (8'he == _T_28[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_4;
      end else if (8'he == _T_25[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_3;
      end else if (8'he == _T_22[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_2;
      end else if (8'he == _T_19[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_1;
      end else if (8'he == _T_15[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_15 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hf == _T_37[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_7;
      end else if (8'hf == _T_34[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_6;
      end else if (8'hf == _T_31[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_5;
      end else if (8'hf == _T_28[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_4;
      end else if (8'hf == _T_25[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_3;
      end else if (8'hf == _T_22[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_2;
      end else if (8'hf == _T_19[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_1;
      end else if (8'hf == _T_15[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_16 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h10 == _T_37[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_7;
      end else if (8'h10 == _T_34[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_6;
      end else if (8'h10 == _T_31[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_5;
      end else if (8'h10 == _T_28[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_4;
      end else if (8'h10 == _T_25[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_3;
      end else if (8'h10 == _T_22[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_2;
      end else if (8'h10 == _T_19[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_1;
      end else if (8'h10 == _T_15[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_17 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h11 == _T_37[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_7;
      end else if (8'h11 == _T_34[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_6;
      end else if (8'h11 == _T_31[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_5;
      end else if (8'h11 == _T_28[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_4;
      end else if (8'h11 == _T_25[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_3;
      end else if (8'h11 == _T_22[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_2;
      end else if (8'h11 == _T_19[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_1;
      end else if (8'h11 == _T_15[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_18 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h12 == _T_37[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_7;
      end else if (8'h12 == _T_34[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_6;
      end else if (8'h12 == _T_31[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_5;
      end else if (8'h12 == _T_28[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_4;
      end else if (8'h12 == _T_25[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_3;
      end else if (8'h12 == _T_22[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_2;
      end else if (8'h12 == _T_19[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_1;
      end else if (8'h12 == _T_15[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_19 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h13 == _T_37[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_7;
      end else if (8'h13 == _T_34[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_6;
      end else if (8'h13 == _T_31[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_5;
      end else if (8'h13 == _T_28[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_4;
      end else if (8'h13 == _T_25[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_3;
      end else if (8'h13 == _T_22[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_2;
      end else if (8'h13 == _T_19[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_1;
      end else if (8'h13 == _T_15[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_20 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h14 == _T_37[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_7;
      end else if (8'h14 == _T_34[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_6;
      end else if (8'h14 == _T_31[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_5;
      end else if (8'h14 == _T_28[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_4;
      end else if (8'h14 == _T_25[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_3;
      end else if (8'h14 == _T_22[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_2;
      end else if (8'h14 == _T_19[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_1;
      end else if (8'h14 == _T_15[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_21 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h15 == _T_37[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_7;
      end else if (8'h15 == _T_34[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_6;
      end else if (8'h15 == _T_31[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_5;
      end else if (8'h15 == _T_28[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_4;
      end else if (8'h15 == _T_25[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_3;
      end else if (8'h15 == _T_22[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_2;
      end else if (8'h15 == _T_19[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_1;
      end else if (8'h15 == _T_15[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_22 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h16 == _T_37[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_7;
      end else if (8'h16 == _T_34[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_6;
      end else if (8'h16 == _T_31[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_5;
      end else if (8'h16 == _T_28[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_4;
      end else if (8'h16 == _T_25[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_3;
      end else if (8'h16 == _T_22[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_2;
      end else if (8'h16 == _T_19[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_1;
      end else if (8'h16 == _T_15[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_23 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h17 == _T_37[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_7;
      end else if (8'h17 == _T_34[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_6;
      end else if (8'h17 == _T_31[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_5;
      end else if (8'h17 == _T_28[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_4;
      end else if (8'h17 == _T_25[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_3;
      end else if (8'h17 == _T_22[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_2;
      end else if (8'h17 == _T_19[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_1;
      end else if (8'h17 == _T_15[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_24 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h18 == _T_37[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_7;
      end else if (8'h18 == _T_34[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_6;
      end else if (8'h18 == _T_31[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_5;
      end else if (8'h18 == _T_28[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_4;
      end else if (8'h18 == _T_25[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_3;
      end else if (8'h18 == _T_22[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_2;
      end else if (8'h18 == _T_19[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_1;
      end else if (8'h18 == _T_15[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_25 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h19 == _T_37[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_7;
      end else if (8'h19 == _T_34[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_6;
      end else if (8'h19 == _T_31[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_5;
      end else if (8'h19 == _T_28[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_4;
      end else if (8'h19 == _T_25[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_3;
      end else if (8'h19 == _T_22[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_2;
      end else if (8'h19 == _T_19[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_1;
      end else if (8'h19 == _T_15[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_26 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1a == _T_37[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_7;
      end else if (8'h1a == _T_34[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_6;
      end else if (8'h1a == _T_31[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_5;
      end else if (8'h1a == _T_28[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_4;
      end else if (8'h1a == _T_25[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_3;
      end else if (8'h1a == _T_22[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_2;
      end else if (8'h1a == _T_19[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_1;
      end else if (8'h1a == _T_15[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_27 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1b == _T_37[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_7;
      end else if (8'h1b == _T_34[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_6;
      end else if (8'h1b == _T_31[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_5;
      end else if (8'h1b == _T_28[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_4;
      end else if (8'h1b == _T_25[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_3;
      end else if (8'h1b == _T_22[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_2;
      end else if (8'h1b == _T_19[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_1;
      end else if (8'h1b == _T_15[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_28 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1c == _T_37[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_7;
      end else if (8'h1c == _T_34[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_6;
      end else if (8'h1c == _T_31[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_5;
      end else if (8'h1c == _T_28[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_4;
      end else if (8'h1c == _T_25[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_3;
      end else if (8'h1c == _T_22[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_2;
      end else if (8'h1c == _T_19[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_1;
      end else if (8'h1c == _T_15[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_29 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1d == _T_37[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_7;
      end else if (8'h1d == _T_34[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_6;
      end else if (8'h1d == _T_31[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_5;
      end else if (8'h1d == _T_28[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_4;
      end else if (8'h1d == _T_25[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_3;
      end else if (8'h1d == _T_22[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_2;
      end else if (8'h1d == _T_19[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_1;
      end else if (8'h1d == _T_15[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_30 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1e == _T_37[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_7;
      end else if (8'h1e == _T_34[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_6;
      end else if (8'h1e == _T_31[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_5;
      end else if (8'h1e == _T_28[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_4;
      end else if (8'h1e == _T_25[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_3;
      end else if (8'h1e == _T_22[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_2;
      end else if (8'h1e == _T_19[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_1;
      end else if (8'h1e == _T_15[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_31 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1f == _T_37[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_7;
      end else if (8'h1f == _T_34[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_6;
      end else if (8'h1f == _T_31[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_5;
      end else if (8'h1f == _T_28[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_4;
      end else if (8'h1f == _T_25[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_3;
      end else if (8'h1f == _T_22[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_2;
      end else if (8'h1f == _T_19[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_1;
      end else if (8'h1f == _T_15[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_32 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h20 == _T_37[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_7;
      end else if (8'h20 == _T_34[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_6;
      end else if (8'h20 == _T_31[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_5;
      end else if (8'h20 == _T_28[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_4;
      end else if (8'h20 == _T_25[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_3;
      end else if (8'h20 == _T_22[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_2;
      end else if (8'h20 == _T_19[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_1;
      end else if (8'h20 == _T_15[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_33 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h21 == _T_37[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_7;
      end else if (8'h21 == _T_34[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_6;
      end else if (8'h21 == _T_31[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_5;
      end else if (8'h21 == _T_28[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_4;
      end else if (8'h21 == _T_25[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_3;
      end else if (8'h21 == _T_22[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_2;
      end else if (8'h21 == _T_19[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_1;
      end else if (8'h21 == _T_15[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_34 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h22 == _T_37[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_7;
      end else if (8'h22 == _T_34[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_6;
      end else if (8'h22 == _T_31[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_5;
      end else if (8'h22 == _T_28[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_4;
      end else if (8'h22 == _T_25[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_3;
      end else if (8'h22 == _T_22[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_2;
      end else if (8'h22 == _T_19[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_1;
      end else if (8'h22 == _T_15[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_35 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h23 == _T_37[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_7;
      end else if (8'h23 == _T_34[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_6;
      end else if (8'h23 == _T_31[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_5;
      end else if (8'h23 == _T_28[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_4;
      end else if (8'h23 == _T_25[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_3;
      end else if (8'h23 == _T_22[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_2;
      end else if (8'h23 == _T_19[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_1;
      end else if (8'h23 == _T_15[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_36 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h24 == _T_37[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_7;
      end else if (8'h24 == _T_34[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_6;
      end else if (8'h24 == _T_31[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_5;
      end else if (8'h24 == _T_28[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_4;
      end else if (8'h24 == _T_25[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_3;
      end else if (8'h24 == _T_22[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_2;
      end else if (8'h24 == _T_19[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_1;
      end else if (8'h24 == _T_15[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_37 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h25 == _T_37[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_7;
      end else if (8'h25 == _T_34[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_6;
      end else if (8'h25 == _T_31[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_5;
      end else if (8'h25 == _T_28[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_4;
      end else if (8'h25 == _T_25[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_3;
      end else if (8'h25 == _T_22[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_2;
      end else if (8'h25 == _T_19[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_1;
      end else if (8'h25 == _T_15[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_38 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h26 == _T_37[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_7;
      end else if (8'h26 == _T_34[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_6;
      end else if (8'h26 == _T_31[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_5;
      end else if (8'h26 == _T_28[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_4;
      end else if (8'h26 == _T_25[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_3;
      end else if (8'h26 == _T_22[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_2;
      end else if (8'h26 == _T_19[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_1;
      end else if (8'h26 == _T_15[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_39 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h27 == _T_37[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_7;
      end else if (8'h27 == _T_34[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_6;
      end else if (8'h27 == _T_31[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_5;
      end else if (8'h27 == _T_28[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_4;
      end else if (8'h27 == _T_25[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_3;
      end else if (8'h27 == _T_22[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_2;
      end else if (8'h27 == _T_19[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_1;
      end else if (8'h27 == _T_15[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_40 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h28 == _T_37[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_7;
      end else if (8'h28 == _T_34[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_6;
      end else if (8'h28 == _T_31[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_5;
      end else if (8'h28 == _T_28[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_4;
      end else if (8'h28 == _T_25[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_3;
      end else if (8'h28 == _T_22[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_2;
      end else if (8'h28 == _T_19[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_1;
      end else if (8'h28 == _T_15[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_41 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h29 == _T_37[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_7;
      end else if (8'h29 == _T_34[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_6;
      end else if (8'h29 == _T_31[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_5;
      end else if (8'h29 == _T_28[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_4;
      end else if (8'h29 == _T_25[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_3;
      end else if (8'h29 == _T_22[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_2;
      end else if (8'h29 == _T_19[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_1;
      end else if (8'h29 == _T_15[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_42 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2a == _T_37[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_7;
      end else if (8'h2a == _T_34[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_6;
      end else if (8'h2a == _T_31[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_5;
      end else if (8'h2a == _T_28[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_4;
      end else if (8'h2a == _T_25[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_3;
      end else if (8'h2a == _T_22[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_2;
      end else if (8'h2a == _T_19[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_1;
      end else if (8'h2a == _T_15[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_43 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2b == _T_37[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_7;
      end else if (8'h2b == _T_34[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_6;
      end else if (8'h2b == _T_31[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_5;
      end else if (8'h2b == _T_28[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_4;
      end else if (8'h2b == _T_25[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_3;
      end else if (8'h2b == _T_22[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_2;
      end else if (8'h2b == _T_19[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_1;
      end else if (8'h2b == _T_15[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_44 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2c == _T_37[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_7;
      end else if (8'h2c == _T_34[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_6;
      end else if (8'h2c == _T_31[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_5;
      end else if (8'h2c == _T_28[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_4;
      end else if (8'h2c == _T_25[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_3;
      end else if (8'h2c == _T_22[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_2;
      end else if (8'h2c == _T_19[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_1;
      end else if (8'h2c == _T_15[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_45 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2d == _T_37[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_7;
      end else if (8'h2d == _T_34[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_6;
      end else if (8'h2d == _T_31[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_5;
      end else if (8'h2d == _T_28[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_4;
      end else if (8'h2d == _T_25[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_3;
      end else if (8'h2d == _T_22[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_2;
      end else if (8'h2d == _T_19[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_1;
      end else if (8'h2d == _T_15[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_46 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2e == _T_37[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_7;
      end else if (8'h2e == _T_34[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_6;
      end else if (8'h2e == _T_31[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_5;
      end else if (8'h2e == _T_28[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_4;
      end else if (8'h2e == _T_25[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_3;
      end else if (8'h2e == _T_22[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_2;
      end else if (8'h2e == _T_19[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_1;
      end else if (8'h2e == _T_15[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_47 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2f == _T_37[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_7;
      end else if (8'h2f == _T_34[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_6;
      end else if (8'h2f == _T_31[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_5;
      end else if (8'h2f == _T_28[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_4;
      end else if (8'h2f == _T_25[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_3;
      end else if (8'h2f == _T_22[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_2;
      end else if (8'h2f == _T_19[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_1;
      end else if (8'h2f == _T_15[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_48 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h30 == _T_37[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_7;
      end else if (8'h30 == _T_34[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_6;
      end else if (8'h30 == _T_31[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_5;
      end else if (8'h30 == _T_28[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_4;
      end else if (8'h30 == _T_25[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_3;
      end else if (8'h30 == _T_22[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_2;
      end else if (8'h30 == _T_19[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_1;
      end else if (8'h30 == _T_15[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_49 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h31 == _T_37[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_7;
      end else if (8'h31 == _T_34[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_6;
      end else if (8'h31 == _T_31[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_5;
      end else if (8'h31 == _T_28[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_4;
      end else if (8'h31 == _T_25[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_3;
      end else if (8'h31 == _T_22[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_2;
      end else if (8'h31 == _T_19[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_1;
      end else if (8'h31 == _T_15[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_50 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h32 == _T_37[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_7;
      end else if (8'h32 == _T_34[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_6;
      end else if (8'h32 == _T_31[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_5;
      end else if (8'h32 == _T_28[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_4;
      end else if (8'h32 == _T_25[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_3;
      end else if (8'h32 == _T_22[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_2;
      end else if (8'h32 == _T_19[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_1;
      end else if (8'h32 == _T_15[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_51 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h33 == _T_37[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_7;
      end else if (8'h33 == _T_34[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_6;
      end else if (8'h33 == _T_31[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_5;
      end else if (8'h33 == _T_28[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_4;
      end else if (8'h33 == _T_25[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_3;
      end else if (8'h33 == _T_22[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_2;
      end else if (8'h33 == _T_19[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_1;
      end else if (8'h33 == _T_15[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_52 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h34 == _T_37[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_7;
      end else if (8'h34 == _T_34[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_6;
      end else if (8'h34 == _T_31[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_5;
      end else if (8'h34 == _T_28[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_4;
      end else if (8'h34 == _T_25[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_3;
      end else if (8'h34 == _T_22[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_2;
      end else if (8'h34 == _T_19[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_1;
      end else if (8'h34 == _T_15[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_53 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h35 == _T_37[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_7;
      end else if (8'h35 == _T_34[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_6;
      end else if (8'h35 == _T_31[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_5;
      end else if (8'h35 == _T_28[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_4;
      end else if (8'h35 == _T_25[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_3;
      end else if (8'h35 == _T_22[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_2;
      end else if (8'h35 == _T_19[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_1;
      end else if (8'h35 == _T_15[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_54 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h36 == _T_37[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_7;
      end else if (8'h36 == _T_34[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_6;
      end else if (8'h36 == _T_31[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_5;
      end else if (8'h36 == _T_28[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_4;
      end else if (8'h36 == _T_25[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_3;
      end else if (8'h36 == _T_22[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_2;
      end else if (8'h36 == _T_19[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_1;
      end else if (8'h36 == _T_15[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_55 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h37 == _T_37[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_7;
      end else if (8'h37 == _T_34[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_6;
      end else if (8'h37 == _T_31[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_5;
      end else if (8'h37 == _T_28[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_4;
      end else if (8'h37 == _T_25[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_3;
      end else if (8'h37 == _T_22[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_2;
      end else if (8'h37 == _T_19[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_1;
      end else if (8'h37 == _T_15[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_56 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h38 == _T_37[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_7;
      end else if (8'h38 == _T_34[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_6;
      end else if (8'h38 == _T_31[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_5;
      end else if (8'h38 == _T_28[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_4;
      end else if (8'h38 == _T_25[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_3;
      end else if (8'h38 == _T_22[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_2;
      end else if (8'h38 == _T_19[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_1;
      end else if (8'h38 == _T_15[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_57 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h39 == _T_37[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_7;
      end else if (8'h39 == _T_34[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_6;
      end else if (8'h39 == _T_31[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_5;
      end else if (8'h39 == _T_28[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_4;
      end else if (8'h39 == _T_25[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_3;
      end else if (8'h39 == _T_22[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_2;
      end else if (8'h39 == _T_19[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_1;
      end else if (8'h39 == _T_15[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_58 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3a == _T_37[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_7;
      end else if (8'h3a == _T_34[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_6;
      end else if (8'h3a == _T_31[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_5;
      end else if (8'h3a == _T_28[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_4;
      end else if (8'h3a == _T_25[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_3;
      end else if (8'h3a == _T_22[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_2;
      end else if (8'h3a == _T_19[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_1;
      end else if (8'h3a == _T_15[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_59 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3b == _T_37[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_7;
      end else if (8'h3b == _T_34[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_6;
      end else if (8'h3b == _T_31[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_5;
      end else if (8'h3b == _T_28[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_4;
      end else if (8'h3b == _T_25[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_3;
      end else if (8'h3b == _T_22[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_2;
      end else if (8'h3b == _T_19[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_1;
      end else if (8'h3b == _T_15[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_60 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3c == _T_37[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_7;
      end else if (8'h3c == _T_34[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_6;
      end else if (8'h3c == _T_31[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_5;
      end else if (8'h3c == _T_28[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_4;
      end else if (8'h3c == _T_25[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_3;
      end else if (8'h3c == _T_22[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_2;
      end else if (8'h3c == _T_19[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_1;
      end else if (8'h3c == _T_15[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_61 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3d == _T_37[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_7;
      end else if (8'h3d == _T_34[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_6;
      end else if (8'h3d == _T_31[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_5;
      end else if (8'h3d == _T_28[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_4;
      end else if (8'h3d == _T_25[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_3;
      end else if (8'h3d == _T_22[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_2;
      end else if (8'h3d == _T_19[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_1;
      end else if (8'h3d == _T_15[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_62 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3e == _T_37[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_7;
      end else if (8'h3e == _T_34[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_6;
      end else if (8'h3e == _T_31[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_5;
      end else if (8'h3e == _T_28[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_4;
      end else if (8'h3e == _T_25[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_3;
      end else if (8'h3e == _T_22[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_2;
      end else if (8'h3e == _T_19[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_1;
      end else if (8'h3e == _T_15[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_63 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3f == _T_37[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_7;
      end else if (8'h3f == _T_34[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_6;
      end else if (8'h3f == _T_31[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_5;
      end else if (8'h3f == _T_28[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_4;
      end else if (8'h3f == _T_25[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_3;
      end else if (8'h3f == _T_22[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_2;
      end else if (8'h3f == _T_19[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_1;
      end else if (8'h3f == _T_15[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_64 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h40 == _T_37[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_7;
      end else if (8'h40 == _T_34[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_6;
      end else if (8'h40 == _T_31[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_5;
      end else if (8'h40 == _T_28[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_4;
      end else if (8'h40 == _T_25[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_3;
      end else if (8'h40 == _T_22[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_2;
      end else if (8'h40 == _T_19[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_1;
      end else if (8'h40 == _T_15[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_65 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h41 == _T_37[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_7;
      end else if (8'h41 == _T_34[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_6;
      end else if (8'h41 == _T_31[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_5;
      end else if (8'h41 == _T_28[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_4;
      end else if (8'h41 == _T_25[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_3;
      end else if (8'h41 == _T_22[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_2;
      end else if (8'h41 == _T_19[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_1;
      end else if (8'h41 == _T_15[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_66 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h42 == _T_37[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_7;
      end else if (8'h42 == _T_34[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_6;
      end else if (8'h42 == _T_31[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_5;
      end else if (8'h42 == _T_28[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_4;
      end else if (8'h42 == _T_25[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_3;
      end else if (8'h42 == _T_22[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_2;
      end else if (8'h42 == _T_19[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_1;
      end else if (8'h42 == _T_15[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_67 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h43 == _T_37[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_7;
      end else if (8'h43 == _T_34[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_6;
      end else if (8'h43 == _T_31[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_5;
      end else if (8'h43 == _T_28[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_4;
      end else if (8'h43 == _T_25[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_3;
      end else if (8'h43 == _T_22[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_2;
      end else if (8'h43 == _T_19[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_1;
      end else if (8'h43 == _T_15[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_68 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h44 == _T_37[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_7;
      end else if (8'h44 == _T_34[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_6;
      end else if (8'h44 == _T_31[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_5;
      end else if (8'h44 == _T_28[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_4;
      end else if (8'h44 == _T_25[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_3;
      end else if (8'h44 == _T_22[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_2;
      end else if (8'h44 == _T_19[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_1;
      end else if (8'h44 == _T_15[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_69 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h45 == _T_37[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_7;
      end else if (8'h45 == _T_34[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_6;
      end else if (8'h45 == _T_31[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_5;
      end else if (8'h45 == _T_28[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_4;
      end else if (8'h45 == _T_25[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_3;
      end else if (8'h45 == _T_22[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_2;
      end else if (8'h45 == _T_19[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_1;
      end else if (8'h45 == _T_15[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_70 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h46 == _T_37[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_7;
      end else if (8'h46 == _T_34[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_6;
      end else if (8'h46 == _T_31[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_5;
      end else if (8'h46 == _T_28[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_4;
      end else if (8'h46 == _T_25[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_3;
      end else if (8'h46 == _T_22[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_2;
      end else if (8'h46 == _T_19[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_1;
      end else if (8'h46 == _T_15[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_71 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h47 == _T_37[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_7;
      end else if (8'h47 == _T_34[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_6;
      end else if (8'h47 == _T_31[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_5;
      end else if (8'h47 == _T_28[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_4;
      end else if (8'h47 == _T_25[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_3;
      end else if (8'h47 == _T_22[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_2;
      end else if (8'h47 == _T_19[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_1;
      end else if (8'h47 == _T_15[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_72 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h48 == _T_37[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_7;
      end else if (8'h48 == _T_34[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_6;
      end else if (8'h48 == _T_31[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_5;
      end else if (8'h48 == _T_28[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_4;
      end else if (8'h48 == _T_25[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_3;
      end else if (8'h48 == _T_22[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_2;
      end else if (8'h48 == _T_19[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_1;
      end else if (8'h48 == _T_15[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_73 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h49 == _T_37[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_7;
      end else if (8'h49 == _T_34[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_6;
      end else if (8'h49 == _T_31[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_5;
      end else if (8'h49 == _T_28[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_4;
      end else if (8'h49 == _T_25[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_3;
      end else if (8'h49 == _T_22[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_2;
      end else if (8'h49 == _T_19[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_1;
      end else if (8'h49 == _T_15[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_74 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4a == _T_37[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_7;
      end else if (8'h4a == _T_34[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_6;
      end else if (8'h4a == _T_31[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_5;
      end else if (8'h4a == _T_28[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_4;
      end else if (8'h4a == _T_25[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_3;
      end else if (8'h4a == _T_22[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_2;
      end else if (8'h4a == _T_19[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_1;
      end else if (8'h4a == _T_15[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_75 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4b == _T_37[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_7;
      end else if (8'h4b == _T_34[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_6;
      end else if (8'h4b == _T_31[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_5;
      end else if (8'h4b == _T_28[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_4;
      end else if (8'h4b == _T_25[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_3;
      end else if (8'h4b == _T_22[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_2;
      end else if (8'h4b == _T_19[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_1;
      end else if (8'h4b == _T_15[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_76 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4c == _T_37[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_7;
      end else if (8'h4c == _T_34[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_6;
      end else if (8'h4c == _T_31[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_5;
      end else if (8'h4c == _T_28[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_4;
      end else if (8'h4c == _T_25[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_3;
      end else if (8'h4c == _T_22[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_2;
      end else if (8'h4c == _T_19[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_1;
      end else if (8'h4c == _T_15[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_77 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4d == _T_37[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_7;
      end else if (8'h4d == _T_34[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_6;
      end else if (8'h4d == _T_31[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_5;
      end else if (8'h4d == _T_28[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_4;
      end else if (8'h4d == _T_25[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_3;
      end else if (8'h4d == _T_22[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_2;
      end else if (8'h4d == _T_19[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_1;
      end else if (8'h4d == _T_15[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_78 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4e == _T_37[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_7;
      end else if (8'h4e == _T_34[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_6;
      end else if (8'h4e == _T_31[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_5;
      end else if (8'h4e == _T_28[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_4;
      end else if (8'h4e == _T_25[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_3;
      end else if (8'h4e == _T_22[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_2;
      end else if (8'h4e == _T_19[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_1;
      end else if (8'h4e == _T_15[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_79 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4f == _T_37[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_7;
      end else if (8'h4f == _T_34[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_6;
      end else if (8'h4f == _T_31[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_5;
      end else if (8'h4f == _T_28[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_4;
      end else if (8'h4f == _T_25[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_3;
      end else if (8'h4f == _T_22[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_2;
      end else if (8'h4f == _T_19[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_1;
      end else if (8'h4f == _T_15[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_80 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h50 == _T_37[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_7;
      end else if (8'h50 == _T_34[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_6;
      end else if (8'h50 == _T_31[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_5;
      end else if (8'h50 == _T_28[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_4;
      end else if (8'h50 == _T_25[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_3;
      end else if (8'h50 == _T_22[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_2;
      end else if (8'h50 == _T_19[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_1;
      end else if (8'h50 == _T_15[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_81 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h51 == _T_37[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_7;
      end else if (8'h51 == _T_34[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_6;
      end else if (8'h51 == _T_31[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_5;
      end else if (8'h51 == _T_28[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_4;
      end else if (8'h51 == _T_25[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_3;
      end else if (8'h51 == _T_22[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_2;
      end else if (8'h51 == _T_19[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_1;
      end else if (8'h51 == _T_15[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_82 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h52 == _T_37[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_7;
      end else if (8'h52 == _T_34[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_6;
      end else if (8'h52 == _T_31[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_5;
      end else if (8'h52 == _T_28[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_4;
      end else if (8'h52 == _T_25[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_3;
      end else if (8'h52 == _T_22[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_2;
      end else if (8'h52 == _T_19[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_1;
      end else if (8'h52 == _T_15[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_83 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h53 == _T_37[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_7;
      end else if (8'h53 == _T_34[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_6;
      end else if (8'h53 == _T_31[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_5;
      end else if (8'h53 == _T_28[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_4;
      end else if (8'h53 == _T_25[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_3;
      end else if (8'h53 == _T_22[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_2;
      end else if (8'h53 == _T_19[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_1;
      end else if (8'h53 == _T_15[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_84 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h54 == _T_37[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_7;
      end else if (8'h54 == _T_34[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_6;
      end else if (8'h54 == _T_31[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_5;
      end else if (8'h54 == _T_28[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_4;
      end else if (8'h54 == _T_25[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_3;
      end else if (8'h54 == _T_22[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_2;
      end else if (8'h54 == _T_19[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_1;
      end else if (8'h54 == _T_15[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_85 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h55 == _T_37[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_7;
      end else if (8'h55 == _T_34[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_6;
      end else if (8'h55 == _T_31[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_5;
      end else if (8'h55 == _T_28[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_4;
      end else if (8'h55 == _T_25[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_3;
      end else if (8'h55 == _T_22[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_2;
      end else if (8'h55 == _T_19[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_1;
      end else if (8'h55 == _T_15[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_86 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h56 == _T_37[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_7;
      end else if (8'h56 == _T_34[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_6;
      end else if (8'h56 == _T_31[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_5;
      end else if (8'h56 == _T_28[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_4;
      end else if (8'h56 == _T_25[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_3;
      end else if (8'h56 == _T_22[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_2;
      end else if (8'h56 == _T_19[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_1;
      end else if (8'h56 == _T_15[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_87 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h57 == _T_37[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_7;
      end else if (8'h57 == _T_34[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_6;
      end else if (8'h57 == _T_31[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_5;
      end else if (8'h57 == _T_28[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_4;
      end else if (8'h57 == _T_25[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_3;
      end else if (8'h57 == _T_22[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_2;
      end else if (8'h57 == _T_19[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_1;
      end else if (8'h57 == _T_15[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_88 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h58 == _T_37[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_7;
      end else if (8'h58 == _T_34[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_6;
      end else if (8'h58 == _T_31[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_5;
      end else if (8'h58 == _T_28[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_4;
      end else if (8'h58 == _T_25[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_3;
      end else if (8'h58 == _T_22[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_2;
      end else if (8'h58 == _T_19[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_1;
      end else if (8'h58 == _T_15[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_89 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h59 == _T_37[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_7;
      end else if (8'h59 == _T_34[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_6;
      end else if (8'h59 == _T_31[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_5;
      end else if (8'h59 == _T_28[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_4;
      end else if (8'h59 == _T_25[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_3;
      end else if (8'h59 == _T_22[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_2;
      end else if (8'h59 == _T_19[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_1;
      end else if (8'h59 == _T_15[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_90 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5a == _T_37[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_7;
      end else if (8'h5a == _T_34[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_6;
      end else if (8'h5a == _T_31[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_5;
      end else if (8'h5a == _T_28[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_4;
      end else if (8'h5a == _T_25[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_3;
      end else if (8'h5a == _T_22[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_2;
      end else if (8'h5a == _T_19[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_1;
      end else if (8'h5a == _T_15[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_91 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5b == _T_37[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_7;
      end else if (8'h5b == _T_34[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_6;
      end else if (8'h5b == _T_31[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_5;
      end else if (8'h5b == _T_28[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_4;
      end else if (8'h5b == _T_25[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_3;
      end else if (8'h5b == _T_22[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_2;
      end else if (8'h5b == _T_19[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_1;
      end else if (8'h5b == _T_15[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_92 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5c == _T_37[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_7;
      end else if (8'h5c == _T_34[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_6;
      end else if (8'h5c == _T_31[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_5;
      end else if (8'h5c == _T_28[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_4;
      end else if (8'h5c == _T_25[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_3;
      end else if (8'h5c == _T_22[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_2;
      end else if (8'h5c == _T_19[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_1;
      end else if (8'h5c == _T_15[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_93 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5d == _T_37[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_7;
      end else if (8'h5d == _T_34[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_6;
      end else if (8'h5d == _T_31[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_5;
      end else if (8'h5d == _T_28[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_4;
      end else if (8'h5d == _T_25[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_3;
      end else if (8'h5d == _T_22[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_2;
      end else if (8'h5d == _T_19[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_1;
      end else if (8'h5d == _T_15[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_94 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5e == _T_37[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_7;
      end else if (8'h5e == _T_34[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_6;
      end else if (8'h5e == _T_31[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_5;
      end else if (8'h5e == _T_28[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_4;
      end else if (8'h5e == _T_25[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_3;
      end else if (8'h5e == _T_22[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_2;
      end else if (8'h5e == _T_19[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_1;
      end else if (8'h5e == _T_15[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_95 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5f == _T_37[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_7;
      end else if (8'h5f == _T_34[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_6;
      end else if (8'h5f == _T_31[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_5;
      end else if (8'h5f == _T_28[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_4;
      end else if (8'h5f == _T_25[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_3;
      end else if (8'h5f == _T_22[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_2;
      end else if (8'h5f == _T_19[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_1;
      end else if (8'h5f == _T_15[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_96 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h60 == _T_37[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_7;
      end else if (8'h60 == _T_34[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_6;
      end else if (8'h60 == _T_31[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_5;
      end else if (8'h60 == _T_28[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_4;
      end else if (8'h60 == _T_25[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_3;
      end else if (8'h60 == _T_22[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_2;
      end else if (8'h60 == _T_19[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_1;
      end else if (8'h60 == _T_15[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_97 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h61 == _T_37[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_7;
      end else if (8'h61 == _T_34[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_6;
      end else if (8'h61 == _T_31[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_5;
      end else if (8'h61 == _T_28[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_4;
      end else if (8'h61 == _T_25[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_3;
      end else if (8'h61 == _T_22[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_2;
      end else if (8'h61 == _T_19[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_1;
      end else if (8'h61 == _T_15[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_98 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h62 == _T_37[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_7;
      end else if (8'h62 == _T_34[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_6;
      end else if (8'h62 == _T_31[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_5;
      end else if (8'h62 == _T_28[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_4;
      end else if (8'h62 == _T_25[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_3;
      end else if (8'h62 == _T_22[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_2;
      end else if (8'h62 == _T_19[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_1;
      end else if (8'h62 == _T_15[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_99 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h63 == _T_37[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_7;
      end else if (8'h63 == _T_34[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_6;
      end else if (8'h63 == _T_31[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_5;
      end else if (8'h63 == _T_28[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_4;
      end else if (8'h63 == _T_25[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_3;
      end else if (8'h63 == _T_22[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_2;
      end else if (8'h63 == _T_19[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_1;
      end else if (8'h63 == _T_15[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_100 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h64 == _T_37[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_7;
      end else if (8'h64 == _T_34[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_6;
      end else if (8'h64 == _T_31[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_5;
      end else if (8'h64 == _T_28[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_4;
      end else if (8'h64 == _T_25[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_3;
      end else if (8'h64 == _T_22[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_2;
      end else if (8'h64 == _T_19[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_1;
      end else if (8'h64 == _T_15[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_101 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h65 == _T_37[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_7;
      end else if (8'h65 == _T_34[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_6;
      end else if (8'h65 == _T_31[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_5;
      end else if (8'h65 == _T_28[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_4;
      end else if (8'h65 == _T_25[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_3;
      end else if (8'h65 == _T_22[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_2;
      end else if (8'h65 == _T_19[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_1;
      end else if (8'h65 == _T_15[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_102 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h66 == _T_37[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_7;
      end else if (8'h66 == _T_34[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_6;
      end else if (8'h66 == _T_31[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_5;
      end else if (8'h66 == _T_28[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_4;
      end else if (8'h66 == _T_25[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_3;
      end else if (8'h66 == _T_22[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_2;
      end else if (8'h66 == _T_19[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_1;
      end else if (8'h66 == _T_15[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_103 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h67 == _T_37[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_7;
      end else if (8'h67 == _T_34[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_6;
      end else if (8'h67 == _T_31[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_5;
      end else if (8'h67 == _T_28[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_4;
      end else if (8'h67 == _T_25[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_3;
      end else if (8'h67 == _T_22[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_2;
      end else if (8'h67 == _T_19[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_1;
      end else if (8'h67 == _T_15[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_104 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h68 == _T_37[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_7;
      end else if (8'h68 == _T_34[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_6;
      end else if (8'h68 == _T_31[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_5;
      end else if (8'h68 == _T_28[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_4;
      end else if (8'h68 == _T_25[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_3;
      end else if (8'h68 == _T_22[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_2;
      end else if (8'h68 == _T_19[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_1;
      end else if (8'h68 == _T_15[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_105 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h69 == _T_37[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_7;
      end else if (8'h69 == _T_34[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_6;
      end else if (8'h69 == _T_31[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_5;
      end else if (8'h69 == _T_28[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_4;
      end else if (8'h69 == _T_25[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_3;
      end else if (8'h69 == _T_22[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_2;
      end else if (8'h69 == _T_19[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_1;
      end else if (8'h69 == _T_15[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_106 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6a == _T_37[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_7;
      end else if (8'h6a == _T_34[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_6;
      end else if (8'h6a == _T_31[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_5;
      end else if (8'h6a == _T_28[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_4;
      end else if (8'h6a == _T_25[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_3;
      end else if (8'h6a == _T_22[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_2;
      end else if (8'h6a == _T_19[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_1;
      end else if (8'h6a == _T_15[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_107 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6b == _T_37[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_7;
      end else if (8'h6b == _T_34[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_6;
      end else if (8'h6b == _T_31[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_5;
      end else if (8'h6b == _T_28[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_4;
      end else if (8'h6b == _T_25[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_3;
      end else if (8'h6b == _T_22[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_2;
      end else if (8'h6b == _T_19[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_1;
      end else if (8'h6b == _T_15[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_108 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6c == _T_37[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_7;
      end else if (8'h6c == _T_34[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_6;
      end else if (8'h6c == _T_31[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_5;
      end else if (8'h6c == _T_28[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_4;
      end else if (8'h6c == _T_25[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_3;
      end else if (8'h6c == _T_22[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_2;
      end else if (8'h6c == _T_19[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_1;
      end else if (8'h6c == _T_15[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_109 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6d == _T_37[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_7;
      end else if (8'h6d == _T_34[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_6;
      end else if (8'h6d == _T_31[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_5;
      end else if (8'h6d == _T_28[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_4;
      end else if (8'h6d == _T_25[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_3;
      end else if (8'h6d == _T_22[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_2;
      end else if (8'h6d == _T_19[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_1;
      end else if (8'h6d == _T_15[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_110 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6e == _T_37[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_7;
      end else if (8'h6e == _T_34[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_6;
      end else if (8'h6e == _T_31[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_5;
      end else if (8'h6e == _T_28[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_4;
      end else if (8'h6e == _T_25[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_3;
      end else if (8'h6e == _T_22[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_2;
      end else if (8'h6e == _T_19[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_1;
      end else if (8'h6e == _T_15[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_111 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6f == _T_37[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_7;
      end else if (8'h6f == _T_34[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_6;
      end else if (8'h6f == _T_31[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_5;
      end else if (8'h6f == _T_28[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_4;
      end else if (8'h6f == _T_25[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_3;
      end else if (8'h6f == _T_22[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_2;
      end else if (8'h6f == _T_19[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_1;
      end else if (8'h6f == _T_15[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_112 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h70 == _T_37[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_7;
      end else if (8'h70 == _T_34[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_6;
      end else if (8'h70 == _T_31[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_5;
      end else if (8'h70 == _T_28[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_4;
      end else if (8'h70 == _T_25[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_3;
      end else if (8'h70 == _T_22[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_2;
      end else if (8'h70 == _T_19[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_1;
      end else if (8'h70 == _T_15[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_113 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h71 == _T_37[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_7;
      end else if (8'h71 == _T_34[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_6;
      end else if (8'h71 == _T_31[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_5;
      end else if (8'h71 == _T_28[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_4;
      end else if (8'h71 == _T_25[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_3;
      end else if (8'h71 == _T_22[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_2;
      end else if (8'h71 == _T_19[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_1;
      end else if (8'h71 == _T_15[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_114 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h72 == _T_37[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_7;
      end else if (8'h72 == _T_34[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_6;
      end else if (8'h72 == _T_31[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_5;
      end else if (8'h72 == _T_28[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_4;
      end else if (8'h72 == _T_25[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_3;
      end else if (8'h72 == _T_22[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_2;
      end else if (8'h72 == _T_19[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_1;
      end else if (8'h72 == _T_15[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_115 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h73 == _T_37[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_7;
      end else if (8'h73 == _T_34[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_6;
      end else if (8'h73 == _T_31[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_5;
      end else if (8'h73 == _T_28[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_4;
      end else if (8'h73 == _T_25[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_3;
      end else if (8'h73 == _T_22[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_2;
      end else if (8'h73 == _T_19[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_1;
      end else if (8'h73 == _T_15[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_116 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h74 == _T_37[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_7;
      end else if (8'h74 == _T_34[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_6;
      end else if (8'h74 == _T_31[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_5;
      end else if (8'h74 == _T_28[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_4;
      end else if (8'h74 == _T_25[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_3;
      end else if (8'h74 == _T_22[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_2;
      end else if (8'h74 == _T_19[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_1;
      end else if (8'h74 == _T_15[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_117 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h75 == _T_37[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_7;
      end else if (8'h75 == _T_34[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_6;
      end else if (8'h75 == _T_31[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_5;
      end else if (8'h75 == _T_28[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_4;
      end else if (8'h75 == _T_25[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_3;
      end else if (8'h75 == _T_22[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_2;
      end else if (8'h75 == _T_19[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_1;
      end else if (8'h75 == _T_15[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_118 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h76 == _T_37[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_7;
      end else if (8'h76 == _T_34[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_6;
      end else if (8'h76 == _T_31[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_5;
      end else if (8'h76 == _T_28[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_4;
      end else if (8'h76 == _T_25[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_3;
      end else if (8'h76 == _T_22[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_2;
      end else if (8'h76 == _T_19[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_1;
      end else if (8'h76 == _T_15[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_119 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h77 == _T_37[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_7;
      end else if (8'h77 == _T_34[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_6;
      end else if (8'h77 == _T_31[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_5;
      end else if (8'h77 == _T_28[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_4;
      end else if (8'h77 == _T_25[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_3;
      end else if (8'h77 == _T_22[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_2;
      end else if (8'h77 == _T_19[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_1;
      end else if (8'h77 == _T_15[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_120 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h78 == _T_37[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_7;
      end else if (8'h78 == _T_34[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_6;
      end else if (8'h78 == _T_31[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_5;
      end else if (8'h78 == _T_28[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_4;
      end else if (8'h78 == _T_25[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_3;
      end else if (8'h78 == _T_22[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_2;
      end else if (8'h78 == _T_19[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_1;
      end else if (8'h78 == _T_15[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_121 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h79 == _T_37[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_7;
      end else if (8'h79 == _T_34[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_6;
      end else if (8'h79 == _T_31[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_5;
      end else if (8'h79 == _T_28[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_4;
      end else if (8'h79 == _T_25[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_3;
      end else if (8'h79 == _T_22[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_2;
      end else if (8'h79 == _T_19[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_1;
      end else if (8'h79 == _T_15[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_122 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7a == _T_37[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_7;
      end else if (8'h7a == _T_34[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_6;
      end else if (8'h7a == _T_31[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_5;
      end else if (8'h7a == _T_28[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_4;
      end else if (8'h7a == _T_25[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_3;
      end else if (8'h7a == _T_22[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_2;
      end else if (8'h7a == _T_19[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_1;
      end else if (8'h7a == _T_15[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_123 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7b == _T_37[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_7;
      end else if (8'h7b == _T_34[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_6;
      end else if (8'h7b == _T_31[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_5;
      end else if (8'h7b == _T_28[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_4;
      end else if (8'h7b == _T_25[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_3;
      end else if (8'h7b == _T_22[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_2;
      end else if (8'h7b == _T_19[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_1;
      end else if (8'h7b == _T_15[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_124 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7c == _T_37[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_7;
      end else if (8'h7c == _T_34[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_6;
      end else if (8'h7c == _T_31[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_5;
      end else if (8'h7c == _T_28[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_4;
      end else if (8'h7c == _T_25[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_3;
      end else if (8'h7c == _T_22[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_2;
      end else if (8'h7c == _T_19[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_1;
      end else if (8'h7c == _T_15[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_125 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7d == _T_37[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_7;
      end else if (8'h7d == _T_34[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_6;
      end else if (8'h7d == _T_31[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_5;
      end else if (8'h7d == _T_28[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_4;
      end else if (8'h7d == _T_25[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_3;
      end else if (8'h7d == _T_22[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_2;
      end else if (8'h7d == _T_19[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_1;
      end else if (8'h7d == _T_15[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_126 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7e == _T_37[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_7;
      end else if (8'h7e == _T_34[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_6;
      end else if (8'h7e == _T_31[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_5;
      end else if (8'h7e == _T_28[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_4;
      end else if (8'h7e == _T_25[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_3;
      end else if (8'h7e == _T_22[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_2;
      end else if (8'h7e == _T_19[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_1;
      end else if (8'h7e == _T_15[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_127 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7f == _T_37[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_7;
      end else if (8'h7f == _T_34[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_6;
      end else if (8'h7f == _T_31[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_5;
      end else if (8'h7f == _T_28[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_4;
      end else if (8'h7f == _T_25[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_3;
      end else if (8'h7f == _T_22[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_2;
      end else if (8'h7f == _T_19[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_1;
      end else if (8'h7f == _T_15[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_128 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h80 == _T_37[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_7;
      end else if (8'h80 == _T_34[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_6;
      end else if (8'h80 == _T_31[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_5;
      end else if (8'h80 == _T_28[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_4;
      end else if (8'h80 == _T_25[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_3;
      end else if (8'h80 == _T_22[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_2;
      end else if (8'h80 == _T_19[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_1;
      end else if (8'h80 == _T_15[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_129 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h81 == _T_37[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_7;
      end else if (8'h81 == _T_34[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_6;
      end else if (8'h81 == _T_31[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_5;
      end else if (8'h81 == _T_28[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_4;
      end else if (8'h81 == _T_25[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_3;
      end else if (8'h81 == _T_22[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_2;
      end else if (8'h81 == _T_19[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_1;
      end else if (8'h81 == _T_15[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_130 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h82 == _T_37[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_7;
      end else if (8'h82 == _T_34[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_6;
      end else if (8'h82 == _T_31[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_5;
      end else if (8'h82 == _T_28[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_4;
      end else if (8'h82 == _T_25[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_3;
      end else if (8'h82 == _T_22[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_2;
      end else if (8'h82 == _T_19[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_1;
      end else if (8'h82 == _T_15[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_131 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h83 == _T_37[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_7;
      end else if (8'h83 == _T_34[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_6;
      end else if (8'h83 == _T_31[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_5;
      end else if (8'h83 == _T_28[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_4;
      end else if (8'h83 == _T_25[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_3;
      end else if (8'h83 == _T_22[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_2;
      end else if (8'h83 == _T_19[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_1;
      end else if (8'h83 == _T_15[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_132 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h84 == _T_37[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_7;
      end else if (8'h84 == _T_34[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_6;
      end else if (8'h84 == _T_31[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_5;
      end else if (8'h84 == _T_28[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_4;
      end else if (8'h84 == _T_25[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_3;
      end else if (8'h84 == _T_22[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_2;
      end else if (8'h84 == _T_19[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_1;
      end else if (8'h84 == _T_15[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_133 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h85 == _T_37[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_7;
      end else if (8'h85 == _T_34[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_6;
      end else if (8'h85 == _T_31[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_5;
      end else if (8'h85 == _T_28[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_4;
      end else if (8'h85 == _T_25[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_3;
      end else if (8'h85 == _T_22[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_2;
      end else if (8'h85 == _T_19[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_1;
      end else if (8'h85 == _T_15[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_134 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h86 == _T_37[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_7;
      end else if (8'h86 == _T_34[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_6;
      end else if (8'h86 == _T_31[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_5;
      end else if (8'h86 == _T_28[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_4;
      end else if (8'h86 == _T_25[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_3;
      end else if (8'h86 == _T_22[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_2;
      end else if (8'h86 == _T_19[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_1;
      end else if (8'h86 == _T_15[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_135 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h87 == _T_37[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_7;
      end else if (8'h87 == _T_34[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_6;
      end else if (8'h87 == _T_31[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_5;
      end else if (8'h87 == _T_28[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_4;
      end else if (8'h87 == _T_25[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_3;
      end else if (8'h87 == _T_22[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_2;
      end else if (8'h87 == _T_19[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_1;
      end else if (8'h87 == _T_15[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_136 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h88 == _T_37[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_7;
      end else if (8'h88 == _T_34[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_6;
      end else if (8'h88 == _T_31[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_5;
      end else if (8'h88 == _T_28[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_4;
      end else if (8'h88 == _T_25[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_3;
      end else if (8'h88 == _T_22[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_2;
      end else if (8'h88 == _T_19[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_1;
      end else if (8'h88 == _T_15[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_137 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h89 == _T_37[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_7;
      end else if (8'h89 == _T_34[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_6;
      end else if (8'h89 == _T_31[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_5;
      end else if (8'h89 == _T_28[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_4;
      end else if (8'h89 == _T_25[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_3;
      end else if (8'h89 == _T_22[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_2;
      end else if (8'h89 == _T_19[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_1;
      end else if (8'h89 == _T_15[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_138 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8a == _T_37[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_7;
      end else if (8'h8a == _T_34[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_6;
      end else if (8'h8a == _T_31[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_5;
      end else if (8'h8a == _T_28[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_4;
      end else if (8'h8a == _T_25[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_3;
      end else if (8'h8a == _T_22[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_2;
      end else if (8'h8a == _T_19[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_1;
      end else if (8'h8a == _T_15[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_139 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8b == _T_37[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_7;
      end else if (8'h8b == _T_34[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_6;
      end else if (8'h8b == _T_31[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_5;
      end else if (8'h8b == _T_28[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_4;
      end else if (8'h8b == _T_25[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_3;
      end else if (8'h8b == _T_22[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_2;
      end else if (8'h8b == _T_19[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_1;
      end else if (8'h8b == _T_15[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_140 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8c == _T_37[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_7;
      end else if (8'h8c == _T_34[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_6;
      end else if (8'h8c == _T_31[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_5;
      end else if (8'h8c == _T_28[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_4;
      end else if (8'h8c == _T_25[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_3;
      end else if (8'h8c == _T_22[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_2;
      end else if (8'h8c == _T_19[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_1;
      end else if (8'h8c == _T_15[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_141 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8d == _T_37[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_7;
      end else if (8'h8d == _T_34[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_6;
      end else if (8'h8d == _T_31[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_5;
      end else if (8'h8d == _T_28[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_4;
      end else if (8'h8d == _T_25[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_3;
      end else if (8'h8d == _T_22[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_2;
      end else if (8'h8d == _T_19[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_1;
      end else if (8'h8d == _T_15[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_142 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8e == _T_37[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_7;
      end else if (8'h8e == _T_34[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_6;
      end else if (8'h8e == _T_31[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_5;
      end else if (8'h8e == _T_28[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_4;
      end else if (8'h8e == _T_25[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_3;
      end else if (8'h8e == _T_22[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_2;
      end else if (8'h8e == _T_19[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_1;
      end else if (8'h8e == _T_15[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_143 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8f == _T_37[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_7;
      end else if (8'h8f == _T_34[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_6;
      end else if (8'h8f == _T_31[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_5;
      end else if (8'h8f == _T_28[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_4;
      end else if (8'h8f == _T_25[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_3;
      end else if (8'h8f == _T_22[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_2;
      end else if (8'h8f == _T_19[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_1;
      end else if (8'h8f == _T_15[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_1_0 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h0 == _T_37[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_7;
      end else if (8'h0 == _T_34[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_6;
      end else if (8'h0 == _T_31[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_5;
      end else if (8'h0 == _T_28[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_4;
      end else if (8'h0 == _T_25[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_3;
      end else if (8'h0 == _T_22[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_2;
      end else if (8'h0 == _T_19[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_1;
      end else if (8'h0 == _T_15[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_1 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1 == _T_37[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_7;
      end else if (8'h1 == _T_34[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_6;
      end else if (8'h1 == _T_31[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_5;
      end else if (8'h1 == _T_28[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_4;
      end else if (8'h1 == _T_25[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_3;
      end else if (8'h1 == _T_22[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_2;
      end else if (8'h1 == _T_19[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_1;
      end else if (8'h1 == _T_15[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_2 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2 == _T_37[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_7;
      end else if (8'h2 == _T_34[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_6;
      end else if (8'h2 == _T_31[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_5;
      end else if (8'h2 == _T_28[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_4;
      end else if (8'h2 == _T_25[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_3;
      end else if (8'h2 == _T_22[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_2;
      end else if (8'h2 == _T_19[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_1;
      end else if (8'h2 == _T_15[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_3 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3 == _T_37[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_7;
      end else if (8'h3 == _T_34[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_6;
      end else if (8'h3 == _T_31[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_5;
      end else if (8'h3 == _T_28[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_4;
      end else if (8'h3 == _T_25[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_3;
      end else if (8'h3 == _T_22[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_2;
      end else if (8'h3 == _T_19[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_1;
      end else if (8'h3 == _T_15[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_4 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4 == _T_37[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_7;
      end else if (8'h4 == _T_34[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_6;
      end else if (8'h4 == _T_31[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_5;
      end else if (8'h4 == _T_28[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_4;
      end else if (8'h4 == _T_25[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_3;
      end else if (8'h4 == _T_22[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_2;
      end else if (8'h4 == _T_19[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_1;
      end else if (8'h4 == _T_15[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_5 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5 == _T_37[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_7;
      end else if (8'h5 == _T_34[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_6;
      end else if (8'h5 == _T_31[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_5;
      end else if (8'h5 == _T_28[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_4;
      end else if (8'h5 == _T_25[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_3;
      end else if (8'h5 == _T_22[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_2;
      end else if (8'h5 == _T_19[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_1;
      end else if (8'h5 == _T_15[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_6 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6 == _T_37[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_7;
      end else if (8'h6 == _T_34[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_6;
      end else if (8'h6 == _T_31[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_5;
      end else if (8'h6 == _T_28[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_4;
      end else if (8'h6 == _T_25[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_3;
      end else if (8'h6 == _T_22[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_2;
      end else if (8'h6 == _T_19[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_1;
      end else if (8'h6 == _T_15[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_7 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7 == _T_37[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_7;
      end else if (8'h7 == _T_34[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_6;
      end else if (8'h7 == _T_31[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_5;
      end else if (8'h7 == _T_28[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_4;
      end else if (8'h7 == _T_25[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_3;
      end else if (8'h7 == _T_22[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_2;
      end else if (8'h7 == _T_19[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_1;
      end else if (8'h7 == _T_15[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_8 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8 == _T_37[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_7;
      end else if (8'h8 == _T_34[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_6;
      end else if (8'h8 == _T_31[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_5;
      end else if (8'h8 == _T_28[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_4;
      end else if (8'h8 == _T_25[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_3;
      end else if (8'h8 == _T_22[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_2;
      end else if (8'h8 == _T_19[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_1;
      end else if (8'h8 == _T_15[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_9 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9 == _T_37[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_7;
      end else if (8'h9 == _T_34[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_6;
      end else if (8'h9 == _T_31[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_5;
      end else if (8'h9 == _T_28[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_4;
      end else if (8'h9 == _T_25[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_3;
      end else if (8'h9 == _T_22[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_2;
      end else if (8'h9 == _T_19[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_1;
      end else if (8'h9 == _T_15[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_10 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha == _T_37[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_7;
      end else if (8'ha == _T_34[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_6;
      end else if (8'ha == _T_31[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_5;
      end else if (8'ha == _T_28[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_4;
      end else if (8'ha == _T_25[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_3;
      end else if (8'ha == _T_22[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_2;
      end else if (8'ha == _T_19[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_1;
      end else if (8'ha == _T_15[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_11 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb == _T_37[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_7;
      end else if (8'hb == _T_34[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_6;
      end else if (8'hb == _T_31[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_5;
      end else if (8'hb == _T_28[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_4;
      end else if (8'hb == _T_25[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_3;
      end else if (8'hb == _T_22[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_2;
      end else if (8'hb == _T_19[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_1;
      end else if (8'hb == _T_15[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_12 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc == _T_37[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_7;
      end else if (8'hc == _T_34[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_6;
      end else if (8'hc == _T_31[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_5;
      end else if (8'hc == _T_28[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_4;
      end else if (8'hc == _T_25[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_3;
      end else if (8'hc == _T_22[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_2;
      end else if (8'hc == _T_19[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_1;
      end else if (8'hc == _T_15[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_13 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd == _T_37[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_7;
      end else if (8'hd == _T_34[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_6;
      end else if (8'hd == _T_31[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_5;
      end else if (8'hd == _T_28[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_4;
      end else if (8'hd == _T_25[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_3;
      end else if (8'hd == _T_22[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_2;
      end else if (8'hd == _T_19[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_1;
      end else if (8'hd == _T_15[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_14 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he == _T_37[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_7;
      end else if (8'he == _T_34[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_6;
      end else if (8'he == _T_31[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_5;
      end else if (8'he == _T_28[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_4;
      end else if (8'he == _T_25[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_3;
      end else if (8'he == _T_22[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_2;
      end else if (8'he == _T_19[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_1;
      end else if (8'he == _T_15[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_15 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf == _T_37[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_7;
      end else if (8'hf == _T_34[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_6;
      end else if (8'hf == _T_31[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_5;
      end else if (8'hf == _T_28[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_4;
      end else if (8'hf == _T_25[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_3;
      end else if (8'hf == _T_22[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_2;
      end else if (8'hf == _T_19[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_1;
      end else if (8'hf == _T_15[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_16 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h10 == _T_37[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_7;
      end else if (8'h10 == _T_34[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_6;
      end else if (8'h10 == _T_31[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_5;
      end else if (8'h10 == _T_28[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_4;
      end else if (8'h10 == _T_25[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_3;
      end else if (8'h10 == _T_22[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_2;
      end else if (8'h10 == _T_19[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_1;
      end else if (8'h10 == _T_15[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_17 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h11 == _T_37[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_7;
      end else if (8'h11 == _T_34[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_6;
      end else if (8'h11 == _T_31[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_5;
      end else if (8'h11 == _T_28[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_4;
      end else if (8'h11 == _T_25[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_3;
      end else if (8'h11 == _T_22[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_2;
      end else if (8'h11 == _T_19[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_1;
      end else if (8'h11 == _T_15[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_18 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h12 == _T_37[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_7;
      end else if (8'h12 == _T_34[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_6;
      end else if (8'h12 == _T_31[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_5;
      end else if (8'h12 == _T_28[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_4;
      end else if (8'h12 == _T_25[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_3;
      end else if (8'h12 == _T_22[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_2;
      end else if (8'h12 == _T_19[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_1;
      end else if (8'h12 == _T_15[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_19 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h13 == _T_37[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_7;
      end else if (8'h13 == _T_34[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_6;
      end else if (8'h13 == _T_31[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_5;
      end else if (8'h13 == _T_28[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_4;
      end else if (8'h13 == _T_25[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_3;
      end else if (8'h13 == _T_22[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_2;
      end else if (8'h13 == _T_19[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_1;
      end else if (8'h13 == _T_15[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_20 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h14 == _T_37[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_7;
      end else if (8'h14 == _T_34[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_6;
      end else if (8'h14 == _T_31[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_5;
      end else if (8'h14 == _T_28[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_4;
      end else if (8'h14 == _T_25[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_3;
      end else if (8'h14 == _T_22[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_2;
      end else if (8'h14 == _T_19[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_1;
      end else if (8'h14 == _T_15[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_21 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h15 == _T_37[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_7;
      end else if (8'h15 == _T_34[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_6;
      end else if (8'h15 == _T_31[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_5;
      end else if (8'h15 == _T_28[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_4;
      end else if (8'h15 == _T_25[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_3;
      end else if (8'h15 == _T_22[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_2;
      end else if (8'h15 == _T_19[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_1;
      end else if (8'h15 == _T_15[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_22 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h16 == _T_37[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_7;
      end else if (8'h16 == _T_34[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_6;
      end else if (8'h16 == _T_31[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_5;
      end else if (8'h16 == _T_28[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_4;
      end else if (8'h16 == _T_25[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_3;
      end else if (8'h16 == _T_22[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_2;
      end else if (8'h16 == _T_19[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_1;
      end else if (8'h16 == _T_15[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_23 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h17 == _T_37[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_7;
      end else if (8'h17 == _T_34[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_6;
      end else if (8'h17 == _T_31[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_5;
      end else if (8'h17 == _T_28[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_4;
      end else if (8'h17 == _T_25[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_3;
      end else if (8'h17 == _T_22[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_2;
      end else if (8'h17 == _T_19[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_1;
      end else if (8'h17 == _T_15[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_24 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h18 == _T_37[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_7;
      end else if (8'h18 == _T_34[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_6;
      end else if (8'h18 == _T_31[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_5;
      end else if (8'h18 == _T_28[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_4;
      end else if (8'h18 == _T_25[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_3;
      end else if (8'h18 == _T_22[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_2;
      end else if (8'h18 == _T_19[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_1;
      end else if (8'h18 == _T_15[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_25 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h19 == _T_37[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_7;
      end else if (8'h19 == _T_34[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_6;
      end else if (8'h19 == _T_31[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_5;
      end else if (8'h19 == _T_28[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_4;
      end else if (8'h19 == _T_25[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_3;
      end else if (8'h19 == _T_22[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_2;
      end else if (8'h19 == _T_19[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_1;
      end else if (8'h19 == _T_15[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_26 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1a == _T_37[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_7;
      end else if (8'h1a == _T_34[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_6;
      end else if (8'h1a == _T_31[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_5;
      end else if (8'h1a == _T_28[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_4;
      end else if (8'h1a == _T_25[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_3;
      end else if (8'h1a == _T_22[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_2;
      end else if (8'h1a == _T_19[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_1;
      end else if (8'h1a == _T_15[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_27 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1b == _T_37[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_7;
      end else if (8'h1b == _T_34[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_6;
      end else if (8'h1b == _T_31[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_5;
      end else if (8'h1b == _T_28[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_4;
      end else if (8'h1b == _T_25[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_3;
      end else if (8'h1b == _T_22[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_2;
      end else if (8'h1b == _T_19[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_1;
      end else if (8'h1b == _T_15[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_28 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1c == _T_37[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_7;
      end else if (8'h1c == _T_34[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_6;
      end else if (8'h1c == _T_31[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_5;
      end else if (8'h1c == _T_28[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_4;
      end else if (8'h1c == _T_25[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_3;
      end else if (8'h1c == _T_22[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_2;
      end else if (8'h1c == _T_19[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_1;
      end else if (8'h1c == _T_15[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_29 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1d == _T_37[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_7;
      end else if (8'h1d == _T_34[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_6;
      end else if (8'h1d == _T_31[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_5;
      end else if (8'h1d == _T_28[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_4;
      end else if (8'h1d == _T_25[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_3;
      end else if (8'h1d == _T_22[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_2;
      end else if (8'h1d == _T_19[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_1;
      end else if (8'h1d == _T_15[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_30 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1e == _T_37[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_7;
      end else if (8'h1e == _T_34[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_6;
      end else if (8'h1e == _T_31[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_5;
      end else if (8'h1e == _T_28[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_4;
      end else if (8'h1e == _T_25[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_3;
      end else if (8'h1e == _T_22[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_2;
      end else if (8'h1e == _T_19[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_1;
      end else if (8'h1e == _T_15[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_31 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1f == _T_37[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_7;
      end else if (8'h1f == _T_34[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_6;
      end else if (8'h1f == _T_31[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_5;
      end else if (8'h1f == _T_28[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_4;
      end else if (8'h1f == _T_25[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_3;
      end else if (8'h1f == _T_22[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_2;
      end else if (8'h1f == _T_19[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_1;
      end else if (8'h1f == _T_15[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_32 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h20 == _T_37[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_7;
      end else if (8'h20 == _T_34[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_6;
      end else if (8'h20 == _T_31[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_5;
      end else if (8'h20 == _T_28[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_4;
      end else if (8'h20 == _T_25[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_3;
      end else if (8'h20 == _T_22[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_2;
      end else if (8'h20 == _T_19[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_1;
      end else if (8'h20 == _T_15[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_33 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h21 == _T_37[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_7;
      end else if (8'h21 == _T_34[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_6;
      end else if (8'h21 == _T_31[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_5;
      end else if (8'h21 == _T_28[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_4;
      end else if (8'h21 == _T_25[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_3;
      end else if (8'h21 == _T_22[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_2;
      end else if (8'h21 == _T_19[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_1;
      end else if (8'h21 == _T_15[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_34 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h22 == _T_37[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_7;
      end else if (8'h22 == _T_34[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_6;
      end else if (8'h22 == _T_31[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_5;
      end else if (8'h22 == _T_28[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_4;
      end else if (8'h22 == _T_25[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_3;
      end else if (8'h22 == _T_22[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_2;
      end else if (8'h22 == _T_19[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_1;
      end else if (8'h22 == _T_15[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_35 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h23 == _T_37[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_7;
      end else if (8'h23 == _T_34[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_6;
      end else if (8'h23 == _T_31[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_5;
      end else if (8'h23 == _T_28[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_4;
      end else if (8'h23 == _T_25[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_3;
      end else if (8'h23 == _T_22[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_2;
      end else if (8'h23 == _T_19[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_1;
      end else if (8'h23 == _T_15[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_36 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h24 == _T_37[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_7;
      end else if (8'h24 == _T_34[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_6;
      end else if (8'h24 == _T_31[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_5;
      end else if (8'h24 == _T_28[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_4;
      end else if (8'h24 == _T_25[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_3;
      end else if (8'h24 == _T_22[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_2;
      end else if (8'h24 == _T_19[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_1;
      end else if (8'h24 == _T_15[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_37 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h25 == _T_37[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_7;
      end else if (8'h25 == _T_34[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_6;
      end else if (8'h25 == _T_31[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_5;
      end else if (8'h25 == _T_28[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_4;
      end else if (8'h25 == _T_25[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_3;
      end else if (8'h25 == _T_22[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_2;
      end else if (8'h25 == _T_19[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_1;
      end else if (8'h25 == _T_15[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_38 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h26 == _T_37[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_7;
      end else if (8'h26 == _T_34[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_6;
      end else if (8'h26 == _T_31[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_5;
      end else if (8'h26 == _T_28[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_4;
      end else if (8'h26 == _T_25[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_3;
      end else if (8'h26 == _T_22[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_2;
      end else if (8'h26 == _T_19[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_1;
      end else if (8'h26 == _T_15[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_39 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h27 == _T_37[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_7;
      end else if (8'h27 == _T_34[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_6;
      end else if (8'h27 == _T_31[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_5;
      end else if (8'h27 == _T_28[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_4;
      end else if (8'h27 == _T_25[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_3;
      end else if (8'h27 == _T_22[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_2;
      end else if (8'h27 == _T_19[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_1;
      end else if (8'h27 == _T_15[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_40 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h28 == _T_37[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_7;
      end else if (8'h28 == _T_34[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_6;
      end else if (8'h28 == _T_31[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_5;
      end else if (8'h28 == _T_28[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_4;
      end else if (8'h28 == _T_25[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_3;
      end else if (8'h28 == _T_22[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_2;
      end else if (8'h28 == _T_19[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_1;
      end else if (8'h28 == _T_15[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_41 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h29 == _T_37[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_7;
      end else if (8'h29 == _T_34[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_6;
      end else if (8'h29 == _T_31[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_5;
      end else if (8'h29 == _T_28[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_4;
      end else if (8'h29 == _T_25[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_3;
      end else if (8'h29 == _T_22[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_2;
      end else if (8'h29 == _T_19[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_1;
      end else if (8'h29 == _T_15[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_42 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2a == _T_37[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_7;
      end else if (8'h2a == _T_34[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_6;
      end else if (8'h2a == _T_31[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_5;
      end else if (8'h2a == _T_28[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_4;
      end else if (8'h2a == _T_25[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_3;
      end else if (8'h2a == _T_22[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_2;
      end else if (8'h2a == _T_19[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_1;
      end else if (8'h2a == _T_15[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_43 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2b == _T_37[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_7;
      end else if (8'h2b == _T_34[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_6;
      end else if (8'h2b == _T_31[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_5;
      end else if (8'h2b == _T_28[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_4;
      end else if (8'h2b == _T_25[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_3;
      end else if (8'h2b == _T_22[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_2;
      end else if (8'h2b == _T_19[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_1;
      end else if (8'h2b == _T_15[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_44 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2c == _T_37[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_7;
      end else if (8'h2c == _T_34[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_6;
      end else if (8'h2c == _T_31[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_5;
      end else if (8'h2c == _T_28[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_4;
      end else if (8'h2c == _T_25[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_3;
      end else if (8'h2c == _T_22[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_2;
      end else if (8'h2c == _T_19[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_1;
      end else if (8'h2c == _T_15[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_45 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2d == _T_37[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_7;
      end else if (8'h2d == _T_34[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_6;
      end else if (8'h2d == _T_31[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_5;
      end else if (8'h2d == _T_28[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_4;
      end else if (8'h2d == _T_25[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_3;
      end else if (8'h2d == _T_22[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_2;
      end else if (8'h2d == _T_19[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_1;
      end else if (8'h2d == _T_15[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_46 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2e == _T_37[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_7;
      end else if (8'h2e == _T_34[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_6;
      end else if (8'h2e == _T_31[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_5;
      end else if (8'h2e == _T_28[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_4;
      end else if (8'h2e == _T_25[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_3;
      end else if (8'h2e == _T_22[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_2;
      end else if (8'h2e == _T_19[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_1;
      end else if (8'h2e == _T_15[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_47 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2f == _T_37[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_7;
      end else if (8'h2f == _T_34[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_6;
      end else if (8'h2f == _T_31[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_5;
      end else if (8'h2f == _T_28[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_4;
      end else if (8'h2f == _T_25[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_3;
      end else if (8'h2f == _T_22[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_2;
      end else if (8'h2f == _T_19[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_1;
      end else if (8'h2f == _T_15[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_48 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h30 == _T_37[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_7;
      end else if (8'h30 == _T_34[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_6;
      end else if (8'h30 == _T_31[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_5;
      end else if (8'h30 == _T_28[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_4;
      end else if (8'h30 == _T_25[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_3;
      end else if (8'h30 == _T_22[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_2;
      end else if (8'h30 == _T_19[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_1;
      end else if (8'h30 == _T_15[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_49 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h31 == _T_37[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_7;
      end else if (8'h31 == _T_34[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_6;
      end else if (8'h31 == _T_31[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_5;
      end else if (8'h31 == _T_28[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_4;
      end else if (8'h31 == _T_25[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_3;
      end else if (8'h31 == _T_22[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_2;
      end else if (8'h31 == _T_19[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_1;
      end else if (8'h31 == _T_15[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_50 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h32 == _T_37[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_7;
      end else if (8'h32 == _T_34[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_6;
      end else if (8'h32 == _T_31[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_5;
      end else if (8'h32 == _T_28[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_4;
      end else if (8'h32 == _T_25[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_3;
      end else if (8'h32 == _T_22[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_2;
      end else if (8'h32 == _T_19[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_1;
      end else if (8'h32 == _T_15[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_51 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h33 == _T_37[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_7;
      end else if (8'h33 == _T_34[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_6;
      end else if (8'h33 == _T_31[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_5;
      end else if (8'h33 == _T_28[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_4;
      end else if (8'h33 == _T_25[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_3;
      end else if (8'h33 == _T_22[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_2;
      end else if (8'h33 == _T_19[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_1;
      end else if (8'h33 == _T_15[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_52 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h34 == _T_37[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_7;
      end else if (8'h34 == _T_34[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_6;
      end else if (8'h34 == _T_31[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_5;
      end else if (8'h34 == _T_28[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_4;
      end else if (8'h34 == _T_25[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_3;
      end else if (8'h34 == _T_22[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_2;
      end else if (8'h34 == _T_19[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_1;
      end else if (8'h34 == _T_15[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_53 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h35 == _T_37[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_7;
      end else if (8'h35 == _T_34[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_6;
      end else if (8'h35 == _T_31[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_5;
      end else if (8'h35 == _T_28[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_4;
      end else if (8'h35 == _T_25[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_3;
      end else if (8'h35 == _T_22[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_2;
      end else if (8'h35 == _T_19[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_1;
      end else if (8'h35 == _T_15[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_54 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h36 == _T_37[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_7;
      end else if (8'h36 == _T_34[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_6;
      end else if (8'h36 == _T_31[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_5;
      end else if (8'h36 == _T_28[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_4;
      end else if (8'h36 == _T_25[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_3;
      end else if (8'h36 == _T_22[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_2;
      end else if (8'h36 == _T_19[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_1;
      end else if (8'h36 == _T_15[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_55 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h37 == _T_37[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_7;
      end else if (8'h37 == _T_34[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_6;
      end else if (8'h37 == _T_31[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_5;
      end else if (8'h37 == _T_28[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_4;
      end else if (8'h37 == _T_25[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_3;
      end else if (8'h37 == _T_22[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_2;
      end else if (8'h37 == _T_19[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_1;
      end else if (8'h37 == _T_15[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_56 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h38 == _T_37[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_7;
      end else if (8'h38 == _T_34[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_6;
      end else if (8'h38 == _T_31[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_5;
      end else if (8'h38 == _T_28[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_4;
      end else if (8'h38 == _T_25[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_3;
      end else if (8'h38 == _T_22[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_2;
      end else if (8'h38 == _T_19[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_1;
      end else if (8'h38 == _T_15[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_57 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h39 == _T_37[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_7;
      end else if (8'h39 == _T_34[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_6;
      end else if (8'h39 == _T_31[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_5;
      end else if (8'h39 == _T_28[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_4;
      end else if (8'h39 == _T_25[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_3;
      end else if (8'h39 == _T_22[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_2;
      end else if (8'h39 == _T_19[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_1;
      end else if (8'h39 == _T_15[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_58 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3a == _T_37[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_7;
      end else if (8'h3a == _T_34[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_6;
      end else if (8'h3a == _T_31[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_5;
      end else if (8'h3a == _T_28[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_4;
      end else if (8'h3a == _T_25[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_3;
      end else if (8'h3a == _T_22[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_2;
      end else if (8'h3a == _T_19[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_1;
      end else if (8'h3a == _T_15[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_59 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3b == _T_37[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_7;
      end else if (8'h3b == _T_34[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_6;
      end else if (8'h3b == _T_31[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_5;
      end else if (8'h3b == _T_28[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_4;
      end else if (8'h3b == _T_25[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_3;
      end else if (8'h3b == _T_22[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_2;
      end else if (8'h3b == _T_19[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_1;
      end else if (8'h3b == _T_15[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_60 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3c == _T_37[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_7;
      end else if (8'h3c == _T_34[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_6;
      end else if (8'h3c == _T_31[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_5;
      end else if (8'h3c == _T_28[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_4;
      end else if (8'h3c == _T_25[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_3;
      end else if (8'h3c == _T_22[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_2;
      end else if (8'h3c == _T_19[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_1;
      end else if (8'h3c == _T_15[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_61 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3d == _T_37[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_7;
      end else if (8'h3d == _T_34[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_6;
      end else if (8'h3d == _T_31[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_5;
      end else if (8'h3d == _T_28[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_4;
      end else if (8'h3d == _T_25[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_3;
      end else if (8'h3d == _T_22[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_2;
      end else if (8'h3d == _T_19[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_1;
      end else if (8'h3d == _T_15[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_62 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3e == _T_37[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_7;
      end else if (8'h3e == _T_34[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_6;
      end else if (8'h3e == _T_31[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_5;
      end else if (8'h3e == _T_28[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_4;
      end else if (8'h3e == _T_25[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_3;
      end else if (8'h3e == _T_22[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_2;
      end else if (8'h3e == _T_19[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_1;
      end else if (8'h3e == _T_15[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_63 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3f == _T_37[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_7;
      end else if (8'h3f == _T_34[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_6;
      end else if (8'h3f == _T_31[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_5;
      end else if (8'h3f == _T_28[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_4;
      end else if (8'h3f == _T_25[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_3;
      end else if (8'h3f == _T_22[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_2;
      end else if (8'h3f == _T_19[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_1;
      end else if (8'h3f == _T_15[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_64 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h40 == _T_37[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_7;
      end else if (8'h40 == _T_34[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_6;
      end else if (8'h40 == _T_31[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_5;
      end else if (8'h40 == _T_28[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_4;
      end else if (8'h40 == _T_25[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_3;
      end else if (8'h40 == _T_22[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_2;
      end else if (8'h40 == _T_19[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_1;
      end else if (8'h40 == _T_15[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_65 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h41 == _T_37[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_7;
      end else if (8'h41 == _T_34[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_6;
      end else if (8'h41 == _T_31[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_5;
      end else if (8'h41 == _T_28[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_4;
      end else if (8'h41 == _T_25[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_3;
      end else if (8'h41 == _T_22[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_2;
      end else if (8'h41 == _T_19[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_1;
      end else if (8'h41 == _T_15[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_66 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h42 == _T_37[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_7;
      end else if (8'h42 == _T_34[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_6;
      end else if (8'h42 == _T_31[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_5;
      end else if (8'h42 == _T_28[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_4;
      end else if (8'h42 == _T_25[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_3;
      end else if (8'h42 == _T_22[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_2;
      end else if (8'h42 == _T_19[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_1;
      end else if (8'h42 == _T_15[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_67 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h43 == _T_37[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_7;
      end else if (8'h43 == _T_34[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_6;
      end else if (8'h43 == _T_31[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_5;
      end else if (8'h43 == _T_28[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_4;
      end else if (8'h43 == _T_25[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_3;
      end else if (8'h43 == _T_22[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_2;
      end else if (8'h43 == _T_19[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_1;
      end else if (8'h43 == _T_15[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_68 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h44 == _T_37[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_7;
      end else if (8'h44 == _T_34[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_6;
      end else if (8'h44 == _T_31[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_5;
      end else if (8'h44 == _T_28[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_4;
      end else if (8'h44 == _T_25[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_3;
      end else if (8'h44 == _T_22[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_2;
      end else if (8'h44 == _T_19[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_1;
      end else if (8'h44 == _T_15[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_69 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h45 == _T_37[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_7;
      end else if (8'h45 == _T_34[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_6;
      end else if (8'h45 == _T_31[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_5;
      end else if (8'h45 == _T_28[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_4;
      end else if (8'h45 == _T_25[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_3;
      end else if (8'h45 == _T_22[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_2;
      end else if (8'h45 == _T_19[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_1;
      end else if (8'h45 == _T_15[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_70 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h46 == _T_37[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_7;
      end else if (8'h46 == _T_34[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_6;
      end else if (8'h46 == _T_31[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_5;
      end else if (8'h46 == _T_28[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_4;
      end else if (8'h46 == _T_25[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_3;
      end else if (8'h46 == _T_22[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_2;
      end else if (8'h46 == _T_19[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_1;
      end else if (8'h46 == _T_15[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_71 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h47 == _T_37[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_7;
      end else if (8'h47 == _T_34[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_6;
      end else if (8'h47 == _T_31[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_5;
      end else if (8'h47 == _T_28[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_4;
      end else if (8'h47 == _T_25[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_3;
      end else if (8'h47 == _T_22[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_2;
      end else if (8'h47 == _T_19[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_1;
      end else if (8'h47 == _T_15[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_72 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h48 == _T_37[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_7;
      end else if (8'h48 == _T_34[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_6;
      end else if (8'h48 == _T_31[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_5;
      end else if (8'h48 == _T_28[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_4;
      end else if (8'h48 == _T_25[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_3;
      end else if (8'h48 == _T_22[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_2;
      end else if (8'h48 == _T_19[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_1;
      end else if (8'h48 == _T_15[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_73 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h49 == _T_37[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_7;
      end else if (8'h49 == _T_34[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_6;
      end else if (8'h49 == _T_31[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_5;
      end else if (8'h49 == _T_28[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_4;
      end else if (8'h49 == _T_25[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_3;
      end else if (8'h49 == _T_22[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_2;
      end else if (8'h49 == _T_19[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_1;
      end else if (8'h49 == _T_15[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_74 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4a == _T_37[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_7;
      end else if (8'h4a == _T_34[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_6;
      end else if (8'h4a == _T_31[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_5;
      end else if (8'h4a == _T_28[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_4;
      end else if (8'h4a == _T_25[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_3;
      end else if (8'h4a == _T_22[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_2;
      end else if (8'h4a == _T_19[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_1;
      end else if (8'h4a == _T_15[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_75 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4b == _T_37[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_7;
      end else if (8'h4b == _T_34[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_6;
      end else if (8'h4b == _T_31[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_5;
      end else if (8'h4b == _T_28[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_4;
      end else if (8'h4b == _T_25[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_3;
      end else if (8'h4b == _T_22[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_2;
      end else if (8'h4b == _T_19[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_1;
      end else if (8'h4b == _T_15[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_76 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4c == _T_37[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_7;
      end else if (8'h4c == _T_34[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_6;
      end else if (8'h4c == _T_31[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_5;
      end else if (8'h4c == _T_28[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_4;
      end else if (8'h4c == _T_25[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_3;
      end else if (8'h4c == _T_22[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_2;
      end else if (8'h4c == _T_19[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_1;
      end else if (8'h4c == _T_15[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_77 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4d == _T_37[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_7;
      end else if (8'h4d == _T_34[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_6;
      end else if (8'h4d == _T_31[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_5;
      end else if (8'h4d == _T_28[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_4;
      end else if (8'h4d == _T_25[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_3;
      end else if (8'h4d == _T_22[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_2;
      end else if (8'h4d == _T_19[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_1;
      end else if (8'h4d == _T_15[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_78 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4e == _T_37[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_7;
      end else if (8'h4e == _T_34[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_6;
      end else if (8'h4e == _T_31[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_5;
      end else if (8'h4e == _T_28[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_4;
      end else if (8'h4e == _T_25[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_3;
      end else if (8'h4e == _T_22[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_2;
      end else if (8'h4e == _T_19[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_1;
      end else if (8'h4e == _T_15[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_79 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4f == _T_37[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_7;
      end else if (8'h4f == _T_34[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_6;
      end else if (8'h4f == _T_31[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_5;
      end else if (8'h4f == _T_28[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_4;
      end else if (8'h4f == _T_25[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_3;
      end else if (8'h4f == _T_22[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_2;
      end else if (8'h4f == _T_19[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_1;
      end else if (8'h4f == _T_15[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_80 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h50 == _T_37[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_7;
      end else if (8'h50 == _T_34[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_6;
      end else if (8'h50 == _T_31[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_5;
      end else if (8'h50 == _T_28[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_4;
      end else if (8'h50 == _T_25[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_3;
      end else if (8'h50 == _T_22[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_2;
      end else if (8'h50 == _T_19[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_1;
      end else if (8'h50 == _T_15[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_81 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h51 == _T_37[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_7;
      end else if (8'h51 == _T_34[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_6;
      end else if (8'h51 == _T_31[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_5;
      end else if (8'h51 == _T_28[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_4;
      end else if (8'h51 == _T_25[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_3;
      end else if (8'h51 == _T_22[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_2;
      end else if (8'h51 == _T_19[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_1;
      end else if (8'h51 == _T_15[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_82 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h52 == _T_37[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_7;
      end else if (8'h52 == _T_34[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_6;
      end else if (8'h52 == _T_31[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_5;
      end else if (8'h52 == _T_28[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_4;
      end else if (8'h52 == _T_25[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_3;
      end else if (8'h52 == _T_22[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_2;
      end else if (8'h52 == _T_19[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_1;
      end else if (8'h52 == _T_15[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_83 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h53 == _T_37[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_7;
      end else if (8'h53 == _T_34[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_6;
      end else if (8'h53 == _T_31[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_5;
      end else if (8'h53 == _T_28[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_4;
      end else if (8'h53 == _T_25[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_3;
      end else if (8'h53 == _T_22[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_2;
      end else if (8'h53 == _T_19[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_1;
      end else if (8'h53 == _T_15[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_84 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h54 == _T_37[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_7;
      end else if (8'h54 == _T_34[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_6;
      end else if (8'h54 == _T_31[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_5;
      end else if (8'h54 == _T_28[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_4;
      end else if (8'h54 == _T_25[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_3;
      end else if (8'h54 == _T_22[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_2;
      end else if (8'h54 == _T_19[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_1;
      end else if (8'h54 == _T_15[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_85 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h55 == _T_37[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_7;
      end else if (8'h55 == _T_34[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_6;
      end else if (8'h55 == _T_31[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_5;
      end else if (8'h55 == _T_28[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_4;
      end else if (8'h55 == _T_25[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_3;
      end else if (8'h55 == _T_22[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_2;
      end else if (8'h55 == _T_19[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_1;
      end else if (8'h55 == _T_15[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_86 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h56 == _T_37[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_7;
      end else if (8'h56 == _T_34[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_6;
      end else if (8'h56 == _T_31[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_5;
      end else if (8'h56 == _T_28[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_4;
      end else if (8'h56 == _T_25[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_3;
      end else if (8'h56 == _T_22[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_2;
      end else if (8'h56 == _T_19[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_1;
      end else if (8'h56 == _T_15[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_87 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h57 == _T_37[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_7;
      end else if (8'h57 == _T_34[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_6;
      end else if (8'h57 == _T_31[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_5;
      end else if (8'h57 == _T_28[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_4;
      end else if (8'h57 == _T_25[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_3;
      end else if (8'h57 == _T_22[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_2;
      end else if (8'h57 == _T_19[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_1;
      end else if (8'h57 == _T_15[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_88 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h58 == _T_37[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_7;
      end else if (8'h58 == _T_34[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_6;
      end else if (8'h58 == _T_31[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_5;
      end else if (8'h58 == _T_28[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_4;
      end else if (8'h58 == _T_25[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_3;
      end else if (8'h58 == _T_22[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_2;
      end else if (8'h58 == _T_19[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_1;
      end else if (8'h58 == _T_15[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_89 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h59 == _T_37[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_7;
      end else if (8'h59 == _T_34[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_6;
      end else if (8'h59 == _T_31[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_5;
      end else if (8'h59 == _T_28[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_4;
      end else if (8'h59 == _T_25[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_3;
      end else if (8'h59 == _T_22[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_2;
      end else if (8'h59 == _T_19[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_1;
      end else if (8'h59 == _T_15[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_90 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5a == _T_37[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_7;
      end else if (8'h5a == _T_34[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_6;
      end else if (8'h5a == _T_31[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_5;
      end else if (8'h5a == _T_28[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_4;
      end else if (8'h5a == _T_25[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_3;
      end else if (8'h5a == _T_22[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_2;
      end else if (8'h5a == _T_19[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_1;
      end else if (8'h5a == _T_15[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_91 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5b == _T_37[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_7;
      end else if (8'h5b == _T_34[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_6;
      end else if (8'h5b == _T_31[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_5;
      end else if (8'h5b == _T_28[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_4;
      end else if (8'h5b == _T_25[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_3;
      end else if (8'h5b == _T_22[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_2;
      end else if (8'h5b == _T_19[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_1;
      end else if (8'h5b == _T_15[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_92 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5c == _T_37[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_7;
      end else if (8'h5c == _T_34[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_6;
      end else if (8'h5c == _T_31[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_5;
      end else if (8'h5c == _T_28[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_4;
      end else if (8'h5c == _T_25[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_3;
      end else if (8'h5c == _T_22[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_2;
      end else if (8'h5c == _T_19[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_1;
      end else if (8'h5c == _T_15[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_93 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5d == _T_37[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_7;
      end else if (8'h5d == _T_34[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_6;
      end else if (8'h5d == _T_31[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_5;
      end else if (8'h5d == _T_28[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_4;
      end else if (8'h5d == _T_25[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_3;
      end else if (8'h5d == _T_22[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_2;
      end else if (8'h5d == _T_19[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_1;
      end else if (8'h5d == _T_15[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_94 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5e == _T_37[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_7;
      end else if (8'h5e == _T_34[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_6;
      end else if (8'h5e == _T_31[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_5;
      end else if (8'h5e == _T_28[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_4;
      end else if (8'h5e == _T_25[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_3;
      end else if (8'h5e == _T_22[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_2;
      end else if (8'h5e == _T_19[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_1;
      end else if (8'h5e == _T_15[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_95 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5f == _T_37[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_7;
      end else if (8'h5f == _T_34[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_6;
      end else if (8'h5f == _T_31[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_5;
      end else if (8'h5f == _T_28[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_4;
      end else if (8'h5f == _T_25[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_3;
      end else if (8'h5f == _T_22[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_2;
      end else if (8'h5f == _T_19[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_1;
      end else if (8'h5f == _T_15[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_96 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h60 == _T_37[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_7;
      end else if (8'h60 == _T_34[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_6;
      end else if (8'h60 == _T_31[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_5;
      end else if (8'h60 == _T_28[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_4;
      end else if (8'h60 == _T_25[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_3;
      end else if (8'h60 == _T_22[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_2;
      end else if (8'h60 == _T_19[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_1;
      end else if (8'h60 == _T_15[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_97 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h61 == _T_37[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_7;
      end else if (8'h61 == _T_34[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_6;
      end else if (8'h61 == _T_31[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_5;
      end else if (8'h61 == _T_28[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_4;
      end else if (8'h61 == _T_25[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_3;
      end else if (8'h61 == _T_22[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_2;
      end else if (8'h61 == _T_19[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_1;
      end else if (8'h61 == _T_15[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_98 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h62 == _T_37[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_7;
      end else if (8'h62 == _T_34[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_6;
      end else if (8'h62 == _T_31[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_5;
      end else if (8'h62 == _T_28[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_4;
      end else if (8'h62 == _T_25[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_3;
      end else if (8'h62 == _T_22[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_2;
      end else if (8'h62 == _T_19[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_1;
      end else if (8'h62 == _T_15[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_99 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h63 == _T_37[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_7;
      end else if (8'h63 == _T_34[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_6;
      end else if (8'h63 == _T_31[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_5;
      end else if (8'h63 == _T_28[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_4;
      end else if (8'h63 == _T_25[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_3;
      end else if (8'h63 == _T_22[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_2;
      end else if (8'h63 == _T_19[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_1;
      end else if (8'h63 == _T_15[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_100 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h64 == _T_37[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_7;
      end else if (8'h64 == _T_34[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_6;
      end else if (8'h64 == _T_31[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_5;
      end else if (8'h64 == _T_28[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_4;
      end else if (8'h64 == _T_25[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_3;
      end else if (8'h64 == _T_22[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_2;
      end else if (8'h64 == _T_19[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_1;
      end else if (8'h64 == _T_15[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_101 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h65 == _T_37[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_7;
      end else if (8'h65 == _T_34[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_6;
      end else if (8'h65 == _T_31[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_5;
      end else if (8'h65 == _T_28[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_4;
      end else if (8'h65 == _T_25[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_3;
      end else if (8'h65 == _T_22[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_2;
      end else if (8'h65 == _T_19[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_1;
      end else if (8'h65 == _T_15[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_102 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h66 == _T_37[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_7;
      end else if (8'h66 == _T_34[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_6;
      end else if (8'h66 == _T_31[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_5;
      end else if (8'h66 == _T_28[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_4;
      end else if (8'h66 == _T_25[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_3;
      end else if (8'h66 == _T_22[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_2;
      end else if (8'h66 == _T_19[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_1;
      end else if (8'h66 == _T_15[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_103 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h67 == _T_37[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_7;
      end else if (8'h67 == _T_34[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_6;
      end else if (8'h67 == _T_31[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_5;
      end else if (8'h67 == _T_28[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_4;
      end else if (8'h67 == _T_25[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_3;
      end else if (8'h67 == _T_22[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_2;
      end else if (8'h67 == _T_19[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_1;
      end else if (8'h67 == _T_15[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_104 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h68 == _T_37[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_7;
      end else if (8'h68 == _T_34[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_6;
      end else if (8'h68 == _T_31[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_5;
      end else if (8'h68 == _T_28[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_4;
      end else if (8'h68 == _T_25[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_3;
      end else if (8'h68 == _T_22[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_2;
      end else if (8'h68 == _T_19[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_1;
      end else if (8'h68 == _T_15[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_105 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h69 == _T_37[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_7;
      end else if (8'h69 == _T_34[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_6;
      end else if (8'h69 == _T_31[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_5;
      end else if (8'h69 == _T_28[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_4;
      end else if (8'h69 == _T_25[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_3;
      end else if (8'h69 == _T_22[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_2;
      end else if (8'h69 == _T_19[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_1;
      end else if (8'h69 == _T_15[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_106 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6a == _T_37[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_7;
      end else if (8'h6a == _T_34[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_6;
      end else if (8'h6a == _T_31[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_5;
      end else if (8'h6a == _T_28[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_4;
      end else if (8'h6a == _T_25[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_3;
      end else if (8'h6a == _T_22[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_2;
      end else if (8'h6a == _T_19[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_1;
      end else if (8'h6a == _T_15[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_107 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6b == _T_37[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_7;
      end else if (8'h6b == _T_34[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_6;
      end else if (8'h6b == _T_31[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_5;
      end else if (8'h6b == _T_28[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_4;
      end else if (8'h6b == _T_25[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_3;
      end else if (8'h6b == _T_22[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_2;
      end else if (8'h6b == _T_19[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_1;
      end else if (8'h6b == _T_15[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_108 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6c == _T_37[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_7;
      end else if (8'h6c == _T_34[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_6;
      end else if (8'h6c == _T_31[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_5;
      end else if (8'h6c == _T_28[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_4;
      end else if (8'h6c == _T_25[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_3;
      end else if (8'h6c == _T_22[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_2;
      end else if (8'h6c == _T_19[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_1;
      end else if (8'h6c == _T_15[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_109 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6d == _T_37[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_7;
      end else if (8'h6d == _T_34[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_6;
      end else if (8'h6d == _T_31[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_5;
      end else if (8'h6d == _T_28[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_4;
      end else if (8'h6d == _T_25[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_3;
      end else if (8'h6d == _T_22[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_2;
      end else if (8'h6d == _T_19[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_1;
      end else if (8'h6d == _T_15[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_110 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6e == _T_37[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_7;
      end else if (8'h6e == _T_34[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_6;
      end else if (8'h6e == _T_31[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_5;
      end else if (8'h6e == _T_28[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_4;
      end else if (8'h6e == _T_25[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_3;
      end else if (8'h6e == _T_22[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_2;
      end else if (8'h6e == _T_19[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_1;
      end else if (8'h6e == _T_15[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_111 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6f == _T_37[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_7;
      end else if (8'h6f == _T_34[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_6;
      end else if (8'h6f == _T_31[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_5;
      end else if (8'h6f == _T_28[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_4;
      end else if (8'h6f == _T_25[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_3;
      end else if (8'h6f == _T_22[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_2;
      end else if (8'h6f == _T_19[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_1;
      end else if (8'h6f == _T_15[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_112 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h70 == _T_37[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_7;
      end else if (8'h70 == _T_34[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_6;
      end else if (8'h70 == _T_31[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_5;
      end else if (8'h70 == _T_28[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_4;
      end else if (8'h70 == _T_25[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_3;
      end else if (8'h70 == _T_22[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_2;
      end else if (8'h70 == _T_19[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_1;
      end else if (8'h70 == _T_15[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_113 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h71 == _T_37[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_7;
      end else if (8'h71 == _T_34[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_6;
      end else if (8'h71 == _T_31[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_5;
      end else if (8'h71 == _T_28[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_4;
      end else if (8'h71 == _T_25[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_3;
      end else if (8'h71 == _T_22[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_2;
      end else if (8'h71 == _T_19[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_1;
      end else if (8'h71 == _T_15[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_114 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h72 == _T_37[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_7;
      end else if (8'h72 == _T_34[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_6;
      end else if (8'h72 == _T_31[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_5;
      end else if (8'h72 == _T_28[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_4;
      end else if (8'h72 == _T_25[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_3;
      end else if (8'h72 == _T_22[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_2;
      end else if (8'h72 == _T_19[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_1;
      end else if (8'h72 == _T_15[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_115 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h73 == _T_37[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_7;
      end else if (8'h73 == _T_34[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_6;
      end else if (8'h73 == _T_31[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_5;
      end else if (8'h73 == _T_28[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_4;
      end else if (8'h73 == _T_25[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_3;
      end else if (8'h73 == _T_22[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_2;
      end else if (8'h73 == _T_19[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_1;
      end else if (8'h73 == _T_15[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_116 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h74 == _T_37[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_7;
      end else if (8'h74 == _T_34[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_6;
      end else if (8'h74 == _T_31[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_5;
      end else if (8'h74 == _T_28[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_4;
      end else if (8'h74 == _T_25[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_3;
      end else if (8'h74 == _T_22[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_2;
      end else if (8'h74 == _T_19[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_1;
      end else if (8'h74 == _T_15[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_117 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h75 == _T_37[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_7;
      end else if (8'h75 == _T_34[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_6;
      end else if (8'h75 == _T_31[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_5;
      end else if (8'h75 == _T_28[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_4;
      end else if (8'h75 == _T_25[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_3;
      end else if (8'h75 == _T_22[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_2;
      end else if (8'h75 == _T_19[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_1;
      end else if (8'h75 == _T_15[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_118 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h76 == _T_37[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_7;
      end else if (8'h76 == _T_34[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_6;
      end else if (8'h76 == _T_31[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_5;
      end else if (8'h76 == _T_28[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_4;
      end else if (8'h76 == _T_25[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_3;
      end else if (8'h76 == _T_22[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_2;
      end else if (8'h76 == _T_19[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_1;
      end else if (8'h76 == _T_15[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_119 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h77 == _T_37[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_7;
      end else if (8'h77 == _T_34[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_6;
      end else if (8'h77 == _T_31[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_5;
      end else if (8'h77 == _T_28[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_4;
      end else if (8'h77 == _T_25[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_3;
      end else if (8'h77 == _T_22[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_2;
      end else if (8'h77 == _T_19[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_1;
      end else if (8'h77 == _T_15[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_120 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h78 == _T_37[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_7;
      end else if (8'h78 == _T_34[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_6;
      end else if (8'h78 == _T_31[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_5;
      end else if (8'h78 == _T_28[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_4;
      end else if (8'h78 == _T_25[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_3;
      end else if (8'h78 == _T_22[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_2;
      end else if (8'h78 == _T_19[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_1;
      end else if (8'h78 == _T_15[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_121 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h79 == _T_37[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_7;
      end else if (8'h79 == _T_34[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_6;
      end else if (8'h79 == _T_31[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_5;
      end else if (8'h79 == _T_28[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_4;
      end else if (8'h79 == _T_25[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_3;
      end else if (8'h79 == _T_22[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_2;
      end else if (8'h79 == _T_19[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_1;
      end else if (8'h79 == _T_15[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_122 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7a == _T_37[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_7;
      end else if (8'h7a == _T_34[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_6;
      end else if (8'h7a == _T_31[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_5;
      end else if (8'h7a == _T_28[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_4;
      end else if (8'h7a == _T_25[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_3;
      end else if (8'h7a == _T_22[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_2;
      end else if (8'h7a == _T_19[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_1;
      end else if (8'h7a == _T_15[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_123 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7b == _T_37[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_7;
      end else if (8'h7b == _T_34[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_6;
      end else if (8'h7b == _T_31[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_5;
      end else if (8'h7b == _T_28[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_4;
      end else if (8'h7b == _T_25[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_3;
      end else if (8'h7b == _T_22[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_2;
      end else if (8'h7b == _T_19[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_1;
      end else if (8'h7b == _T_15[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_124 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7c == _T_37[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_7;
      end else if (8'h7c == _T_34[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_6;
      end else if (8'h7c == _T_31[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_5;
      end else if (8'h7c == _T_28[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_4;
      end else if (8'h7c == _T_25[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_3;
      end else if (8'h7c == _T_22[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_2;
      end else if (8'h7c == _T_19[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_1;
      end else if (8'h7c == _T_15[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_125 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7d == _T_37[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_7;
      end else if (8'h7d == _T_34[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_6;
      end else if (8'h7d == _T_31[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_5;
      end else if (8'h7d == _T_28[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_4;
      end else if (8'h7d == _T_25[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_3;
      end else if (8'h7d == _T_22[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_2;
      end else if (8'h7d == _T_19[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_1;
      end else if (8'h7d == _T_15[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_126 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7e == _T_37[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_7;
      end else if (8'h7e == _T_34[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_6;
      end else if (8'h7e == _T_31[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_5;
      end else if (8'h7e == _T_28[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_4;
      end else if (8'h7e == _T_25[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_3;
      end else if (8'h7e == _T_22[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_2;
      end else if (8'h7e == _T_19[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_1;
      end else if (8'h7e == _T_15[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_127 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7f == _T_37[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_7;
      end else if (8'h7f == _T_34[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_6;
      end else if (8'h7f == _T_31[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_5;
      end else if (8'h7f == _T_28[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_4;
      end else if (8'h7f == _T_25[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_3;
      end else if (8'h7f == _T_22[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_2;
      end else if (8'h7f == _T_19[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_1;
      end else if (8'h7f == _T_15[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_128 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h80 == _T_37[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_7;
      end else if (8'h80 == _T_34[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_6;
      end else if (8'h80 == _T_31[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_5;
      end else if (8'h80 == _T_28[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_4;
      end else if (8'h80 == _T_25[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_3;
      end else if (8'h80 == _T_22[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_2;
      end else if (8'h80 == _T_19[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_1;
      end else if (8'h80 == _T_15[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_129 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h81 == _T_37[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_7;
      end else if (8'h81 == _T_34[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_6;
      end else if (8'h81 == _T_31[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_5;
      end else if (8'h81 == _T_28[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_4;
      end else if (8'h81 == _T_25[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_3;
      end else if (8'h81 == _T_22[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_2;
      end else if (8'h81 == _T_19[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_1;
      end else if (8'h81 == _T_15[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_130 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h82 == _T_37[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_7;
      end else if (8'h82 == _T_34[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_6;
      end else if (8'h82 == _T_31[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_5;
      end else if (8'h82 == _T_28[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_4;
      end else if (8'h82 == _T_25[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_3;
      end else if (8'h82 == _T_22[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_2;
      end else if (8'h82 == _T_19[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_1;
      end else if (8'h82 == _T_15[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_131 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h83 == _T_37[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_7;
      end else if (8'h83 == _T_34[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_6;
      end else if (8'h83 == _T_31[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_5;
      end else if (8'h83 == _T_28[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_4;
      end else if (8'h83 == _T_25[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_3;
      end else if (8'h83 == _T_22[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_2;
      end else if (8'h83 == _T_19[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_1;
      end else if (8'h83 == _T_15[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_132 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h84 == _T_37[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_7;
      end else if (8'h84 == _T_34[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_6;
      end else if (8'h84 == _T_31[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_5;
      end else if (8'h84 == _T_28[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_4;
      end else if (8'h84 == _T_25[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_3;
      end else if (8'h84 == _T_22[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_2;
      end else if (8'h84 == _T_19[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_1;
      end else if (8'h84 == _T_15[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_133 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h85 == _T_37[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_7;
      end else if (8'h85 == _T_34[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_6;
      end else if (8'h85 == _T_31[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_5;
      end else if (8'h85 == _T_28[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_4;
      end else if (8'h85 == _T_25[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_3;
      end else if (8'h85 == _T_22[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_2;
      end else if (8'h85 == _T_19[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_1;
      end else if (8'h85 == _T_15[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_134 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h86 == _T_37[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_7;
      end else if (8'h86 == _T_34[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_6;
      end else if (8'h86 == _T_31[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_5;
      end else if (8'h86 == _T_28[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_4;
      end else if (8'h86 == _T_25[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_3;
      end else if (8'h86 == _T_22[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_2;
      end else if (8'h86 == _T_19[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_1;
      end else if (8'h86 == _T_15[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_135 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h87 == _T_37[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_7;
      end else if (8'h87 == _T_34[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_6;
      end else if (8'h87 == _T_31[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_5;
      end else if (8'h87 == _T_28[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_4;
      end else if (8'h87 == _T_25[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_3;
      end else if (8'h87 == _T_22[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_2;
      end else if (8'h87 == _T_19[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_1;
      end else if (8'h87 == _T_15[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_136 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h88 == _T_37[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_7;
      end else if (8'h88 == _T_34[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_6;
      end else if (8'h88 == _T_31[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_5;
      end else if (8'h88 == _T_28[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_4;
      end else if (8'h88 == _T_25[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_3;
      end else if (8'h88 == _T_22[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_2;
      end else if (8'h88 == _T_19[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_1;
      end else if (8'h88 == _T_15[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_137 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h89 == _T_37[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_7;
      end else if (8'h89 == _T_34[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_6;
      end else if (8'h89 == _T_31[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_5;
      end else if (8'h89 == _T_28[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_4;
      end else if (8'h89 == _T_25[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_3;
      end else if (8'h89 == _T_22[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_2;
      end else if (8'h89 == _T_19[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_1;
      end else if (8'h89 == _T_15[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_138 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8a == _T_37[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_7;
      end else if (8'h8a == _T_34[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_6;
      end else if (8'h8a == _T_31[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_5;
      end else if (8'h8a == _T_28[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_4;
      end else if (8'h8a == _T_25[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_3;
      end else if (8'h8a == _T_22[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_2;
      end else if (8'h8a == _T_19[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_1;
      end else if (8'h8a == _T_15[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_139 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8b == _T_37[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_7;
      end else if (8'h8b == _T_34[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_6;
      end else if (8'h8b == _T_31[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_5;
      end else if (8'h8b == _T_28[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_4;
      end else if (8'h8b == _T_25[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_3;
      end else if (8'h8b == _T_22[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_2;
      end else if (8'h8b == _T_19[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_1;
      end else if (8'h8b == _T_15[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_140 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8c == _T_37[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_7;
      end else if (8'h8c == _T_34[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_6;
      end else if (8'h8c == _T_31[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_5;
      end else if (8'h8c == _T_28[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_4;
      end else if (8'h8c == _T_25[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_3;
      end else if (8'h8c == _T_22[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_2;
      end else if (8'h8c == _T_19[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_1;
      end else if (8'h8c == _T_15[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_141 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8d == _T_37[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_7;
      end else if (8'h8d == _T_34[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_6;
      end else if (8'h8d == _T_31[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_5;
      end else if (8'h8d == _T_28[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_4;
      end else if (8'h8d == _T_25[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_3;
      end else if (8'h8d == _T_22[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_2;
      end else if (8'h8d == _T_19[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_1;
      end else if (8'h8d == _T_15[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_142 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8e == _T_37[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_7;
      end else if (8'h8e == _T_34[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_6;
      end else if (8'h8e == _T_31[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_5;
      end else if (8'h8e == _T_28[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_4;
      end else if (8'h8e == _T_25[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_3;
      end else if (8'h8e == _T_22[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_2;
      end else if (8'h8e == _T_19[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_1;
      end else if (8'h8e == _T_15[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_143 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8f == _T_37[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_7;
      end else if (8'h8f == _T_34[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_6;
      end else if (8'h8f == _T_31[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_5;
      end else if (8'h8f == _T_28[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_4;
      end else if (8'h8f == _T_25[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_3;
      end else if (8'h8f == _T_22[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_2;
      end else if (8'h8f == _T_19[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_1;
      end else if (8'h8f == _T_15[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_2_0 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h0 == _T_37[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_7;
      end else if (8'h0 == _T_34[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_6;
      end else if (8'h0 == _T_31[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_5;
      end else if (8'h0 == _T_28[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_4;
      end else if (8'h0 == _T_25[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_3;
      end else if (8'h0 == _T_22[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_2;
      end else if (8'h0 == _T_19[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_1;
      end else if (8'h0 == _T_15[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_1 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1 == _T_37[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_7;
      end else if (8'h1 == _T_34[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_6;
      end else if (8'h1 == _T_31[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_5;
      end else if (8'h1 == _T_28[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_4;
      end else if (8'h1 == _T_25[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_3;
      end else if (8'h1 == _T_22[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_2;
      end else if (8'h1 == _T_19[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_1;
      end else if (8'h1 == _T_15[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_2 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2 == _T_37[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_7;
      end else if (8'h2 == _T_34[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_6;
      end else if (8'h2 == _T_31[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_5;
      end else if (8'h2 == _T_28[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_4;
      end else if (8'h2 == _T_25[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_3;
      end else if (8'h2 == _T_22[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_2;
      end else if (8'h2 == _T_19[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_1;
      end else if (8'h2 == _T_15[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_3 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3 == _T_37[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_7;
      end else if (8'h3 == _T_34[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_6;
      end else if (8'h3 == _T_31[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_5;
      end else if (8'h3 == _T_28[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_4;
      end else if (8'h3 == _T_25[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_3;
      end else if (8'h3 == _T_22[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_2;
      end else if (8'h3 == _T_19[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_1;
      end else if (8'h3 == _T_15[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_4 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4 == _T_37[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_7;
      end else if (8'h4 == _T_34[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_6;
      end else if (8'h4 == _T_31[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_5;
      end else if (8'h4 == _T_28[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_4;
      end else if (8'h4 == _T_25[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_3;
      end else if (8'h4 == _T_22[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_2;
      end else if (8'h4 == _T_19[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_1;
      end else if (8'h4 == _T_15[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_5 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5 == _T_37[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_7;
      end else if (8'h5 == _T_34[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_6;
      end else if (8'h5 == _T_31[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_5;
      end else if (8'h5 == _T_28[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_4;
      end else if (8'h5 == _T_25[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_3;
      end else if (8'h5 == _T_22[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_2;
      end else if (8'h5 == _T_19[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_1;
      end else if (8'h5 == _T_15[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_6 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6 == _T_37[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_7;
      end else if (8'h6 == _T_34[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_6;
      end else if (8'h6 == _T_31[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_5;
      end else if (8'h6 == _T_28[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_4;
      end else if (8'h6 == _T_25[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_3;
      end else if (8'h6 == _T_22[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_2;
      end else if (8'h6 == _T_19[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_1;
      end else if (8'h6 == _T_15[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_7 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7 == _T_37[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_7;
      end else if (8'h7 == _T_34[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_6;
      end else if (8'h7 == _T_31[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_5;
      end else if (8'h7 == _T_28[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_4;
      end else if (8'h7 == _T_25[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_3;
      end else if (8'h7 == _T_22[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_2;
      end else if (8'h7 == _T_19[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_1;
      end else if (8'h7 == _T_15[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_8 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8 == _T_37[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_7;
      end else if (8'h8 == _T_34[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_6;
      end else if (8'h8 == _T_31[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_5;
      end else if (8'h8 == _T_28[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_4;
      end else if (8'h8 == _T_25[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_3;
      end else if (8'h8 == _T_22[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_2;
      end else if (8'h8 == _T_19[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_1;
      end else if (8'h8 == _T_15[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_9 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9 == _T_37[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_7;
      end else if (8'h9 == _T_34[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_6;
      end else if (8'h9 == _T_31[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_5;
      end else if (8'h9 == _T_28[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_4;
      end else if (8'h9 == _T_25[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_3;
      end else if (8'h9 == _T_22[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_2;
      end else if (8'h9 == _T_19[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_1;
      end else if (8'h9 == _T_15[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_10 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha == _T_37[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_7;
      end else if (8'ha == _T_34[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_6;
      end else if (8'ha == _T_31[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_5;
      end else if (8'ha == _T_28[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_4;
      end else if (8'ha == _T_25[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_3;
      end else if (8'ha == _T_22[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_2;
      end else if (8'ha == _T_19[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_1;
      end else if (8'ha == _T_15[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_11 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb == _T_37[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_7;
      end else if (8'hb == _T_34[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_6;
      end else if (8'hb == _T_31[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_5;
      end else if (8'hb == _T_28[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_4;
      end else if (8'hb == _T_25[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_3;
      end else if (8'hb == _T_22[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_2;
      end else if (8'hb == _T_19[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_1;
      end else if (8'hb == _T_15[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_12 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc == _T_37[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_7;
      end else if (8'hc == _T_34[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_6;
      end else if (8'hc == _T_31[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_5;
      end else if (8'hc == _T_28[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_4;
      end else if (8'hc == _T_25[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_3;
      end else if (8'hc == _T_22[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_2;
      end else if (8'hc == _T_19[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_1;
      end else if (8'hc == _T_15[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_13 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd == _T_37[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_7;
      end else if (8'hd == _T_34[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_6;
      end else if (8'hd == _T_31[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_5;
      end else if (8'hd == _T_28[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_4;
      end else if (8'hd == _T_25[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_3;
      end else if (8'hd == _T_22[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_2;
      end else if (8'hd == _T_19[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_1;
      end else if (8'hd == _T_15[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_14 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he == _T_37[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_7;
      end else if (8'he == _T_34[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_6;
      end else if (8'he == _T_31[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_5;
      end else if (8'he == _T_28[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_4;
      end else if (8'he == _T_25[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_3;
      end else if (8'he == _T_22[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_2;
      end else if (8'he == _T_19[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_1;
      end else if (8'he == _T_15[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_15 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf == _T_37[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_7;
      end else if (8'hf == _T_34[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_6;
      end else if (8'hf == _T_31[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_5;
      end else if (8'hf == _T_28[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_4;
      end else if (8'hf == _T_25[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_3;
      end else if (8'hf == _T_22[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_2;
      end else if (8'hf == _T_19[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_1;
      end else if (8'hf == _T_15[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_16 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h10 == _T_37[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_7;
      end else if (8'h10 == _T_34[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_6;
      end else if (8'h10 == _T_31[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_5;
      end else if (8'h10 == _T_28[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_4;
      end else if (8'h10 == _T_25[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_3;
      end else if (8'h10 == _T_22[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_2;
      end else if (8'h10 == _T_19[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_1;
      end else if (8'h10 == _T_15[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_17 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h11 == _T_37[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_7;
      end else if (8'h11 == _T_34[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_6;
      end else if (8'h11 == _T_31[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_5;
      end else if (8'h11 == _T_28[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_4;
      end else if (8'h11 == _T_25[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_3;
      end else if (8'h11 == _T_22[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_2;
      end else if (8'h11 == _T_19[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_1;
      end else if (8'h11 == _T_15[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_18 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h12 == _T_37[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_7;
      end else if (8'h12 == _T_34[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_6;
      end else if (8'h12 == _T_31[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_5;
      end else if (8'h12 == _T_28[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_4;
      end else if (8'h12 == _T_25[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_3;
      end else if (8'h12 == _T_22[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_2;
      end else if (8'h12 == _T_19[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_1;
      end else if (8'h12 == _T_15[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_19 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h13 == _T_37[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_7;
      end else if (8'h13 == _T_34[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_6;
      end else if (8'h13 == _T_31[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_5;
      end else if (8'h13 == _T_28[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_4;
      end else if (8'h13 == _T_25[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_3;
      end else if (8'h13 == _T_22[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_2;
      end else if (8'h13 == _T_19[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_1;
      end else if (8'h13 == _T_15[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_20 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h14 == _T_37[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_7;
      end else if (8'h14 == _T_34[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_6;
      end else if (8'h14 == _T_31[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_5;
      end else if (8'h14 == _T_28[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_4;
      end else if (8'h14 == _T_25[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_3;
      end else if (8'h14 == _T_22[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_2;
      end else if (8'h14 == _T_19[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_1;
      end else if (8'h14 == _T_15[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_21 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h15 == _T_37[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_7;
      end else if (8'h15 == _T_34[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_6;
      end else if (8'h15 == _T_31[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_5;
      end else if (8'h15 == _T_28[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_4;
      end else if (8'h15 == _T_25[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_3;
      end else if (8'h15 == _T_22[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_2;
      end else if (8'h15 == _T_19[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_1;
      end else if (8'h15 == _T_15[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_22 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h16 == _T_37[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_7;
      end else if (8'h16 == _T_34[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_6;
      end else if (8'h16 == _T_31[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_5;
      end else if (8'h16 == _T_28[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_4;
      end else if (8'h16 == _T_25[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_3;
      end else if (8'h16 == _T_22[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_2;
      end else if (8'h16 == _T_19[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_1;
      end else if (8'h16 == _T_15[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_23 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h17 == _T_37[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_7;
      end else if (8'h17 == _T_34[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_6;
      end else if (8'h17 == _T_31[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_5;
      end else if (8'h17 == _T_28[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_4;
      end else if (8'h17 == _T_25[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_3;
      end else if (8'h17 == _T_22[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_2;
      end else if (8'h17 == _T_19[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_1;
      end else if (8'h17 == _T_15[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_24 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h18 == _T_37[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_7;
      end else if (8'h18 == _T_34[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_6;
      end else if (8'h18 == _T_31[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_5;
      end else if (8'h18 == _T_28[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_4;
      end else if (8'h18 == _T_25[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_3;
      end else if (8'h18 == _T_22[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_2;
      end else if (8'h18 == _T_19[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_1;
      end else if (8'h18 == _T_15[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_25 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h19 == _T_37[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_7;
      end else if (8'h19 == _T_34[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_6;
      end else if (8'h19 == _T_31[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_5;
      end else if (8'h19 == _T_28[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_4;
      end else if (8'h19 == _T_25[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_3;
      end else if (8'h19 == _T_22[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_2;
      end else if (8'h19 == _T_19[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_1;
      end else if (8'h19 == _T_15[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_26 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1a == _T_37[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_7;
      end else if (8'h1a == _T_34[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_6;
      end else if (8'h1a == _T_31[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_5;
      end else if (8'h1a == _T_28[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_4;
      end else if (8'h1a == _T_25[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_3;
      end else if (8'h1a == _T_22[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_2;
      end else if (8'h1a == _T_19[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_1;
      end else if (8'h1a == _T_15[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_27 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1b == _T_37[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_7;
      end else if (8'h1b == _T_34[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_6;
      end else if (8'h1b == _T_31[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_5;
      end else if (8'h1b == _T_28[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_4;
      end else if (8'h1b == _T_25[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_3;
      end else if (8'h1b == _T_22[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_2;
      end else if (8'h1b == _T_19[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_1;
      end else if (8'h1b == _T_15[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_28 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1c == _T_37[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_7;
      end else if (8'h1c == _T_34[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_6;
      end else if (8'h1c == _T_31[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_5;
      end else if (8'h1c == _T_28[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_4;
      end else if (8'h1c == _T_25[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_3;
      end else if (8'h1c == _T_22[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_2;
      end else if (8'h1c == _T_19[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_1;
      end else if (8'h1c == _T_15[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_29 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1d == _T_37[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_7;
      end else if (8'h1d == _T_34[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_6;
      end else if (8'h1d == _T_31[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_5;
      end else if (8'h1d == _T_28[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_4;
      end else if (8'h1d == _T_25[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_3;
      end else if (8'h1d == _T_22[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_2;
      end else if (8'h1d == _T_19[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_1;
      end else if (8'h1d == _T_15[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_30 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1e == _T_37[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_7;
      end else if (8'h1e == _T_34[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_6;
      end else if (8'h1e == _T_31[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_5;
      end else if (8'h1e == _T_28[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_4;
      end else if (8'h1e == _T_25[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_3;
      end else if (8'h1e == _T_22[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_2;
      end else if (8'h1e == _T_19[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_1;
      end else if (8'h1e == _T_15[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_31 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1f == _T_37[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_7;
      end else if (8'h1f == _T_34[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_6;
      end else if (8'h1f == _T_31[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_5;
      end else if (8'h1f == _T_28[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_4;
      end else if (8'h1f == _T_25[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_3;
      end else if (8'h1f == _T_22[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_2;
      end else if (8'h1f == _T_19[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_1;
      end else if (8'h1f == _T_15[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_32 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h20 == _T_37[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_7;
      end else if (8'h20 == _T_34[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_6;
      end else if (8'h20 == _T_31[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_5;
      end else if (8'h20 == _T_28[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_4;
      end else if (8'h20 == _T_25[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_3;
      end else if (8'h20 == _T_22[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_2;
      end else if (8'h20 == _T_19[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_1;
      end else if (8'h20 == _T_15[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_33 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h21 == _T_37[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_7;
      end else if (8'h21 == _T_34[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_6;
      end else if (8'h21 == _T_31[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_5;
      end else if (8'h21 == _T_28[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_4;
      end else if (8'h21 == _T_25[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_3;
      end else if (8'h21 == _T_22[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_2;
      end else if (8'h21 == _T_19[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_1;
      end else if (8'h21 == _T_15[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_34 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h22 == _T_37[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_7;
      end else if (8'h22 == _T_34[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_6;
      end else if (8'h22 == _T_31[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_5;
      end else if (8'h22 == _T_28[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_4;
      end else if (8'h22 == _T_25[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_3;
      end else if (8'h22 == _T_22[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_2;
      end else if (8'h22 == _T_19[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_1;
      end else if (8'h22 == _T_15[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_35 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h23 == _T_37[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_7;
      end else if (8'h23 == _T_34[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_6;
      end else if (8'h23 == _T_31[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_5;
      end else if (8'h23 == _T_28[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_4;
      end else if (8'h23 == _T_25[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_3;
      end else if (8'h23 == _T_22[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_2;
      end else if (8'h23 == _T_19[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_1;
      end else if (8'h23 == _T_15[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_36 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h24 == _T_37[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_7;
      end else if (8'h24 == _T_34[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_6;
      end else if (8'h24 == _T_31[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_5;
      end else if (8'h24 == _T_28[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_4;
      end else if (8'h24 == _T_25[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_3;
      end else if (8'h24 == _T_22[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_2;
      end else if (8'h24 == _T_19[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_1;
      end else if (8'h24 == _T_15[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_37 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h25 == _T_37[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_7;
      end else if (8'h25 == _T_34[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_6;
      end else if (8'h25 == _T_31[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_5;
      end else if (8'h25 == _T_28[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_4;
      end else if (8'h25 == _T_25[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_3;
      end else if (8'h25 == _T_22[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_2;
      end else if (8'h25 == _T_19[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_1;
      end else if (8'h25 == _T_15[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_38 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h26 == _T_37[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_7;
      end else if (8'h26 == _T_34[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_6;
      end else if (8'h26 == _T_31[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_5;
      end else if (8'h26 == _T_28[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_4;
      end else if (8'h26 == _T_25[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_3;
      end else if (8'h26 == _T_22[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_2;
      end else if (8'h26 == _T_19[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_1;
      end else if (8'h26 == _T_15[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_39 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h27 == _T_37[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_7;
      end else if (8'h27 == _T_34[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_6;
      end else if (8'h27 == _T_31[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_5;
      end else if (8'h27 == _T_28[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_4;
      end else if (8'h27 == _T_25[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_3;
      end else if (8'h27 == _T_22[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_2;
      end else if (8'h27 == _T_19[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_1;
      end else if (8'h27 == _T_15[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_40 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h28 == _T_37[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_7;
      end else if (8'h28 == _T_34[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_6;
      end else if (8'h28 == _T_31[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_5;
      end else if (8'h28 == _T_28[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_4;
      end else if (8'h28 == _T_25[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_3;
      end else if (8'h28 == _T_22[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_2;
      end else if (8'h28 == _T_19[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_1;
      end else if (8'h28 == _T_15[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_41 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h29 == _T_37[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_7;
      end else if (8'h29 == _T_34[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_6;
      end else if (8'h29 == _T_31[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_5;
      end else if (8'h29 == _T_28[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_4;
      end else if (8'h29 == _T_25[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_3;
      end else if (8'h29 == _T_22[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_2;
      end else if (8'h29 == _T_19[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_1;
      end else if (8'h29 == _T_15[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_42 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2a == _T_37[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_7;
      end else if (8'h2a == _T_34[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_6;
      end else if (8'h2a == _T_31[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_5;
      end else if (8'h2a == _T_28[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_4;
      end else if (8'h2a == _T_25[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_3;
      end else if (8'h2a == _T_22[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_2;
      end else if (8'h2a == _T_19[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_1;
      end else if (8'h2a == _T_15[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_43 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2b == _T_37[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_7;
      end else if (8'h2b == _T_34[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_6;
      end else if (8'h2b == _T_31[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_5;
      end else if (8'h2b == _T_28[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_4;
      end else if (8'h2b == _T_25[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_3;
      end else if (8'h2b == _T_22[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_2;
      end else if (8'h2b == _T_19[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_1;
      end else if (8'h2b == _T_15[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_44 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2c == _T_37[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_7;
      end else if (8'h2c == _T_34[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_6;
      end else if (8'h2c == _T_31[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_5;
      end else if (8'h2c == _T_28[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_4;
      end else if (8'h2c == _T_25[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_3;
      end else if (8'h2c == _T_22[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_2;
      end else if (8'h2c == _T_19[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_1;
      end else if (8'h2c == _T_15[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_45 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2d == _T_37[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_7;
      end else if (8'h2d == _T_34[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_6;
      end else if (8'h2d == _T_31[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_5;
      end else if (8'h2d == _T_28[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_4;
      end else if (8'h2d == _T_25[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_3;
      end else if (8'h2d == _T_22[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_2;
      end else if (8'h2d == _T_19[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_1;
      end else if (8'h2d == _T_15[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_46 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2e == _T_37[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_7;
      end else if (8'h2e == _T_34[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_6;
      end else if (8'h2e == _T_31[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_5;
      end else if (8'h2e == _T_28[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_4;
      end else if (8'h2e == _T_25[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_3;
      end else if (8'h2e == _T_22[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_2;
      end else if (8'h2e == _T_19[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_1;
      end else if (8'h2e == _T_15[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_47 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2f == _T_37[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_7;
      end else if (8'h2f == _T_34[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_6;
      end else if (8'h2f == _T_31[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_5;
      end else if (8'h2f == _T_28[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_4;
      end else if (8'h2f == _T_25[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_3;
      end else if (8'h2f == _T_22[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_2;
      end else if (8'h2f == _T_19[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_1;
      end else if (8'h2f == _T_15[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_48 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h30 == _T_37[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_7;
      end else if (8'h30 == _T_34[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_6;
      end else if (8'h30 == _T_31[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_5;
      end else if (8'h30 == _T_28[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_4;
      end else if (8'h30 == _T_25[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_3;
      end else if (8'h30 == _T_22[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_2;
      end else if (8'h30 == _T_19[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_1;
      end else if (8'h30 == _T_15[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_49 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h31 == _T_37[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_7;
      end else if (8'h31 == _T_34[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_6;
      end else if (8'h31 == _T_31[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_5;
      end else if (8'h31 == _T_28[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_4;
      end else if (8'h31 == _T_25[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_3;
      end else if (8'h31 == _T_22[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_2;
      end else if (8'h31 == _T_19[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_1;
      end else if (8'h31 == _T_15[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_50 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h32 == _T_37[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_7;
      end else if (8'h32 == _T_34[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_6;
      end else if (8'h32 == _T_31[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_5;
      end else if (8'h32 == _T_28[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_4;
      end else if (8'h32 == _T_25[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_3;
      end else if (8'h32 == _T_22[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_2;
      end else if (8'h32 == _T_19[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_1;
      end else if (8'h32 == _T_15[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_51 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h33 == _T_37[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_7;
      end else if (8'h33 == _T_34[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_6;
      end else if (8'h33 == _T_31[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_5;
      end else if (8'h33 == _T_28[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_4;
      end else if (8'h33 == _T_25[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_3;
      end else if (8'h33 == _T_22[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_2;
      end else if (8'h33 == _T_19[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_1;
      end else if (8'h33 == _T_15[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_52 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h34 == _T_37[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_7;
      end else if (8'h34 == _T_34[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_6;
      end else if (8'h34 == _T_31[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_5;
      end else if (8'h34 == _T_28[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_4;
      end else if (8'h34 == _T_25[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_3;
      end else if (8'h34 == _T_22[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_2;
      end else if (8'h34 == _T_19[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_1;
      end else if (8'h34 == _T_15[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_53 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h35 == _T_37[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_7;
      end else if (8'h35 == _T_34[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_6;
      end else if (8'h35 == _T_31[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_5;
      end else if (8'h35 == _T_28[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_4;
      end else if (8'h35 == _T_25[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_3;
      end else if (8'h35 == _T_22[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_2;
      end else if (8'h35 == _T_19[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_1;
      end else if (8'h35 == _T_15[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_54 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h36 == _T_37[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_7;
      end else if (8'h36 == _T_34[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_6;
      end else if (8'h36 == _T_31[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_5;
      end else if (8'h36 == _T_28[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_4;
      end else if (8'h36 == _T_25[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_3;
      end else if (8'h36 == _T_22[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_2;
      end else if (8'h36 == _T_19[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_1;
      end else if (8'h36 == _T_15[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_55 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h37 == _T_37[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_7;
      end else if (8'h37 == _T_34[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_6;
      end else if (8'h37 == _T_31[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_5;
      end else if (8'h37 == _T_28[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_4;
      end else if (8'h37 == _T_25[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_3;
      end else if (8'h37 == _T_22[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_2;
      end else if (8'h37 == _T_19[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_1;
      end else if (8'h37 == _T_15[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_56 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h38 == _T_37[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_7;
      end else if (8'h38 == _T_34[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_6;
      end else if (8'h38 == _T_31[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_5;
      end else if (8'h38 == _T_28[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_4;
      end else if (8'h38 == _T_25[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_3;
      end else if (8'h38 == _T_22[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_2;
      end else if (8'h38 == _T_19[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_1;
      end else if (8'h38 == _T_15[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_57 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h39 == _T_37[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_7;
      end else if (8'h39 == _T_34[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_6;
      end else if (8'h39 == _T_31[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_5;
      end else if (8'h39 == _T_28[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_4;
      end else if (8'h39 == _T_25[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_3;
      end else if (8'h39 == _T_22[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_2;
      end else if (8'h39 == _T_19[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_1;
      end else if (8'h39 == _T_15[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_58 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3a == _T_37[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_7;
      end else if (8'h3a == _T_34[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_6;
      end else if (8'h3a == _T_31[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_5;
      end else if (8'h3a == _T_28[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_4;
      end else if (8'h3a == _T_25[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_3;
      end else if (8'h3a == _T_22[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_2;
      end else if (8'h3a == _T_19[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_1;
      end else if (8'h3a == _T_15[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_59 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3b == _T_37[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_7;
      end else if (8'h3b == _T_34[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_6;
      end else if (8'h3b == _T_31[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_5;
      end else if (8'h3b == _T_28[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_4;
      end else if (8'h3b == _T_25[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_3;
      end else if (8'h3b == _T_22[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_2;
      end else if (8'h3b == _T_19[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_1;
      end else if (8'h3b == _T_15[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_60 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3c == _T_37[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_7;
      end else if (8'h3c == _T_34[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_6;
      end else if (8'h3c == _T_31[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_5;
      end else if (8'h3c == _T_28[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_4;
      end else if (8'h3c == _T_25[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_3;
      end else if (8'h3c == _T_22[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_2;
      end else if (8'h3c == _T_19[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_1;
      end else if (8'h3c == _T_15[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_61 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3d == _T_37[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_7;
      end else if (8'h3d == _T_34[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_6;
      end else if (8'h3d == _T_31[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_5;
      end else if (8'h3d == _T_28[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_4;
      end else if (8'h3d == _T_25[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_3;
      end else if (8'h3d == _T_22[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_2;
      end else if (8'h3d == _T_19[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_1;
      end else if (8'h3d == _T_15[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_62 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3e == _T_37[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_7;
      end else if (8'h3e == _T_34[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_6;
      end else if (8'h3e == _T_31[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_5;
      end else if (8'h3e == _T_28[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_4;
      end else if (8'h3e == _T_25[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_3;
      end else if (8'h3e == _T_22[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_2;
      end else if (8'h3e == _T_19[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_1;
      end else if (8'h3e == _T_15[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_63 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3f == _T_37[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_7;
      end else if (8'h3f == _T_34[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_6;
      end else if (8'h3f == _T_31[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_5;
      end else if (8'h3f == _T_28[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_4;
      end else if (8'h3f == _T_25[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_3;
      end else if (8'h3f == _T_22[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_2;
      end else if (8'h3f == _T_19[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_1;
      end else if (8'h3f == _T_15[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_64 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h40 == _T_37[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_7;
      end else if (8'h40 == _T_34[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_6;
      end else if (8'h40 == _T_31[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_5;
      end else if (8'h40 == _T_28[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_4;
      end else if (8'h40 == _T_25[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_3;
      end else if (8'h40 == _T_22[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_2;
      end else if (8'h40 == _T_19[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_1;
      end else if (8'h40 == _T_15[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_65 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h41 == _T_37[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_7;
      end else if (8'h41 == _T_34[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_6;
      end else if (8'h41 == _T_31[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_5;
      end else if (8'h41 == _T_28[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_4;
      end else if (8'h41 == _T_25[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_3;
      end else if (8'h41 == _T_22[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_2;
      end else if (8'h41 == _T_19[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_1;
      end else if (8'h41 == _T_15[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_66 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h42 == _T_37[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_7;
      end else if (8'h42 == _T_34[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_6;
      end else if (8'h42 == _T_31[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_5;
      end else if (8'h42 == _T_28[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_4;
      end else if (8'h42 == _T_25[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_3;
      end else if (8'h42 == _T_22[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_2;
      end else if (8'h42 == _T_19[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_1;
      end else if (8'h42 == _T_15[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_67 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h43 == _T_37[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_7;
      end else if (8'h43 == _T_34[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_6;
      end else if (8'h43 == _T_31[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_5;
      end else if (8'h43 == _T_28[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_4;
      end else if (8'h43 == _T_25[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_3;
      end else if (8'h43 == _T_22[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_2;
      end else if (8'h43 == _T_19[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_1;
      end else if (8'h43 == _T_15[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_68 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h44 == _T_37[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_7;
      end else if (8'h44 == _T_34[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_6;
      end else if (8'h44 == _T_31[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_5;
      end else if (8'h44 == _T_28[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_4;
      end else if (8'h44 == _T_25[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_3;
      end else if (8'h44 == _T_22[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_2;
      end else if (8'h44 == _T_19[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_1;
      end else if (8'h44 == _T_15[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_69 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h45 == _T_37[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_7;
      end else if (8'h45 == _T_34[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_6;
      end else if (8'h45 == _T_31[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_5;
      end else if (8'h45 == _T_28[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_4;
      end else if (8'h45 == _T_25[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_3;
      end else if (8'h45 == _T_22[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_2;
      end else if (8'h45 == _T_19[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_1;
      end else if (8'h45 == _T_15[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_70 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h46 == _T_37[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_7;
      end else if (8'h46 == _T_34[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_6;
      end else if (8'h46 == _T_31[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_5;
      end else if (8'h46 == _T_28[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_4;
      end else if (8'h46 == _T_25[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_3;
      end else if (8'h46 == _T_22[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_2;
      end else if (8'h46 == _T_19[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_1;
      end else if (8'h46 == _T_15[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_71 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h47 == _T_37[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_7;
      end else if (8'h47 == _T_34[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_6;
      end else if (8'h47 == _T_31[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_5;
      end else if (8'h47 == _T_28[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_4;
      end else if (8'h47 == _T_25[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_3;
      end else if (8'h47 == _T_22[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_2;
      end else if (8'h47 == _T_19[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_1;
      end else if (8'h47 == _T_15[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_72 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h48 == _T_37[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_7;
      end else if (8'h48 == _T_34[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_6;
      end else if (8'h48 == _T_31[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_5;
      end else if (8'h48 == _T_28[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_4;
      end else if (8'h48 == _T_25[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_3;
      end else if (8'h48 == _T_22[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_2;
      end else if (8'h48 == _T_19[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_1;
      end else if (8'h48 == _T_15[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_73 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h49 == _T_37[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_7;
      end else if (8'h49 == _T_34[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_6;
      end else if (8'h49 == _T_31[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_5;
      end else if (8'h49 == _T_28[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_4;
      end else if (8'h49 == _T_25[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_3;
      end else if (8'h49 == _T_22[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_2;
      end else if (8'h49 == _T_19[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_1;
      end else if (8'h49 == _T_15[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_74 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4a == _T_37[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_7;
      end else if (8'h4a == _T_34[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_6;
      end else if (8'h4a == _T_31[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_5;
      end else if (8'h4a == _T_28[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_4;
      end else if (8'h4a == _T_25[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_3;
      end else if (8'h4a == _T_22[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_2;
      end else if (8'h4a == _T_19[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_1;
      end else if (8'h4a == _T_15[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_75 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4b == _T_37[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_7;
      end else if (8'h4b == _T_34[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_6;
      end else if (8'h4b == _T_31[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_5;
      end else if (8'h4b == _T_28[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_4;
      end else if (8'h4b == _T_25[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_3;
      end else if (8'h4b == _T_22[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_2;
      end else if (8'h4b == _T_19[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_1;
      end else if (8'h4b == _T_15[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_76 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4c == _T_37[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_7;
      end else if (8'h4c == _T_34[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_6;
      end else if (8'h4c == _T_31[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_5;
      end else if (8'h4c == _T_28[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_4;
      end else if (8'h4c == _T_25[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_3;
      end else if (8'h4c == _T_22[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_2;
      end else if (8'h4c == _T_19[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_1;
      end else if (8'h4c == _T_15[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_77 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4d == _T_37[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_7;
      end else if (8'h4d == _T_34[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_6;
      end else if (8'h4d == _T_31[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_5;
      end else if (8'h4d == _T_28[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_4;
      end else if (8'h4d == _T_25[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_3;
      end else if (8'h4d == _T_22[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_2;
      end else if (8'h4d == _T_19[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_1;
      end else if (8'h4d == _T_15[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_78 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4e == _T_37[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_7;
      end else if (8'h4e == _T_34[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_6;
      end else if (8'h4e == _T_31[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_5;
      end else if (8'h4e == _T_28[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_4;
      end else if (8'h4e == _T_25[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_3;
      end else if (8'h4e == _T_22[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_2;
      end else if (8'h4e == _T_19[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_1;
      end else if (8'h4e == _T_15[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_79 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4f == _T_37[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_7;
      end else if (8'h4f == _T_34[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_6;
      end else if (8'h4f == _T_31[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_5;
      end else if (8'h4f == _T_28[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_4;
      end else if (8'h4f == _T_25[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_3;
      end else if (8'h4f == _T_22[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_2;
      end else if (8'h4f == _T_19[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_1;
      end else if (8'h4f == _T_15[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_80 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h50 == _T_37[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_7;
      end else if (8'h50 == _T_34[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_6;
      end else if (8'h50 == _T_31[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_5;
      end else if (8'h50 == _T_28[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_4;
      end else if (8'h50 == _T_25[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_3;
      end else if (8'h50 == _T_22[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_2;
      end else if (8'h50 == _T_19[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_1;
      end else if (8'h50 == _T_15[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_81 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h51 == _T_37[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_7;
      end else if (8'h51 == _T_34[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_6;
      end else if (8'h51 == _T_31[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_5;
      end else if (8'h51 == _T_28[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_4;
      end else if (8'h51 == _T_25[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_3;
      end else if (8'h51 == _T_22[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_2;
      end else if (8'h51 == _T_19[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_1;
      end else if (8'h51 == _T_15[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_82 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h52 == _T_37[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_7;
      end else if (8'h52 == _T_34[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_6;
      end else if (8'h52 == _T_31[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_5;
      end else if (8'h52 == _T_28[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_4;
      end else if (8'h52 == _T_25[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_3;
      end else if (8'h52 == _T_22[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_2;
      end else if (8'h52 == _T_19[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_1;
      end else if (8'h52 == _T_15[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_83 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h53 == _T_37[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_7;
      end else if (8'h53 == _T_34[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_6;
      end else if (8'h53 == _T_31[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_5;
      end else if (8'h53 == _T_28[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_4;
      end else if (8'h53 == _T_25[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_3;
      end else if (8'h53 == _T_22[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_2;
      end else if (8'h53 == _T_19[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_1;
      end else if (8'h53 == _T_15[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_84 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h54 == _T_37[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_7;
      end else if (8'h54 == _T_34[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_6;
      end else if (8'h54 == _T_31[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_5;
      end else if (8'h54 == _T_28[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_4;
      end else if (8'h54 == _T_25[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_3;
      end else if (8'h54 == _T_22[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_2;
      end else if (8'h54 == _T_19[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_1;
      end else if (8'h54 == _T_15[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_85 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h55 == _T_37[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_7;
      end else if (8'h55 == _T_34[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_6;
      end else if (8'h55 == _T_31[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_5;
      end else if (8'h55 == _T_28[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_4;
      end else if (8'h55 == _T_25[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_3;
      end else if (8'h55 == _T_22[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_2;
      end else if (8'h55 == _T_19[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_1;
      end else if (8'h55 == _T_15[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_86 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h56 == _T_37[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_7;
      end else if (8'h56 == _T_34[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_6;
      end else if (8'h56 == _T_31[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_5;
      end else if (8'h56 == _T_28[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_4;
      end else if (8'h56 == _T_25[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_3;
      end else if (8'h56 == _T_22[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_2;
      end else if (8'h56 == _T_19[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_1;
      end else if (8'h56 == _T_15[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_87 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h57 == _T_37[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_7;
      end else if (8'h57 == _T_34[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_6;
      end else if (8'h57 == _T_31[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_5;
      end else if (8'h57 == _T_28[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_4;
      end else if (8'h57 == _T_25[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_3;
      end else if (8'h57 == _T_22[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_2;
      end else if (8'h57 == _T_19[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_1;
      end else if (8'h57 == _T_15[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_88 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h58 == _T_37[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_7;
      end else if (8'h58 == _T_34[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_6;
      end else if (8'h58 == _T_31[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_5;
      end else if (8'h58 == _T_28[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_4;
      end else if (8'h58 == _T_25[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_3;
      end else if (8'h58 == _T_22[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_2;
      end else if (8'h58 == _T_19[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_1;
      end else if (8'h58 == _T_15[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_89 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h59 == _T_37[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_7;
      end else if (8'h59 == _T_34[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_6;
      end else if (8'h59 == _T_31[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_5;
      end else if (8'h59 == _T_28[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_4;
      end else if (8'h59 == _T_25[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_3;
      end else if (8'h59 == _T_22[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_2;
      end else if (8'h59 == _T_19[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_1;
      end else if (8'h59 == _T_15[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_90 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5a == _T_37[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_7;
      end else if (8'h5a == _T_34[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_6;
      end else if (8'h5a == _T_31[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_5;
      end else if (8'h5a == _T_28[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_4;
      end else if (8'h5a == _T_25[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_3;
      end else if (8'h5a == _T_22[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_2;
      end else if (8'h5a == _T_19[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_1;
      end else if (8'h5a == _T_15[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_91 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5b == _T_37[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_7;
      end else if (8'h5b == _T_34[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_6;
      end else if (8'h5b == _T_31[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_5;
      end else if (8'h5b == _T_28[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_4;
      end else if (8'h5b == _T_25[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_3;
      end else if (8'h5b == _T_22[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_2;
      end else if (8'h5b == _T_19[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_1;
      end else if (8'h5b == _T_15[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_92 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5c == _T_37[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_7;
      end else if (8'h5c == _T_34[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_6;
      end else if (8'h5c == _T_31[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_5;
      end else if (8'h5c == _T_28[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_4;
      end else if (8'h5c == _T_25[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_3;
      end else if (8'h5c == _T_22[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_2;
      end else if (8'h5c == _T_19[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_1;
      end else if (8'h5c == _T_15[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_93 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5d == _T_37[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_7;
      end else if (8'h5d == _T_34[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_6;
      end else if (8'h5d == _T_31[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_5;
      end else if (8'h5d == _T_28[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_4;
      end else if (8'h5d == _T_25[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_3;
      end else if (8'h5d == _T_22[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_2;
      end else if (8'h5d == _T_19[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_1;
      end else if (8'h5d == _T_15[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_94 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5e == _T_37[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_7;
      end else if (8'h5e == _T_34[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_6;
      end else if (8'h5e == _T_31[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_5;
      end else if (8'h5e == _T_28[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_4;
      end else if (8'h5e == _T_25[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_3;
      end else if (8'h5e == _T_22[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_2;
      end else if (8'h5e == _T_19[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_1;
      end else if (8'h5e == _T_15[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_95 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5f == _T_37[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_7;
      end else if (8'h5f == _T_34[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_6;
      end else if (8'h5f == _T_31[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_5;
      end else if (8'h5f == _T_28[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_4;
      end else if (8'h5f == _T_25[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_3;
      end else if (8'h5f == _T_22[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_2;
      end else if (8'h5f == _T_19[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_1;
      end else if (8'h5f == _T_15[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_96 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h60 == _T_37[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_7;
      end else if (8'h60 == _T_34[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_6;
      end else if (8'h60 == _T_31[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_5;
      end else if (8'h60 == _T_28[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_4;
      end else if (8'h60 == _T_25[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_3;
      end else if (8'h60 == _T_22[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_2;
      end else if (8'h60 == _T_19[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_1;
      end else if (8'h60 == _T_15[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_97 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h61 == _T_37[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_7;
      end else if (8'h61 == _T_34[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_6;
      end else if (8'h61 == _T_31[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_5;
      end else if (8'h61 == _T_28[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_4;
      end else if (8'h61 == _T_25[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_3;
      end else if (8'h61 == _T_22[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_2;
      end else if (8'h61 == _T_19[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_1;
      end else if (8'h61 == _T_15[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_98 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h62 == _T_37[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_7;
      end else if (8'h62 == _T_34[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_6;
      end else if (8'h62 == _T_31[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_5;
      end else if (8'h62 == _T_28[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_4;
      end else if (8'h62 == _T_25[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_3;
      end else if (8'h62 == _T_22[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_2;
      end else if (8'h62 == _T_19[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_1;
      end else if (8'h62 == _T_15[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_99 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h63 == _T_37[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_7;
      end else if (8'h63 == _T_34[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_6;
      end else if (8'h63 == _T_31[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_5;
      end else if (8'h63 == _T_28[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_4;
      end else if (8'h63 == _T_25[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_3;
      end else if (8'h63 == _T_22[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_2;
      end else if (8'h63 == _T_19[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_1;
      end else if (8'h63 == _T_15[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_100 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h64 == _T_37[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_7;
      end else if (8'h64 == _T_34[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_6;
      end else if (8'h64 == _T_31[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_5;
      end else if (8'h64 == _T_28[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_4;
      end else if (8'h64 == _T_25[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_3;
      end else if (8'h64 == _T_22[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_2;
      end else if (8'h64 == _T_19[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_1;
      end else if (8'h64 == _T_15[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_101 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h65 == _T_37[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_7;
      end else if (8'h65 == _T_34[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_6;
      end else if (8'h65 == _T_31[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_5;
      end else if (8'h65 == _T_28[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_4;
      end else if (8'h65 == _T_25[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_3;
      end else if (8'h65 == _T_22[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_2;
      end else if (8'h65 == _T_19[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_1;
      end else if (8'h65 == _T_15[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_102 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h66 == _T_37[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_7;
      end else if (8'h66 == _T_34[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_6;
      end else if (8'h66 == _T_31[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_5;
      end else if (8'h66 == _T_28[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_4;
      end else if (8'h66 == _T_25[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_3;
      end else if (8'h66 == _T_22[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_2;
      end else if (8'h66 == _T_19[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_1;
      end else if (8'h66 == _T_15[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_103 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h67 == _T_37[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_7;
      end else if (8'h67 == _T_34[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_6;
      end else if (8'h67 == _T_31[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_5;
      end else if (8'h67 == _T_28[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_4;
      end else if (8'h67 == _T_25[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_3;
      end else if (8'h67 == _T_22[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_2;
      end else if (8'h67 == _T_19[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_1;
      end else if (8'h67 == _T_15[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_104 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h68 == _T_37[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_7;
      end else if (8'h68 == _T_34[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_6;
      end else if (8'h68 == _T_31[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_5;
      end else if (8'h68 == _T_28[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_4;
      end else if (8'h68 == _T_25[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_3;
      end else if (8'h68 == _T_22[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_2;
      end else if (8'h68 == _T_19[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_1;
      end else if (8'h68 == _T_15[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_105 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h69 == _T_37[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_7;
      end else if (8'h69 == _T_34[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_6;
      end else if (8'h69 == _T_31[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_5;
      end else if (8'h69 == _T_28[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_4;
      end else if (8'h69 == _T_25[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_3;
      end else if (8'h69 == _T_22[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_2;
      end else if (8'h69 == _T_19[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_1;
      end else if (8'h69 == _T_15[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_106 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6a == _T_37[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_7;
      end else if (8'h6a == _T_34[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_6;
      end else if (8'h6a == _T_31[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_5;
      end else if (8'h6a == _T_28[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_4;
      end else if (8'h6a == _T_25[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_3;
      end else if (8'h6a == _T_22[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_2;
      end else if (8'h6a == _T_19[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_1;
      end else if (8'h6a == _T_15[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_107 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6b == _T_37[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_7;
      end else if (8'h6b == _T_34[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_6;
      end else if (8'h6b == _T_31[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_5;
      end else if (8'h6b == _T_28[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_4;
      end else if (8'h6b == _T_25[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_3;
      end else if (8'h6b == _T_22[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_2;
      end else if (8'h6b == _T_19[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_1;
      end else if (8'h6b == _T_15[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_108 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6c == _T_37[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_7;
      end else if (8'h6c == _T_34[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_6;
      end else if (8'h6c == _T_31[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_5;
      end else if (8'h6c == _T_28[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_4;
      end else if (8'h6c == _T_25[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_3;
      end else if (8'h6c == _T_22[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_2;
      end else if (8'h6c == _T_19[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_1;
      end else if (8'h6c == _T_15[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_109 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6d == _T_37[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_7;
      end else if (8'h6d == _T_34[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_6;
      end else if (8'h6d == _T_31[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_5;
      end else if (8'h6d == _T_28[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_4;
      end else if (8'h6d == _T_25[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_3;
      end else if (8'h6d == _T_22[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_2;
      end else if (8'h6d == _T_19[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_1;
      end else if (8'h6d == _T_15[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_110 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6e == _T_37[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_7;
      end else if (8'h6e == _T_34[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_6;
      end else if (8'h6e == _T_31[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_5;
      end else if (8'h6e == _T_28[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_4;
      end else if (8'h6e == _T_25[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_3;
      end else if (8'h6e == _T_22[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_2;
      end else if (8'h6e == _T_19[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_1;
      end else if (8'h6e == _T_15[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_111 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6f == _T_37[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_7;
      end else if (8'h6f == _T_34[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_6;
      end else if (8'h6f == _T_31[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_5;
      end else if (8'h6f == _T_28[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_4;
      end else if (8'h6f == _T_25[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_3;
      end else if (8'h6f == _T_22[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_2;
      end else if (8'h6f == _T_19[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_1;
      end else if (8'h6f == _T_15[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_112 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h70 == _T_37[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_7;
      end else if (8'h70 == _T_34[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_6;
      end else if (8'h70 == _T_31[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_5;
      end else if (8'h70 == _T_28[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_4;
      end else if (8'h70 == _T_25[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_3;
      end else if (8'h70 == _T_22[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_2;
      end else if (8'h70 == _T_19[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_1;
      end else if (8'h70 == _T_15[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_113 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h71 == _T_37[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_7;
      end else if (8'h71 == _T_34[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_6;
      end else if (8'h71 == _T_31[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_5;
      end else if (8'h71 == _T_28[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_4;
      end else if (8'h71 == _T_25[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_3;
      end else if (8'h71 == _T_22[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_2;
      end else if (8'h71 == _T_19[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_1;
      end else if (8'h71 == _T_15[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_114 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h72 == _T_37[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_7;
      end else if (8'h72 == _T_34[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_6;
      end else if (8'h72 == _T_31[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_5;
      end else if (8'h72 == _T_28[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_4;
      end else if (8'h72 == _T_25[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_3;
      end else if (8'h72 == _T_22[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_2;
      end else if (8'h72 == _T_19[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_1;
      end else if (8'h72 == _T_15[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_115 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h73 == _T_37[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_7;
      end else if (8'h73 == _T_34[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_6;
      end else if (8'h73 == _T_31[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_5;
      end else if (8'h73 == _T_28[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_4;
      end else if (8'h73 == _T_25[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_3;
      end else if (8'h73 == _T_22[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_2;
      end else if (8'h73 == _T_19[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_1;
      end else if (8'h73 == _T_15[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_116 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h74 == _T_37[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_7;
      end else if (8'h74 == _T_34[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_6;
      end else if (8'h74 == _T_31[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_5;
      end else if (8'h74 == _T_28[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_4;
      end else if (8'h74 == _T_25[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_3;
      end else if (8'h74 == _T_22[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_2;
      end else if (8'h74 == _T_19[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_1;
      end else if (8'h74 == _T_15[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_117 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h75 == _T_37[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_7;
      end else if (8'h75 == _T_34[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_6;
      end else if (8'h75 == _T_31[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_5;
      end else if (8'h75 == _T_28[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_4;
      end else if (8'h75 == _T_25[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_3;
      end else if (8'h75 == _T_22[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_2;
      end else if (8'h75 == _T_19[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_1;
      end else if (8'h75 == _T_15[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_118 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h76 == _T_37[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_7;
      end else if (8'h76 == _T_34[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_6;
      end else if (8'h76 == _T_31[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_5;
      end else if (8'h76 == _T_28[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_4;
      end else if (8'h76 == _T_25[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_3;
      end else if (8'h76 == _T_22[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_2;
      end else if (8'h76 == _T_19[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_1;
      end else if (8'h76 == _T_15[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_119 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h77 == _T_37[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_7;
      end else if (8'h77 == _T_34[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_6;
      end else if (8'h77 == _T_31[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_5;
      end else if (8'h77 == _T_28[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_4;
      end else if (8'h77 == _T_25[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_3;
      end else if (8'h77 == _T_22[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_2;
      end else if (8'h77 == _T_19[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_1;
      end else if (8'h77 == _T_15[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_120 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h78 == _T_37[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_7;
      end else if (8'h78 == _T_34[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_6;
      end else if (8'h78 == _T_31[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_5;
      end else if (8'h78 == _T_28[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_4;
      end else if (8'h78 == _T_25[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_3;
      end else if (8'h78 == _T_22[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_2;
      end else if (8'h78 == _T_19[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_1;
      end else if (8'h78 == _T_15[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_121 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h79 == _T_37[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_7;
      end else if (8'h79 == _T_34[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_6;
      end else if (8'h79 == _T_31[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_5;
      end else if (8'h79 == _T_28[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_4;
      end else if (8'h79 == _T_25[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_3;
      end else if (8'h79 == _T_22[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_2;
      end else if (8'h79 == _T_19[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_1;
      end else if (8'h79 == _T_15[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_122 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7a == _T_37[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_7;
      end else if (8'h7a == _T_34[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_6;
      end else if (8'h7a == _T_31[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_5;
      end else if (8'h7a == _T_28[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_4;
      end else if (8'h7a == _T_25[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_3;
      end else if (8'h7a == _T_22[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_2;
      end else if (8'h7a == _T_19[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_1;
      end else if (8'h7a == _T_15[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_123 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7b == _T_37[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_7;
      end else if (8'h7b == _T_34[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_6;
      end else if (8'h7b == _T_31[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_5;
      end else if (8'h7b == _T_28[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_4;
      end else if (8'h7b == _T_25[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_3;
      end else if (8'h7b == _T_22[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_2;
      end else if (8'h7b == _T_19[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_1;
      end else if (8'h7b == _T_15[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_124 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7c == _T_37[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_7;
      end else if (8'h7c == _T_34[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_6;
      end else if (8'h7c == _T_31[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_5;
      end else if (8'h7c == _T_28[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_4;
      end else if (8'h7c == _T_25[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_3;
      end else if (8'h7c == _T_22[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_2;
      end else if (8'h7c == _T_19[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_1;
      end else if (8'h7c == _T_15[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_125 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7d == _T_37[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_7;
      end else if (8'h7d == _T_34[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_6;
      end else if (8'h7d == _T_31[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_5;
      end else if (8'h7d == _T_28[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_4;
      end else if (8'h7d == _T_25[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_3;
      end else if (8'h7d == _T_22[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_2;
      end else if (8'h7d == _T_19[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_1;
      end else if (8'h7d == _T_15[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_126 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7e == _T_37[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_7;
      end else if (8'h7e == _T_34[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_6;
      end else if (8'h7e == _T_31[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_5;
      end else if (8'h7e == _T_28[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_4;
      end else if (8'h7e == _T_25[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_3;
      end else if (8'h7e == _T_22[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_2;
      end else if (8'h7e == _T_19[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_1;
      end else if (8'h7e == _T_15[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_127 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7f == _T_37[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_7;
      end else if (8'h7f == _T_34[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_6;
      end else if (8'h7f == _T_31[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_5;
      end else if (8'h7f == _T_28[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_4;
      end else if (8'h7f == _T_25[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_3;
      end else if (8'h7f == _T_22[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_2;
      end else if (8'h7f == _T_19[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_1;
      end else if (8'h7f == _T_15[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_128 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h80 == _T_37[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_7;
      end else if (8'h80 == _T_34[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_6;
      end else if (8'h80 == _T_31[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_5;
      end else if (8'h80 == _T_28[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_4;
      end else if (8'h80 == _T_25[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_3;
      end else if (8'h80 == _T_22[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_2;
      end else if (8'h80 == _T_19[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_1;
      end else if (8'h80 == _T_15[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_129 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h81 == _T_37[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_7;
      end else if (8'h81 == _T_34[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_6;
      end else if (8'h81 == _T_31[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_5;
      end else if (8'h81 == _T_28[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_4;
      end else if (8'h81 == _T_25[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_3;
      end else if (8'h81 == _T_22[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_2;
      end else if (8'h81 == _T_19[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_1;
      end else if (8'h81 == _T_15[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_130 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h82 == _T_37[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_7;
      end else if (8'h82 == _T_34[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_6;
      end else if (8'h82 == _T_31[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_5;
      end else if (8'h82 == _T_28[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_4;
      end else if (8'h82 == _T_25[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_3;
      end else if (8'h82 == _T_22[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_2;
      end else if (8'h82 == _T_19[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_1;
      end else if (8'h82 == _T_15[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_131 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h83 == _T_37[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_7;
      end else if (8'h83 == _T_34[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_6;
      end else if (8'h83 == _T_31[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_5;
      end else if (8'h83 == _T_28[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_4;
      end else if (8'h83 == _T_25[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_3;
      end else if (8'h83 == _T_22[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_2;
      end else if (8'h83 == _T_19[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_1;
      end else if (8'h83 == _T_15[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_132 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h84 == _T_37[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_7;
      end else if (8'h84 == _T_34[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_6;
      end else if (8'h84 == _T_31[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_5;
      end else if (8'h84 == _T_28[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_4;
      end else if (8'h84 == _T_25[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_3;
      end else if (8'h84 == _T_22[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_2;
      end else if (8'h84 == _T_19[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_1;
      end else if (8'h84 == _T_15[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_133 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h85 == _T_37[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_7;
      end else if (8'h85 == _T_34[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_6;
      end else if (8'h85 == _T_31[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_5;
      end else if (8'h85 == _T_28[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_4;
      end else if (8'h85 == _T_25[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_3;
      end else if (8'h85 == _T_22[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_2;
      end else if (8'h85 == _T_19[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_1;
      end else if (8'h85 == _T_15[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_134 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h86 == _T_37[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_7;
      end else if (8'h86 == _T_34[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_6;
      end else if (8'h86 == _T_31[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_5;
      end else if (8'h86 == _T_28[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_4;
      end else if (8'h86 == _T_25[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_3;
      end else if (8'h86 == _T_22[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_2;
      end else if (8'h86 == _T_19[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_1;
      end else if (8'h86 == _T_15[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_135 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h87 == _T_37[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_7;
      end else if (8'h87 == _T_34[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_6;
      end else if (8'h87 == _T_31[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_5;
      end else if (8'h87 == _T_28[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_4;
      end else if (8'h87 == _T_25[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_3;
      end else if (8'h87 == _T_22[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_2;
      end else if (8'h87 == _T_19[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_1;
      end else if (8'h87 == _T_15[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_136 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h88 == _T_37[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_7;
      end else if (8'h88 == _T_34[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_6;
      end else if (8'h88 == _T_31[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_5;
      end else if (8'h88 == _T_28[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_4;
      end else if (8'h88 == _T_25[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_3;
      end else if (8'h88 == _T_22[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_2;
      end else if (8'h88 == _T_19[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_1;
      end else if (8'h88 == _T_15[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_137 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h89 == _T_37[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_7;
      end else if (8'h89 == _T_34[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_6;
      end else if (8'h89 == _T_31[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_5;
      end else if (8'h89 == _T_28[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_4;
      end else if (8'h89 == _T_25[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_3;
      end else if (8'h89 == _T_22[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_2;
      end else if (8'h89 == _T_19[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_1;
      end else if (8'h89 == _T_15[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_138 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8a == _T_37[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_7;
      end else if (8'h8a == _T_34[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_6;
      end else if (8'h8a == _T_31[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_5;
      end else if (8'h8a == _T_28[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_4;
      end else if (8'h8a == _T_25[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_3;
      end else if (8'h8a == _T_22[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_2;
      end else if (8'h8a == _T_19[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_1;
      end else if (8'h8a == _T_15[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_139 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8b == _T_37[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_7;
      end else if (8'h8b == _T_34[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_6;
      end else if (8'h8b == _T_31[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_5;
      end else if (8'h8b == _T_28[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_4;
      end else if (8'h8b == _T_25[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_3;
      end else if (8'h8b == _T_22[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_2;
      end else if (8'h8b == _T_19[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_1;
      end else if (8'h8b == _T_15[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_140 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8c == _T_37[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_7;
      end else if (8'h8c == _T_34[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_6;
      end else if (8'h8c == _T_31[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_5;
      end else if (8'h8c == _T_28[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_4;
      end else if (8'h8c == _T_25[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_3;
      end else if (8'h8c == _T_22[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_2;
      end else if (8'h8c == _T_19[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_1;
      end else if (8'h8c == _T_15[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_141 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8d == _T_37[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_7;
      end else if (8'h8d == _T_34[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_6;
      end else if (8'h8d == _T_31[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_5;
      end else if (8'h8d == _T_28[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_4;
      end else if (8'h8d == _T_25[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_3;
      end else if (8'h8d == _T_22[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_2;
      end else if (8'h8d == _T_19[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_1;
      end else if (8'h8d == _T_15[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_142 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8e == _T_37[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_7;
      end else if (8'h8e == _T_34[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_6;
      end else if (8'h8e == _T_31[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_5;
      end else if (8'h8e == _T_28[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_4;
      end else if (8'h8e == _T_25[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_3;
      end else if (8'h8e == _T_22[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_2;
      end else if (8'h8e == _T_19[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_1;
      end else if (8'h8e == _T_15[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_143 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8f == _T_37[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_7;
      end else if (8'h8f == _T_34[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_6;
      end else if (8'h8f == _T_31[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_5;
      end else if (8'h8f == _T_28[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_4;
      end else if (8'h8f == _T_25[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_3;
      end else if (8'h8f == _T_22[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_2;
      end else if (8'h8f == _T_19[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_1;
      end else if (8'h8f == _T_15[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      pixelIndex <= 32'h0;
    end else if (io_valid_in) begin
      if (_T_90) begin
        pixelIndex <= 32'h0;
      end else begin
        pixelIndex <= _T_88;
      end
    end
  end
endmodule
module ImageProcessing(
  input         clock,
  input         reset,
  input  [5:0]  io_SPI_filterIndex,
  input         io_SPI_invert,
  input         io_SPI_distort,
  input  [10:0] io_rowIndex,
  input  [10:0] io_colIndex,
  output [3:0]  io_pixelVal_out_0,
  output [3:0]  io_pixelVal_out_1,
  output [3:0]  io_pixelVal_out_2
);
  wire  filter_clock; // @[ImageProcessing.scala 23:22]
  wire  filter_reset; // @[ImageProcessing.scala 23:22]
  wire [5:0] filter_io_SPI_filterIndex; // @[ImageProcessing.scala 23:22]
  wire  filter_io_SPI_distort; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_0; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_1; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_2; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_3; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_4; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_5; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_6; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_7; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_0; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_1; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_2; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_3; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_4; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_5; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_6; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_7; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_0; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_1; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_2; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_3; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_4; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_5; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_6; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_7; // @[ImageProcessing.scala 23:22]
  wire  filter_io_valid_out; // @[ImageProcessing.scala 23:22]
  wire  videoBuffer_clock; // @[ImageProcessing.scala 24:27]
  wire  videoBuffer_reset; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_0; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_1; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_2; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_3; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_4; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_5; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_6; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_7; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_0; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_1; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_2; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_3; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_4; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_5; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_6; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_7; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_0; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_1; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_2; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_3; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_4; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_5; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_6; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_7; // @[ImageProcessing.scala 24:27]
  wire  videoBuffer_io_valid_in; // @[ImageProcessing.scala 24:27]
  wire [10:0] videoBuffer_io_rowIndex; // @[ImageProcessing.scala 24:27]
  wire [10:0] videoBuffer_io_colIndex; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_out_0; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_out_1; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_out_2; // @[ImageProcessing.scala 24:27]
  Filter filter ( // @[ImageProcessing.scala 23:22]
    .clock(filter_clock),
    .reset(filter_reset),
    .io_SPI_filterIndex(filter_io_SPI_filterIndex),
    .io_SPI_distort(filter_io_SPI_distort),
    .io_pixelVal_out_0_0(filter_io_pixelVal_out_0_0),
    .io_pixelVal_out_0_1(filter_io_pixelVal_out_0_1),
    .io_pixelVal_out_0_2(filter_io_pixelVal_out_0_2),
    .io_pixelVal_out_0_3(filter_io_pixelVal_out_0_3),
    .io_pixelVal_out_0_4(filter_io_pixelVal_out_0_4),
    .io_pixelVal_out_0_5(filter_io_pixelVal_out_0_5),
    .io_pixelVal_out_0_6(filter_io_pixelVal_out_0_6),
    .io_pixelVal_out_0_7(filter_io_pixelVal_out_0_7),
    .io_pixelVal_out_1_0(filter_io_pixelVal_out_1_0),
    .io_pixelVal_out_1_1(filter_io_pixelVal_out_1_1),
    .io_pixelVal_out_1_2(filter_io_pixelVal_out_1_2),
    .io_pixelVal_out_1_3(filter_io_pixelVal_out_1_3),
    .io_pixelVal_out_1_4(filter_io_pixelVal_out_1_4),
    .io_pixelVal_out_1_5(filter_io_pixelVal_out_1_5),
    .io_pixelVal_out_1_6(filter_io_pixelVal_out_1_6),
    .io_pixelVal_out_1_7(filter_io_pixelVal_out_1_7),
    .io_pixelVal_out_2_0(filter_io_pixelVal_out_2_0),
    .io_pixelVal_out_2_1(filter_io_pixelVal_out_2_1),
    .io_pixelVal_out_2_2(filter_io_pixelVal_out_2_2),
    .io_pixelVal_out_2_3(filter_io_pixelVal_out_2_3),
    .io_pixelVal_out_2_4(filter_io_pixelVal_out_2_4),
    .io_pixelVal_out_2_5(filter_io_pixelVal_out_2_5),
    .io_pixelVal_out_2_6(filter_io_pixelVal_out_2_6),
    .io_pixelVal_out_2_7(filter_io_pixelVal_out_2_7),
    .io_valid_out(filter_io_valid_out)
  );
  VideoBuffer videoBuffer ( // @[ImageProcessing.scala 24:27]
    .clock(videoBuffer_clock),
    .reset(videoBuffer_reset),
    .io_pixelVal_in_0_0(videoBuffer_io_pixelVal_in_0_0),
    .io_pixelVal_in_0_1(videoBuffer_io_pixelVal_in_0_1),
    .io_pixelVal_in_0_2(videoBuffer_io_pixelVal_in_0_2),
    .io_pixelVal_in_0_3(videoBuffer_io_pixelVal_in_0_3),
    .io_pixelVal_in_0_4(videoBuffer_io_pixelVal_in_0_4),
    .io_pixelVal_in_0_5(videoBuffer_io_pixelVal_in_0_5),
    .io_pixelVal_in_0_6(videoBuffer_io_pixelVal_in_0_6),
    .io_pixelVal_in_0_7(videoBuffer_io_pixelVal_in_0_7),
    .io_pixelVal_in_1_0(videoBuffer_io_pixelVal_in_1_0),
    .io_pixelVal_in_1_1(videoBuffer_io_pixelVal_in_1_1),
    .io_pixelVal_in_1_2(videoBuffer_io_pixelVal_in_1_2),
    .io_pixelVal_in_1_3(videoBuffer_io_pixelVal_in_1_3),
    .io_pixelVal_in_1_4(videoBuffer_io_pixelVal_in_1_4),
    .io_pixelVal_in_1_5(videoBuffer_io_pixelVal_in_1_5),
    .io_pixelVal_in_1_6(videoBuffer_io_pixelVal_in_1_6),
    .io_pixelVal_in_1_7(videoBuffer_io_pixelVal_in_1_7),
    .io_pixelVal_in_2_0(videoBuffer_io_pixelVal_in_2_0),
    .io_pixelVal_in_2_1(videoBuffer_io_pixelVal_in_2_1),
    .io_pixelVal_in_2_2(videoBuffer_io_pixelVal_in_2_2),
    .io_pixelVal_in_2_3(videoBuffer_io_pixelVal_in_2_3),
    .io_pixelVal_in_2_4(videoBuffer_io_pixelVal_in_2_4),
    .io_pixelVal_in_2_5(videoBuffer_io_pixelVal_in_2_5),
    .io_pixelVal_in_2_6(videoBuffer_io_pixelVal_in_2_6),
    .io_pixelVal_in_2_7(videoBuffer_io_pixelVal_in_2_7),
    .io_valid_in(videoBuffer_io_valid_in),
    .io_rowIndex(videoBuffer_io_rowIndex),
    .io_colIndex(videoBuffer_io_colIndex),
    .io_pixelVal_out_0(videoBuffer_io_pixelVal_out_0),
    .io_pixelVal_out_1(videoBuffer_io_pixelVal_out_1),
    .io_pixelVal_out_2(videoBuffer_io_pixelVal_out_2)
  );
  assign io_pixelVal_out_0 = videoBuffer_io_pixelVal_out_0; // @[ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25]
  assign io_pixelVal_out_1 = videoBuffer_io_pixelVal_out_1; // @[ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25]
  assign io_pixelVal_out_2 = videoBuffer_io_pixelVal_out_2; // @[ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25]
  assign filter_clock = clock;
  assign filter_reset = reset;
  assign filter_io_SPI_filterIndex = io_SPI_filterIndex; // @[ImageProcessing.scala 29:29]
  assign filter_io_SPI_distort = io_SPI_distort; // @[ImageProcessing.scala 31:29]
  assign videoBuffer_clock = clock;
  assign videoBuffer_reset = reset;
  assign videoBuffer_io_pixelVal_in_0_0 = filter_io_pixelVal_out_0_0; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_1 = filter_io_pixelVal_out_0_1; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_2 = filter_io_pixelVal_out_0_2; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_3 = filter_io_pixelVal_out_0_3; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_4 = filter_io_pixelVal_out_0_4; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_5 = filter_io_pixelVal_out_0_5; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_6 = filter_io_pixelVal_out_0_6; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_7 = filter_io_pixelVal_out_0_7; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_0 = filter_io_pixelVal_out_1_0; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_1 = filter_io_pixelVal_out_1_1; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_2 = filter_io_pixelVal_out_1_2; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_3 = filter_io_pixelVal_out_1_3; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_4 = filter_io_pixelVal_out_1_4; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_5 = filter_io_pixelVal_out_1_5; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_6 = filter_io_pixelVal_out_1_6; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_7 = filter_io_pixelVal_out_1_7; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_0 = filter_io_pixelVal_out_2_0; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_1 = filter_io_pixelVal_out_2_1; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_2 = filter_io_pixelVal_out_2_2; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_3 = filter_io_pixelVal_out_2_3; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_4 = filter_io_pixelVal_out_2_4; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_5 = filter_io_pixelVal_out_2_5; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_6 = filter_io_pixelVal_out_2_6; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_7 = filter_io_pixelVal_out_2_7; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_valid_in = filter_io_valid_out; // @[ImageProcessing.scala 39:27]
  assign videoBuffer_io_rowIndex = io_rowIndex; // @[ImageProcessing.scala 26:27]
  assign videoBuffer_io_colIndex = io_colIndex; // @[ImageProcessing.scala 27:27]
endmodule
