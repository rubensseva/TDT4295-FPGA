module DotProd(
  input        clock,
  input        reset,
  input  [7:0] io_dataInA,
  input  [7:0] io_dataInB,
  output [8:0] io_dataOut,
  output       io_outputValid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] countVal; // @[Counter.scala 29:33]
  wire  countReset = countVal == 4'h8; // @[Counter.scala 38:24]
  wire [3:0] _T_2 = countVal + 4'h1; // @[Counter.scala 39:22]
  reg [8:0] accumulator; // @[DotProd.scala 19:28]
  wire [15:0] product = $signed(io_dataInA) * $signed(io_dataInB); // @[DotProd.scala 20:35]
  wire [15:0] _GEN_5 = {{7{accumulator[8]}},accumulator}; // @[DotProd.scala 21:30]
  wire [15:0] _T_6 = $signed(_GEN_5) + $signed(product); // @[DotProd.scala 21:30]
  wire  _T_11 = ~reset; // @[DotProd.scala 29:11]
  wire [15:0] _GEN_4 = countReset ? $signed(16'sh0) : $signed(_T_6); // @[DotProd.scala 25:20]
  assign io_dataOut = _T_6[8:0]; // @[DotProd.scala 23:14]
  assign io_outputValid = countVal == 4'h8; // @[DotProd.scala 26:20 DotProd.scala 31:20]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  countVal = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  accumulator = _RAND_1[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      countVal <= 4'h0;
    end else if (countReset) begin
      countVal <= 4'h0;
    end else begin
      countVal <= _T_2;
    end
    if (reset) begin
      accumulator <= 9'sh0;
    end else begin
      accumulator <= _GEN_4[8:0];
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (countReset & _T_11) begin
          $fwrite(32'h80000002,"VALOUTidghspdolgnfgkln\n"); // @[DotProd.scala 29:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module KernelConvolution(
  input        clock,
  input        reset,
  input  [4:0] io_kernelVal_in,
  input  [3:0] io_pixelVal_in_0,
  input  [3:0] io_pixelVal_in_1,
  input  [3:0] io_pixelVal_in_2,
  input  [3:0] io_pixelVal_in_3,
  input  [3:0] io_pixelVal_in_4,
  input  [3:0] io_pixelVal_in_5,
  input  [3:0] io_pixelVal_in_6,
  input  [3:0] io_pixelVal_in_7,
  output [8:0] io_pixelVal_out_0,
  output [8:0] io_pixelVal_out_1,
  output [8:0] io_pixelVal_out_2,
  output [8:0] io_pixelVal_out_3,
  output [8:0] io_pixelVal_out_4,
  output [8:0] io_pixelVal_out_5,
  output [8:0] io_pixelVal_out_6,
  output [8:0] io_pixelVal_out_7,
  output       io_valid_out
);
  wire  DotProd_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_1_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_1_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_1_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_1_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_1_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_1_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_2_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_2_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_2_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_2_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_2_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_2_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_3_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_3_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_3_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_3_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_3_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_3_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_4_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_4_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_4_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_4_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_4_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_4_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_5_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_5_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_5_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_5_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_5_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_5_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_6_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_6_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_6_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_6_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_6_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_6_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_7_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_7_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_7_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_7_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_7_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_7_io_outputValid; // @[KernelConvolution.scala 21:58]
  DotProd DotProd ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_clock),
    .reset(DotProd_reset),
    .io_dataInA(DotProd_io_dataInA),
    .io_dataInB(DotProd_io_dataInB),
    .io_dataOut(DotProd_io_dataOut),
    .io_outputValid(DotProd_io_outputValid)
  );
  DotProd DotProd_1 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_1_clock),
    .reset(DotProd_1_reset),
    .io_dataInA(DotProd_1_io_dataInA),
    .io_dataInB(DotProd_1_io_dataInB),
    .io_dataOut(DotProd_1_io_dataOut),
    .io_outputValid(DotProd_1_io_outputValid)
  );
  DotProd DotProd_2 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_2_clock),
    .reset(DotProd_2_reset),
    .io_dataInA(DotProd_2_io_dataInA),
    .io_dataInB(DotProd_2_io_dataInB),
    .io_dataOut(DotProd_2_io_dataOut),
    .io_outputValid(DotProd_2_io_outputValid)
  );
  DotProd DotProd_3 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_3_clock),
    .reset(DotProd_3_reset),
    .io_dataInA(DotProd_3_io_dataInA),
    .io_dataInB(DotProd_3_io_dataInB),
    .io_dataOut(DotProd_3_io_dataOut),
    .io_outputValid(DotProd_3_io_outputValid)
  );
  DotProd DotProd_4 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_4_clock),
    .reset(DotProd_4_reset),
    .io_dataInA(DotProd_4_io_dataInA),
    .io_dataInB(DotProd_4_io_dataInB),
    .io_dataOut(DotProd_4_io_dataOut),
    .io_outputValid(DotProd_4_io_outputValid)
  );
  DotProd DotProd_5 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_5_clock),
    .reset(DotProd_5_reset),
    .io_dataInA(DotProd_5_io_dataInA),
    .io_dataInB(DotProd_5_io_dataInB),
    .io_dataOut(DotProd_5_io_dataOut),
    .io_outputValid(DotProd_5_io_outputValid)
  );
  DotProd DotProd_6 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_6_clock),
    .reset(DotProd_6_reset),
    .io_dataInA(DotProd_6_io_dataInA),
    .io_dataInB(DotProd_6_io_dataInB),
    .io_dataOut(DotProd_6_io_dataOut),
    .io_outputValid(DotProd_6_io_outputValid)
  );
  DotProd DotProd_7 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_7_clock),
    .reset(DotProd_7_reset),
    .io_dataInA(DotProd_7_io_dataInA),
    .io_dataInB(DotProd_7_io_dataInB),
    .io_dataOut(DotProd_7_io_dataOut),
    .io_outputValid(DotProd_7_io_outputValid)
  );
  assign io_pixelVal_out_0 = DotProd_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_1 = DotProd_1_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_2 = DotProd_2_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_3 = DotProd_3_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_4 = DotProd_4_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_5 = DotProd_5_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_6 = DotProd_6_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_7 = DotProd_7_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_valid_out = DotProd_io_outputValid; // @[KernelConvolution.scala 35:30]
  assign DotProd_clock = clock;
  assign DotProd_reset = reset;
  assign DotProd_io_dataInA = {{4'd0}, io_pixelVal_in_0}; // @[KernelConvolution.scala 21:32]
  assign DotProd_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_1_clock = clock;
  assign DotProd_1_reset = reset;
  assign DotProd_1_io_dataInA = {{4'd0}, io_pixelVal_in_1}; // @[KernelConvolution.scala 21:32]
  assign DotProd_1_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_2_clock = clock;
  assign DotProd_2_reset = reset;
  assign DotProd_2_io_dataInA = {{4'd0}, io_pixelVal_in_2}; // @[KernelConvolution.scala 21:32]
  assign DotProd_2_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_3_clock = clock;
  assign DotProd_3_reset = reset;
  assign DotProd_3_io_dataInA = {{4'd0}, io_pixelVal_in_3}; // @[KernelConvolution.scala 21:32]
  assign DotProd_3_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_4_clock = clock;
  assign DotProd_4_reset = reset;
  assign DotProd_4_io_dataInA = {{4'd0}, io_pixelVal_in_4}; // @[KernelConvolution.scala 21:32]
  assign DotProd_4_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_5_clock = clock;
  assign DotProd_5_reset = reset;
  assign DotProd_5_io_dataInA = {{4'd0}, io_pixelVal_in_5}; // @[KernelConvolution.scala 21:32]
  assign DotProd_5_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_6_clock = clock;
  assign DotProd_6_reset = reset;
  assign DotProd_6_io_dataInA = {{4'd0}, io_pixelVal_in_6}; // @[KernelConvolution.scala 21:32]
  assign DotProd_6_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_7_clock = clock;
  assign DotProd_7_reset = reset;
  assign DotProd_7_io_dataInA = {{4'd0}, io_pixelVal_in_7}; // @[KernelConvolution.scala 21:32]
  assign DotProd_7_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
endmodule
module Filter(
  input        clock,
  input        reset,
  input  [5:0] io_SPI_filterIndex,
  input        io_SPI_distort,
  output [3:0] io_pixelVal_out_0_0,
  output [3:0] io_pixelVal_out_0_1,
  output [3:0] io_pixelVal_out_0_2,
  output [3:0] io_pixelVal_out_0_3,
  output [3:0] io_pixelVal_out_0_4,
  output [3:0] io_pixelVal_out_0_5,
  output [3:0] io_pixelVal_out_0_6,
  output [3:0] io_pixelVal_out_0_7,
  output [3:0] io_pixelVal_out_1_0,
  output [3:0] io_pixelVal_out_1_1,
  output [3:0] io_pixelVal_out_1_2,
  output [3:0] io_pixelVal_out_1_3,
  output [3:0] io_pixelVal_out_1_4,
  output [3:0] io_pixelVal_out_1_5,
  output [3:0] io_pixelVal_out_1_6,
  output [3:0] io_pixelVal_out_1_7,
  output [3:0] io_pixelVal_out_2_0,
  output [3:0] io_pixelVal_out_2_1,
  output [3:0] io_pixelVal_out_2_2,
  output [3:0] io_pixelVal_out_2_3,
  output [3:0] io_pixelVal_out_2_4,
  output [3:0] io_pixelVal_out_2_5,
  output [3:0] io_pixelVal_out_2_6,
  output [3:0] io_pixelVal_out_2_7,
  output       io_valid_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  KernelConvolution_clock; // @[Filter.scala 142:36]
  wire  KernelConvolution_reset; // @[Filter.scala 142:36]
  wire [4:0] KernelConvolution_io_kernelVal_in; // @[Filter.scala 142:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_0; // @[Filter.scala 142:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_1; // @[Filter.scala 142:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_2; // @[Filter.scala 142:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_3; // @[Filter.scala 142:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_4; // @[Filter.scala 142:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_5; // @[Filter.scala 142:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_6; // @[Filter.scala 142:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_7; // @[Filter.scala 142:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_0; // @[Filter.scala 142:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_1; // @[Filter.scala 142:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_2; // @[Filter.scala 142:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_3; // @[Filter.scala 142:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_4; // @[Filter.scala 142:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_5; // @[Filter.scala 142:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_6; // @[Filter.scala 142:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_7; // @[Filter.scala 142:36]
  wire  KernelConvolution_io_valid_out; // @[Filter.scala 142:36]
  wire  KernelConvolution_1_clock; // @[Filter.scala 143:36]
  wire  KernelConvolution_1_reset; // @[Filter.scala 143:36]
  wire [4:0] KernelConvolution_1_io_kernelVal_in; // @[Filter.scala 143:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_0; // @[Filter.scala 143:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_1; // @[Filter.scala 143:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_2; // @[Filter.scala 143:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_3; // @[Filter.scala 143:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_4; // @[Filter.scala 143:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_5; // @[Filter.scala 143:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_6; // @[Filter.scala 143:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_7; // @[Filter.scala 143:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_0; // @[Filter.scala 143:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_1; // @[Filter.scala 143:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_2; // @[Filter.scala 143:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_3; // @[Filter.scala 143:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_4; // @[Filter.scala 143:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_5; // @[Filter.scala 143:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_6; // @[Filter.scala 143:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_7; // @[Filter.scala 143:36]
  wire  KernelConvolution_1_io_valid_out; // @[Filter.scala 143:36]
  wire  KernelConvolution_2_clock; // @[Filter.scala 144:36]
  wire  KernelConvolution_2_reset; // @[Filter.scala 144:36]
  wire [4:0] KernelConvolution_2_io_kernelVal_in; // @[Filter.scala 144:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_0; // @[Filter.scala 144:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_1; // @[Filter.scala 144:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_2; // @[Filter.scala 144:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_3; // @[Filter.scala 144:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_4; // @[Filter.scala 144:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_5; // @[Filter.scala 144:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_6; // @[Filter.scala 144:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_7; // @[Filter.scala 144:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_0; // @[Filter.scala 144:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_1; // @[Filter.scala 144:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_2; // @[Filter.scala 144:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_3; // @[Filter.scala 144:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_4; // @[Filter.scala 144:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_5; // @[Filter.scala 144:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_6; // @[Filter.scala 144:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_7; // @[Filter.scala 144:36]
  wire  KernelConvolution_2_io_valid_out; // @[Filter.scala 144:36]
  reg [3:0] kernelCounter; // @[Counter.scala 29:33]
  wire  kernelCountReset = kernelCounter == 4'h8; // @[Counter.scala 38:24]
  wire [3:0] _T_14 = kernelCounter + 4'h1; // @[Counter.scala 39:22]
  wire  _GEN_18683 = 3'h0 == io_SPI_filterIndex[2:0]; // @[Filter.scala 150:41]
  wire  _GEN_18684 = 4'h4 == kernelCounter; // @[Filter.scala 150:41]
  wire [4:0] _GEN_7 = _GEN_18683 & _GEN_18684 ? $signed(5'sh1) : $signed(5'sh0); // @[Filter.scala 150:41]
  wire  _GEN_18686 = 4'h5 == kernelCounter; // @[Filter.scala 150:41]
  wire [4:0] _GEN_8 = _GEN_18683 & _GEN_18686 ? $signed(5'sh0) : $signed(_GEN_7); // @[Filter.scala 150:41]
  wire  _GEN_18688 = 4'h6 == kernelCounter; // @[Filter.scala 150:41]
  wire [4:0] _GEN_9 = _GEN_18683 & _GEN_18688 ? $signed(5'sh0) : $signed(_GEN_8); // @[Filter.scala 150:41]
  wire  _GEN_18690 = 4'h7 == kernelCounter; // @[Filter.scala 150:41]
  wire [4:0] _GEN_10 = _GEN_18683 & _GEN_18690 ? $signed(5'sh0) : $signed(_GEN_9); // @[Filter.scala 150:41]
  wire  _GEN_18692 = 4'h8 == kernelCounter; // @[Filter.scala 150:41]
  wire [4:0] _GEN_11 = _GEN_18683 & _GEN_18692 ? $signed(5'sh0) : $signed(_GEN_10); // @[Filter.scala 150:41]
  wire  _GEN_18693 = 3'h1 == io_SPI_filterIndex[2:0]; // @[Filter.scala 150:41]
  wire  _GEN_18694 = 4'h0 == kernelCounter; // @[Filter.scala 150:41]
  wire [4:0] _GEN_12 = _GEN_18693 & _GEN_18694 ? $signed(5'sh1) : $signed(_GEN_11); // @[Filter.scala 150:41]
  wire  _GEN_18696 = 4'h1 == kernelCounter; // @[Filter.scala 150:41]
  wire [4:0] _GEN_13 = _GEN_18693 & _GEN_18696 ? $signed(5'sh1) : $signed(_GEN_12); // @[Filter.scala 150:41]
  wire  _GEN_18698 = 4'h2 == kernelCounter; // @[Filter.scala 150:41]
  wire [4:0] _GEN_14 = _GEN_18693 & _GEN_18698 ? $signed(5'sh1) : $signed(_GEN_13); // @[Filter.scala 150:41]
  wire  _GEN_18700 = 4'h3 == kernelCounter; // @[Filter.scala 150:41]
  wire [4:0] _GEN_15 = _GEN_18693 & _GEN_18700 ? $signed(5'sh1) : $signed(_GEN_14); // @[Filter.scala 150:41]
  wire [4:0] _GEN_16 = _GEN_18693 & _GEN_18684 ? $signed(5'sh1) : $signed(_GEN_15); // @[Filter.scala 150:41]
  wire [4:0] _GEN_17 = _GEN_18693 & _GEN_18686 ? $signed(5'sh1) : $signed(_GEN_16); // @[Filter.scala 150:41]
  wire [4:0] _GEN_18 = _GEN_18693 & _GEN_18688 ? $signed(5'sh1) : $signed(_GEN_17); // @[Filter.scala 150:41]
  wire [4:0] _GEN_19 = _GEN_18693 & _GEN_18690 ? $signed(5'sh1) : $signed(_GEN_18); // @[Filter.scala 150:41]
  wire [4:0] _GEN_20 = _GEN_18693 & _GEN_18692 ? $signed(5'sh1) : $signed(_GEN_19); // @[Filter.scala 150:41]
  wire  _GEN_18711 = 3'h2 == io_SPI_filterIndex[2:0]; // @[Filter.scala 150:41]
  wire [4:0] _GEN_21 = _GEN_18711 & _GEN_18694 ? $signed(5'sh1) : $signed(_GEN_20); // @[Filter.scala 150:41]
  wire [4:0] _GEN_22 = _GEN_18711 & _GEN_18696 ? $signed(5'sh2) : $signed(_GEN_21); // @[Filter.scala 150:41]
  wire [4:0] _GEN_23 = _GEN_18711 & _GEN_18698 ? $signed(5'sh1) : $signed(_GEN_22); // @[Filter.scala 150:41]
  wire [4:0] _GEN_24 = _GEN_18711 & _GEN_18700 ? $signed(5'sh2) : $signed(_GEN_23); // @[Filter.scala 150:41]
  wire [4:0] _GEN_25 = _GEN_18711 & _GEN_18684 ? $signed(5'sh4) : $signed(_GEN_24); // @[Filter.scala 150:41]
  wire [4:0] _GEN_26 = _GEN_18711 & _GEN_18686 ? $signed(5'sh2) : $signed(_GEN_25); // @[Filter.scala 150:41]
  wire [4:0] _GEN_27 = _GEN_18711 & _GEN_18688 ? $signed(5'sh1) : $signed(_GEN_26); // @[Filter.scala 150:41]
  wire [4:0] _GEN_28 = _GEN_18711 & _GEN_18690 ? $signed(5'sh2) : $signed(_GEN_27); // @[Filter.scala 150:41]
  wire [4:0] _GEN_29 = _GEN_18711 & _GEN_18692 ? $signed(5'sh1) : $signed(_GEN_28); // @[Filter.scala 150:41]
  wire  _GEN_18729 = 3'h3 == io_SPI_filterIndex[2:0]; // @[Filter.scala 150:41]
  wire [4:0] _GEN_30 = _GEN_18729 & _GEN_18694 ? $signed(5'sh0) : $signed(_GEN_29); // @[Filter.scala 150:41]
  wire [4:0] _GEN_31 = _GEN_18729 & _GEN_18696 ? $signed(-5'sh1) : $signed(_GEN_30); // @[Filter.scala 150:41]
  wire [4:0] _GEN_32 = _GEN_18729 & _GEN_18698 ? $signed(5'sh0) : $signed(_GEN_31); // @[Filter.scala 150:41]
  wire [4:0] _GEN_33 = _GEN_18729 & _GEN_18700 ? $signed(-5'sh1) : $signed(_GEN_32); // @[Filter.scala 150:41]
  wire [4:0] _GEN_34 = _GEN_18729 & _GEN_18684 ? $signed(5'sh4) : $signed(_GEN_33); // @[Filter.scala 150:41]
  wire [4:0] _GEN_35 = _GEN_18729 & _GEN_18686 ? $signed(-5'sh1) : $signed(_GEN_34); // @[Filter.scala 150:41]
  wire [4:0] _GEN_36 = _GEN_18729 & _GEN_18688 ? $signed(5'sh0) : $signed(_GEN_35); // @[Filter.scala 150:41]
  wire [4:0] _GEN_37 = _GEN_18729 & _GEN_18690 ? $signed(-5'sh1) : $signed(_GEN_36); // @[Filter.scala 150:41]
  wire [4:0] _GEN_38 = _GEN_18729 & _GEN_18692 ? $signed(5'sh0) : $signed(_GEN_37); // @[Filter.scala 150:41]
  wire  _GEN_18747 = 3'h4 == io_SPI_filterIndex[2:0]; // @[Filter.scala 150:41]
  wire [4:0] _GEN_39 = _GEN_18747 & _GEN_18694 ? $signed(-5'sh1) : $signed(_GEN_38); // @[Filter.scala 150:41]
  wire [4:0] _GEN_40 = _GEN_18747 & _GEN_18696 ? $signed(-5'sh1) : $signed(_GEN_39); // @[Filter.scala 150:41]
  wire [4:0] _GEN_41 = _GEN_18747 & _GEN_18698 ? $signed(-5'sh1) : $signed(_GEN_40); // @[Filter.scala 150:41]
  wire [4:0] _GEN_42 = _GEN_18747 & _GEN_18700 ? $signed(-5'sh1) : $signed(_GEN_41); // @[Filter.scala 150:41]
  wire [4:0] _GEN_43 = _GEN_18747 & _GEN_18684 ? $signed(5'sh8) : $signed(_GEN_42); // @[Filter.scala 150:41]
  wire [4:0] _GEN_44 = _GEN_18747 & _GEN_18686 ? $signed(-5'sh1) : $signed(_GEN_43); // @[Filter.scala 150:41]
  wire [4:0] _GEN_45 = _GEN_18747 & _GEN_18688 ? $signed(-5'sh1) : $signed(_GEN_44); // @[Filter.scala 150:41]
  wire [4:0] _GEN_46 = _GEN_18747 & _GEN_18690 ? $signed(-5'sh1) : $signed(_GEN_45); // @[Filter.scala 150:41]
  wire [4:0] _GEN_47 = _GEN_18747 & _GEN_18692 ? $signed(-5'sh1) : $signed(_GEN_46); // @[Filter.scala 150:41]
  wire  _GEN_18765 = 3'h5 == io_SPI_filterIndex[2:0]; // @[Filter.scala 150:41]
  wire [4:0] _GEN_48 = _GEN_18765 & _GEN_18694 ? $signed(5'sh0) : $signed(_GEN_47); // @[Filter.scala 150:41]
  wire [4:0] _GEN_49 = _GEN_18765 & _GEN_18696 ? $signed(-5'sh1) : $signed(_GEN_48); // @[Filter.scala 150:41]
  wire [4:0] _GEN_50 = _GEN_18765 & _GEN_18698 ? $signed(5'sh0) : $signed(_GEN_49); // @[Filter.scala 150:41]
  wire [4:0] _GEN_51 = _GEN_18765 & _GEN_18700 ? $signed(-5'sh1) : $signed(_GEN_50); // @[Filter.scala 150:41]
  wire [4:0] _GEN_52 = _GEN_18765 & _GEN_18684 ? $signed(5'sh5) : $signed(_GEN_51); // @[Filter.scala 150:41]
  wire [4:0] _GEN_53 = _GEN_18765 & _GEN_18686 ? $signed(-5'sh1) : $signed(_GEN_52); // @[Filter.scala 150:41]
  wire [4:0] _GEN_54 = _GEN_18765 & _GEN_18688 ? $signed(5'sh0) : $signed(_GEN_53); // @[Filter.scala 150:41]
  wire [4:0] _GEN_55 = _GEN_18765 & _GEN_18690 ? $signed(-5'sh1) : $signed(_GEN_54); // @[Filter.scala 150:41]
  reg [1:0] imageCounterX; // @[Counter.scala 29:33]
  wire  imageCounterXReset = imageCounterX == 2'h2; // @[Counter.scala 38:24]
  wire [1:0] _T_20 = imageCounterX + 2'h1; // @[Counter.scala 39:22]
  reg [1:0] imageCounterY; // @[Counter.scala 29:33]
  wire  _T_21 = imageCounterY == 2'h2; // @[Counter.scala 38:24]
  wire [1:0] _T_23 = imageCounterY + 2'h1; // @[Counter.scala 39:22]
  reg [31:0] pixelIndex; // @[Filter.scala 155:31]
  wire [32:0] _T_24 = {{1'd0}, pixelIndex}; // @[Filter.scala 158:31]
  wire [31:0] _GEN_0 = _T_24[31:0] % 32'h10; // @[Filter.scala 158:38]
  wire [4:0] _T_26 = _GEN_0[4:0]; // @[Filter.scala 158:38]
  wire [4:0] _GEN_18983 = {{3'd0}, imageCounterX}; // @[Filter.scala 158:53]
  wire [4:0] _T_28 = _T_26 + _GEN_18983; // @[Filter.scala 158:53]
  wire [4:0] _T_30 = _T_28 - 5'h1; // @[Filter.scala 158:69]
  wire [31:0] _T_33 = _T_24[31:0] / 32'h10; // @[Filter.scala 159:38]
  wire [31:0] _GEN_18984 = {{30'd0}, imageCounterY}; // @[Filter.scala 159:53]
  wire [31:0] _T_35 = _T_33 + _GEN_18984; // @[Filter.scala 159:53]
  wire [31:0] _T_37 = _T_35 - 32'h1; // @[Filter.scala 159:69]
  wire  _T_39 = _T_30 >= 5'h10; // @[Filter.scala 162:31]
  wire  _T_43 = _T_37 >= 32'hc; // @[Filter.scala 162:63]
  wire  _T_44 = _T_39 | _T_43; // @[Filter.scala 162:58]
  wire [36:0] _T_45 = _T_37 * 32'h10; // @[Filter.scala 165:66]
  wire [36:0] _GEN_18985 = {{32'd0}, _T_30}; // @[Filter.scala 165:81]
  wire [36:0] _T_47 = _T_45 + _GEN_18985; // @[Filter.scala 165:81]
  wire [3:0] _GEN_179 = 8'h8 == _T_47[7:0] ? 4'h0 : 4'hf; // @[Filter.scala 165:86]
  wire [3:0] _GEN_180 = 8'h9 == _T_47[7:0] ? 4'h0 : _GEN_179; // @[Filter.scala 165:86]
  wire [3:0] _GEN_181 = 8'ha == _T_47[7:0] ? 4'h0 : _GEN_180; // @[Filter.scala 165:86]
  wire [3:0] _GEN_182 = 8'hb == _T_47[7:0] ? 4'h0 : _GEN_181; // @[Filter.scala 165:86]
  wire [3:0] _GEN_183 = 8'hc == _T_47[7:0] ? 4'h0 : _GEN_182; // @[Filter.scala 165:86]
  wire [3:0] _GEN_184 = 8'hd == _T_47[7:0] ? 4'h0 : _GEN_183; // @[Filter.scala 165:86]
  wire [3:0] _GEN_185 = 8'he == _T_47[7:0] ? 4'h0 : _GEN_184; // @[Filter.scala 165:86]
  wire [3:0] _GEN_186 = 8'hf == _T_47[7:0] ? 4'h0 : _GEN_185; // @[Filter.scala 165:86]
  wire [3:0] _GEN_187 = 8'h10 == _T_47[7:0] ? 4'hf : _GEN_186; // @[Filter.scala 165:86]
  wire [3:0] _GEN_188 = 8'h11 == _T_47[7:0] ? 4'hf : _GEN_187; // @[Filter.scala 165:86]
  wire [3:0] _GEN_189 = 8'h12 == _T_47[7:0] ? 4'hf : _GEN_188; // @[Filter.scala 165:86]
  wire [3:0] _GEN_190 = 8'h13 == _T_47[7:0] ? 4'hf : _GEN_189; // @[Filter.scala 165:86]
  wire [3:0] _GEN_191 = 8'h14 == _T_47[7:0] ? 4'hf : _GEN_190; // @[Filter.scala 165:86]
  wire [3:0] _GEN_192 = 8'h15 == _T_47[7:0] ? 4'hf : _GEN_191; // @[Filter.scala 165:86]
  wire [3:0] _GEN_193 = 8'h16 == _T_47[7:0] ? 4'hf : _GEN_192; // @[Filter.scala 165:86]
  wire [3:0] _GEN_194 = 8'h17 == _T_47[7:0] ? 4'hf : _GEN_193; // @[Filter.scala 165:86]
  wire [3:0] _GEN_195 = 8'h18 == _T_47[7:0] ? 4'h0 : _GEN_194; // @[Filter.scala 165:86]
  wire [3:0] _GEN_196 = 8'h19 == _T_47[7:0] ? 4'h0 : _GEN_195; // @[Filter.scala 165:86]
  wire [3:0] _GEN_197 = 8'h1a == _T_47[7:0] ? 4'h0 : _GEN_196; // @[Filter.scala 165:86]
  wire [3:0] _GEN_198 = 8'h1b == _T_47[7:0] ? 4'h0 : _GEN_197; // @[Filter.scala 165:86]
  wire [3:0] _GEN_199 = 8'h1c == _T_47[7:0] ? 4'h0 : _GEN_198; // @[Filter.scala 165:86]
  wire [3:0] _GEN_200 = 8'h1d == _T_47[7:0] ? 4'h0 : _GEN_199; // @[Filter.scala 165:86]
  wire [3:0] _GEN_201 = 8'h1e == _T_47[7:0] ? 4'h0 : _GEN_200; // @[Filter.scala 165:86]
  wire [3:0] _GEN_202 = 8'h1f == _T_47[7:0] ? 4'h0 : _GEN_201; // @[Filter.scala 165:86]
  wire [3:0] _GEN_203 = 8'h20 == _T_47[7:0] ? 4'hf : _GEN_202; // @[Filter.scala 165:86]
  wire [3:0] _GEN_204 = 8'h21 == _T_47[7:0] ? 4'hf : _GEN_203; // @[Filter.scala 165:86]
  wire [3:0] _GEN_205 = 8'h22 == _T_47[7:0] ? 4'hf : _GEN_204; // @[Filter.scala 165:86]
  wire [3:0] _GEN_206 = 8'h23 == _T_47[7:0] ? 4'hf : _GEN_205; // @[Filter.scala 165:86]
  wire [3:0] _GEN_207 = 8'h24 == _T_47[7:0] ? 4'hf : _GEN_206; // @[Filter.scala 165:86]
  wire [3:0] _GEN_208 = 8'h25 == _T_47[7:0] ? 4'hf : _GEN_207; // @[Filter.scala 165:86]
  wire [3:0] _GEN_209 = 8'h26 == _T_47[7:0] ? 4'hf : _GEN_208; // @[Filter.scala 165:86]
  wire [3:0] _GEN_210 = 8'h27 == _T_47[7:0] ? 4'hf : _GEN_209; // @[Filter.scala 165:86]
  wire [3:0] _GEN_211 = 8'h28 == _T_47[7:0] ? 4'h0 : _GEN_210; // @[Filter.scala 165:86]
  wire [3:0] _GEN_212 = 8'h29 == _T_47[7:0] ? 4'h0 : _GEN_211; // @[Filter.scala 165:86]
  wire [3:0] _GEN_213 = 8'h2a == _T_47[7:0] ? 4'h0 : _GEN_212; // @[Filter.scala 165:86]
  wire [3:0] _GEN_214 = 8'h2b == _T_47[7:0] ? 4'h0 : _GEN_213; // @[Filter.scala 165:86]
  wire [3:0] _GEN_215 = 8'h2c == _T_47[7:0] ? 4'h0 : _GEN_214; // @[Filter.scala 165:86]
  wire [3:0] _GEN_216 = 8'h2d == _T_47[7:0] ? 4'h0 : _GEN_215; // @[Filter.scala 165:86]
  wire [3:0] _GEN_217 = 8'h2e == _T_47[7:0] ? 4'h0 : _GEN_216; // @[Filter.scala 165:86]
  wire [3:0] _GEN_218 = 8'h2f == _T_47[7:0] ? 4'h0 : _GEN_217; // @[Filter.scala 165:86]
  wire [3:0] _GEN_219 = 8'h30 == _T_47[7:0] ? 4'hf : _GEN_218; // @[Filter.scala 165:86]
  wire [3:0] _GEN_220 = 8'h31 == _T_47[7:0] ? 4'hf : _GEN_219; // @[Filter.scala 165:86]
  wire [3:0] _GEN_221 = 8'h32 == _T_47[7:0] ? 4'hf : _GEN_220; // @[Filter.scala 165:86]
  wire [3:0] _GEN_222 = 8'h33 == _T_47[7:0] ? 4'hf : _GEN_221; // @[Filter.scala 165:86]
  wire [3:0] _GEN_223 = 8'h34 == _T_47[7:0] ? 4'hf : _GEN_222; // @[Filter.scala 165:86]
  wire [3:0] _GEN_224 = 8'h35 == _T_47[7:0] ? 4'hf : _GEN_223; // @[Filter.scala 165:86]
  wire [3:0] _GEN_225 = 8'h36 == _T_47[7:0] ? 4'hf : _GEN_224; // @[Filter.scala 165:86]
  wire [3:0] _GEN_226 = 8'h37 == _T_47[7:0] ? 4'hf : _GEN_225; // @[Filter.scala 165:86]
  wire [3:0] _GEN_227 = 8'h38 == _T_47[7:0] ? 4'h0 : _GEN_226; // @[Filter.scala 165:86]
  wire [3:0] _GEN_228 = 8'h39 == _T_47[7:0] ? 4'h0 : _GEN_227; // @[Filter.scala 165:86]
  wire [3:0] _GEN_229 = 8'h3a == _T_47[7:0] ? 4'h0 : _GEN_228; // @[Filter.scala 165:86]
  wire [3:0] _GEN_230 = 8'h3b == _T_47[7:0] ? 4'h0 : _GEN_229; // @[Filter.scala 165:86]
  wire [3:0] _GEN_231 = 8'h3c == _T_47[7:0] ? 4'h0 : _GEN_230; // @[Filter.scala 165:86]
  wire [3:0] _GEN_232 = 8'h3d == _T_47[7:0] ? 4'h0 : _GEN_231; // @[Filter.scala 165:86]
  wire [3:0] _GEN_233 = 8'h3e == _T_47[7:0] ? 4'h0 : _GEN_232; // @[Filter.scala 165:86]
  wire [3:0] _GEN_234 = 8'h3f == _T_47[7:0] ? 4'h0 : _GEN_233; // @[Filter.scala 165:86]
  wire [3:0] _GEN_235 = 8'h40 == _T_47[7:0] ? 4'hf : _GEN_234; // @[Filter.scala 165:86]
  wire [3:0] _GEN_236 = 8'h41 == _T_47[7:0] ? 4'hf : _GEN_235; // @[Filter.scala 165:86]
  wire [3:0] _GEN_237 = 8'h42 == _T_47[7:0] ? 4'hf : _GEN_236; // @[Filter.scala 165:86]
  wire [3:0] _GEN_238 = 8'h43 == _T_47[7:0] ? 4'hf : _GEN_237; // @[Filter.scala 165:86]
  wire [3:0] _GEN_239 = 8'h44 == _T_47[7:0] ? 4'hf : _GEN_238; // @[Filter.scala 165:86]
  wire [3:0] _GEN_240 = 8'h45 == _T_47[7:0] ? 4'hf : _GEN_239; // @[Filter.scala 165:86]
  wire [3:0] _GEN_241 = 8'h46 == _T_47[7:0] ? 4'hf : _GEN_240; // @[Filter.scala 165:86]
  wire [3:0] _GEN_242 = 8'h47 == _T_47[7:0] ? 4'hf : _GEN_241; // @[Filter.scala 165:86]
  wire [3:0] _GEN_243 = 8'h48 == _T_47[7:0] ? 4'h0 : _GEN_242; // @[Filter.scala 165:86]
  wire [3:0] _GEN_244 = 8'h49 == _T_47[7:0] ? 4'h0 : _GEN_243; // @[Filter.scala 165:86]
  wire [3:0] _GEN_245 = 8'h4a == _T_47[7:0] ? 4'h0 : _GEN_244; // @[Filter.scala 165:86]
  wire [3:0] _GEN_246 = 8'h4b == _T_47[7:0] ? 4'h0 : _GEN_245; // @[Filter.scala 165:86]
  wire [3:0] _GEN_247 = 8'h4c == _T_47[7:0] ? 4'h0 : _GEN_246; // @[Filter.scala 165:86]
  wire [3:0] _GEN_248 = 8'h4d == _T_47[7:0] ? 4'h0 : _GEN_247; // @[Filter.scala 165:86]
  wire [3:0] _GEN_249 = 8'h4e == _T_47[7:0] ? 4'h0 : _GEN_248; // @[Filter.scala 165:86]
  wire [3:0] _GEN_250 = 8'h4f == _T_47[7:0] ? 4'h0 : _GEN_249; // @[Filter.scala 165:86]
  wire [3:0] _GEN_251 = 8'h50 == _T_47[7:0] ? 4'hf : _GEN_250; // @[Filter.scala 165:86]
  wire [3:0] _GEN_252 = 8'h51 == _T_47[7:0] ? 4'hf : _GEN_251; // @[Filter.scala 165:86]
  wire [3:0] _GEN_253 = 8'h52 == _T_47[7:0] ? 4'hf : _GEN_252; // @[Filter.scala 165:86]
  wire [3:0] _GEN_254 = 8'h53 == _T_47[7:0] ? 4'hf : _GEN_253; // @[Filter.scala 165:86]
  wire [3:0] _GEN_255 = 8'h54 == _T_47[7:0] ? 4'hf : _GEN_254; // @[Filter.scala 165:86]
  wire [3:0] _GEN_256 = 8'h55 == _T_47[7:0] ? 4'hf : _GEN_255; // @[Filter.scala 165:86]
  wire [3:0] _GEN_257 = 8'h56 == _T_47[7:0] ? 4'hf : _GEN_256; // @[Filter.scala 165:86]
  wire [3:0] _GEN_258 = 8'h57 == _T_47[7:0] ? 4'hf : _GEN_257; // @[Filter.scala 165:86]
  wire [3:0] _GEN_259 = 8'h58 == _T_47[7:0] ? 4'h0 : _GEN_258; // @[Filter.scala 165:86]
  wire [3:0] _GEN_260 = 8'h59 == _T_47[7:0] ? 4'h0 : _GEN_259; // @[Filter.scala 165:86]
  wire [3:0] _GEN_261 = 8'h5a == _T_47[7:0] ? 4'h0 : _GEN_260; // @[Filter.scala 165:86]
  wire [3:0] _GEN_262 = 8'h5b == _T_47[7:0] ? 4'h0 : _GEN_261; // @[Filter.scala 165:86]
  wire [3:0] _GEN_263 = 8'h5c == _T_47[7:0] ? 4'h0 : _GEN_262; // @[Filter.scala 165:86]
  wire [3:0] _GEN_264 = 8'h5d == _T_47[7:0] ? 4'h0 : _GEN_263; // @[Filter.scala 165:86]
  wire [3:0] _GEN_265 = 8'h5e == _T_47[7:0] ? 4'h0 : _GEN_264; // @[Filter.scala 165:86]
  wire [3:0] _GEN_266 = 8'h5f == _T_47[7:0] ? 4'h0 : _GEN_265; // @[Filter.scala 165:86]
  wire [3:0] _GEN_267 = 8'h60 == _T_47[7:0] ? 4'h0 : _GEN_266; // @[Filter.scala 165:86]
  wire [3:0] _GEN_268 = 8'h61 == _T_47[7:0] ? 4'h0 : _GEN_267; // @[Filter.scala 165:86]
  wire [3:0] _GEN_269 = 8'h62 == _T_47[7:0] ? 4'h0 : _GEN_268; // @[Filter.scala 165:86]
  wire [3:0] _GEN_270 = 8'h63 == _T_47[7:0] ? 4'h0 : _GEN_269; // @[Filter.scala 165:86]
  wire [3:0] _GEN_271 = 8'h64 == _T_47[7:0] ? 4'h0 : _GEN_270; // @[Filter.scala 165:86]
  wire [3:0] _GEN_272 = 8'h65 == _T_47[7:0] ? 4'h0 : _GEN_271; // @[Filter.scala 165:86]
  wire [3:0] _GEN_273 = 8'h66 == _T_47[7:0] ? 4'h0 : _GEN_272; // @[Filter.scala 165:86]
  wire [3:0] _GEN_274 = 8'h67 == _T_47[7:0] ? 4'h0 : _GEN_273; // @[Filter.scala 165:86]
  wire [3:0] _GEN_275 = 8'h68 == _T_47[7:0] ? 4'hf : _GEN_274; // @[Filter.scala 165:86]
  wire [3:0] _GEN_276 = 8'h69 == _T_47[7:0] ? 4'hf : _GEN_275; // @[Filter.scala 165:86]
  wire [3:0] _GEN_277 = 8'h6a == _T_47[7:0] ? 4'hf : _GEN_276; // @[Filter.scala 165:86]
  wire [3:0] _GEN_278 = 8'h6b == _T_47[7:0] ? 4'hf : _GEN_277; // @[Filter.scala 165:86]
  wire [3:0] _GEN_279 = 8'h6c == _T_47[7:0] ? 4'hf : _GEN_278; // @[Filter.scala 165:86]
  wire [3:0] _GEN_280 = 8'h6d == _T_47[7:0] ? 4'hf : _GEN_279; // @[Filter.scala 165:86]
  wire [3:0] _GEN_281 = 8'h6e == _T_47[7:0] ? 4'hf : _GEN_280; // @[Filter.scala 165:86]
  wire [3:0] _GEN_282 = 8'h6f == _T_47[7:0] ? 4'hf : _GEN_281; // @[Filter.scala 165:86]
  wire [3:0] _GEN_283 = 8'h70 == _T_47[7:0] ? 4'h0 : _GEN_282; // @[Filter.scala 165:86]
  wire [3:0] _GEN_284 = 8'h71 == _T_47[7:0] ? 4'h0 : _GEN_283; // @[Filter.scala 165:86]
  wire [3:0] _GEN_285 = 8'h72 == _T_47[7:0] ? 4'h0 : _GEN_284; // @[Filter.scala 165:86]
  wire [3:0] _GEN_286 = 8'h73 == _T_47[7:0] ? 4'h0 : _GEN_285; // @[Filter.scala 165:86]
  wire [3:0] _GEN_287 = 8'h74 == _T_47[7:0] ? 4'h0 : _GEN_286; // @[Filter.scala 165:86]
  wire [3:0] _GEN_288 = 8'h75 == _T_47[7:0] ? 4'h0 : _GEN_287; // @[Filter.scala 165:86]
  wire [3:0] _GEN_289 = 8'h76 == _T_47[7:0] ? 4'h0 : _GEN_288; // @[Filter.scala 165:86]
  wire [3:0] _GEN_290 = 8'h77 == _T_47[7:0] ? 4'h0 : _GEN_289; // @[Filter.scala 165:86]
  wire [3:0] _GEN_291 = 8'h78 == _T_47[7:0] ? 4'hf : _GEN_290; // @[Filter.scala 165:86]
  wire [3:0] _GEN_292 = 8'h79 == _T_47[7:0] ? 4'hf : _GEN_291; // @[Filter.scala 165:86]
  wire [3:0] _GEN_293 = 8'h7a == _T_47[7:0] ? 4'hf : _GEN_292; // @[Filter.scala 165:86]
  wire [3:0] _GEN_294 = 8'h7b == _T_47[7:0] ? 4'hf : _GEN_293; // @[Filter.scala 165:86]
  wire [3:0] _GEN_295 = 8'h7c == _T_47[7:0] ? 4'hf : _GEN_294; // @[Filter.scala 165:86]
  wire [3:0] _GEN_296 = 8'h7d == _T_47[7:0] ? 4'hf : _GEN_295; // @[Filter.scala 165:86]
  wire [3:0] _GEN_297 = 8'h7e == _T_47[7:0] ? 4'hf : _GEN_296; // @[Filter.scala 165:86]
  wire [3:0] _GEN_298 = 8'h7f == _T_47[7:0] ? 4'hf : _GEN_297; // @[Filter.scala 165:86]
  wire [3:0] _GEN_299 = 8'h80 == _T_47[7:0] ? 4'h0 : _GEN_298; // @[Filter.scala 165:86]
  wire [3:0] _GEN_300 = 8'h81 == _T_47[7:0] ? 4'h0 : _GEN_299; // @[Filter.scala 165:86]
  wire [3:0] _GEN_301 = 8'h82 == _T_47[7:0] ? 4'h0 : _GEN_300; // @[Filter.scala 165:86]
  wire [3:0] _GEN_302 = 8'h83 == _T_47[7:0] ? 4'h0 : _GEN_301; // @[Filter.scala 165:86]
  wire [3:0] _GEN_303 = 8'h84 == _T_47[7:0] ? 4'h0 : _GEN_302; // @[Filter.scala 165:86]
  wire [3:0] _GEN_304 = 8'h85 == _T_47[7:0] ? 4'h0 : _GEN_303; // @[Filter.scala 165:86]
  wire [3:0] _GEN_305 = 8'h86 == _T_47[7:0] ? 4'h0 : _GEN_304; // @[Filter.scala 165:86]
  wire [3:0] _GEN_306 = 8'h87 == _T_47[7:0] ? 4'h0 : _GEN_305; // @[Filter.scala 165:86]
  wire [3:0] _GEN_307 = 8'h88 == _T_47[7:0] ? 4'hf : _GEN_306; // @[Filter.scala 165:86]
  wire [3:0] _GEN_308 = 8'h89 == _T_47[7:0] ? 4'hf : _GEN_307; // @[Filter.scala 165:86]
  wire [3:0] _GEN_309 = 8'h8a == _T_47[7:0] ? 4'hf : _GEN_308; // @[Filter.scala 165:86]
  wire [3:0] _GEN_310 = 8'h8b == _T_47[7:0] ? 4'hf : _GEN_309; // @[Filter.scala 165:86]
  wire [3:0] _GEN_311 = 8'h8c == _T_47[7:0] ? 4'hf : _GEN_310; // @[Filter.scala 165:86]
  wire [3:0] _GEN_312 = 8'h8d == _T_47[7:0] ? 4'hf : _GEN_311; // @[Filter.scala 165:86]
  wire [3:0] _GEN_313 = 8'h8e == _T_47[7:0] ? 4'hf : _GEN_312; // @[Filter.scala 165:86]
  wire [3:0] _GEN_314 = 8'h8f == _T_47[7:0] ? 4'hf : _GEN_313; // @[Filter.scala 165:86]
  wire [3:0] _GEN_315 = 8'h90 == _T_47[7:0] ? 4'h0 : _GEN_314; // @[Filter.scala 165:86]
  wire [3:0] _GEN_316 = 8'h91 == _T_47[7:0] ? 4'h0 : _GEN_315; // @[Filter.scala 165:86]
  wire [3:0] _GEN_317 = 8'h92 == _T_47[7:0] ? 4'h0 : _GEN_316; // @[Filter.scala 165:86]
  wire [3:0] _GEN_318 = 8'h93 == _T_47[7:0] ? 4'h0 : _GEN_317; // @[Filter.scala 165:86]
  wire [3:0] _GEN_319 = 8'h94 == _T_47[7:0] ? 4'h0 : _GEN_318; // @[Filter.scala 165:86]
  wire [3:0] _GEN_320 = 8'h95 == _T_47[7:0] ? 4'h0 : _GEN_319; // @[Filter.scala 165:86]
  wire [3:0] _GEN_321 = 8'h96 == _T_47[7:0] ? 4'h0 : _GEN_320; // @[Filter.scala 165:86]
  wire [3:0] _GEN_322 = 8'h97 == _T_47[7:0] ? 4'h0 : _GEN_321; // @[Filter.scala 165:86]
  wire [3:0] _GEN_323 = 8'h98 == _T_47[7:0] ? 4'hf : _GEN_322; // @[Filter.scala 165:86]
  wire [3:0] _GEN_324 = 8'h99 == _T_47[7:0] ? 4'hf : _GEN_323; // @[Filter.scala 165:86]
  wire [3:0] _GEN_325 = 8'h9a == _T_47[7:0] ? 4'hf : _GEN_324; // @[Filter.scala 165:86]
  wire [3:0] _GEN_326 = 8'h9b == _T_47[7:0] ? 4'hf : _GEN_325; // @[Filter.scala 165:86]
  wire [3:0] _GEN_327 = 8'h9c == _T_47[7:0] ? 4'hf : _GEN_326; // @[Filter.scala 165:86]
  wire [3:0] _GEN_328 = 8'h9d == _T_47[7:0] ? 4'hf : _GEN_327; // @[Filter.scala 165:86]
  wire [3:0] _GEN_329 = 8'h9e == _T_47[7:0] ? 4'hf : _GEN_328; // @[Filter.scala 165:86]
  wire [3:0] _GEN_330 = 8'h9f == _T_47[7:0] ? 4'hf : _GEN_329; // @[Filter.scala 165:86]
  wire [3:0] _GEN_331 = 8'ha0 == _T_47[7:0] ? 4'h0 : _GEN_330; // @[Filter.scala 165:86]
  wire [3:0] _GEN_332 = 8'ha1 == _T_47[7:0] ? 4'h0 : _GEN_331; // @[Filter.scala 165:86]
  wire [3:0] _GEN_333 = 8'ha2 == _T_47[7:0] ? 4'h0 : _GEN_332; // @[Filter.scala 165:86]
  wire [3:0] _GEN_334 = 8'ha3 == _T_47[7:0] ? 4'h0 : _GEN_333; // @[Filter.scala 165:86]
  wire [3:0] _GEN_335 = 8'ha4 == _T_47[7:0] ? 4'h0 : _GEN_334; // @[Filter.scala 165:86]
  wire [3:0] _GEN_336 = 8'ha5 == _T_47[7:0] ? 4'h0 : _GEN_335; // @[Filter.scala 165:86]
  wire [3:0] _GEN_337 = 8'ha6 == _T_47[7:0] ? 4'h0 : _GEN_336; // @[Filter.scala 165:86]
  wire [3:0] _GEN_338 = 8'ha7 == _T_47[7:0] ? 4'h0 : _GEN_337; // @[Filter.scala 165:86]
  wire [3:0] _GEN_339 = 8'ha8 == _T_47[7:0] ? 4'hf : _GEN_338; // @[Filter.scala 165:86]
  wire [3:0] _GEN_340 = 8'ha9 == _T_47[7:0] ? 4'hf : _GEN_339; // @[Filter.scala 165:86]
  wire [3:0] _GEN_341 = 8'haa == _T_47[7:0] ? 4'hf : _GEN_340; // @[Filter.scala 165:86]
  wire [3:0] _GEN_342 = 8'hab == _T_47[7:0] ? 4'hf : _GEN_341; // @[Filter.scala 165:86]
  wire [3:0] _GEN_343 = 8'hac == _T_47[7:0] ? 4'hf : _GEN_342; // @[Filter.scala 165:86]
  wire [3:0] _GEN_344 = 8'had == _T_47[7:0] ? 4'hf : _GEN_343; // @[Filter.scala 165:86]
  wire [3:0] _GEN_345 = 8'hae == _T_47[7:0] ? 4'hf : _GEN_344; // @[Filter.scala 165:86]
  wire [3:0] _GEN_346 = 8'haf == _T_47[7:0] ? 4'hf : _GEN_345; // @[Filter.scala 165:86]
  wire [3:0] _GEN_347 = 8'hb0 == _T_47[7:0] ? 4'h0 : _GEN_346; // @[Filter.scala 165:86]
  wire [3:0] _GEN_348 = 8'hb1 == _T_47[7:0] ? 4'h0 : _GEN_347; // @[Filter.scala 165:86]
  wire [3:0] _GEN_349 = 8'hb2 == _T_47[7:0] ? 4'h0 : _GEN_348; // @[Filter.scala 165:86]
  wire [3:0] _GEN_350 = 8'hb3 == _T_47[7:0] ? 4'h0 : _GEN_349; // @[Filter.scala 165:86]
  wire [3:0] _GEN_351 = 8'hb4 == _T_47[7:0] ? 4'h0 : _GEN_350; // @[Filter.scala 165:86]
  wire [3:0] _GEN_352 = 8'hb5 == _T_47[7:0] ? 4'h0 : _GEN_351; // @[Filter.scala 165:86]
  wire [3:0] _GEN_353 = 8'hb6 == _T_47[7:0] ? 4'h0 : _GEN_352; // @[Filter.scala 165:86]
  wire [3:0] _GEN_354 = 8'hb7 == _T_47[7:0] ? 4'h0 : _GEN_353; // @[Filter.scala 165:86]
  wire [3:0] _GEN_355 = 8'hb8 == _T_47[7:0] ? 4'hf : _GEN_354; // @[Filter.scala 165:86]
  wire [3:0] _GEN_356 = 8'hb9 == _T_47[7:0] ? 4'hf : _GEN_355; // @[Filter.scala 165:86]
  wire [3:0] _GEN_357 = 8'hba == _T_47[7:0] ? 4'hf : _GEN_356; // @[Filter.scala 165:86]
  wire [3:0] _GEN_358 = 8'hbb == _T_47[7:0] ? 4'hf : _GEN_357; // @[Filter.scala 165:86]
  wire [3:0] _GEN_359 = 8'hbc == _T_47[7:0] ? 4'hf : _GEN_358; // @[Filter.scala 165:86]
  wire [3:0] _GEN_360 = 8'hbd == _T_47[7:0] ? 4'hf : _GEN_359; // @[Filter.scala 165:86]
  wire [3:0] _GEN_361 = 8'hbe == _T_47[7:0] ? 4'hf : _GEN_360; // @[Filter.scala 165:86]
  wire [3:0] _GEN_362 = 8'hbf == _T_47[7:0] ? 4'hf : _GEN_361; // @[Filter.scala 165:86]
  wire [4:0] _GEN_18986 = {{1'd0}, _GEN_362}; // @[Filter.scala 165:86]
  wire [8:0] _T_49 = _GEN_18986 * 5'h14; // @[Filter.scala 165:86]
  wire [3:0] _GEN_459 = 8'h60 == _T_47[7:0] ? 4'hf : 4'h0; // @[Filter.scala 165:126]
  wire [3:0] _GEN_460 = 8'h61 == _T_47[7:0] ? 4'hf : _GEN_459; // @[Filter.scala 165:126]
  wire [3:0] _GEN_461 = 8'h62 == _T_47[7:0] ? 4'hf : _GEN_460; // @[Filter.scala 165:126]
  wire [3:0] _GEN_462 = 8'h63 == _T_47[7:0] ? 4'hf : _GEN_461; // @[Filter.scala 165:126]
  wire [3:0] _GEN_463 = 8'h64 == _T_47[7:0] ? 4'hf : _GEN_462; // @[Filter.scala 165:126]
  wire [3:0] _GEN_464 = 8'h65 == _T_47[7:0] ? 4'hf : _GEN_463; // @[Filter.scala 165:126]
  wire [3:0] _GEN_465 = 8'h66 == _T_47[7:0] ? 4'hf : _GEN_464; // @[Filter.scala 165:126]
  wire [3:0] _GEN_466 = 8'h67 == _T_47[7:0] ? 4'hf : _GEN_465; // @[Filter.scala 165:126]
  wire [3:0] _GEN_467 = 8'h68 == _T_47[7:0] ? 4'hf : _GEN_466; // @[Filter.scala 165:126]
  wire [3:0] _GEN_468 = 8'h69 == _T_47[7:0] ? 4'hf : _GEN_467; // @[Filter.scala 165:126]
  wire [3:0] _GEN_469 = 8'h6a == _T_47[7:0] ? 4'hf : _GEN_468; // @[Filter.scala 165:126]
  wire [3:0] _GEN_470 = 8'h6b == _T_47[7:0] ? 4'hf : _GEN_469; // @[Filter.scala 165:126]
  wire [3:0] _GEN_471 = 8'h6c == _T_47[7:0] ? 4'hf : _GEN_470; // @[Filter.scala 165:126]
  wire [3:0] _GEN_472 = 8'h6d == _T_47[7:0] ? 4'hf : _GEN_471; // @[Filter.scala 165:126]
  wire [3:0] _GEN_473 = 8'h6e == _T_47[7:0] ? 4'hf : _GEN_472; // @[Filter.scala 165:126]
  wire [3:0] _GEN_474 = 8'h6f == _T_47[7:0] ? 4'hf : _GEN_473; // @[Filter.scala 165:126]
  wire [3:0] _GEN_475 = 8'h70 == _T_47[7:0] ? 4'hf : _GEN_474; // @[Filter.scala 165:126]
  wire [3:0] _GEN_476 = 8'h71 == _T_47[7:0] ? 4'hf : _GEN_475; // @[Filter.scala 165:126]
  wire [3:0] _GEN_477 = 8'h72 == _T_47[7:0] ? 4'hf : _GEN_476; // @[Filter.scala 165:126]
  wire [3:0] _GEN_478 = 8'h73 == _T_47[7:0] ? 4'hf : _GEN_477; // @[Filter.scala 165:126]
  wire [3:0] _GEN_479 = 8'h74 == _T_47[7:0] ? 4'hf : _GEN_478; // @[Filter.scala 165:126]
  wire [3:0] _GEN_480 = 8'h75 == _T_47[7:0] ? 4'hf : _GEN_479; // @[Filter.scala 165:126]
  wire [3:0] _GEN_481 = 8'h76 == _T_47[7:0] ? 4'hf : _GEN_480; // @[Filter.scala 165:126]
  wire [3:0] _GEN_482 = 8'h77 == _T_47[7:0] ? 4'hf : _GEN_481; // @[Filter.scala 165:126]
  wire [3:0] _GEN_483 = 8'h78 == _T_47[7:0] ? 4'hf : _GEN_482; // @[Filter.scala 165:126]
  wire [3:0] _GEN_484 = 8'h79 == _T_47[7:0] ? 4'hf : _GEN_483; // @[Filter.scala 165:126]
  wire [3:0] _GEN_485 = 8'h7a == _T_47[7:0] ? 4'hf : _GEN_484; // @[Filter.scala 165:126]
  wire [3:0] _GEN_486 = 8'h7b == _T_47[7:0] ? 4'hf : _GEN_485; // @[Filter.scala 165:126]
  wire [3:0] _GEN_487 = 8'h7c == _T_47[7:0] ? 4'hf : _GEN_486; // @[Filter.scala 165:126]
  wire [3:0] _GEN_488 = 8'h7d == _T_47[7:0] ? 4'hf : _GEN_487; // @[Filter.scala 165:126]
  wire [3:0] _GEN_489 = 8'h7e == _T_47[7:0] ? 4'hf : _GEN_488; // @[Filter.scala 165:126]
  wire [3:0] _GEN_490 = 8'h7f == _T_47[7:0] ? 4'hf : _GEN_489; // @[Filter.scala 165:126]
  wire [3:0] _GEN_491 = 8'h80 == _T_47[7:0] ? 4'hf : _GEN_490; // @[Filter.scala 165:126]
  wire [3:0] _GEN_492 = 8'h81 == _T_47[7:0] ? 4'hf : _GEN_491; // @[Filter.scala 165:126]
  wire [3:0] _GEN_493 = 8'h82 == _T_47[7:0] ? 4'hf : _GEN_492; // @[Filter.scala 165:126]
  wire [3:0] _GEN_494 = 8'h83 == _T_47[7:0] ? 4'hf : _GEN_493; // @[Filter.scala 165:126]
  wire [3:0] _GEN_495 = 8'h84 == _T_47[7:0] ? 4'hf : _GEN_494; // @[Filter.scala 165:126]
  wire [3:0] _GEN_496 = 8'h85 == _T_47[7:0] ? 4'hf : _GEN_495; // @[Filter.scala 165:126]
  wire [3:0] _GEN_497 = 8'h86 == _T_47[7:0] ? 4'hf : _GEN_496; // @[Filter.scala 165:126]
  wire [3:0] _GEN_498 = 8'h87 == _T_47[7:0] ? 4'hf : _GEN_497; // @[Filter.scala 165:126]
  wire [3:0] _GEN_499 = 8'h88 == _T_47[7:0] ? 4'hf : _GEN_498; // @[Filter.scala 165:126]
  wire [3:0] _GEN_500 = 8'h89 == _T_47[7:0] ? 4'hf : _GEN_499; // @[Filter.scala 165:126]
  wire [3:0] _GEN_501 = 8'h8a == _T_47[7:0] ? 4'hf : _GEN_500; // @[Filter.scala 165:126]
  wire [3:0] _GEN_502 = 8'h8b == _T_47[7:0] ? 4'hf : _GEN_501; // @[Filter.scala 165:126]
  wire [3:0] _GEN_503 = 8'h8c == _T_47[7:0] ? 4'hf : _GEN_502; // @[Filter.scala 165:126]
  wire [3:0] _GEN_504 = 8'h8d == _T_47[7:0] ? 4'hf : _GEN_503; // @[Filter.scala 165:126]
  wire [3:0] _GEN_505 = 8'h8e == _T_47[7:0] ? 4'hf : _GEN_504; // @[Filter.scala 165:126]
  wire [3:0] _GEN_506 = 8'h8f == _T_47[7:0] ? 4'hf : _GEN_505; // @[Filter.scala 165:126]
  wire [3:0] _GEN_507 = 8'h90 == _T_47[7:0] ? 4'hf : _GEN_506; // @[Filter.scala 165:126]
  wire [3:0] _GEN_508 = 8'h91 == _T_47[7:0] ? 4'hf : _GEN_507; // @[Filter.scala 165:126]
  wire [3:0] _GEN_509 = 8'h92 == _T_47[7:0] ? 4'hf : _GEN_508; // @[Filter.scala 165:126]
  wire [3:0] _GEN_510 = 8'h93 == _T_47[7:0] ? 4'hf : _GEN_509; // @[Filter.scala 165:126]
  wire [3:0] _GEN_511 = 8'h94 == _T_47[7:0] ? 4'hf : _GEN_510; // @[Filter.scala 165:126]
  wire [3:0] _GEN_512 = 8'h95 == _T_47[7:0] ? 4'hf : _GEN_511; // @[Filter.scala 165:126]
  wire [3:0] _GEN_513 = 8'h96 == _T_47[7:0] ? 4'hf : _GEN_512; // @[Filter.scala 165:126]
  wire [3:0] _GEN_514 = 8'h97 == _T_47[7:0] ? 4'hf : _GEN_513; // @[Filter.scala 165:126]
  wire [3:0] _GEN_515 = 8'h98 == _T_47[7:0] ? 4'hf : _GEN_514; // @[Filter.scala 165:126]
  wire [3:0] _GEN_516 = 8'h99 == _T_47[7:0] ? 4'hf : _GEN_515; // @[Filter.scala 165:126]
  wire [3:0] _GEN_517 = 8'h9a == _T_47[7:0] ? 4'hf : _GEN_516; // @[Filter.scala 165:126]
  wire [3:0] _GEN_518 = 8'h9b == _T_47[7:0] ? 4'hf : _GEN_517; // @[Filter.scala 165:126]
  wire [3:0] _GEN_519 = 8'h9c == _T_47[7:0] ? 4'hf : _GEN_518; // @[Filter.scala 165:126]
  wire [3:0] _GEN_520 = 8'h9d == _T_47[7:0] ? 4'hf : _GEN_519; // @[Filter.scala 165:126]
  wire [3:0] _GEN_521 = 8'h9e == _T_47[7:0] ? 4'hf : _GEN_520; // @[Filter.scala 165:126]
  wire [3:0] _GEN_522 = 8'h9f == _T_47[7:0] ? 4'hf : _GEN_521; // @[Filter.scala 165:126]
  wire [3:0] _GEN_523 = 8'ha0 == _T_47[7:0] ? 4'hf : _GEN_522; // @[Filter.scala 165:126]
  wire [3:0] _GEN_524 = 8'ha1 == _T_47[7:0] ? 4'hf : _GEN_523; // @[Filter.scala 165:126]
  wire [3:0] _GEN_525 = 8'ha2 == _T_47[7:0] ? 4'hf : _GEN_524; // @[Filter.scala 165:126]
  wire [3:0] _GEN_526 = 8'ha3 == _T_47[7:0] ? 4'hf : _GEN_525; // @[Filter.scala 165:126]
  wire [3:0] _GEN_527 = 8'ha4 == _T_47[7:0] ? 4'hf : _GEN_526; // @[Filter.scala 165:126]
  wire [3:0] _GEN_528 = 8'ha5 == _T_47[7:0] ? 4'hf : _GEN_527; // @[Filter.scala 165:126]
  wire [3:0] _GEN_529 = 8'ha6 == _T_47[7:0] ? 4'hf : _GEN_528; // @[Filter.scala 165:126]
  wire [3:0] _GEN_530 = 8'ha7 == _T_47[7:0] ? 4'hf : _GEN_529; // @[Filter.scala 165:126]
  wire [3:0] _GEN_531 = 8'ha8 == _T_47[7:0] ? 4'hf : _GEN_530; // @[Filter.scala 165:126]
  wire [3:0] _GEN_532 = 8'ha9 == _T_47[7:0] ? 4'hf : _GEN_531; // @[Filter.scala 165:126]
  wire [3:0] _GEN_533 = 8'haa == _T_47[7:0] ? 4'hf : _GEN_532; // @[Filter.scala 165:126]
  wire [3:0] _GEN_534 = 8'hab == _T_47[7:0] ? 4'hf : _GEN_533; // @[Filter.scala 165:126]
  wire [3:0] _GEN_535 = 8'hac == _T_47[7:0] ? 4'hf : _GEN_534; // @[Filter.scala 165:126]
  wire [3:0] _GEN_536 = 8'had == _T_47[7:0] ? 4'hf : _GEN_535; // @[Filter.scala 165:126]
  wire [3:0] _GEN_537 = 8'hae == _T_47[7:0] ? 4'hf : _GEN_536; // @[Filter.scala 165:126]
  wire [3:0] _GEN_538 = 8'haf == _T_47[7:0] ? 4'hf : _GEN_537; // @[Filter.scala 165:126]
  wire [3:0] _GEN_539 = 8'hb0 == _T_47[7:0] ? 4'hf : _GEN_538; // @[Filter.scala 165:126]
  wire [3:0] _GEN_540 = 8'hb1 == _T_47[7:0] ? 4'hf : _GEN_539; // @[Filter.scala 165:126]
  wire [3:0] _GEN_541 = 8'hb2 == _T_47[7:0] ? 4'hf : _GEN_540; // @[Filter.scala 165:126]
  wire [3:0] _GEN_542 = 8'hb3 == _T_47[7:0] ? 4'hf : _GEN_541; // @[Filter.scala 165:126]
  wire [3:0] _GEN_543 = 8'hb4 == _T_47[7:0] ? 4'hf : _GEN_542; // @[Filter.scala 165:126]
  wire [3:0] _GEN_544 = 8'hb5 == _T_47[7:0] ? 4'hf : _GEN_543; // @[Filter.scala 165:126]
  wire [3:0] _GEN_545 = 8'hb6 == _T_47[7:0] ? 4'hf : _GEN_544; // @[Filter.scala 165:126]
  wire [3:0] _GEN_546 = 8'hb7 == _T_47[7:0] ? 4'hf : _GEN_545; // @[Filter.scala 165:126]
  wire [3:0] _GEN_547 = 8'hb8 == _T_47[7:0] ? 4'hf : _GEN_546; // @[Filter.scala 165:126]
  wire [3:0] _GEN_548 = 8'hb9 == _T_47[7:0] ? 4'hf : _GEN_547; // @[Filter.scala 165:126]
  wire [3:0] _GEN_549 = 8'hba == _T_47[7:0] ? 4'hf : _GEN_548; // @[Filter.scala 165:126]
  wire [3:0] _GEN_550 = 8'hbb == _T_47[7:0] ? 4'hf : _GEN_549; // @[Filter.scala 165:126]
  wire [3:0] _GEN_551 = 8'hbc == _T_47[7:0] ? 4'hf : _GEN_550; // @[Filter.scala 165:126]
  wire [3:0] _GEN_552 = 8'hbd == _T_47[7:0] ? 4'hf : _GEN_551; // @[Filter.scala 165:126]
  wire [3:0] _GEN_553 = 8'hbe == _T_47[7:0] ? 4'hf : _GEN_552; // @[Filter.scala 165:126]
  wire [3:0] _GEN_554 = 8'hbf == _T_47[7:0] ? 4'hf : _GEN_553; // @[Filter.scala 165:126]
  wire [6:0] _GEN_18988 = {{3'd0}, _GEN_554}; // @[Filter.scala 165:126]
  wire [10:0] _T_54 = _GEN_18988 * 7'h46; // @[Filter.scala 165:126]
  wire [10:0] _GEN_18989 = {{2'd0}, _T_49}; // @[Filter.scala 165:93]
  wire [10:0] _T_56 = _GEN_18989 + _T_54; // @[Filter.scala 165:93]
  wire [3:0] _GEN_563 = 8'h8 == _T_47[7:0] ? 4'hf : 4'h0; // @[Filter.scala 165:166]
  wire [3:0] _GEN_564 = 8'h9 == _T_47[7:0] ? 4'hf : _GEN_563; // @[Filter.scala 165:166]
  wire [3:0] _GEN_565 = 8'ha == _T_47[7:0] ? 4'hf : _GEN_564; // @[Filter.scala 165:166]
  wire [3:0] _GEN_566 = 8'hb == _T_47[7:0] ? 4'hf : _GEN_565; // @[Filter.scala 165:166]
  wire [3:0] _GEN_567 = 8'hc == _T_47[7:0] ? 4'hf : _GEN_566; // @[Filter.scala 165:166]
  wire [3:0] _GEN_568 = 8'hd == _T_47[7:0] ? 4'hf : _GEN_567; // @[Filter.scala 165:166]
  wire [3:0] _GEN_569 = 8'he == _T_47[7:0] ? 4'hf : _GEN_568; // @[Filter.scala 165:166]
  wire [3:0] _GEN_570 = 8'hf == _T_47[7:0] ? 4'hf : _GEN_569; // @[Filter.scala 165:166]
  wire [3:0] _GEN_571 = 8'h10 == _T_47[7:0] ? 4'h0 : _GEN_570; // @[Filter.scala 165:166]
  wire [3:0] _GEN_572 = 8'h11 == _T_47[7:0] ? 4'h0 : _GEN_571; // @[Filter.scala 165:166]
  wire [3:0] _GEN_573 = 8'h12 == _T_47[7:0] ? 4'h0 : _GEN_572; // @[Filter.scala 165:166]
  wire [3:0] _GEN_574 = 8'h13 == _T_47[7:0] ? 4'h0 : _GEN_573; // @[Filter.scala 165:166]
  wire [3:0] _GEN_575 = 8'h14 == _T_47[7:0] ? 4'h0 : _GEN_574; // @[Filter.scala 165:166]
  wire [3:0] _GEN_576 = 8'h15 == _T_47[7:0] ? 4'h0 : _GEN_575; // @[Filter.scala 165:166]
  wire [3:0] _GEN_577 = 8'h16 == _T_47[7:0] ? 4'h0 : _GEN_576; // @[Filter.scala 165:166]
  wire [3:0] _GEN_578 = 8'h17 == _T_47[7:0] ? 4'h0 : _GEN_577; // @[Filter.scala 165:166]
  wire [3:0] _GEN_579 = 8'h18 == _T_47[7:0] ? 4'hf : _GEN_578; // @[Filter.scala 165:166]
  wire [3:0] _GEN_580 = 8'h19 == _T_47[7:0] ? 4'hf : _GEN_579; // @[Filter.scala 165:166]
  wire [3:0] _GEN_581 = 8'h1a == _T_47[7:0] ? 4'hf : _GEN_580; // @[Filter.scala 165:166]
  wire [3:0] _GEN_582 = 8'h1b == _T_47[7:0] ? 4'hf : _GEN_581; // @[Filter.scala 165:166]
  wire [3:0] _GEN_583 = 8'h1c == _T_47[7:0] ? 4'hf : _GEN_582; // @[Filter.scala 165:166]
  wire [3:0] _GEN_584 = 8'h1d == _T_47[7:0] ? 4'hf : _GEN_583; // @[Filter.scala 165:166]
  wire [3:0] _GEN_585 = 8'h1e == _T_47[7:0] ? 4'hf : _GEN_584; // @[Filter.scala 165:166]
  wire [3:0] _GEN_586 = 8'h1f == _T_47[7:0] ? 4'hf : _GEN_585; // @[Filter.scala 165:166]
  wire [3:0] _GEN_587 = 8'h20 == _T_47[7:0] ? 4'h0 : _GEN_586; // @[Filter.scala 165:166]
  wire [3:0] _GEN_588 = 8'h21 == _T_47[7:0] ? 4'h0 : _GEN_587; // @[Filter.scala 165:166]
  wire [3:0] _GEN_589 = 8'h22 == _T_47[7:0] ? 4'h0 : _GEN_588; // @[Filter.scala 165:166]
  wire [3:0] _GEN_590 = 8'h23 == _T_47[7:0] ? 4'h0 : _GEN_589; // @[Filter.scala 165:166]
  wire [3:0] _GEN_591 = 8'h24 == _T_47[7:0] ? 4'h0 : _GEN_590; // @[Filter.scala 165:166]
  wire [3:0] _GEN_592 = 8'h25 == _T_47[7:0] ? 4'h0 : _GEN_591; // @[Filter.scala 165:166]
  wire [3:0] _GEN_593 = 8'h26 == _T_47[7:0] ? 4'h0 : _GEN_592; // @[Filter.scala 165:166]
  wire [3:0] _GEN_594 = 8'h27 == _T_47[7:0] ? 4'h0 : _GEN_593; // @[Filter.scala 165:166]
  wire [3:0] _GEN_595 = 8'h28 == _T_47[7:0] ? 4'hf : _GEN_594; // @[Filter.scala 165:166]
  wire [3:0] _GEN_596 = 8'h29 == _T_47[7:0] ? 4'hf : _GEN_595; // @[Filter.scala 165:166]
  wire [3:0] _GEN_597 = 8'h2a == _T_47[7:0] ? 4'hf : _GEN_596; // @[Filter.scala 165:166]
  wire [3:0] _GEN_598 = 8'h2b == _T_47[7:0] ? 4'hf : _GEN_597; // @[Filter.scala 165:166]
  wire [3:0] _GEN_599 = 8'h2c == _T_47[7:0] ? 4'hf : _GEN_598; // @[Filter.scala 165:166]
  wire [3:0] _GEN_600 = 8'h2d == _T_47[7:0] ? 4'hf : _GEN_599; // @[Filter.scala 165:166]
  wire [3:0] _GEN_601 = 8'h2e == _T_47[7:0] ? 4'hf : _GEN_600; // @[Filter.scala 165:166]
  wire [3:0] _GEN_602 = 8'h2f == _T_47[7:0] ? 4'hf : _GEN_601; // @[Filter.scala 165:166]
  wire [3:0] _GEN_603 = 8'h30 == _T_47[7:0] ? 4'h0 : _GEN_602; // @[Filter.scala 165:166]
  wire [3:0] _GEN_604 = 8'h31 == _T_47[7:0] ? 4'h0 : _GEN_603; // @[Filter.scala 165:166]
  wire [3:0] _GEN_605 = 8'h32 == _T_47[7:0] ? 4'h0 : _GEN_604; // @[Filter.scala 165:166]
  wire [3:0] _GEN_606 = 8'h33 == _T_47[7:0] ? 4'h0 : _GEN_605; // @[Filter.scala 165:166]
  wire [3:0] _GEN_607 = 8'h34 == _T_47[7:0] ? 4'h0 : _GEN_606; // @[Filter.scala 165:166]
  wire [3:0] _GEN_608 = 8'h35 == _T_47[7:0] ? 4'h0 : _GEN_607; // @[Filter.scala 165:166]
  wire [3:0] _GEN_609 = 8'h36 == _T_47[7:0] ? 4'h0 : _GEN_608; // @[Filter.scala 165:166]
  wire [3:0] _GEN_610 = 8'h37 == _T_47[7:0] ? 4'h0 : _GEN_609; // @[Filter.scala 165:166]
  wire [3:0] _GEN_611 = 8'h38 == _T_47[7:0] ? 4'hf : _GEN_610; // @[Filter.scala 165:166]
  wire [3:0] _GEN_612 = 8'h39 == _T_47[7:0] ? 4'hf : _GEN_611; // @[Filter.scala 165:166]
  wire [3:0] _GEN_613 = 8'h3a == _T_47[7:0] ? 4'hf : _GEN_612; // @[Filter.scala 165:166]
  wire [3:0] _GEN_614 = 8'h3b == _T_47[7:0] ? 4'hf : _GEN_613; // @[Filter.scala 165:166]
  wire [3:0] _GEN_615 = 8'h3c == _T_47[7:0] ? 4'hf : _GEN_614; // @[Filter.scala 165:166]
  wire [3:0] _GEN_616 = 8'h3d == _T_47[7:0] ? 4'hf : _GEN_615; // @[Filter.scala 165:166]
  wire [3:0] _GEN_617 = 8'h3e == _T_47[7:0] ? 4'hf : _GEN_616; // @[Filter.scala 165:166]
  wire [3:0] _GEN_618 = 8'h3f == _T_47[7:0] ? 4'hf : _GEN_617; // @[Filter.scala 165:166]
  wire [3:0] _GEN_619 = 8'h40 == _T_47[7:0] ? 4'h0 : _GEN_618; // @[Filter.scala 165:166]
  wire [3:0] _GEN_620 = 8'h41 == _T_47[7:0] ? 4'h0 : _GEN_619; // @[Filter.scala 165:166]
  wire [3:0] _GEN_621 = 8'h42 == _T_47[7:0] ? 4'h0 : _GEN_620; // @[Filter.scala 165:166]
  wire [3:0] _GEN_622 = 8'h43 == _T_47[7:0] ? 4'h0 : _GEN_621; // @[Filter.scala 165:166]
  wire [3:0] _GEN_623 = 8'h44 == _T_47[7:0] ? 4'h0 : _GEN_622; // @[Filter.scala 165:166]
  wire [3:0] _GEN_624 = 8'h45 == _T_47[7:0] ? 4'h0 : _GEN_623; // @[Filter.scala 165:166]
  wire [3:0] _GEN_625 = 8'h46 == _T_47[7:0] ? 4'h0 : _GEN_624; // @[Filter.scala 165:166]
  wire [3:0] _GEN_626 = 8'h47 == _T_47[7:0] ? 4'h0 : _GEN_625; // @[Filter.scala 165:166]
  wire [3:0] _GEN_627 = 8'h48 == _T_47[7:0] ? 4'hf : _GEN_626; // @[Filter.scala 165:166]
  wire [3:0] _GEN_628 = 8'h49 == _T_47[7:0] ? 4'hf : _GEN_627; // @[Filter.scala 165:166]
  wire [3:0] _GEN_629 = 8'h4a == _T_47[7:0] ? 4'hf : _GEN_628; // @[Filter.scala 165:166]
  wire [3:0] _GEN_630 = 8'h4b == _T_47[7:0] ? 4'hf : _GEN_629; // @[Filter.scala 165:166]
  wire [3:0] _GEN_631 = 8'h4c == _T_47[7:0] ? 4'hf : _GEN_630; // @[Filter.scala 165:166]
  wire [3:0] _GEN_632 = 8'h4d == _T_47[7:0] ? 4'hf : _GEN_631; // @[Filter.scala 165:166]
  wire [3:0] _GEN_633 = 8'h4e == _T_47[7:0] ? 4'hf : _GEN_632; // @[Filter.scala 165:166]
  wire [3:0] _GEN_634 = 8'h4f == _T_47[7:0] ? 4'hf : _GEN_633; // @[Filter.scala 165:166]
  wire [3:0] _GEN_635 = 8'h50 == _T_47[7:0] ? 4'h0 : _GEN_634; // @[Filter.scala 165:166]
  wire [3:0] _GEN_636 = 8'h51 == _T_47[7:0] ? 4'h0 : _GEN_635; // @[Filter.scala 165:166]
  wire [3:0] _GEN_637 = 8'h52 == _T_47[7:0] ? 4'h0 : _GEN_636; // @[Filter.scala 165:166]
  wire [3:0] _GEN_638 = 8'h53 == _T_47[7:0] ? 4'h0 : _GEN_637; // @[Filter.scala 165:166]
  wire [3:0] _GEN_639 = 8'h54 == _T_47[7:0] ? 4'h0 : _GEN_638; // @[Filter.scala 165:166]
  wire [3:0] _GEN_640 = 8'h55 == _T_47[7:0] ? 4'h0 : _GEN_639; // @[Filter.scala 165:166]
  wire [3:0] _GEN_641 = 8'h56 == _T_47[7:0] ? 4'h0 : _GEN_640; // @[Filter.scala 165:166]
  wire [3:0] _GEN_642 = 8'h57 == _T_47[7:0] ? 4'h0 : _GEN_641; // @[Filter.scala 165:166]
  wire [3:0] _GEN_643 = 8'h58 == _T_47[7:0] ? 4'hf : _GEN_642; // @[Filter.scala 165:166]
  wire [3:0] _GEN_644 = 8'h59 == _T_47[7:0] ? 4'hf : _GEN_643; // @[Filter.scala 165:166]
  wire [3:0] _GEN_645 = 8'h5a == _T_47[7:0] ? 4'hf : _GEN_644; // @[Filter.scala 165:166]
  wire [3:0] _GEN_646 = 8'h5b == _T_47[7:0] ? 4'hf : _GEN_645; // @[Filter.scala 165:166]
  wire [3:0] _GEN_647 = 8'h5c == _T_47[7:0] ? 4'hf : _GEN_646; // @[Filter.scala 165:166]
  wire [3:0] _GEN_648 = 8'h5d == _T_47[7:0] ? 4'hf : _GEN_647; // @[Filter.scala 165:166]
  wire [3:0] _GEN_649 = 8'h5e == _T_47[7:0] ? 4'hf : _GEN_648; // @[Filter.scala 165:166]
  wire [3:0] _GEN_650 = 8'h5f == _T_47[7:0] ? 4'hf : _GEN_649; // @[Filter.scala 165:166]
  wire [3:0] _GEN_651 = 8'h60 == _T_47[7:0] ? 4'h0 : _GEN_650; // @[Filter.scala 165:166]
  wire [3:0] _GEN_652 = 8'h61 == _T_47[7:0] ? 4'h0 : _GEN_651; // @[Filter.scala 165:166]
  wire [3:0] _GEN_653 = 8'h62 == _T_47[7:0] ? 4'h0 : _GEN_652; // @[Filter.scala 165:166]
  wire [3:0] _GEN_654 = 8'h63 == _T_47[7:0] ? 4'h0 : _GEN_653; // @[Filter.scala 165:166]
  wire [3:0] _GEN_655 = 8'h64 == _T_47[7:0] ? 4'h0 : _GEN_654; // @[Filter.scala 165:166]
  wire [3:0] _GEN_656 = 8'h65 == _T_47[7:0] ? 4'h0 : _GEN_655; // @[Filter.scala 165:166]
  wire [3:0] _GEN_657 = 8'h66 == _T_47[7:0] ? 4'h0 : _GEN_656; // @[Filter.scala 165:166]
  wire [3:0] _GEN_658 = 8'h67 == _T_47[7:0] ? 4'h0 : _GEN_657; // @[Filter.scala 165:166]
  wire [3:0] _GEN_659 = 8'h68 == _T_47[7:0] ? 4'hf : _GEN_658; // @[Filter.scala 165:166]
  wire [3:0] _GEN_660 = 8'h69 == _T_47[7:0] ? 4'hf : _GEN_659; // @[Filter.scala 165:166]
  wire [3:0] _GEN_661 = 8'h6a == _T_47[7:0] ? 4'hf : _GEN_660; // @[Filter.scala 165:166]
  wire [3:0] _GEN_662 = 8'h6b == _T_47[7:0] ? 4'hf : _GEN_661; // @[Filter.scala 165:166]
  wire [3:0] _GEN_663 = 8'h6c == _T_47[7:0] ? 4'hf : _GEN_662; // @[Filter.scala 165:166]
  wire [3:0] _GEN_664 = 8'h6d == _T_47[7:0] ? 4'hf : _GEN_663; // @[Filter.scala 165:166]
  wire [3:0] _GEN_665 = 8'h6e == _T_47[7:0] ? 4'hf : _GEN_664; // @[Filter.scala 165:166]
  wire [3:0] _GEN_666 = 8'h6f == _T_47[7:0] ? 4'hf : _GEN_665; // @[Filter.scala 165:166]
  wire [3:0] _GEN_667 = 8'h70 == _T_47[7:0] ? 4'h0 : _GEN_666; // @[Filter.scala 165:166]
  wire [3:0] _GEN_668 = 8'h71 == _T_47[7:0] ? 4'h0 : _GEN_667; // @[Filter.scala 165:166]
  wire [3:0] _GEN_669 = 8'h72 == _T_47[7:0] ? 4'h0 : _GEN_668; // @[Filter.scala 165:166]
  wire [3:0] _GEN_670 = 8'h73 == _T_47[7:0] ? 4'h0 : _GEN_669; // @[Filter.scala 165:166]
  wire [3:0] _GEN_671 = 8'h74 == _T_47[7:0] ? 4'h0 : _GEN_670; // @[Filter.scala 165:166]
  wire [3:0] _GEN_672 = 8'h75 == _T_47[7:0] ? 4'h0 : _GEN_671; // @[Filter.scala 165:166]
  wire [3:0] _GEN_673 = 8'h76 == _T_47[7:0] ? 4'h0 : _GEN_672; // @[Filter.scala 165:166]
  wire [3:0] _GEN_674 = 8'h77 == _T_47[7:0] ? 4'h0 : _GEN_673; // @[Filter.scala 165:166]
  wire [3:0] _GEN_675 = 8'h78 == _T_47[7:0] ? 4'hf : _GEN_674; // @[Filter.scala 165:166]
  wire [3:0] _GEN_676 = 8'h79 == _T_47[7:0] ? 4'hf : _GEN_675; // @[Filter.scala 165:166]
  wire [3:0] _GEN_677 = 8'h7a == _T_47[7:0] ? 4'hf : _GEN_676; // @[Filter.scala 165:166]
  wire [3:0] _GEN_678 = 8'h7b == _T_47[7:0] ? 4'hf : _GEN_677; // @[Filter.scala 165:166]
  wire [3:0] _GEN_679 = 8'h7c == _T_47[7:0] ? 4'hf : _GEN_678; // @[Filter.scala 165:166]
  wire [3:0] _GEN_680 = 8'h7d == _T_47[7:0] ? 4'hf : _GEN_679; // @[Filter.scala 165:166]
  wire [3:0] _GEN_681 = 8'h7e == _T_47[7:0] ? 4'hf : _GEN_680; // @[Filter.scala 165:166]
  wire [3:0] _GEN_682 = 8'h7f == _T_47[7:0] ? 4'hf : _GEN_681; // @[Filter.scala 165:166]
  wire [3:0] _GEN_683 = 8'h80 == _T_47[7:0] ? 4'h0 : _GEN_682; // @[Filter.scala 165:166]
  wire [3:0] _GEN_684 = 8'h81 == _T_47[7:0] ? 4'h0 : _GEN_683; // @[Filter.scala 165:166]
  wire [3:0] _GEN_685 = 8'h82 == _T_47[7:0] ? 4'h0 : _GEN_684; // @[Filter.scala 165:166]
  wire [3:0] _GEN_686 = 8'h83 == _T_47[7:0] ? 4'h0 : _GEN_685; // @[Filter.scala 165:166]
  wire [3:0] _GEN_687 = 8'h84 == _T_47[7:0] ? 4'h0 : _GEN_686; // @[Filter.scala 165:166]
  wire [3:0] _GEN_688 = 8'h85 == _T_47[7:0] ? 4'h0 : _GEN_687; // @[Filter.scala 165:166]
  wire [3:0] _GEN_689 = 8'h86 == _T_47[7:0] ? 4'h0 : _GEN_688; // @[Filter.scala 165:166]
  wire [3:0] _GEN_690 = 8'h87 == _T_47[7:0] ? 4'h0 : _GEN_689; // @[Filter.scala 165:166]
  wire [3:0] _GEN_691 = 8'h88 == _T_47[7:0] ? 4'hf : _GEN_690; // @[Filter.scala 165:166]
  wire [3:0] _GEN_692 = 8'h89 == _T_47[7:0] ? 4'hf : _GEN_691; // @[Filter.scala 165:166]
  wire [3:0] _GEN_693 = 8'h8a == _T_47[7:0] ? 4'hf : _GEN_692; // @[Filter.scala 165:166]
  wire [3:0] _GEN_694 = 8'h8b == _T_47[7:0] ? 4'hf : _GEN_693; // @[Filter.scala 165:166]
  wire [3:0] _GEN_695 = 8'h8c == _T_47[7:0] ? 4'hf : _GEN_694; // @[Filter.scala 165:166]
  wire [3:0] _GEN_696 = 8'h8d == _T_47[7:0] ? 4'hf : _GEN_695; // @[Filter.scala 165:166]
  wire [3:0] _GEN_697 = 8'h8e == _T_47[7:0] ? 4'hf : _GEN_696; // @[Filter.scala 165:166]
  wire [3:0] _GEN_698 = 8'h8f == _T_47[7:0] ? 4'hf : _GEN_697; // @[Filter.scala 165:166]
  wire [3:0] _GEN_699 = 8'h90 == _T_47[7:0] ? 4'h0 : _GEN_698; // @[Filter.scala 165:166]
  wire [3:0] _GEN_700 = 8'h91 == _T_47[7:0] ? 4'h0 : _GEN_699; // @[Filter.scala 165:166]
  wire [3:0] _GEN_701 = 8'h92 == _T_47[7:0] ? 4'h0 : _GEN_700; // @[Filter.scala 165:166]
  wire [3:0] _GEN_702 = 8'h93 == _T_47[7:0] ? 4'h0 : _GEN_701; // @[Filter.scala 165:166]
  wire [3:0] _GEN_703 = 8'h94 == _T_47[7:0] ? 4'h0 : _GEN_702; // @[Filter.scala 165:166]
  wire [3:0] _GEN_704 = 8'h95 == _T_47[7:0] ? 4'h0 : _GEN_703; // @[Filter.scala 165:166]
  wire [3:0] _GEN_705 = 8'h96 == _T_47[7:0] ? 4'h0 : _GEN_704; // @[Filter.scala 165:166]
  wire [3:0] _GEN_706 = 8'h97 == _T_47[7:0] ? 4'h0 : _GEN_705; // @[Filter.scala 165:166]
  wire [3:0] _GEN_707 = 8'h98 == _T_47[7:0] ? 4'hf : _GEN_706; // @[Filter.scala 165:166]
  wire [3:0] _GEN_708 = 8'h99 == _T_47[7:0] ? 4'hf : _GEN_707; // @[Filter.scala 165:166]
  wire [3:0] _GEN_709 = 8'h9a == _T_47[7:0] ? 4'hf : _GEN_708; // @[Filter.scala 165:166]
  wire [3:0] _GEN_710 = 8'h9b == _T_47[7:0] ? 4'hf : _GEN_709; // @[Filter.scala 165:166]
  wire [3:0] _GEN_711 = 8'h9c == _T_47[7:0] ? 4'hf : _GEN_710; // @[Filter.scala 165:166]
  wire [3:0] _GEN_712 = 8'h9d == _T_47[7:0] ? 4'hf : _GEN_711; // @[Filter.scala 165:166]
  wire [3:0] _GEN_713 = 8'h9e == _T_47[7:0] ? 4'hf : _GEN_712; // @[Filter.scala 165:166]
  wire [3:0] _GEN_714 = 8'h9f == _T_47[7:0] ? 4'hf : _GEN_713; // @[Filter.scala 165:166]
  wire [3:0] _GEN_715 = 8'ha0 == _T_47[7:0] ? 4'h0 : _GEN_714; // @[Filter.scala 165:166]
  wire [3:0] _GEN_716 = 8'ha1 == _T_47[7:0] ? 4'h0 : _GEN_715; // @[Filter.scala 165:166]
  wire [3:0] _GEN_717 = 8'ha2 == _T_47[7:0] ? 4'h0 : _GEN_716; // @[Filter.scala 165:166]
  wire [3:0] _GEN_718 = 8'ha3 == _T_47[7:0] ? 4'h0 : _GEN_717; // @[Filter.scala 165:166]
  wire [3:0] _GEN_719 = 8'ha4 == _T_47[7:0] ? 4'h0 : _GEN_718; // @[Filter.scala 165:166]
  wire [3:0] _GEN_720 = 8'ha5 == _T_47[7:0] ? 4'h0 : _GEN_719; // @[Filter.scala 165:166]
  wire [3:0] _GEN_721 = 8'ha6 == _T_47[7:0] ? 4'h0 : _GEN_720; // @[Filter.scala 165:166]
  wire [3:0] _GEN_722 = 8'ha7 == _T_47[7:0] ? 4'h0 : _GEN_721; // @[Filter.scala 165:166]
  wire [3:0] _GEN_723 = 8'ha8 == _T_47[7:0] ? 4'hf : _GEN_722; // @[Filter.scala 165:166]
  wire [3:0] _GEN_724 = 8'ha9 == _T_47[7:0] ? 4'hf : _GEN_723; // @[Filter.scala 165:166]
  wire [3:0] _GEN_725 = 8'haa == _T_47[7:0] ? 4'hf : _GEN_724; // @[Filter.scala 165:166]
  wire [3:0] _GEN_726 = 8'hab == _T_47[7:0] ? 4'hf : _GEN_725; // @[Filter.scala 165:166]
  wire [3:0] _GEN_727 = 8'hac == _T_47[7:0] ? 4'hf : _GEN_726; // @[Filter.scala 165:166]
  wire [3:0] _GEN_728 = 8'had == _T_47[7:0] ? 4'hf : _GEN_727; // @[Filter.scala 165:166]
  wire [3:0] _GEN_729 = 8'hae == _T_47[7:0] ? 4'hf : _GEN_728; // @[Filter.scala 165:166]
  wire [3:0] _GEN_730 = 8'haf == _T_47[7:0] ? 4'hf : _GEN_729; // @[Filter.scala 165:166]
  wire [3:0] _GEN_731 = 8'hb0 == _T_47[7:0] ? 4'h0 : _GEN_730; // @[Filter.scala 165:166]
  wire [3:0] _GEN_732 = 8'hb1 == _T_47[7:0] ? 4'h0 : _GEN_731; // @[Filter.scala 165:166]
  wire [3:0] _GEN_733 = 8'hb2 == _T_47[7:0] ? 4'h0 : _GEN_732; // @[Filter.scala 165:166]
  wire [3:0] _GEN_734 = 8'hb3 == _T_47[7:0] ? 4'h0 : _GEN_733; // @[Filter.scala 165:166]
  wire [3:0] _GEN_735 = 8'hb4 == _T_47[7:0] ? 4'h0 : _GEN_734; // @[Filter.scala 165:166]
  wire [3:0] _GEN_736 = 8'hb5 == _T_47[7:0] ? 4'h0 : _GEN_735; // @[Filter.scala 165:166]
  wire [3:0] _GEN_737 = 8'hb6 == _T_47[7:0] ? 4'h0 : _GEN_736; // @[Filter.scala 165:166]
  wire [3:0] _GEN_738 = 8'hb7 == _T_47[7:0] ? 4'h0 : _GEN_737; // @[Filter.scala 165:166]
  wire [3:0] _GEN_739 = 8'hb8 == _T_47[7:0] ? 4'hf : _GEN_738; // @[Filter.scala 165:166]
  wire [3:0] _GEN_740 = 8'hb9 == _T_47[7:0] ? 4'hf : _GEN_739; // @[Filter.scala 165:166]
  wire [3:0] _GEN_741 = 8'hba == _T_47[7:0] ? 4'hf : _GEN_740; // @[Filter.scala 165:166]
  wire [3:0] _GEN_742 = 8'hbb == _T_47[7:0] ? 4'hf : _GEN_741; // @[Filter.scala 165:166]
  wire [3:0] _GEN_743 = 8'hbc == _T_47[7:0] ? 4'hf : _GEN_742; // @[Filter.scala 165:166]
  wire [3:0] _GEN_744 = 8'hbd == _T_47[7:0] ? 4'hf : _GEN_743; // @[Filter.scala 165:166]
  wire [3:0] _GEN_745 = 8'hbe == _T_47[7:0] ? 4'hf : _GEN_744; // @[Filter.scala 165:166]
  wire [3:0] _GEN_746 = 8'hbf == _T_47[7:0] ? 4'hf : _GEN_745; // @[Filter.scala 165:166]
  wire [7:0] _T_61 = _GEN_746 * 4'ha; // @[Filter.scala 165:166]
  wire [10:0] _GEN_18991 = {{3'd0}, _T_61}; // @[Filter.scala 165:133]
  wire [10:0] _T_63 = _T_56 + _GEN_18991; // @[Filter.scala 165:133]
  wire [10:0] _T_64 = _T_63 / 11'h64; // @[Filter.scala 165:174]
  wire [10:0] _GEN_939 = io_SPI_distort ? _T_64 : {{7'd0}, _GEN_362}; // @[Filter.scala 164:35]
  wire [10:0] _GEN_940 = _T_44 ? 11'h0 : _GEN_939; // @[Filter.scala 162:80]
  wire [10:0] _GEN_1709 = io_SPI_distort ? _T_64 : {{7'd0}, _GEN_554}; // @[Filter.scala 164:35]
  wire [10:0] _GEN_1710 = _T_44 ? 11'h0 : _GEN_1709; // @[Filter.scala 162:80]
  wire [10:0] _GEN_2479 = io_SPI_distort ? _T_64 : {{7'd0}, _GEN_746}; // @[Filter.scala 164:35]
  wire [10:0] _GEN_2480 = _T_44 ? 11'h0 : _GEN_2479; // @[Filter.scala 162:80]
  wire [31:0] _T_132 = pixelIndex + 32'h1; // @[Filter.scala 158:31]
  wire [31:0] _GEN_1 = _T_132 % 32'h10; // @[Filter.scala 158:38]
  wire [4:0] _T_133 = _GEN_1[4:0]; // @[Filter.scala 158:38]
  wire [4:0] _T_135 = _T_133 + _GEN_18983; // @[Filter.scala 158:53]
  wire [4:0] _T_137 = _T_135 - 5'h1; // @[Filter.scala 158:69]
  wire [31:0] _T_140 = _T_132 / 32'h10; // @[Filter.scala 159:38]
  wire [31:0] _T_142 = _T_140 + _GEN_18984; // @[Filter.scala 159:53]
  wire [31:0] _T_144 = _T_142 - 32'h1; // @[Filter.scala 159:69]
  wire  _T_146 = _T_137 >= 5'h10; // @[Filter.scala 162:31]
  wire  _T_150 = _T_144 >= 32'hc; // @[Filter.scala 162:63]
  wire  _T_151 = _T_146 | _T_150; // @[Filter.scala 162:58]
  wire [36:0] _T_152 = _T_144 * 32'h10; // @[Filter.scala 165:66]
  wire [36:0] _GEN_19011 = {{32'd0}, _T_137}; // @[Filter.scala 165:81]
  wire [36:0] _T_154 = _T_152 + _GEN_19011; // @[Filter.scala 165:81]
  wire [3:0] _GEN_2489 = 8'h8 == _T_154[7:0] ? 4'h0 : 4'hf; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2490 = 8'h9 == _T_154[7:0] ? 4'h0 : _GEN_2489; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2491 = 8'ha == _T_154[7:0] ? 4'h0 : _GEN_2490; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2492 = 8'hb == _T_154[7:0] ? 4'h0 : _GEN_2491; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2493 = 8'hc == _T_154[7:0] ? 4'h0 : _GEN_2492; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2494 = 8'hd == _T_154[7:0] ? 4'h0 : _GEN_2493; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2495 = 8'he == _T_154[7:0] ? 4'h0 : _GEN_2494; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2496 = 8'hf == _T_154[7:0] ? 4'h0 : _GEN_2495; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2497 = 8'h10 == _T_154[7:0] ? 4'hf : _GEN_2496; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2498 = 8'h11 == _T_154[7:0] ? 4'hf : _GEN_2497; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2499 = 8'h12 == _T_154[7:0] ? 4'hf : _GEN_2498; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2500 = 8'h13 == _T_154[7:0] ? 4'hf : _GEN_2499; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2501 = 8'h14 == _T_154[7:0] ? 4'hf : _GEN_2500; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2502 = 8'h15 == _T_154[7:0] ? 4'hf : _GEN_2501; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2503 = 8'h16 == _T_154[7:0] ? 4'hf : _GEN_2502; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2504 = 8'h17 == _T_154[7:0] ? 4'hf : _GEN_2503; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2505 = 8'h18 == _T_154[7:0] ? 4'h0 : _GEN_2504; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2506 = 8'h19 == _T_154[7:0] ? 4'h0 : _GEN_2505; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2507 = 8'h1a == _T_154[7:0] ? 4'h0 : _GEN_2506; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2508 = 8'h1b == _T_154[7:0] ? 4'h0 : _GEN_2507; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2509 = 8'h1c == _T_154[7:0] ? 4'h0 : _GEN_2508; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2510 = 8'h1d == _T_154[7:0] ? 4'h0 : _GEN_2509; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2511 = 8'h1e == _T_154[7:0] ? 4'h0 : _GEN_2510; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2512 = 8'h1f == _T_154[7:0] ? 4'h0 : _GEN_2511; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2513 = 8'h20 == _T_154[7:0] ? 4'hf : _GEN_2512; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2514 = 8'h21 == _T_154[7:0] ? 4'hf : _GEN_2513; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2515 = 8'h22 == _T_154[7:0] ? 4'hf : _GEN_2514; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2516 = 8'h23 == _T_154[7:0] ? 4'hf : _GEN_2515; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2517 = 8'h24 == _T_154[7:0] ? 4'hf : _GEN_2516; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2518 = 8'h25 == _T_154[7:0] ? 4'hf : _GEN_2517; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2519 = 8'h26 == _T_154[7:0] ? 4'hf : _GEN_2518; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2520 = 8'h27 == _T_154[7:0] ? 4'hf : _GEN_2519; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2521 = 8'h28 == _T_154[7:0] ? 4'h0 : _GEN_2520; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2522 = 8'h29 == _T_154[7:0] ? 4'h0 : _GEN_2521; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2523 = 8'h2a == _T_154[7:0] ? 4'h0 : _GEN_2522; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2524 = 8'h2b == _T_154[7:0] ? 4'h0 : _GEN_2523; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2525 = 8'h2c == _T_154[7:0] ? 4'h0 : _GEN_2524; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2526 = 8'h2d == _T_154[7:0] ? 4'h0 : _GEN_2525; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2527 = 8'h2e == _T_154[7:0] ? 4'h0 : _GEN_2526; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2528 = 8'h2f == _T_154[7:0] ? 4'h0 : _GEN_2527; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2529 = 8'h30 == _T_154[7:0] ? 4'hf : _GEN_2528; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2530 = 8'h31 == _T_154[7:0] ? 4'hf : _GEN_2529; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2531 = 8'h32 == _T_154[7:0] ? 4'hf : _GEN_2530; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2532 = 8'h33 == _T_154[7:0] ? 4'hf : _GEN_2531; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2533 = 8'h34 == _T_154[7:0] ? 4'hf : _GEN_2532; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2534 = 8'h35 == _T_154[7:0] ? 4'hf : _GEN_2533; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2535 = 8'h36 == _T_154[7:0] ? 4'hf : _GEN_2534; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2536 = 8'h37 == _T_154[7:0] ? 4'hf : _GEN_2535; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2537 = 8'h38 == _T_154[7:0] ? 4'h0 : _GEN_2536; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2538 = 8'h39 == _T_154[7:0] ? 4'h0 : _GEN_2537; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2539 = 8'h3a == _T_154[7:0] ? 4'h0 : _GEN_2538; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2540 = 8'h3b == _T_154[7:0] ? 4'h0 : _GEN_2539; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2541 = 8'h3c == _T_154[7:0] ? 4'h0 : _GEN_2540; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2542 = 8'h3d == _T_154[7:0] ? 4'h0 : _GEN_2541; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2543 = 8'h3e == _T_154[7:0] ? 4'h0 : _GEN_2542; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2544 = 8'h3f == _T_154[7:0] ? 4'h0 : _GEN_2543; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2545 = 8'h40 == _T_154[7:0] ? 4'hf : _GEN_2544; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2546 = 8'h41 == _T_154[7:0] ? 4'hf : _GEN_2545; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2547 = 8'h42 == _T_154[7:0] ? 4'hf : _GEN_2546; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2548 = 8'h43 == _T_154[7:0] ? 4'hf : _GEN_2547; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2549 = 8'h44 == _T_154[7:0] ? 4'hf : _GEN_2548; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2550 = 8'h45 == _T_154[7:0] ? 4'hf : _GEN_2549; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2551 = 8'h46 == _T_154[7:0] ? 4'hf : _GEN_2550; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2552 = 8'h47 == _T_154[7:0] ? 4'hf : _GEN_2551; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2553 = 8'h48 == _T_154[7:0] ? 4'h0 : _GEN_2552; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2554 = 8'h49 == _T_154[7:0] ? 4'h0 : _GEN_2553; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2555 = 8'h4a == _T_154[7:0] ? 4'h0 : _GEN_2554; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2556 = 8'h4b == _T_154[7:0] ? 4'h0 : _GEN_2555; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2557 = 8'h4c == _T_154[7:0] ? 4'h0 : _GEN_2556; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2558 = 8'h4d == _T_154[7:0] ? 4'h0 : _GEN_2557; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2559 = 8'h4e == _T_154[7:0] ? 4'h0 : _GEN_2558; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2560 = 8'h4f == _T_154[7:0] ? 4'h0 : _GEN_2559; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2561 = 8'h50 == _T_154[7:0] ? 4'hf : _GEN_2560; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2562 = 8'h51 == _T_154[7:0] ? 4'hf : _GEN_2561; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2563 = 8'h52 == _T_154[7:0] ? 4'hf : _GEN_2562; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2564 = 8'h53 == _T_154[7:0] ? 4'hf : _GEN_2563; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2565 = 8'h54 == _T_154[7:0] ? 4'hf : _GEN_2564; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2566 = 8'h55 == _T_154[7:0] ? 4'hf : _GEN_2565; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2567 = 8'h56 == _T_154[7:0] ? 4'hf : _GEN_2566; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2568 = 8'h57 == _T_154[7:0] ? 4'hf : _GEN_2567; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2569 = 8'h58 == _T_154[7:0] ? 4'h0 : _GEN_2568; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2570 = 8'h59 == _T_154[7:0] ? 4'h0 : _GEN_2569; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2571 = 8'h5a == _T_154[7:0] ? 4'h0 : _GEN_2570; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2572 = 8'h5b == _T_154[7:0] ? 4'h0 : _GEN_2571; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2573 = 8'h5c == _T_154[7:0] ? 4'h0 : _GEN_2572; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2574 = 8'h5d == _T_154[7:0] ? 4'h0 : _GEN_2573; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2575 = 8'h5e == _T_154[7:0] ? 4'h0 : _GEN_2574; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2576 = 8'h5f == _T_154[7:0] ? 4'h0 : _GEN_2575; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2577 = 8'h60 == _T_154[7:0] ? 4'h0 : _GEN_2576; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2578 = 8'h61 == _T_154[7:0] ? 4'h0 : _GEN_2577; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2579 = 8'h62 == _T_154[7:0] ? 4'h0 : _GEN_2578; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2580 = 8'h63 == _T_154[7:0] ? 4'h0 : _GEN_2579; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2581 = 8'h64 == _T_154[7:0] ? 4'h0 : _GEN_2580; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2582 = 8'h65 == _T_154[7:0] ? 4'h0 : _GEN_2581; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2583 = 8'h66 == _T_154[7:0] ? 4'h0 : _GEN_2582; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2584 = 8'h67 == _T_154[7:0] ? 4'h0 : _GEN_2583; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2585 = 8'h68 == _T_154[7:0] ? 4'hf : _GEN_2584; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2586 = 8'h69 == _T_154[7:0] ? 4'hf : _GEN_2585; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2587 = 8'h6a == _T_154[7:0] ? 4'hf : _GEN_2586; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2588 = 8'h6b == _T_154[7:0] ? 4'hf : _GEN_2587; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2589 = 8'h6c == _T_154[7:0] ? 4'hf : _GEN_2588; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2590 = 8'h6d == _T_154[7:0] ? 4'hf : _GEN_2589; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2591 = 8'h6e == _T_154[7:0] ? 4'hf : _GEN_2590; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2592 = 8'h6f == _T_154[7:0] ? 4'hf : _GEN_2591; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2593 = 8'h70 == _T_154[7:0] ? 4'h0 : _GEN_2592; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2594 = 8'h71 == _T_154[7:0] ? 4'h0 : _GEN_2593; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2595 = 8'h72 == _T_154[7:0] ? 4'h0 : _GEN_2594; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2596 = 8'h73 == _T_154[7:0] ? 4'h0 : _GEN_2595; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2597 = 8'h74 == _T_154[7:0] ? 4'h0 : _GEN_2596; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2598 = 8'h75 == _T_154[7:0] ? 4'h0 : _GEN_2597; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2599 = 8'h76 == _T_154[7:0] ? 4'h0 : _GEN_2598; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2600 = 8'h77 == _T_154[7:0] ? 4'h0 : _GEN_2599; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2601 = 8'h78 == _T_154[7:0] ? 4'hf : _GEN_2600; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2602 = 8'h79 == _T_154[7:0] ? 4'hf : _GEN_2601; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2603 = 8'h7a == _T_154[7:0] ? 4'hf : _GEN_2602; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2604 = 8'h7b == _T_154[7:0] ? 4'hf : _GEN_2603; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2605 = 8'h7c == _T_154[7:0] ? 4'hf : _GEN_2604; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2606 = 8'h7d == _T_154[7:0] ? 4'hf : _GEN_2605; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2607 = 8'h7e == _T_154[7:0] ? 4'hf : _GEN_2606; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2608 = 8'h7f == _T_154[7:0] ? 4'hf : _GEN_2607; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2609 = 8'h80 == _T_154[7:0] ? 4'h0 : _GEN_2608; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2610 = 8'h81 == _T_154[7:0] ? 4'h0 : _GEN_2609; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2611 = 8'h82 == _T_154[7:0] ? 4'h0 : _GEN_2610; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2612 = 8'h83 == _T_154[7:0] ? 4'h0 : _GEN_2611; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2613 = 8'h84 == _T_154[7:0] ? 4'h0 : _GEN_2612; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2614 = 8'h85 == _T_154[7:0] ? 4'h0 : _GEN_2613; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2615 = 8'h86 == _T_154[7:0] ? 4'h0 : _GEN_2614; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2616 = 8'h87 == _T_154[7:0] ? 4'h0 : _GEN_2615; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2617 = 8'h88 == _T_154[7:0] ? 4'hf : _GEN_2616; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2618 = 8'h89 == _T_154[7:0] ? 4'hf : _GEN_2617; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2619 = 8'h8a == _T_154[7:0] ? 4'hf : _GEN_2618; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2620 = 8'h8b == _T_154[7:0] ? 4'hf : _GEN_2619; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2621 = 8'h8c == _T_154[7:0] ? 4'hf : _GEN_2620; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2622 = 8'h8d == _T_154[7:0] ? 4'hf : _GEN_2621; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2623 = 8'h8e == _T_154[7:0] ? 4'hf : _GEN_2622; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2624 = 8'h8f == _T_154[7:0] ? 4'hf : _GEN_2623; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2625 = 8'h90 == _T_154[7:0] ? 4'h0 : _GEN_2624; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2626 = 8'h91 == _T_154[7:0] ? 4'h0 : _GEN_2625; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2627 = 8'h92 == _T_154[7:0] ? 4'h0 : _GEN_2626; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2628 = 8'h93 == _T_154[7:0] ? 4'h0 : _GEN_2627; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2629 = 8'h94 == _T_154[7:0] ? 4'h0 : _GEN_2628; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2630 = 8'h95 == _T_154[7:0] ? 4'h0 : _GEN_2629; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2631 = 8'h96 == _T_154[7:0] ? 4'h0 : _GEN_2630; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2632 = 8'h97 == _T_154[7:0] ? 4'h0 : _GEN_2631; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2633 = 8'h98 == _T_154[7:0] ? 4'hf : _GEN_2632; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2634 = 8'h99 == _T_154[7:0] ? 4'hf : _GEN_2633; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2635 = 8'h9a == _T_154[7:0] ? 4'hf : _GEN_2634; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2636 = 8'h9b == _T_154[7:0] ? 4'hf : _GEN_2635; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2637 = 8'h9c == _T_154[7:0] ? 4'hf : _GEN_2636; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2638 = 8'h9d == _T_154[7:0] ? 4'hf : _GEN_2637; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2639 = 8'h9e == _T_154[7:0] ? 4'hf : _GEN_2638; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2640 = 8'h9f == _T_154[7:0] ? 4'hf : _GEN_2639; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2641 = 8'ha0 == _T_154[7:0] ? 4'h0 : _GEN_2640; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2642 = 8'ha1 == _T_154[7:0] ? 4'h0 : _GEN_2641; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2643 = 8'ha2 == _T_154[7:0] ? 4'h0 : _GEN_2642; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2644 = 8'ha3 == _T_154[7:0] ? 4'h0 : _GEN_2643; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2645 = 8'ha4 == _T_154[7:0] ? 4'h0 : _GEN_2644; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2646 = 8'ha5 == _T_154[7:0] ? 4'h0 : _GEN_2645; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2647 = 8'ha6 == _T_154[7:0] ? 4'h0 : _GEN_2646; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2648 = 8'ha7 == _T_154[7:0] ? 4'h0 : _GEN_2647; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2649 = 8'ha8 == _T_154[7:0] ? 4'hf : _GEN_2648; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2650 = 8'ha9 == _T_154[7:0] ? 4'hf : _GEN_2649; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2651 = 8'haa == _T_154[7:0] ? 4'hf : _GEN_2650; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2652 = 8'hab == _T_154[7:0] ? 4'hf : _GEN_2651; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2653 = 8'hac == _T_154[7:0] ? 4'hf : _GEN_2652; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2654 = 8'had == _T_154[7:0] ? 4'hf : _GEN_2653; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2655 = 8'hae == _T_154[7:0] ? 4'hf : _GEN_2654; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2656 = 8'haf == _T_154[7:0] ? 4'hf : _GEN_2655; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2657 = 8'hb0 == _T_154[7:0] ? 4'h0 : _GEN_2656; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2658 = 8'hb1 == _T_154[7:0] ? 4'h0 : _GEN_2657; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2659 = 8'hb2 == _T_154[7:0] ? 4'h0 : _GEN_2658; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2660 = 8'hb3 == _T_154[7:0] ? 4'h0 : _GEN_2659; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2661 = 8'hb4 == _T_154[7:0] ? 4'h0 : _GEN_2660; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2662 = 8'hb5 == _T_154[7:0] ? 4'h0 : _GEN_2661; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2663 = 8'hb6 == _T_154[7:0] ? 4'h0 : _GEN_2662; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2664 = 8'hb7 == _T_154[7:0] ? 4'h0 : _GEN_2663; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2665 = 8'hb8 == _T_154[7:0] ? 4'hf : _GEN_2664; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2666 = 8'hb9 == _T_154[7:0] ? 4'hf : _GEN_2665; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2667 = 8'hba == _T_154[7:0] ? 4'hf : _GEN_2666; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2668 = 8'hbb == _T_154[7:0] ? 4'hf : _GEN_2667; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2669 = 8'hbc == _T_154[7:0] ? 4'hf : _GEN_2668; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2670 = 8'hbd == _T_154[7:0] ? 4'hf : _GEN_2669; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2671 = 8'hbe == _T_154[7:0] ? 4'hf : _GEN_2670; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2672 = 8'hbf == _T_154[7:0] ? 4'hf : _GEN_2671; // @[Filter.scala 165:86]
  wire [4:0] _GEN_19012 = {{1'd0}, _GEN_2672}; // @[Filter.scala 165:86]
  wire [8:0] _T_156 = _GEN_19012 * 5'h14; // @[Filter.scala 165:86]
  wire [3:0] _GEN_2769 = 8'h60 == _T_154[7:0] ? 4'hf : 4'h0; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2770 = 8'h61 == _T_154[7:0] ? 4'hf : _GEN_2769; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2771 = 8'h62 == _T_154[7:0] ? 4'hf : _GEN_2770; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2772 = 8'h63 == _T_154[7:0] ? 4'hf : _GEN_2771; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2773 = 8'h64 == _T_154[7:0] ? 4'hf : _GEN_2772; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2774 = 8'h65 == _T_154[7:0] ? 4'hf : _GEN_2773; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2775 = 8'h66 == _T_154[7:0] ? 4'hf : _GEN_2774; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2776 = 8'h67 == _T_154[7:0] ? 4'hf : _GEN_2775; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2777 = 8'h68 == _T_154[7:0] ? 4'hf : _GEN_2776; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2778 = 8'h69 == _T_154[7:0] ? 4'hf : _GEN_2777; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2779 = 8'h6a == _T_154[7:0] ? 4'hf : _GEN_2778; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2780 = 8'h6b == _T_154[7:0] ? 4'hf : _GEN_2779; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2781 = 8'h6c == _T_154[7:0] ? 4'hf : _GEN_2780; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2782 = 8'h6d == _T_154[7:0] ? 4'hf : _GEN_2781; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2783 = 8'h6e == _T_154[7:0] ? 4'hf : _GEN_2782; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2784 = 8'h6f == _T_154[7:0] ? 4'hf : _GEN_2783; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2785 = 8'h70 == _T_154[7:0] ? 4'hf : _GEN_2784; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2786 = 8'h71 == _T_154[7:0] ? 4'hf : _GEN_2785; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2787 = 8'h72 == _T_154[7:0] ? 4'hf : _GEN_2786; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2788 = 8'h73 == _T_154[7:0] ? 4'hf : _GEN_2787; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2789 = 8'h74 == _T_154[7:0] ? 4'hf : _GEN_2788; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2790 = 8'h75 == _T_154[7:0] ? 4'hf : _GEN_2789; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2791 = 8'h76 == _T_154[7:0] ? 4'hf : _GEN_2790; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2792 = 8'h77 == _T_154[7:0] ? 4'hf : _GEN_2791; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2793 = 8'h78 == _T_154[7:0] ? 4'hf : _GEN_2792; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2794 = 8'h79 == _T_154[7:0] ? 4'hf : _GEN_2793; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2795 = 8'h7a == _T_154[7:0] ? 4'hf : _GEN_2794; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2796 = 8'h7b == _T_154[7:0] ? 4'hf : _GEN_2795; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2797 = 8'h7c == _T_154[7:0] ? 4'hf : _GEN_2796; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2798 = 8'h7d == _T_154[7:0] ? 4'hf : _GEN_2797; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2799 = 8'h7e == _T_154[7:0] ? 4'hf : _GEN_2798; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2800 = 8'h7f == _T_154[7:0] ? 4'hf : _GEN_2799; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2801 = 8'h80 == _T_154[7:0] ? 4'hf : _GEN_2800; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2802 = 8'h81 == _T_154[7:0] ? 4'hf : _GEN_2801; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2803 = 8'h82 == _T_154[7:0] ? 4'hf : _GEN_2802; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2804 = 8'h83 == _T_154[7:0] ? 4'hf : _GEN_2803; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2805 = 8'h84 == _T_154[7:0] ? 4'hf : _GEN_2804; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2806 = 8'h85 == _T_154[7:0] ? 4'hf : _GEN_2805; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2807 = 8'h86 == _T_154[7:0] ? 4'hf : _GEN_2806; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2808 = 8'h87 == _T_154[7:0] ? 4'hf : _GEN_2807; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2809 = 8'h88 == _T_154[7:0] ? 4'hf : _GEN_2808; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2810 = 8'h89 == _T_154[7:0] ? 4'hf : _GEN_2809; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2811 = 8'h8a == _T_154[7:0] ? 4'hf : _GEN_2810; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2812 = 8'h8b == _T_154[7:0] ? 4'hf : _GEN_2811; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2813 = 8'h8c == _T_154[7:0] ? 4'hf : _GEN_2812; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2814 = 8'h8d == _T_154[7:0] ? 4'hf : _GEN_2813; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2815 = 8'h8e == _T_154[7:0] ? 4'hf : _GEN_2814; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2816 = 8'h8f == _T_154[7:0] ? 4'hf : _GEN_2815; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2817 = 8'h90 == _T_154[7:0] ? 4'hf : _GEN_2816; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2818 = 8'h91 == _T_154[7:0] ? 4'hf : _GEN_2817; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2819 = 8'h92 == _T_154[7:0] ? 4'hf : _GEN_2818; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2820 = 8'h93 == _T_154[7:0] ? 4'hf : _GEN_2819; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2821 = 8'h94 == _T_154[7:0] ? 4'hf : _GEN_2820; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2822 = 8'h95 == _T_154[7:0] ? 4'hf : _GEN_2821; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2823 = 8'h96 == _T_154[7:0] ? 4'hf : _GEN_2822; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2824 = 8'h97 == _T_154[7:0] ? 4'hf : _GEN_2823; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2825 = 8'h98 == _T_154[7:0] ? 4'hf : _GEN_2824; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2826 = 8'h99 == _T_154[7:0] ? 4'hf : _GEN_2825; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2827 = 8'h9a == _T_154[7:0] ? 4'hf : _GEN_2826; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2828 = 8'h9b == _T_154[7:0] ? 4'hf : _GEN_2827; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2829 = 8'h9c == _T_154[7:0] ? 4'hf : _GEN_2828; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2830 = 8'h9d == _T_154[7:0] ? 4'hf : _GEN_2829; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2831 = 8'h9e == _T_154[7:0] ? 4'hf : _GEN_2830; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2832 = 8'h9f == _T_154[7:0] ? 4'hf : _GEN_2831; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2833 = 8'ha0 == _T_154[7:0] ? 4'hf : _GEN_2832; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2834 = 8'ha1 == _T_154[7:0] ? 4'hf : _GEN_2833; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2835 = 8'ha2 == _T_154[7:0] ? 4'hf : _GEN_2834; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2836 = 8'ha3 == _T_154[7:0] ? 4'hf : _GEN_2835; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2837 = 8'ha4 == _T_154[7:0] ? 4'hf : _GEN_2836; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2838 = 8'ha5 == _T_154[7:0] ? 4'hf : _GEN_2837; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2839 = 8'ha6 == _T_154[7:0] ? 4'hf : _GEN_2838; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2840 = 8'ha7 == _T_154[7:0] ? 4'hf : _GEN_2839; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2841 = 8'ha8 == _T_154[7:0] ? 4'hf : _GEN_2840; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2842 = 8'ha9 == _T_154[7:0] ? 4'hf : _GEN_2841; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2843 = 8'haa == _T_154[7:0] ? 4'hf : _GEN_2842; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2844 = 8'hab == _T_154[7:0] ? 4'hf : _GEN_2843; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2845 = 8'hac == _T_154[7:0] ? 4'hf : _GEN_2844; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2846 = 8'had == _T_154[7:0] ? 4'hf : _GEN_2845; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2847 = 8'hae == _T_154[7:0] ? 4'hf : _GEN_2846; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2848 = 8'haf == _T_154[7:0] ? 4'hf : _GEN_2847; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2849 = 8'hb0 == _T_154[7:0] ? 4'hf : _GEN_2848; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2850 = 8'hb1 == _T_154[7:0] ? 4'hf : _GEN_2849; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2851 = 8'hb2 == _T_154[7:0] ? 4'hf : _GEN_2850; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2852 = 8'hb3 == _T_154[7:0] ? 4'hf : _GEN_2851; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2853 = 8'hb4 == _T_154[7:0] ? 4'hf : _GEN_2852; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2854 = 8'hb5 == _T_154[7:0] ? 4'hf : _GEN_2853; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2855 = 8'hb6 == _T_154[7:0] ? 4'hf : _GEN_2854; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2856 = 8'hb7 == _T_154[7:0] ? 4'hf : _GEN_2855; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2857 = 8'hb8 == _T_154[7:0] ? 4'hf : _GEN_2856; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2858 = 8'hb9 == _T_154[7:0] ? 4'hf : _GEN_2857; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2859 = 8'hba == _T_154[7:0] ? 4'hf : _GEN_2858; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2860 = 8'hbb == _T_154[7:0] ? 4'hf : _GEN_2859; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2861 = 8'hbc == _T_154[7:0] ? 4'hf : _GEN_2860; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2862 = 8'hbd == _T_154[7:0] ? 4'hf : _GEN_2861; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2863 = 8'hbe == _T_154[7:0] ? 4'hf : _GEN_2862; // @[Filter.scala 165:126]
  wire [3:0] _GEN_2864 = 8'hbf == _T_154[7:0] ? 4'hf : _GEN_2863; // @[Filter.scala 165:126]
  wire [6:0] _GEN_19014 = {{3'd0}, _GEN_2864}; // @[Filter.scala 165:126]
  wire [10:0] _T_161 = _GEN_19014 * 7'h46; // @[Filter.scala 165:126]
  wire [10:0] _GEN_19015 = {{2'd0}, _T_156}; // @[Filter.scala 165:93]
  wire [10:0] _T_163 = _GEN_19015 + _T_161; // @[Filter.scala 165:93]
  wire [3:0] _GEN_2873 = 8'h8 == _T_154[7:0] ? 4'hf : 4'h0; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2874 = 8'h9 == _T_154[7:0] ? 4'hf : _GEN_2873; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2875 = 8'ha == _T_154[7:0] ? 4'hf : _GEN_2874; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2876 = 8'hb == _T_154[7:0] ? 4'hf : _GEN_2875; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2877 = 8'hc == _T_154[7:0] ? 4'hf : _GEN_2876; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2878 = 8'hd == _T_154[7:0] ? 4'hf : _GEN_2877; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2879 = 8'he == _T_154[7:0] ? 4'hf : _GEN_2878; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2880 = 8'hf == _T_154[7:0] ? 4'hf : _GEN_2879; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2881 = 8'h10 == _T_154[7:0] ? 4'h0 : _GEN_2880; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2882 = 8'h11 == _T_154[7:0] ? 4'h0 : _GEN_2881; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2883 = 8'h12 == _T_154[7:0] ? 4'h0 : _GEN_2882; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2884 = 8'h13 == _T_154[7:0] ? 4'h0 : _GEN_2883; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2885 = 8'h14 == _T_154[7:0] ? 4'h0 : _GEN_2884; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2886 = 8'h15 == _T_154[7:0] ? 4'h0 : _GEN_2885; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2887 = 8'h16 == _T_154[7:0] ? 4'h0 : _GEN_2886; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2888 = 8'h17 == _T_154[7:0] ? 4'h0 : _GEN_2887; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2889 = 8'h18 == _T_154[7:0] ? 4'hf : _GEN_2888; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2890 = 8'h19 == _T_154[7:0] ? 4'hf : _GEN_2889; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2891 = 8'h1a == _T_154[7:0] ? 4'hf : _GEN_2890; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2892 = 8'h1b == _T_154[7:0] ? 4'hf : _GEN_2891; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2893 = 8'h1c == _T_154[7:0] ? 4'hf : _GEN_2892; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2894 = 8'h1d == _T_154[7:0] ? 4'hf : _GEN_2893; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2895 = 8'h1e == _T_154[7:0] ? 4'hf : _GEN_2894; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2896 = 8'h1f == _T_154[7:0] ? 4'hf : _GEN_2895; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2897 = 8'h20 == _T_154[7:0] ? 4'h0 : _GEN_2896; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2898 = 8'h21 == _T_154[7:0] ? 4'h0 : _GEN_2897; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2899 = 8'h22 == _T_154[7:0] ? 4'h0 : _GEN_2898; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2900 = 8'h23 == _T_154[7:0] ? 4'h0 : _GEN_2899; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2901 = 8'h24 == _T_154[7:0] ? 4'h0 : _GEN_2900; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2902 = 8'h25 == _T_154[7:0] ? 4'h0 : _GEN_2901; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2903 = 8'h26 == _T_154[7:0] ? 4'h0 : _GEN_2902; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2904 = 8'h27 == _T_154[7:0] ? 4'h0 : _GEN_2903; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2905 = 8'h28 == _T_154[7:0] ? 4'hf : _GEN_2904; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2906 = 8'h29 == _T_154[7:0] ? 4'hf : _GEN_2905; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2907 = 8'h2a == _T_154[7:0] ? 4'hf : _GEN_2906; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2908 = 8'h2b == _T_154[7:0] ? 4'hf : _GEN_2907; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2909 = 8'h2c == _T_154[7:0] ? 4'hf : _GEN_2908; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2910 = 8'h2d == _T_154[7:0] ? 4'hf : _GEN_2909; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2911 = 8'h2e == _T_154[7:0] ? 4'hf : _GEN_2910; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2912 = 8'h2f == _T_154[7:0] ? 4'hf : _GEN_2911; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2913 = 8'h30 == _T_154[7:0] ? 4'h0 : _GEN_2912; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2914 = 8'h31 == _T_154[7:0] ? 4'h0 : _GEN_2913; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2915 = 8'h32 == _T_154[7:0] ? 4'h0 : _GEN_2914; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2916 = 8'h33 == _T_154[7:0] ? 4'h0 : _GEN_2915; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2917 = 8'h34 == _T_154[7:0] ? 4'h0 : _GEN_2916; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2918 = 8'h35 == _T_154[7:0] ? 4'h0 : _GEN_2917; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2919 = 8'h36 == _T_154[7:0] ? 4'h0 : _GEN_2918; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2920 = 8'h37 == _T_154[7:0] ? 4'h0 : _GEN_2919; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2921 = 8'h38 == _T_154[7:0] ? 4'hf : _GEN_2920; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2922 = 8'h39 == _T_154[7:0] ? 4'hf : _GEN_2921; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2923 = 8'h3a == _T_154[7:0] ? 4'hf : _GEN_2922; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2924 = 8'h3b == _T_154[7:0] ? 4'hf : _GEN_2923; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2925 = 8'h3c == _T_154[7:0] ? 4'hf : _GEN_2924; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2926 = 8'h3d == _T_154[7:0] ? 4'hf : _GEN_2925; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2927 = 8'h3e == _T_154[7:0] ? 4'hf : _GEN_2926; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2928 = 8'h3f == _T_154[7:0] ? 4'hf : _GEN_2927; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2929 = 8'h40 == _T_154[7:0] ? 4'h0 : _GEN_2928; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2930 = 8'h41 == _T_154[7:0] ? 4'h0 : _GEN_2929; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2931 = 8'h42 == _T_154[7:0] ? 4'h0 : _GEN_2930; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2932 = 8'h43 == _T_154[7:0] ? 4'h0 : _GEN_2931; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2933 = 8'h44 == _T_154[7:0] ? 4'h0 : _GEN_2932; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2934 = 8'h45 == _T_154[7:0] ? 4'h0 : _GEN_2933; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2935 = 8'h46 == _T_154[7:0] ? 4'h0 : _GEN_2934; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2936 = 8'h47 == _T_154[7:0] ? 4'h0 : _GEN_2935; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2937 = 8'h48 == _T_154[7:0] ? 4'hf : _GEN_2936; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2938 = 8'h49 == _T_154[7:0] ? 4'hf : _GEN_2937; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2939 = 8'h4a == _T_154[7:0] ? 4'hf : _GEN_2938; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2940 = 8'h4b == _T_154[7:0] ? 4'hf : _GEN_2939; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2941 = 8'h4c == _T_154[7:0] ? 4'hf : _GEN_2940; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2942 = 8'h4d == _T_154[7:0] ? 4'hf : _GEN_2941; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2943 = 8'h4e == _T_154[7:0] ? 4'hf : _GEN_2942; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2944 = 8'h4f == _T_154[7:0] ? 4'hf : _GEN_2943; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2945 = 8'h50 == _T_154[7:0] ? 4'h0 : _GEN_2944; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2946 = 8'h51 == _T_154[7:0] ? 4'h0 : _GEN_2945; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2947 = 8'h52 == _T_154[7:0] ? 4'h0 : _GEN_2946; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2948 = 8'h53 == _T_154[7:0] ? 4'h0 : _GEN_2947; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2949 = 8'h54 == _T_154[7:0] ? 4'h0 : _GEN_2948; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2950 = 8'h55 == _T_154[7:0] ? 4'h0 : _GEN_2949; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2951 = 8'h56 == _T_154[7:0] ? 4'h0 : _GEN_2950; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2952 = 8'h57 == _T_154[7:0] ? 4'h0 : _GEN_2951; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2953 = 8'h58 == _T_154[7:0] ? 4'hf : _GEN_2952; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2954 = 8'h59 == _T_154[7:0] ? 4'hf : _GEN_2953; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2955 = 8'h5a == _T_154[7:0] ? 4'hf : _GEN_2954; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2956 = 8'h5b == _T_154[7:0] ? 4'hf : _GEN_2955; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2957 = 8'h5c == _T_154[7:0] ? 4'hf : _GEN_2956; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2958 = 8'h5d == _T_154[7:0] ? 4'hf : _GEN_2957; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2959 = 8'h5e == _T_154[7:0] ? 4'hf : _GEN_2958; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2960 = 8'h5f == _T_154[7:0] ? 4'hf : _GEN_2959; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2961 = 8'h60 == _T_154[7:0] ? 4'h0 : _GEN_2960; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2962 = 8'h61 == _T_154[7:0] ? 4'h0 : _GEN_2961; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2963 = 8'h62 == _T_154[7:0] ? 4'h0 : _GEN_2962; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2964 = 8'h63 == _T_154[7:0] ? 4'h0 : _GEN_2963; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2965 = 8'h64 == _T_154[7:0] ? 4'h0 : _GEN_2964; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2966 = 8'h65 == _T_154[7:0] ? 4'h0 : _GEN_2965; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2967 = 8'h66 == _T_154[7:0] ? 4'h0 : _GEN_2966; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2968 = 8'h67 == _T_154[7:0] ? 4'h0 : _GEN_2967; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2969 = 8'h68 == _T_154[7:0] ? 4'hf : _GEN_2968; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2970 = 8'h69 == _T_154[7:0] ? 4'hf : _GEN_2969; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2971 = 8'h6a == _T_154[7:0] ? 4'hf : _GEN_2970; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2972 = 8'h6b == _T_154[7:0] ? 4'hf : _GEN_2971; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2973 = 8'h6c == _T_154[7:0] ? 4'hf : _GEN_2972; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2974 = 8'h6d == _T_154[7:0] ? 4'hf : _GEN_2973; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2975 = 8'h6e == _T_154[7:0] ? 4'hf : _GEN_2974; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2976 = 8'h6f == _T_154[7:0] ? 4'hf : _GEN_2975; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2977 = 8'h70 == _T_154[7:0] ? 4'h0 : _GEN_2976; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2978 = 8'h71 == _T_154[7:0] ? 4'h0 : _GEN_2977; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2979 = 8'h72 == _T_154[7:0] ? 4'h0 : _GEN_2978; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2980 = 8'h73 == _T_154[7:0] ? 4'h0 : _GEN_2979; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2981 = 8'h74 == _T_154[7:0] ? 4'h0 : _GEN_2980; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2982 = 8'h75 == _T_154[7:0] ? 4'h0 : _GEN_2981; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2983 = 8'h76 == _T_154[7:0] ? 4'h0 : _GEN_2982; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2984 = 8'h77 == _T_154[7:0] ? 4'h0 : _GEN_2983; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2985 = 8'h78 == _T_154[7:0] ? 4'hf : _GEN_2984; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2986 = 8'h79 == _T_154[7:0] ? 4'hf : _GEN_2985; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2987 = 8'h7a == _T_154[7:0] ? 4'hf : _GEN_2986; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2988 = 8'h7b == _T_154[7:0] ? 4'hf : _GEN_2987; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2989 = 8'h7c == _T_154[7:0] ? 4'hf : _GEN_2988; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2990 = 8'h7d == _T_154[7:0] ? 4'hf : _GEN_2989; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2991 = 8'h7e == _T_154[7:0] ? 4'hf : _GEN_2990; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2992 = 8'h7f == _T_154[7:0] ? 4'hf : _GEN_2991; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2993 = 8'h80 == _T_154[7:0] ? 4'h0 : _GEN_2992; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2994 = 8'h81 == _T_154[7:0] ? 4'h0 : _GEN_2993; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2995 = 8'h82 == _T_154[7:0] ? 4'h0 : _GEN_2994; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2996 = 8'h83 == _T_154[7:0] ? 4'h0 : _GEN_2995; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2997 = 8'h84 == _T_154[7:0] ? 4'h0 : _GEN_2996; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2998 = 8'h85 == _T_154[7:0] ? 4'h0 : _GEN_2997; // @[Filter.scala 165:166]
  wire [3:0] _GEN_2999 = 8'h86 == _T_154[7:0] ? 4'h0 : _GEN_2998; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3000 = 8'h87 == _T_154[7:0] ? 4'h0 : _GEN_2999; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3001 = 8'h88 == _T_154[7:0] ? 4'hf : _GEN_3000; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3002 = 8'h89 == _T_154[7:0] ? 4'hf : _GEN_3001; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3003 = 8'h8a == _T_154[7:0] ? 4'hf : _GEN_3002; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3004 = 8'h8b == _T_154[7:0] ? 4'hf : _GEN_3003; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3005 = 8'h8c == _T_154[7:0] ? 4'hf : _GEN_3004; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3006 = 8'h8d == _T_154[7:0] ? 4'hf : _GEN_3005; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3007 = 8'h8e == _T_154[7:0] ? 4'hf : _GEN_3006; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3008 = 8'h8f == _T_154[7:0] ? 4'hf : _GEN_3007; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3009 = 8'h90 == _T_154[7:0] ? 4'h0 : _GEN_3008; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3010 = 8'h91 == _T_154[7:0] ? 4'h0 : _GEN_3009; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3011 = 8'h92 == _T_154[7:0] ? 4'h0 : _GEN_3010; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3012 = 8'h93 == _T_154[7:0] ? 4'h0 : _GEN_3011; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3013 = 8'h94 == _T_154[7:0] ? 4'h0 : _GEN_3012; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3014 = 8'h95 == _T_154[7:0] ? 4'h0 : _GEN_3013; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3015 = 8'h96 == _T_154[7:0] ? 4'h0 : _GEN_3014; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3016 = 8'h97 == _T_154[7:0] ? 4'h0 : _GEN_3015; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3017 = 8'h98 == _T_154[7:0] ? 4'hf : _GEN_3016; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3018 = 8'h99 == _T_154[7:0] ? 4'hf : _GEN_3017; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3019 = 8'h9a == _T_154[7:0] ? 4'hf : _GEN_3018; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3020 = 8'h9b == _T_154[7:0] ? 4'hf : _GEN_3019; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3021 = 8'h9c == _T_154[7:0] ? 4'hf : _GEN_3020; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3022 = 8'h9d == _T_154[7:0] ? 4'hf : _GEN_3021; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3023 = 8'h9e == _T_154[7:0] ? 4'hf : _GEN_3022; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3024 = 8'h9f == _T_154[7:0] ? 4'hf : _GEN_3023; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3025 = 8'ha0 == _T_154[7:0] ? 4'h0 : _GEN_3024; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3026 = 8'ha1 == _T_154[7:0] ? 4'h0 : _GEN_3025; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3027 = 8'ha2 == _T_154[7:0] ? 4'h0 : _GEN_3026; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3028 = 8'ha3 == _T_154[7:0] ? 4'h0 : _GEN_3027; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3029 = 8'ha4 == _T_154[7:0] ? 4'h0 : _GEN_3028; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3030 = 8'ha5 == _T_154[7:0] ? 4'h0 : _GEN_3029; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3031 = 8'ha6 == _T_154[7:0] ? 4'h0 : _GEN_3030; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3032 = 8'ha7 == _T_154[7:0] ? 4'h0 : _GEN_3031; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3033 = 8'ha8 == _T_154[7:0] ? 4'hf : _GEN_3032; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3034 = 8'ha9 == _T_154[7:0] ? 4'hf : _GEN_3033; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3035 = 8'haa == _T_154[7:0] ? 4'hf : _GEN_3034; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3036 = 8'hab == _T_154[7:0] ? 4'hf : _GEN_3035; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3037 = 8'hac == _T_154[7:0] ? 4'hf : _GEN_3036; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3038 = 8'had == _T_154[7:0] ? 4'hf : _GEN_3037; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3039 = 8'hae == _T_154[7:0] ? 4'hf : _GEN_3038; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3040 = 8'haf == _T_154[7:0] ? 4'hf : _GEN_3039; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3041 = 8'hb0 == _T_154[7:0] ? 4'h0 : _GEN_3040; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3042 = 8'hb1 == _T_154[7:0] ? 4'h0 : _GEN_3041; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3043 = 8'hb2 == _T_154[7:0] ? 4'h0 : _GEN_3042; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3044 = 8'hb3 == _T_154[7:0] ? 4'h0 : _GEN_3043; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3045 = 8'hb4 == _T_154[7:0] ? 4'h0 : _GEN_3044; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3046 = 8'hb5 == _T_154[7:0] ? 4'h0 : _GEN_3045; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3047 = 8'hb6 == _T_154[7:0] ? 4'h0 : _GEN_3046; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3048 = 8'hb7 == _T_154[7:0] ? 4'h0 : _GEN_3047; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3049 = 8'hb8 == _T_154[7:0] ? 4'hf : _GEN_3048; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3050 = 8'hb9 == _T_154[7:0] ? 4'hf : _GEN_3049; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3051 = 8'hba == _T_154[7:0] ? 4'hf : _GEN_3050; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3052 = 8'hbb == _T_154[7:0] ? 4'hf : _GEN_3051; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3053 = 8'hbc == _T_154[7:0] ? 4'hf : _GEN_3052; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3054 = 8'hbd == _T_154[7:0] ? 4'hf : _GEN_3053; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3055 = 8'hbe == _T_154[7:0] ? 4'hf : _GEN_3054; // @[Filter.scala 165:166]
  wire [3:0] _GEN_3056 = 8'hbf == _T_154[7:0] ? 4'hf : _GEN_3055; // @[Filter.scala 165:166]
  wire [7:0] _T_168 = _GEN_3056 * 4'ha; // @[Filter.scala 165:166]
  wire [10:0] _GEN_19017 = {{3'd0}, _T_168}; // @[Filter.scala 165:133]
  wire [10:0] _T_170 = _T_163 + _GEN_19017; // @[Filter.scala 165:133]
  wire [10:0] _T_171 = _T_170 / 11'h64; // @[Filter.scala 165:174]
  wire [10:0] _GEN_3249 = io_SPI_distort ? _T_171 : {{7'd0}, _GEN_2672}; // @[Filter.scala 164:35]
  wire [10:0] _GEN_3250 = _T_151 ? 11'h0 : _GEN_3249; // @[Filter.scala 162:80]
  wire [10:0] _GEN_4019 = io_SPI_distort ? _T_171 : {{7'd0}, _GEN_2864}; // @[Filter.scala 164:35]
  wire [10:0] _GEN_4020 = _T_151 ? 11'h0 : _GEN_4019; // @[Filter.scala 162:80]
  wire [10:0] _GEN_4789 = io_SPI_distort ? _T_171 : {{7'd0}, _GEN_3056}; // @[Filter.scala 164:35]
  wire [10:0] _GEN_4790 = _T_151 ? 11'h0 : _GEN_4789; // @[Filter.scala 162:80]
  wire [31:0] _T_239 = pixelIndex + 32'h2; // @[Filter.scala 158:31]
  wire [31:0] _GEN_2 = _T_239 % 32'h10; // @[Filter.scala 158:38]
  wire [4:0] _T_240 = _GEN_2[4:0]; // @[Filter.scala 158:38]
  wire [4:0] _T_242 = _T_240 + _GEN_18983; // @[Filter.scala 158:53]
  wire [4:0] _T_244 = _T_242 - 5'h1; // @[Filter.scala 158:69]
  wire [31:0] _T_247 = _T_239 / 32'h10; // @[Filter.scala 159:38]
  wire [31:0] _T_249 = _T_247 + _GEN_18984; // @[Filter.scala 159:53]
  wire [31:0] _T_251 = _T_249 - 32'h1; // @[Filter.scala 159:69]
  wire  _T_253 = _T_244 >= 5'h10; // @[Filter.scala 162:31]
  wire  _T_257 = _T_251 >= 32'hc; // @[Filter.scala 162:63]
  wire  _T_258 = _T_253 | _T_257; // @[Filter.scala 162:58]
  wire [36:0] _T_259 = _T_251 * 32'h10; // @[Filter.scala 165:66]
  wire [36:0] _GEN_19037 = {{32'd0}, _T_244}; // @[Filter.scala 165:81]
  wire [36:0] _T_261 = _T_259 + _GEN_19037; // @[Filter.scala 165:81]
  wire [3:0] _GEN_4799 = 8'h8 == _T_261[7:0] ? 4'h0 : 4'hf; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4800 = 8'h9 == _T_261[7:0] ? 4'h0 : _GEN_4799; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4801 = 8'ha == _T_261[7:0] ? 4'h0 : _GEN_4800; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4802 = 8'hb == _T_261[7:0] ? 4'h0 : _GEN_4801; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4803 = 8'hc == _T_261[7:0] ? 4'h0 : _GEN_4802; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4804 = 8'hd == _T_261[7:0] ? 4'h0 : _GEN_4803; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4805 = 8'he == _T_261[7:0] ? 4'h0 : _GEN_4804; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4806 = 8'hf == _T_261[7:0] ? 4'h0 : _GEN_4805; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4807 = 8'h10 == _T_261[7:0] ? 4'hf : _GEN_4806; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4808 = 8'h11 == _T_261[7:0] ? 4'hf : _GEN_4807; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4809 = 8'h12 == _T_261[7:0] ? 4'hf : _GEN_4808; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4810 = 8'h13 == _T_261[7:0] ? 4'hf : _GEN_4809; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4811 = 8'h14 == _T_261[7:0] ? 4'hf : _GEN_4810; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4812 = 8'h15 == _T_261[7:0] ? 4'hf : _GEN_4811; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4813 = 8'h16 == _T_261[7:0] ? 4'hf : _GEN_4812; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4814 = 8'h17 == _T_261[7:0] ? 4'hf : _GEN_4813; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4815 = 8'h18 == _T_261[7:0] ? 4'h0 : _GEN_4814; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4816 = 8'h19 == _T_261[7:0] ? 4'h0 : _GEN_4815; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4817 = 8'h1a == _T_261[7:0] ? 4'h0 : _GEN_4816; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4818 = 8'h1b == _T_261[7:0] ? 4'h0 : _GEN_4817; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4819 = 8'h1c == _T_261[7:0] ? 4'h0 : _GEN_4818; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4820 = 8'h1d == _T_261[7:0] ? 4'h0 : _GEN_4819; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4821 = 8'h1e == _T_261[7:0] ? 4'h0 : _GEN_4820; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4822 = 8'h1f == _T_261[7:0] ? 4'h0 : _GEN_4821; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4823 = 8'h20 == _T_261[7:0] ? 4'hf : _GEN_4822; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4824 = 8'h21 == _T_261[7:0] ? 4'hf : _GEN_4823; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4825 = 8'h22 == _T_261[7:0] ? 4'hf : _GEN_4824; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4826 = 8'h23 == _T_261[7:0] ? 4'hf : _GEN_4825; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4827 = 8'h24 == _T_261[7:0] ? 4'hf : _GEN_4826; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4828 = 8'h25 == _T_261[7:0] ? 4'hf : _GEN_4827; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4829 = 8'h26 == _T_261[7:0] ? 4'hf : _GEN_4828; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4830 = 8'h27 == _T_261[7:0] ? 4'hf : _GEN_4829; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4831 = 8'h28 == _T_261[7:0] ? 4'h0 : _GEN_4830; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4832 = 8'h29 == _T_261[7:0] ? 4'h0 : _GEN_4831; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4833 = 8'h2a == _T_261[7:0] ? 4'h0 : _GEN_4832; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4834 = 8'h2b == _T_261[7:0] ? 4'h0 : _GEN_4833; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4835 = 8'h2c == _T_261[7:0] ? 4'h0 : _GEN_4834; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4836 = 8'h2d == _T_261[7:0] ? 4'h0 : _GEN_4835; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4837 = 8'h2e == _T_261[7:0] ? 4'h0 : _GEN_4836; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4838 = 8'h2f == _T_261[7:0] ? 4'h0 : _GEN_4837; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4839 = 8'h30 == _T_261[7:0] ? 4'hf : _GEN_4838; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4840 = 8'h31 == _T_261[7:0] ? 4'hf : _GEN_4839; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4841 = 8'h32 == _T_261[7:0] ? 4'hf : _GEN_4840; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4842 = 8'h33 == _T_261[7:0] ? 4'hf : _GEN_4841; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4843 = 8'h34 == _T_261[7:0] ? 4'hf : _GEN_4842; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4844 = 8'h35 == _T_261[7:0] ? 4'hf : _GEN_4843; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4845 = 8'h36 == _T_261[7:0] ? 4'hf : _GEN_4844; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4846 = 8'h37 == _T_261[7:0] ? 4'hf : _GEN_4845; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4847 = 8'h38 == _T_261[7:0] ? 4'h0 : _GEN_4846; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4848 = 8'h39 == _T_261[7:0] ? 4'h0 : _GEN_4847; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4849 = 8'h3a == _T_261[7:0] ? 4'h0 : _GEN_4848; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4850 = 8'h3b == _T_261[7:0] ? 4'h0 : _GEN_4849; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4851 = 8'h3c == _T_261[7:0] ? 4'h0 : _GEN_4850; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4852 = 8'h3d == _T_261[7:0] ? 4'h0 : _GEN_4851; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4853 = 8'h3e == _T_261[7:0] ? 4'h0 : _GEN_4852; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4854 = 8'h3f == _T_261[7:0] ? 4'h0 : _GEN_4853; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4855 = 8'h40 == _T_261[7:0] ? 4'hf : _GEN_4854; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4856 = 8'h41 == _T_261[7:0] ? 4'hf : _GEN_4855; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4857 = 8'h42 == _T_261[7:0] ? 4'hf : _GEN_4856; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4858 = 8'h43 == _T_261[7:0] ? 4'hf : _GEN_4857; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4859 = 8'h44 == _T_261[7:0] ? 4'hf : _GEN_4858; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4860 = 8'h45 == _T_261[7:0] ? 4'hf : _GEN_4859; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4861 = 8'h46 == _T_261[7:0] ? 4'hf : _GEN_4860; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4862 = 8'h47 == _T_261[7:0] ? 4'hf : _GEN_4861; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4863 = 8'h48 == _T_261[7:0] ? 4'h0 : _GEN_4862; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4864 = 8'h49 == _T_261[7:0] ? 4'h0 : _GEN_4863; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4865 = 8'h4a == _T_261[7:0] ? 4'h0 : _GEN_4864; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4866 = 8'h4b == _T_261[7:0] ? 4'h0 : _GEN_4865; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4867 = 8'h4c == _T_261[7:0] ? 4'h0 : _GEN_4866; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4868 = 8'h4d == _T_261[7:0] ? 4'h0 : _GEN_4867; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4869 = 8'h4e == _T_261[7:0] ? 4'h0 : _GEN_4868; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4870 = 8'h4f == _T_261[7:0] ? 4'h0 : _GEN_4869; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4871 = 8'h50 == _T_261[7:0] ? 4'hf : _GEN_4870; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4872 = 8'h51 == _T_261[7:0] ? 4'hf : _GEN_4871; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4873 = 8'h52 == _T_261[7:0] ? 4'hf : _GEN_4872; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4874 = 8'h53 == _T_261[7:0] ? 4'hf : _GEN_4873; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4875 = 8'h54 == _T_261[7:0] ? 4'hf : _GEN_4874; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4876 = 8'h55 == _T_261[7:0] ? 4'hf : _GEN_4875; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4877 = 8'h56 == _T_261[7:0] ? 4'hf : _GEN_4876; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4878 = 8'h57 == _T_261[7:0] ? 4'hf : _GEN_4877; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4879 = 8'h58 == _T_261[7:0] ? 4'h0 : _GEN_4878; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4880 = 8'h59 == _T_261[7:0] ? 4'h0 : _GEN_4879; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4881 = 8'h5a == _T_261[7:0] ? 4'h0 : _GEN_4880; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4882 = 8'h5b == _T_261[7:0] ? 4'h0 : _GEN_4881; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4883 = 8'h5c == _T_261[7:0] ? 4'h0 : _GEN_4882; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4884 = 8'h5d == _T_261[7:0] ? 4'h0 : _GEN_4883; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4885 = 8'h5e == _T_261[7:0] ? 4'h0 : _GEN_4884; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4886 = 8'h5f == _T_261[7:0] ? 4'h0 : _GEN_4885; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4887 = 8'h60 == _T_261[7:0] ? 4'h0 : _GEN_4886; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4888 = 8'h61 == _T_261[7:0] ? 4'h0 : _GEN_4887; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4889 = 8'h62 == _T_261[7:0] ? 4'h0 : _GEN_4888; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4890 = 8'h63 == _T_261[7:0] ? 4'h0 : _GEN_4889; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4891 = 8'h64 == _T_261[7:0] ? 4'h0 : _GEN_4890; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4892 = 8'h65 == _T_261[7:0] ? 4'h0 : _GEN_4891; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4893 = 8'h66 == _T_261[7:0] ? 4'h0 : _GEN_4892; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4894 = 8'h67 == _T_261[7:0] ? 4'h0 : _GEN_4893; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4895 = 8'h68 == _T_261[7:0] ? 4'hf : _GEN_4894; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4896 = 8'h69 == _T_261[7:0] ? 4'hf : _GEN_4895; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4897 = 8'h6a == _T_261[7:0] ? 4'hf : _GEN_4896; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4898 = 8'h6b == _T_261[7:0] ? 4'hf : _GEN_4897; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4899 = 8'h6c == _T_261[7:0] ? 4'hf : _GEN_4898; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4900 = 8'h6d == _T_261[7:0] ? 4'hf : _GEN_4899; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4901 = 8'h6e == _T_261[7:0] ? 4'hf : _GEN_4900; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4902 = 8'h6f == _T_261[7:0] ? 4'hf : _GEN_4901; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4903 = 8'h70 == _T_261[7:0] ? 4'h0 : _GEN_4902; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4904 = 8'h71 == _T_261[7:0] ? 4'h0 : _GEN_4903; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4905 = 8'h72 == _T_261[7:0] ? 4'h0 : _GEN_4904; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4906 = 8'h73 == _T_261[7:0] ? 4'h0 : _GEN_4905; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4907 = 8'h74 == _T_261[7:0] ? 4'h0 : _GEN_4906; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4908 = 8'h75 == _T_261[7:0] ? 4'h0 : _GEN_4907; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4909 = 8'h76 == _T_261[7:0] ? 4'h0 : _GEN_4908; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4910 = 8'h77 == _T_261[7:0] ? 4'h0 : _GEN_4909; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4911 = 8'h78 == _T_261[7:0] ? 4'hf : _GEN_4910; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4912 = 8'h79 == _T_261[7:0] ? 4'hf : _GEN_4911; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4913 = 8'h7a == _T_261[7:0] ? 4'hf : _GEN_4912; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4914 = 8'h7b == _T_261[7:0] ? 4'hf : _GEN_4913; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4915 = 8'h7c == _T_261[7:0] ? 4'hf : _GEN_4914; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4916 = 8'h7d == _T_261[7:0] ? 4'hf : _GEN_4915; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4917 = 8'h7e == _T_261[7:0] ? 4'hf : _GEN_4916; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4918 = 8'h7f == _T_261[7:0] ? 4'hf : _GEN_4917; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4919 = 8'h80 == _T_261[7:0] ? 4'h0 : _GEN_4918; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4920 = 8'h81 == _T_261[7:0] ? 4'h0 : _GEN_4919; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4921 = 8'h82 == _T_261[7:0] ? 4'h0 : _GEN_4920; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4922 = 8'h83 == _T_261[7:0] ? 4'h0 : _GEN_4921; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4923 = 8'h84 == _T_261[7:0] ? 4'h0 : _GEN_4922; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4924 = 8'h85 == _T_261[7:0] ? 4'h0 : _GEN_4923; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4925 = 8'h86 == _T_261[7:0] ? 4'h0 : _GEN_4924; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4926 = 8'h87 == _T_261[7:0] ? 4'h0 : _GEN_4925; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4927 = 8'h88 == _T_261[7:0] ? 4'hf : _GEN_4926; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4928 = 8'h89 == _T_261[7:0] ? 4'hf : _GEN_4927; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4929 = 8'h8a == _T_261[7:0] ? 4'hf : _GEN_4928; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4930 = 8'h8b == _T_261[7:0] ? 4'hf : _GEN_4929; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4931 = 8'h8c == _T_261[7:0] ? 4'hf : _GEN_4930; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4932 = 8'h8d == _T_261[7:0] ? 4'hf : _GEN_4931; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4933 = 8'h8e == _T_261[7:0] ? 4'hf : _GEN_4932; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4934 = 8'h8f == _T_261[7:0] ? 4'hf : _GEN_4933; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4935 = 8'h90 == _T_261[7:0] ? 4'h0 : _GEN_4934; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4936 = 8'h91 == _T_261[7:0] ? 4'h0 : _GEN_4935; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4937 = 8'h92 == _T_261[7:0] ? 4'h0 : _GEN_4936; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4938 = 8'h93 == _T_261[7:0] ? 4'h0 : _GEN_4937; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4939 = 8'h94 == _T_261[7:0] ? 4'h0 : _GEN_4938; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4940 = 8'h95 == _T_261[7:0] ? 4'h0 : _GEN_4939; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4941 = 8'h96 == _T_261[7:0] ? 4'h0 : _GEN_4940; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4942 = 8'h97 == _T_261[7:0] ? 4'h0 : _GEN_4941; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4943 = 8'h98 == _T_261[7:0] ? 4'hf : _GEN_4942; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4944 = 8'h99 == _T_261[7:0] ? 4'hf : _GEN_4943; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4945 = 8'h9a == _T_261[7:0] ? 4'hf : _GEN_4944; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4946 = 8'h9b == _T_261[7:0] ? 4'hf : _GEN_4945; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4947 = 8'h9c == _T_261[7:0] ? 4'hf : _GEN_4946; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4948 = 8'h9d == _T_261[7:0] ? 4'hf : _GEN_4947; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4949 = 8'h9e == _T_261[7:0] ? 4'hf : _GEN_4948; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4950 = 8'h9f == _T_261[7:0] ? 4'hf : _GEN_4949; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4951 = 8'ha0 == _T_261[7:0] ? 4'h0 : _GEN_4950; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4952 = 8'ha1 == _T_261[7:0] ? 4'h0 : _GEN_4951; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4953 = 8'ha2 == _T_261[7:0] ? 4'h0 : _GEN_4952; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4954 = 8'ha3 == _T_261[7:0] ? 4'h0 : _GEN_4953; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4955 = 8'ha4 == _T_261[7:0] ? 4'h0 : _GEN_4954; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4956 = 8'ha5 == _T_261[7:0] ? 4'h0 : _GEN_4955; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4957 = 8'ha6 == _T_261[7:0] ? 4'h0 : _GEN_4956; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4958 = 8'ha7 == _T_261[7:0] ? 4'h0 : _GEN_4957; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4959 = 8'ha8 == _T_261[7:0] ? 4'hf : _GEN_4958; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4960 = 8'ha9 == _T_261[7:0] ? 4'hf : _GEN_4959; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4961 = 8'haa == _T_261[7:0] ? 4'hf : _GEN_4960; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4962 = 8'hab == _T_261[7:0] ? 4'hf : _GEN_4961; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4963 = 8'hac == _T_261[7:0] ? 4'hf : _GEN_4962; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4964 = 8'had == _T_261[7:0] ? 4'hf : _GEN_4963; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4965 = 8'hae == _T_261[7:0] ? 4'hf : _GEN_4964; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4966 = 8'haf == _T_261[7:0] ? 4'hf : _GEN_4965; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4967 = 8'hb0 == _T_261[7:0] ? 4'h0 : _GEN_4966; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4968 = 8'hb1 == _T_261[7:0] ? 4'h0 : _GEN_4967; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4969 = 8'hb2 == _T_261[7:0] ? 4'h0 : _GEN_4968; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4970 = 8'hb3 == _T_261[7:0] ? 4'h0 : _GEN_4969; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4971 = 8'hb4 == _T_261[7:0] ? 4'h0 : _GEN_4970; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4972 = 8'hb5 == _T_261[7:0] ? 4'h0 : _GEN_4971; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4973 = 8'hb6 == _T_261[7:0] ? 4'h0 : _GEN_4972; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4974 = 8'hb7 == _T_261[7:0] ? 4'h0 : _GEN_4973; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4975 = 8'hb8 == _T_261[7:0] ? 4'hf : _GEN_4974; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4976 = 8'hb9 == _T_261[7:0] ? 4'hf : _GEN_4975; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4977 = 8'hba == _T_261[7:0] ? 4'hf : _GEN_4976; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4978 = 8'hbb == _T_261[7:0] ? 4'hf : _GEN_4977; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4979 = 8'hbc == _T_261[7:0] ? 4'hf : _GEN_4978; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4980 = 8'hbd == _T_261[7:0] ? 4'hf : _GEN_4979; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4981 = 8'hbe == _T_261[7:0] ? 4'hf : _GEN_4980; // @[Filter.scala 165:86]
  wire [3:0] _GEN_4982 = 8'hbf == _T_261[7:0] ? 4'hf : _GEN_4981; // @[Filter.scala 165:86]
  wire [4:0] _GEN_19038 = {{1'd0}, _GEN_4982}; // @[Filter.scala 165:86]
  wire [8:0] _T_263 = _GEN_19038 * 5'h14; // @[Filter.scala 165:86]
  wire [3:0] _GEN_5079 = 8'h60 == _T_261[7:0] ? 4'hf : 4'h0; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5080 = 8'h61 == _T_261[7:0] ? 4'hf : _GEN_5079; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5081 = 8'h62 == _T_261[7:0] ? 4'hf : _GEN_5080; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5082 = 8'h63 == _T_261[7:0] ? 4'hf : _GEN_5081; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5083 = 8'h64 == _T_261[7:0] ? 4'hf : _GEN_5082; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5084 = 8'h65 == _T_261[7:0] ? 4'hf : _GEN_5083; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5085 = 8'h66 == _T_261[7:0] ? 4'hf : _GEN_5084; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5086 = 8'h67 == _T_261[7:0] ? 4'hf : _GEN_5085; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5087 = 8'h68 == _T_261[7:0] ? 4'hf : _GEN_5086; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5088 = 8'h69 == _T_261[7:0] ? 4'hf : _GEN_5087; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5089 = 8'h6a == _T_261[7:0] ? 4'hf : _GEN_5088; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5090 = 8'h6b == _T_261[7:0] ? 4'hf : _GEN_5089; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5091 = 8'h6c == _T_261[7:0] ? 4'hf : _GEN_5090; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5092 = 8'h6d == _T_261[7:0] ? 4'hf : _GEN_5091; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5093 = 8'h6e == _T_261[7:0] ? 4'hf : _GEN_5092; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5094 = 8'h6f == _T_261[7:0] ? 4'hf : _GEN_5093; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5095 = 8'h70 == _T_261[7:0] ? 4'hf : _GEN_5094; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5096 = 8'h71 == _T_261[7:0] ? 4'hf : _GEN_5095; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5097 = 8'h72 == _T_261[7:0] ? 4'hf : _GEN_5096; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5098 = 8'h73 == _T_261[7:0] ? 4'hf : _GEN_5097; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5099 = 8'h74 == _T_261[7:0] ? 4'hf : _GEN_5098; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5100 = 8'h75 == _T_261[7:0] ? 4'hf : _GEN_5099; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5101 = 8'h76 == _T_261[7:0] ? 4'hf : _GEN_5100; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5102 = 8'h77 == _T_261[7:0] ? 4'hf : _GEN_5101; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5103 = 8'h78 == _T_261[7:0] ? 4'hf : _GEN_5102; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5104 = 8'h79 == _T_261[7:0] ? 4'hf : _GEN_5103; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5105 = 8'h7a == _T_261[7:0] ? 4'hf : _GEN_5104; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5106 = 8'h7b == _T_261[7:0] ? 4'hf : _GEN_5105; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5107 = 8'h7c == _T_261[7:0] ? 4'hf : _GEN_5106; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5108 = 8'h7d == _T_261[7:0] ? 4'hf : _GEN_5107; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5109 = 8'h7e == _T_261[7:0] ? 4'hf : _GEN_5108; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5110 = 8'h7f == _T_261[7:0] ? 4'hf : _GEN_5109; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5111 = 8'h80 == _T_261[7:0] ? 4'hf : _GEN_5110; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5112 = 8'h81 == _T_261[7:0] ? 4'hf : _GEN_5111; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5113 = 8'h82 == _T_261[7:0] ? 4'hf : _GEN_5112; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5114 = 8'h83 == _T_261[7:0] ? 4'hf : _GEN_5113; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5115 = 8'h84 == _T_261[7:0] ? 4'hf : _GEN_5114; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5116 = 8'h85 == _T_261[7:0] ? 4'hf : _GEN_5115; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5117 = 8'h86 == _T_261[7:0] ? 4'hf : _GEN_5116; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5118 = 8'h87 == _T_261[7:0] ? 4'hf : _GEN_5117; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5119 = 8'h88 == _T_261[7:0] ? 4'hf : _GEN_5118; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5120 = 8'h89 == _T_261[7:0] ? 4'hf : _GEN_5119; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5121 = 8'h8a == _T_261[7:0] ? 4'hf : _GEN_5120; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5122 = 8'h8b == _T_261[7:0] ? 4'hf : _GEN_5121; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5123 = 8'h8c == _T_261[7:0] ? 4'hf : _GEN_5122; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5124 = 8'h8d == _T_261[7:0] ? 4'hf : _GEN_5123; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5125 = 8'h8e == _T_261[7:0] ? 4'hf : _GEN_5124; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5126 = 8'h8f == _T_261[7:0] ? 4'hf : _GEN_5125; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5127 = 8'h90 == _T_261[7:0] ? 4'hf : _GEN_5126; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5128 = 8'h91 == _T_261[7:0] ? 4'hf : _GEN_5127; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5129 = 8'h92 == _T_261[7:0] ? 4'hf : _GEN_5128; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5130 = 8'h93 == _T_261[7:0] ? 4'hf : _GEN_5129; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5131 = 8'h94 == _T_261[7:0] ? 4'hf : _GEN_5130; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5132 = 8'h95 == _T_261[7:0] ? 4'hf : _GEN_5131; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5133 = 8'h96 == _T_261[7:0] ? 4'hf : _GEN_5132; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5134 = 8'h97 == _T_261[7:0] ? 4'hf : _GEN_5133; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5135 = 8'h98 == _T_261[7:0] ? 4'hf : _GEN_5134; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5136 = 8'h99 == _T_261[7:0] ? 4'hf : _GEN_5135; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5137 = 8'h9a == _T_261[7:0] ? 4'hf : _GEN_5136; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5138 = 8'h9b == _T_261[7:0] ? 4'hf : _GEN_5137; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5139 = 8'h9c == _T_261[7:0] ? 4'hf : _GEN_5138; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5140 = 8'h9d == _T_261[7:0] ? 4'hf : _GEN_5139; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5141 = 8'h9e == _T_261[7:0] ? 4'hf : _GEN_5140; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5142 = 8'h9f == _T_261[7:0] ? 4'hf : _GEN_5141; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5143 = 8'ha0 == _T_261[7:0] ? 4'hf : _GEN_5142; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5144 = 8'ha1 == _T_261[7:0] ? 4'hf : _GEN_5143; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5145 = 8'ha2 == _T_261[7:0] ? 4'hf : _GEN_5144; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5146 = 8'ha3 == _T_261[7:0] ? 4'hf : _GEN_5145; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5147 = 8'ha4 == _T_261[7:0] ? 4'hf : _GEN_5146; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5148 = 8'ha5 == _T_261[7:0] ? 4'hf : _GEN_5147; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5149 = 8'ha6 == _T_261[7:0] ? 4'hf : _GEN_5148; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5150 = 8'ha7 == _T_261[7:0] ? 4'hf : _GEN_5149; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5151 = 8'ha8 == _T_261[7:0] ? 4'hf : _GEN_5150; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5152 = 8'ha9 == _T_261[7:0] ? 4'hf : _GEN_5151; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5153 = 8'haa == _T_261[7:0] ? 4'hf : _GEN_5152; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5154 = 8'hab == _T_261[7:0] ? 4'hf : _GEN_5153; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5155 = 8'hac == _T_261[7:0] ? 4'hf : _GEN_5154; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5156 = 8'had == _T_261[7:0] ? 4'hf : _GEN_5155; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5157 = 8'hae == _T_261[7:0] ? 4'hf : _GEN_5156; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5158 = 8'haf == _T_261[7:0] ? 4'hf : _GEN_5157; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5159 = 8'hb0 == _T_261[7:0] ? 4'hf : _GEN_5158; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5160 = 8'hb1 == _T_261[7:0] ? 4'hf : _GEN_5159; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5161 = 8'hb2 == _T_261[7:0] ? 4'hf : _GEN_5160; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5162 = 8'hb3 == _T_261[7:0] ? 4'hf : _GEN_5161; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5163 = 8'hb4 == _T_261[7:0] ? 4'hf : _GEN_5162; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5164 = 8'hb5 == _T_261[7:0] ? 4'hf : _GEN_5163; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5165 = 8'hb6 == _T_261[7:0] ? 4'hf : _GEN_5164; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5166 = 8'hb7 == _T_261[7:0] ? 4'hf : _GEN_5165; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5167 = 8'hb8 == _T_261[7:0] ? 4'hf : _GEN_5166; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5168 = 8'hb9 == _T_261[7:0] ? 4'hf : _GEN_5167; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5169 = 8'hba == _T_261[7:0] ? 4'hf : _GEN_5168; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5170 = 8'hbb == _T_261[7:0] ? 4'hf : _GEN_5169; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5171 = 8'hbc == _T_261[7:0] ? 4'hf : _GEN_5170; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5172 = 8'hbd == _T_261[7:0] ? 4'hf : _GEN_5171; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5173 = 8'hbe == _T_261[7:0] ? 4'hf : _GEN_5172; // @[Filter.scala 165:126]
  wire [3:0] _GEN_5174 = 8'hbf == _T_261[7:0] ? 4'hf : _GEN_5173; // @[Filter.scala 165:126]
  wire [6:0] _GEN_19040 = {{3'd0}, _GEN_5174}; // @[Filter.scala 165:126]
  wire [10:0] _T_268 = _GEN_19040 * 7'h46; // @[Filter.scala 165:126]
  wire [10:0] _GEN_19041 = {{2'd0}, _T_263}; // @[Filter.scala 165:93]
  wire [10:0] _T_270 = _GEN_19041 + _T_268; // @[Filter.scala 165:93]
  wire [3:0] _GEN_5183 = 8'h8 == _T_261[7:0] ? 4'hf : 4'h0; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5184 = 8'h9 == _T_261[7:0] ? 4'hf : _GEN_5183; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5185 = 8'ha == _T_261[7:0] ? 4'hf : _GEN_5184; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5186 = 8'hb == _T_261[7:0] ? 4'hf : _GEN_5185; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5187 = 8'hc == _T_261[7:0] ? 4'hf : _GEN_5186; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5188 = 8'hd == _T_261[7:0] ? 4'hf : _GEN_5187; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5189 = 8'he == _T_261[7:0] ? 4'hf : _GEN_5188; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5190 = 8'hf == _T_261[7:0] ? 4'hf : _GEN_5189; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5191 = 8'h10 == _T_261[7:0] ? 4'h0 : _GEN_5190; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5192 = 8'h11 == _T_261[7:0] ? 4'h0 : _GEN_5191; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5193 = 8'h12 == _T_261[7:0] ? 4'h0 : _GEN_5192; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5194 = 8'h13 == _T_261[7:0] ? 4'h0 : _GEN_5193; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5195 = 8'h14 == _T_261[7:0] ? 4'h0 : _GEN_5194; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5196 = 8'h15 == _T_261[7:0] ? 4'h0 : _GEN_5195; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5197 = 8'h16 == _T_261[7:0] ? 4'h0 : _GEN_5196; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5198 = 8'h17 == _T_261[7:0] ? 4'h0 : _GEN_5197; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5199 = 8'h18 == _T_261[7:0] ? 4'hf : _GEN_5198; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5200 = 8'h19 == _T_261[7:0] ? 4'hf : _GEN_5199; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5201 = 8'h1a == _T_261[7:0] ? 4'hf : _GEN_5200; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5202 = 8'h1b == _T_261[7:0] ? 4'hf : _GEN_5201; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5203 = 8'h1c == _T_261[7:0] ? 4'hf : _GEN_5202; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5204 = 8'h1d == _T_261[7:0] ? 4'hf : _GEN_5203; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5205 = 8'h1e == _T_261[7:0] ? 4'hf : _GEN_5204; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5206 = 8'h1f == _T_261[7:0] ? 4'hf : _GEN_5205; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5207 = 8'h20 == _T_261[7:0] ? 4'h0 : _GEN_5206; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5208 = 8'h21 == _T_261[7:0] ? 4'h0 : _GEN_5207; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5209 = 8'h22 == _T_261[7:0] ? 4'h0 : _GEN_5208; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5210 = 8'h23 == _T_261[7:0] ? 4'h0 : _GEN_5209; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5211 = 8'h24 == _T_261[7:0] ? 4'h0 : _GEN_5210; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5212 = 8'h25 == _T_261[7:0] ? 4'h0 : _GEN_5211; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5213 = 8'h26 == _T_261[7:0] ? 4'h0 : _GEN_5212; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5214 = 8'h27 == _T_261[7:0] ? 4'h0 : _GEN_5213; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5215 = 8'h28 == _T_261[7:0] ? 4'hf : _GEN_5214; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5216 = 8'h29 == _T_261[7:0] ? 4'hf : _GEN_5215; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5217 = 8'h2a == _T_261[7:0] ? 4'hf : _GEN_5216; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5218 = 8'h2b == _T_261[7:0] ? 4'hf : _GEN_5217; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5219 = 8'h2c == _T_261[7:0] ? 4'hf : _GEN_5218; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5220 = 8'h2d == _T_261[7:0] ? 4'hf : _GEN_5219; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5221 = 8'h2e == _T_261[7:0] ? 4'hf : _GEN_5220; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5222 = 8'h2f == _T_261[7:0] ? 4'hf : _GEN_5221; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5223 = 8'h30 == _T_261[7:0] ? 4'h0 : _GEN_5222; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5224 = 8'h31 == _T_261[7:0] ? 4'h0 : _GEN_5223; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5225 = 8'h32 == _T_261[7:0] ? 4'h0 : _GEN_5224; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5226 = 8'h33 == _T_261[7:0] ? 4'h0 : _GEN_5225; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5227 = 8'h34 == _T_261[7:0] ? 4'h0 : _GEN_5226; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5228 = 8'h35 == _T_261[7:0] ? 4'h0 : _GEN_5227; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5229 = 8'h36 == _T_261[7:0] ? 4'h0 : _GEN_5228; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5230 = 8'h37 == _T_261[7:0] ? 4'h0 : _GEN_5229; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5231 = 8'h38 == _T_261[7:0] ? 4'hf : _GEN_5230; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5232 = 8'h39 == _T_261[7:0] ? 4'hf : _GEN_5231; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5233 = 8'h3a == _T_261[7:0] ? 4'hf : _GEN_5232; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5234 = 8'h3b == _T_261[7:0] ? 4'hf : _GEN_5233; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5235 = 8'h3c == _T_261[7:0] ? 4'hf : _GEN_5234; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5236 = 8'h3d == _T_261[7:0] ? 4'hf : _GEN_5235; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5237 = 8'h3e == _T_261[7:0] ? 4'hf : _GEN_5236; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5238 = 8'h3f == _T_261[7:0] ? 4'hf : _GEN_5237; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5239 = 8'h40 == _T_261[7:0] ? 4'h0 : _GEN_5238; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5240 = 8'h41 == _T_261[7:0] ? 4'h0 : _GEN_5239; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5241 = 8'h42 == _T_261[7:0] ? 4'h0 : _GEN_5240; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5242 = 8'h43 == _T_261[7:0] ? 4'h0 : _GEN_5241; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5243 = 8'h44 == _T_261[7:0] ? 4'h0 : _GEN_5242; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5244 = 8'h45 == _T_261[7:0] ? 4'h0 : _GEN_5243; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5245 = 8'h46 == _T_261[7:0] ? 4'h0 : _GEN_5244; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5246 = 8'h47 == _T_261[7:0] ? 4'h0 : _GEN_5245; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5247 = 8'h48 == _T_261[7:0] ? 4'hf : _GEN_5246; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5248 = 8'h49 == _T_261[7:0] ? 4'hf : _GEN_5247; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5249 = 8'h4a == _T_261[7:0] ? 4'hf : _GEN_5248; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5250 = 8'h4b == _T_261[7:0] ? 4'hf : _GEN_5249; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5251 = 8'h4c == _T_261[7:0] ? 4'hf : _GEN_5250; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5252 = 8'h4d == _T_261[7:0] ? 4'hf : _GEN_5251; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5253 = 8'h4e == _T_261[7:0] ? 4'hf : _GEN_5252; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5254 = 8'h4f == _T_261[7:0] ? 4'hf : _GEN_5253; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5255 = 8'h50 == _T_261[7:0] ? 4'h0 : _GEN_5254; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5256 = 8'h51 == _T_261[7:0] ? 4'h0 : _GEN_5255; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5257 = 8'h52 == _T_261[7:0] ? 4'h0 : _GEN_5256; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5258 = 8'h53 == _T_261[7:0] ? 4'h0 : _GEN_5257; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5259 = 8'h54 == _T_261[7:0] ? 4'h0 : _GEN_5258; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5260 = 8'h55 == _T_261[7:0] ? 4'h0 : _GEN_5259; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5261 = 8'h56 == _T_261[7:0] ? 4'h0 : _GEN_5260; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5262 = 8'h57 == _T_261[7:0] ? 4'h0 : _GEN_5261; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5263 = 8'h58 == _T_261[7:0] ? 4'hf : _GEN_5262; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5264 = 8'h59 == _T_261[7:0] ? 4'hf : _GEN_5263; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5265 = 8'h5a == _T_261[7:0] ? 4'hf : _GEN_5264; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5266 = 8'h5b == _T_261[7:0] ? 4'hf : _GEN_5265; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5267 = 8'h5c == _T_261[7:0] ? 4'hf : _GEN_5266; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5268 = 8'h5d == _T_261[7:0] ? 4'hf : _GEN_5267; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5269 = 8'h5e == _T_261[7:0] ? 4'hf : _GEN_5268; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5270 = 8'h5f == _T_261[7:0] ? 4'hf : _GEN_5269; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5271 = 8'h60 == _T_261[7:0] ? 4'h0 : _GEN_5270; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5272 = 8'h61 == _T_261[7:0] ? 4'h0 : _GEN_5271; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5273 = 8'h62 == _T_261[7:0] ? 4'h0 : _GEN_5272; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5274 = 8'h63 == _T_261[7:0] ? 4'h0 : _GEN_5273; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5275 = 8'h64 == _T_261[7:0] ? 4'h0 : _GEN_5274; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5276 = 8'h65 == _T_261[7:0] ? 4'h0 : _GEN_5275; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5277 = 8'h66 == _T_261[7:0] ? 4'h0 : _GEN_5276; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5278 = 8'h67 == _T_261[7:0] ? 4'h0 : _GEN_5277; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5279 = 8'h68 == _T_261[7:0] ? 4'hf : _GEN_5278; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5280 = 8'h69 == _T_261[7:0] ? 4'hf : _GEN_5279; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5281 = 8'h6a == _T_261[7:0] ? 4'hf : _GEN_5280; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5282 = 8'h6b == _T_261[7:0] ? 4'hf : _GEN_5281; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5283 = 8'h6c == _T_261[7:0] ? 4'hf : _GEN_5282; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5284 = 8'h6d == _T_261[7:0] ? 4'hf : _GEN_5283; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5285 = 8'h6e == _T_261[7:0] ? 4'hf : _GEN_5284; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5286 = 8'h6f == _T_261[7:0] ? 4'hf : _GEN_5285; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5287 = 8'h70 == _T_261[7:0] ? 4'h0 : _GEN_5286; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5288 = 8'h71 == _T_261[7:0] ? 4'h0 : _GEN_5287; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5289 = 8'h72 == _T_261[7:0] ? 4'h0 : _GEN_5288; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5290 = 8'h73 == _T_261[7:0] ? 4'h0 : _GEN_5289; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5291 = 8'h74 == _T_261[7:0] ? 4'h0 : _GEN_5290; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5292 = 8'h75 == _T_261[7:0] ? 4'h0 : _GEN_5291; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5293 = 8'h76 == _T_261[7:0] ? 4'h0 : _GEN_5292; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5294 = 8'h77 == _T_261[7:0] ? 4'h0 : _GEN_5293; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5295 = 8'h78 == _T_261[7:0] ? 4'hf : _GEN_5294; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5296 = 8'h79 == _T_261[7:0] ? 4'hf : _GEN_5295; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5297 = 8'h7a == _T_261[7:0] ? 4'hf : _GEN_5296; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5298 = 8'h7b == _T_261[7:0] ? 4'hf : _GEN_5297; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5299 = 8'h7c == _T_261[7:0] ? 4'hf : _GEN_5298; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5300 = 8'h7d == _T_261[7:0] ? 4'hf : _GEN_5299; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5301 = 8'h7e == _T_261[7:0] ? 4'hf : _GEN_5300; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5302 = 8'h7f == _T_261[7:0] ? 4'hf : _GEN_5301; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5303 = 8'h80 == _T_261[7:0] ? 4'h0 : _GEN_5302; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5304 = 8'h81 == _T_261[7:0] ? 4'h0 : _GEN_5303; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5305 = 8'h82 == _T_261[7:0] ? 4'h0 : _GEN_5304; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5306 = 8'h83 == _T_261[7:0] ? 4'h0 : _GEN_5305; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5307 = 8'h84 == _T_261[7:0] ? 4'h0 : _GEN_5306; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5308 = 8'h85 == _T_261[7:0] ? 4'h0 : _GEN_5307; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5309 = 8'h86 == _T_261[7:0] ? 4'h0 : _GEN_5308; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5310 = 8'h87 == _T_261[7:0] ? 4'h0 : _GEN_5309; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5311 = 8'h88 == _T_261[7:0] ? 4'hf : _GEN_5310; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5312 = 8'h89 == _T_261[7:0] ? 4'hf : _GEN_5311; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5313 = 8'h8a == _T_261[7:0] ? 4'hf : _GEN_5312; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5314 = 8'h8b == _T_261[7:0] ? 4'hf : _GEN_5313; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5315 = 8'h8c == _T_261[7:0] ? 4'hf : _GEN_5314; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5316 = 8'h8d == _T_261[7:0] ? 4'hf : _GEN_5315; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5317 = 8'h8e == _T_261[7:0] ? 4'hf : _GEN_5316; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5318 = 8'h8f == _T_261[7:0] ? 4'hf : _GEN_5317; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5319 = 8'h90 == _T_261[7:0] ? 4'h0 : _GEN_5318; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5320 = 8'h91 == _T_261[7:0] ? 4'h0 : _GEN_5319; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5321 = 8'h92 == _T_261[7:0] ? 4'h0 : _GEN_5320; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5322 = 8'h93 == _T_261[7:0] ? 4'h0 : _GEN_5321; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5323 = 8'h94 == _T_261[7:0] ? 4'h0 : _GEN_5322; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5324 = 8'h95 == _T_261[7:0] ? 4'h0 : _GEN_5323; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5325 = 8'h96 == _T_261[7:0] ? 4'h0 : _GEN_5324; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5326 = 8'h97 == _T_261[7:0] ? 4'h0 : _GEN_5325; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5327 = 8'h98 == _T_261[7:0] ? 4'hf : _GEN_5326; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5328 = 8'h99 == _T_261[7:0] ? 4'hf : _GEN_5327; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5329 = 8'h9a == _T_261[7:0] ? 4'hf : _GEN_5328; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5330 = 8'h9b == _T_261[7:0] ? 4'hf : _GEN_5329; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5331 = 8'h9c == _T_261[7:0] ? 4'hf : _GEN_5330; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5332 = 8'h9d == _T_261[7:0] ? 4'hf : _GEN_5331; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5333 = 8'h9e == _T_261[7:0] ? 4'hf : _GEN_5332; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5334 = 8'h9f == _T_261[7:0] ? 4'hf : _GEN_5333; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5335 = 8'ha0 == _T_261[7:0] ? 4'h0 : _GEN_5334; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5336 = 8'ha1 == _T_261[7:0] ? 4'h0 : _GEN_5335; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5337 = 8'ha2 == _T_261[7:0] ? 4'h0 : _GEN_5336; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5338 = 8'ha3 == _T_261[7:0] ? 4'h0 : _GEN_5337; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5339 = 8'ha4 == _T_261[7:0] ? 4'h0 : _GEN_5338; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5340 = 8'ha5 == _T_261[7:0] ? 4'h0 : _GEN_5339; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5341 = 8'ha6 == _T_261[7:0] ? 4'h0 : _GEN_5340; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5342 = 8'ha7 == _T_261[7:0] ? 4'h0 : _GEN_5341; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5343 = 8'ha8 == _T_261[7:0] ? 4'hf : _GEN_5342; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5344 = 8'ha9 == _T_261[7:0] ? 4'hf : _GEN_5343; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5345 = 8'haa == _T_261[7:0] ? 4'hf : _GEN_5344; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5346 = 8'hab == _T_261[7:0] ? 4'hf : _GEN_5345; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5347 = 8'hac == _T_261[7:0] ? 4'hf : _GEN_5346; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5348 = 8'had == _T_261[7:0] ? 4'hf : _GEN_5347; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5349 = 8'hae == _T_261[7:0] ? 4'hf : _GEN_5348; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5350 = 8'haf == _T_261[7:0] ? 4'hf : _GEN_5349; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5351 = 8'hb0 == _T_261[7:0] ? 4'h0 : _GEN_5350; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5352 = 8'hb1 == _T_261[7:0] ? 4'h0 : _GEN_5351; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5353 = 8'hb2 == _T_261[7:0] ? 4'h0 : _GEN_5352; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5354 = 8'hb3 == _T_261[7:0] ? 4'h0 : _GEN_5353; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5355 = 8'hb4 == _T_261[7:0] ? 4'h0 : _GEN_5354; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5356 = 8'hb5 == _T_261[7:0] ? 4'h0 : _GEN_5355; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5357 = 8'hb6 == _T_261[7:0] ? 4'h0 : _GEN_5356; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5358 = 8'hb7 == _T_261[7:0] ? 4'h0 : _GEN_5357; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5359 = 8'hb8 == _T_261[7:0] ? 4'hf : _GEN_5358; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5360 = 8'hb9 == _T_261[7:0] ? 4'hf : _GEN_5359; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5361 = 8'hba == _T_261[7:0] ? 4'hf : _GEN_5360; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5362 = 8'hbb == _T_261[7:0] ? 4'hf : _GEN_5361; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5363 = 8'hbc == _T_261[7:0] ? 4'hf : _GEN_5362; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5364 = 8'hbd == _T_261[7:0] ? 4'hf : _GEN_5363; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5365 = 8'hbe == _T_261[7:0] ? 4'hf : _GEN_5364; // @[Filter.scala 165:166]
  wire [3:0] _GEN_5366 = 8'hbf == _T_261[7:0] ? 4'hf : _GEN_5365; // @[Filter.scala 165:166]
  wire [7:0] _T_275 = _GEN_5366 * 4'ha; // @[Filter.scala 165:166]
  wire [10:0] _GEN_19043 = {{3'd0}, _T_275}; // @[Filter.scala 165:133]
  wire [10:0] _T_277 = _T_270 + _GEN_19043; // @[Filter.scala 165:133]
  wire [10:0] _T_278 = _T_277 / 11'h64; // @[Filter.scala 165:174]
  wire [10:0] _GEN_5559 = io_SPI_distort ? _T_278 : {{7'd0}, _GEN_4982}; // @[Filter.scala 164:35]
  wire [10:0] _GEN_5560 = _T_258 ? 11'h0 : _GEN_5559; // @[Filter.scala 162:80]
  wire [10:0] _GEN_6329 = io_SPI_distort ? _T_278 : {{7'd0}, _GEN_5174}; // @[Filter.scala 164:35]
  wire [10:0] _GEN_6330 = _T_258 ? 11'h0 : _GEN_6329; // @[Filter.scala 162:80]
  wire [10:0] _GEN_7099 = io_SPI_distort ? _T_278 : {{7'd0}, _GEN_5366}; // @[Filter.scala 164:35]
  wire [10:0] _GEN_7100 = _T_258 ? 11'h0 : _GEN_7099; // @[Filter.scala 162:80]
  wire [31:0] _T_346 = pixelIndex + 32'h3; // @[Filter.scala 158:31]
  wire [31:0] _GEN_3 = _T_346 % 32'h10; // @[Filter.scala 158:38]
  wire [4:0] _T_347 = _GEN_3[4:0]; // @[Filter.scala 158:38]
  wire [4:0] _T_349 = _T_347 + _GEN_18983; // @[Filter.scala 158:53]
  wire [4:0] _T_351 = _T_349 - 5'h1; // @[Filter.scala 158:69]
  wire [31:0] _T_354 = _T_346 / 32'h10; // @[Filter.scala 159:38]
  wire [31:0] _T_356 = _T_354 + _GEN_18984; // @[Filter.scala 159:53]
  wire [31:0] _T_358 = _T_356 - 32'h1; // @[Filter.scala 159:69]
  wire  _T_360 = _T_351 >= 5'h10; // @[Filter.scala 162:31]
  wire  _T_364 = _T_358 >= 32'hc; // @[Filter.scala 162:63]
  wire  _T_365 = _T_360 | _T_364; // @[Filter.scala 162:58]
  wire [36:0] _T_366 = _T_358 * 32'h10; // @[Filter.scala 165:66]
  wire [36:0] _GEN_19063 = {{32'd0}, _T_351}; // @[Filter.scala 165:81]
  wire [36:0] _T_368 = _T_366 + _GEN_19063; // @[Filter.scala 165:81]
  wire [3:0] _GEN_7109 = 8'h8 == _T_368[7:0] ? 4'h0 : 4'hf; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7110 = 8'h9 == _T_368[7:0] ? 4'h0 : _GEN_7109; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7111 = 8'ha == _T_368[7:0] ? 4'h0 : _GEN_7110; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7112 = 8'hb == _T_368[7:0] ? 4'h0 : _GEN_7111; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7113 = 8'hc == _T_368[7:0] ? 4'h0 : _GEN_7112; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7114 = 8'hd == _T_368[7:0] ? 4'h0 : _GEN_7113; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7115 = 8'he == _T_368[7:0] ? 4'h0 : _GEN_7114; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7116 = 8'hf == _T_368[7:0] ? 4'h0 : _GEN_7115; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7117 = 8'h10 == _T_368[7:0] ? 4'hf : _GEN_7116; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7118 = 8'h11 == _T_368[7:0] ? 4'hf : _GEN_7117; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7119 = 8'h12 == _T_368[7:0] ? 4'hf : _GEN_7118; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7120 = 8'h13 == _T_368[7:0] ? 4'hf : _GEN_7119; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7121 = 8'h14 == _T_368[7:0] ? 4'hf : _GEN_7120; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7122 = 8'h15 == _T_368[7:0] ? 4'hf : _GEN_7121; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7123 = 8'h16 == _T_368[7:0] ? 4'hf : _GEN_7122; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7124 = 8'h17 == _T_368[7:0] ? 4'hf : _GEN_7123; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7125 = 8'h18 == _T_368[7:0] ? 4'h0 : _GEN_7124; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7126 = 8'h19 == _T_368[7:0] ? 4'h0 : _GEN_7125; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7127 = 8'h1a == _T_368[7:0] ? 4'h0 : _GEN_7126; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7128 = 8'h1b == _T_368[7:0] ? 4'h0 : _GEN_7127; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7129 = 8'h1c == _T_368[7:0] ? 4'h0 : _GEN_7128; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7130 = 8'h1d == _T_368[7:0] ? 4'h0 : _GEN_7129; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7131 = 8'h1e == _T_368[7:0] ? 4'h0 : _GEN_7130; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7132 = 8'h1f == _T_368[7:0] ? 4'h0 : _GEN_7131; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7133 = 8'h20 == _T_368[7:0] ? 4'hf : _GEN_7132; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7134 = 8'h21 == _T_368[7:0] ? 4'hf : _GEN_7133; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7135 = 8'h22 == _T_368[7:0] ? 4'hf : _GEN_7134; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7136 = 8'h23 == _T_368[7:0] ? 4'hf : _GEN_7135; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7137 = 8'h24 == _T_368[7:0] ? 4'hf : _GEN_7136; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7138 = 8'h25 == _T_368[7:0] ? 4'hf : _GEN_7137; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7139 = 8'h26 == _T_368[7:0] ? 4'hf : _GEN_7138; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7140 = 8'h27 == _T_368[7:0] ? 4'hf : _GEN_7139; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7141 = 8'h28 == _T_368[7:0] ? 4'h0 : _GEN_7140; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7142 = 8'h29 == _T_368[7:0] ? 4'h0 : _GEN_7141; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7143 = 8'h2a == _T_368[7:0] ? 4'h0 : _GEN_7142; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7144 = 8'h2b == _T_368[7:0] ? 4'h0 : _GEN_7143; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7145 = 8'h2c == _T_368[7:0] ? 4'h0 : _GEN_7144; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7146 = 8'h2d == _T_368[7:0] ? 4'h0 : _GEN_7145; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7147 = 8'h2e == _T_368[7:0] ? 4'h0 : _GEN_7146; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7148 = 8'h2f == _T_368[7:0] ? 4'h0 : _GEN_7147; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7149 = 8'h30 == _T_368[7:0] ? 4'hf : _GEN_7148; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7150 = 8'h31 == _T_368[7:0] ? 4'hf : _GEN_7149; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7151 = 8'h32 == _T_368[7:0] ? 4'hf : _GEN_7150; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7152 = 8'h33 == _T_368[7:0] ? 4'hf : _GEN_7151; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7153 = 8'h34 == _T_368[7:0] ? 4'hf : _GEN_7152; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7154 = 8'h35 == _T_368[7:0] ? 4'hf : _GEN_7153; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7155 = 8'h36 == _T_368[7:0] ? 4'hf : _GEN_7154; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7156 = 8'h37 == _T_368[7:0] ? 4'hf : _GEN_7155; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7157 = 8'h38 == _T_368[7:0] ? 4'h0 : _GEN_7156; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7158 = 8'h39 == _T_368[7:0] ? 4'h0 : _GEN_7157; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7159 = 8'h3a == _T_368[7:0] ? 4'h0 : _GEN_7158; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7160 = 8'h3b == _T_368[7:0] ? 4'h0 : _GEN_7159; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7161 = 8'h3c == _T_368[7:0] ? 4'h0 : _GEN_7160; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7162 = 8'h3d == _T_368[7:0] ? 4'h0 : _GEN_7161; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7163 = 8'h3e == _T_368[7:0] ? 4'h0 : _GEN_7162; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7164 = 8'h3f == _T_368[7:0] ? 4'h0 : _GEN_7163; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7165 = 8'h40 == _T_368[7:0] ? 4'hf : _GEN_7164; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7166 = 8'h41 == _T_368[7:0] ? 4'hf : _GEN_7165; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7167 = 8'h42 == _T_368[7:0] ? 4'hf : _GEN_7166; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7168 = 8'h43 == _T_368[7:0] ? 4'hf : _GEN_7167; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7169 = 8'h44 == _T_368[7:0] ? 4'hf : _GEN_7168; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7170 = 8'h45 == _T_368[7:0] ? 4'hf : _GEN_7169; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7171 = 8'h46 == _T_368[7:0] ? 4'hf : _GEN_7170; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7172 = 8'h47 == _T_368[7:0] ? 4'hf : _GEN_7171; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7173 = 8'h48 == _T_368[7:0] ? 4'h0 : _GEN_7172; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7174 = 8'h49 == _T_368[7:0] ? 4'h0 : _GEN_7173; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7175 = 8'h4a == _T_368[7:0] ? 4'h0 : _GEN_7174; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7176 = 8'h4b == _T_368[7:0] ? 4'h0 : _GEN_7175; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7177 = 8'h4c == _T_368[7:0] ? 4'h0 : _GEN_7176; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7178 = 8'h4d == _T_368[7:0] ? 4'h0 : _GEN_7177; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7179 = 8'h4e == _T_368[7:0] ? 4'h0 : _GEN_7178; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7180 = 8'h4f == _T_368[7:0] ? 4'h0 : _GEN_7179; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7181 = 8'h50 == _T_368[7:0] ? 4'hf : _GEN_7180; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7182 = 8'h51 == _T_368[7:0] ? 4'hf : _GEN_7181; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7183 = 8'h52 == _T_368[7:0] ? 4'hf : _GEN_7182; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7184 = 8'h53 == _T_368[7:0] ? 4'hf : _GEN_7183; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7185 = 8'h54 == _T_368[7:0] ? 4'hf : _GEN_7184; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7186 = 8'h55 == _T_368[7:0] ? 4'hf : _GEN_7185; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7187 = 8'h56 == _T_368[7:0] ? 4'hf : _GEN_7186; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7188 = 8'h57 == _T_368[7:0] ? 4'hf : _GEN_7187; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7189 = 8'h58 == _T_368[7:0] ? 4'h0 : _GEN_7188; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7190 = 8'h59 == _T_368[7:0] ? 4'h0 : _GEN_7189; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7191 = 8'h5a == _T_368[7:0] ? 4'h0 : _GEN_7190; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7192 = 8'h5b == _T_368[7:0] ? 4'h0 : _GEN_7191; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7193 = 8'h5c == _T_368[7:0] ? 4'h0 : _GEN_7192; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7194 = 8'h5d == _T_368[7:0] ? 4'h0 : _GEN_7193; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7195 = 8'h5e == _T_368[7:0] ? 4'h0 : _GEN_7194; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7196 = 8'h5f == _T_368[7:0] ? 4'h0 : _GEN_7195; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7197 = 8'h60 == _T_368[7:0] ? 4'h0 : _GEN_7196; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7198 = 8'h61 == _T_368[7:0] ? 4'h0 : _GEN_7197; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7199 = 8'h62 == _T_368[7:0] ? 4'h0 : _GEN_7198; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7200 = 8'h63 == _T_368[7:0] ? 4'h0 : _GEN_7199; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7201 = 8'h64 == _T_368[7:0] ? 4'h0 : _GEN_7200; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7202 = 8'h65 == _T_368[7:0] ? 4'h0 : _GEN_7201; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7203 = 8'h66 == _T_368[7:0] ? 4'h0 : _GEN_7202; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7204 = 8'h67 == _T_368[7:0] ? 4'h0 : _GEN_7203; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7205 = 8'h68 == _T_368[7:0] ? 4'hf : _GEN_7204; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7206 = 8'h69 == _T_368[7:0] ? 4'hf : _GEN_7205; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7207 = 8'h6a == _T_368[7:0] ? 4'hf : _GEN_7206; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7208 = 8'h6b == _T_368[7:0] ? 4'hf : _GEN_7207; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7209 = 8'h6c == _T_368[7:0] ? 4'hf : _GEN_7208; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7210 = 8'h6d == _T_368[7:0] ? 4'hf : _GEN_7209; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7211 = 8'h6e == _T_368[7:0] ? 4'hf : _GEN_7210; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7212 = 8'h6f == _T_368[7:0] ? 4'hf : _GEN_7211; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7213 = 8'h70 == _T_368[7:0] ? 4'h0 : _GEN_7212; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7214 = 8'h71 == _T_368[7:0] ? 4'h0 : _GEN_7213; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7215 = 8'h72 == _T_368[7:0] ? 4'h0 : _GEN_7214; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7216 = 8'h73 == _T_368[7:0] ? 4'h0 : _GEN_7215; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7217 = 8'h74 == _T_368[7:0] ? 4'h0 : _GEN_7216; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7218 = 8'h75 == _T_368[7:0] ? 4'h0 : _GEN_7217; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7219 = 8'h76 == _T_368[7:0] ? 4'h0 : _GEN_7218; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7220 = 8'h77 == _T_368[7:0] ? 4'h0 : _GEN_7219; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7221 = 8'h78 == _T_368[7:0] ? 4'hf : _GEN_7220; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7222 = 8'h79 == _T_368[7:0] ? 4'hf : _GEN_7221; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7223 = 8'h7a == _T_368[7:0] ? 4'hf : _GEN_7222; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7224 = 8'h7b == _T_368[7:0] ? 4'hf : _GEN_7223; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7225 = 8'h7c == _T_368[7:0] ? 4'hf : _GEN_7224; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7226 = 8'h7d == _T_368[7:0] ? 4'hf : _GEN_7225; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7227 = 8'h7e == _T_368[7:0] ? 4'hf : _GEN_7226; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7228 = 8'h7f == _T_368[7:0] ? 4'hf : _GEN_7227; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7229 = 8'h80 == _T_368[7:0] ? 4'h0 : _GEN_7228; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7230 = 8'h81 == _T_368[7:0] ? 4'h0 : _GEN_7229; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7231 = 8'h82 == _T_368[7:0] ? 4'h0 : _GEN_7230; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7232 = 8'h83 == _T_368[7:0] ? 4'h0 : _GEN_7231; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7233 = 8'h84 == _T_368[7:0] ? 4'h0 : _GEN_7232; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7234 = 8'h85 == _T_368[7:0] ? 4'h0 : _GEN_7233; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7235 = 8'h86 == _T_368[7:0] ? 4'h0 : _GEN_7234; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7236 = 8'h87 == _T_368[7:0] ? 4'h0 : _GEN_7235; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7237 = 8'h88 == _T_368[7:0] ? 4'hf : _GEN_7236; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7238 = 8'h89 == _T_368[7:0] ? 4'hf : _GEN_7237; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7239 = 8'h8a == _T_368[7:0] ? 4'hf : _GEN_7238; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7240 = 8'h8b == _T_368[7:0] ? 4'hf : _GEN_7239; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7241 = 8'h8c == _T_368[7:0] ? 4'hf : _GEN_7240; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7242 = 8'h8d == _T_368[7:0] ? 4'hf : _GEN_7241; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7243 = 8'h8e == _T_368[7:0] ? 4'hf : _GEN_7242; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7244 = 8'h8f == _T_368[7:0] ? 4'hf : _GEN_7243; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7245 = 8'h90 == _T_368[7:0] ? 4'h0 : _GEN_7244; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7246 = 8'h91 == _T_368[7:0] ? 4'h0 : _GEN_7245; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7247 = 8'h92 == _T_368[7:0] ? 4'h0 : _GEN_7246; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7248 = 8'h93 == _T_368[7:0] ? 4'h0 : _GEN_7247; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7249 = 8'h94 == _T_368[7:0] ? 4'h0 : _GEN_7248; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7250 = 8'h95 == _T_368[7:0] ? 4'h0 : _GEN_7249; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7251 = 8'h96 == _T_368[7:0] ? 4'h0 : _GEN_7250; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7252 = 8'h97 == _T_368[7:0] ? 4'h0 : _GEN_7251; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7253 = 8'h98 == _T_368[7:0] ? 4'hf : _GEN_7252; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7254 = 8'h99 == _T_368[7:0] ? 4'hf : _GEN_7253; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7255 = 8'h9a == _T_368[7:0] ? 4'hf : _GEN_7254; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7256 = 8'h9b == _T_368[7:0] ? 4'hf : _GEN_7255; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7257 = 8'h9c == _T_368[7:0] ? 4'hf : _GEN_7256; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7258 = 8'h9d == _T_368[7:0] ? 4'hf : _GEN_7257; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7259 = 8'h9e == _T_368[7:0] ? 4'hf : _GEN_7258; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7260 = 8'h9f == _T_368[7:0] ? 4'hf : _GEN_7259; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7261 = 8'ha0 == _T_368[7:0] ? 4'h0 : _GEN_7260; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7262 = 8'ha1 == _T_368[7:0] ? 4'h0 : _GEN_7261; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7263 = 8'ha2 == _T_368[7:0] ? 4'h0 : _GEN_7262; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7264 = 8'ha3 == _T_368[7:0] ? 4'h0 : _GEN_7263; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7265 = 8'ha4 == _T_368[7:0] ? 4'h0 : _GEN_7264; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7266 = 8'ha5 == _T_368[7:0] ? 4'h0 : _GEN_7265; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7267 = 8'ha6 == _T_368[7:0] ? 4'h0 : _GEN_7266; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7268 = 8'ha7 == _T_368[7:0] ? 4'h0 : _GEN_7267; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7269 = 8'ha8 == _T_368[7:0] ? 4'hf : _GEN_7268; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7270 = 8'ha9 == _T_368[7:0] ? 4'hf : _GEN_7269; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7271 = 8'haa == _T_368[7:0] ? 4'hf : _GEN_7270; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7272 = 8'hab == _T_368[7:0] ? 4'hf : _GEN_7271; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7273 = 8'hac == _T_368[7:0] ? 4'hf : _GEN_7272; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7274 = 8'had == _T_368[7:0] ? 4'hf : _GEN_7273; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7275 = 8'hae == _T_368[7:0] ? 4'hf : _GEN_7274; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7276 = 8'haf == _T_368[7:0] ? 4'hf : _GEN_7275; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7277 = 8'hb0 == _T_368[7:0] ? 4'h0 : _GEN_7276; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7278 = 8'hb1 == _T_368[7:0] ? 4'h0 : _GEN_7277; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7279 = 8'hb2 == _T_368[7:0] ? 4'h0 : _GEN_7278; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7280 = 8'hb3 == _T_368[7:0] ? 4'h0 : _GEN_7279; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7281 = 8'hb4 == _T_368[7:0] ? 4'h0 : _GEN_7280; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7282 = 8'hb5 == _T_368[7:0] ? 4'h0 : _GEN_7281; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7283 = 8'hb6 == _T_368[7:0] ? 4'h0 : _GEN_7282; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7284 = 8'hb7 == _T_368[7:0] ? 4'h0 : _GEN_7283; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7285 = 8'hb8 == _T_368[7:0] ? 4'hf : _GEN_7284; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7286 = 8'hb9 == _T_368[7:0] ? 4'hf : _GEN_7285; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7287 = 8'hba == _T_368[7:0] ? 4'hf : _GEN_7286; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7288 = 8'hbb == _T_368[7:0] ? 4'hf : _GEN_7287; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7289 = 8'hbc == _T_368[7:0] ? 4'hf : _GEN_7288; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7290 = 8'hbd == _T_368[7:0] ? 4'hf : _GEN_7289; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7291 = 8'hbe == _T_368[7:0] ? 4'hf : _GEN_7290; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7292 = 8'hbf == _T_368[7:0] ? 4'hf : _GEN_7291; // @[Filter.scala 165:86]
  wire [4:0] _GEN_19064 = {{1'd0}, _GEN_7292}; // @[Filter.scala 165:86]
  wire [8:0] _T_370 = _GEN_19064 * 5'h14; // @[Filter.scala 165:86]
  wire [3:0] _GEN_7389 = 8'h60 == _T_368[7:0] ? 4'hf : 4'h0; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7390 = 8'h61 == _T_368[7:0] ? 4'hf : _GEN_7389; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7391 = 8'h62 == _T_368[7:0] ? 4'hf : _GEN_7390; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7392 = 8'h63 == _T_368[7:0] ? 4'hf : _GEN_7391; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7393 = 8'h64 == _T_368[7:0] ? 4'hf : _GEN_7392; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7394 = 8'h65 == _T_368[7:0] ? 4'hf : _GEN_7393; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7395 = 8'h66 == _T_368[7:0] ? 4'hf : _GEN_7394; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7396 = 8'h67 == _T_368[7:0] ? 4'hf : _GEN_7395; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7397 = 8'h68 == _T_368[7:0] ? 4'hf : _GEN_7396; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7398 = 8'h69 == _T_368[7:0] ? 4'hf : _GEN_7397; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7399 = 8'h6a == _T_368[7:0] ? 4'hf : _GEN_7398; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7400 = 8'h6b == _T_368[7:0] ? 4'hf : _GEN_7399; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7401 = 8'h6c == _T_368[7:0] ? 4'hf : _GEN_7400; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7402 = 8'h6d == _T_368[7:0] ? 4'hf : _GEN_7401; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7403 = 8'h6e == _T_368[7:0] ? 4'hf : _GEN_7402; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7404 = 8'h6f == _T_368[7:0] ? 4'hf : _GEN_7403; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7405 = 8'h70 == _T_368[7:0] ? 4'hf : _GEN_7404; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7406 = 8'h71 == _T_368[7:0] ? 4'hf : _GEN_7405; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7407 = 8'h72 == _T_368[7:0] ? 4'hf : _GEN_7406; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7408 = 8'h73 == _T_368[7:0] ? 4'hf : _GEN_7407; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7409 = 8'h74 == _T_368[7:0] ? 4'hf : _GEN_7408; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7410 = 8'h75 == _T_368[7:0] ? 4'hf : _GEN_7409; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7411 = 8'h76 == _T_368[7:0] ? 4'hf : _GEN_7410; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7412 = 8'h77 == _T_368[7:0] ? 4'hf : _GEN_7411; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7413 = 8'h78 == _T_368[7:0] ? 4'hf : _GEN_7412; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7414 = 8'h79 == _T_368[7:0] ? 4'hf : _GEN_7413; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7415 = 8'h7a == _T_368[7:0] ? 4'hf : _GEN_7414; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7416 = 8'h7b == _T_368[7:0] ? 4'hf : _GEN_7415; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7417 = 8'h7c == _T_368[7:0] ? 4'hf : _GEN_7416; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7418 = 8'h7d == _T_368[7:0] ? 4'hf : _GEN_7417; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7419 = 8'h7e == _T_368[7:0] ? 4'hf : _GEN_7418; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7420 = 8'h7f == _T_368[7:0] ? 4'hf : _GEN_7419; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7421 = 8'h80 == _T_368[7:0] ? 4'hf : _GEN_7420; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7422 = 8'h81 == _T_368[7:0] ? 4'hf : _GEN_7421; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7423 = 8'h82 == _T_368[7:0] ? 4'hf : _GEN_7422; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7424 = 8'h83 == _T_368[7:0] ? 4'hf : _GEN_7423; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7425 = 8'h84 == _T_368[7:0] ? 4'hf : _GEN_7424; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7426 = 8'h85 == _T_368[7:0] ? 4'hf : _GEN_7425; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7427 = 8'h86 == _T_368[7:0] ? 4'hf : _GEN_7426; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7428 = 8'h87 == _T_368[7:0] ? 4'hf : _GEN_7427; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7429 = 8'h88 == _T_368[7:0] ? 4'hf : _GEN_7428; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7430 = 8'h89 == _T_368[7:0] ? 4'hf : _GEN_7429; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7431 = 8'h8a == _T_368[7:0] ? 4'hf : _GEN_7430; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7432 = 8'h8b == _T_368[7:0] ? 4'hf : _GEN_7431; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7433 = 8'h8c == _T_368[7:0] ? 4'hf : _GEN_7432; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7434 = 8'h8d == _T_368[7:0] ? 4'hf : _GEN_7433; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7435 = 8'h8e == _T_368[7:0] ? 4'hf : _GEN_7434; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7436 = 8'h8f == _T_368[7:0] ? 4'hf : _GEN_7435; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7437 = 8'h90 == _T_368[7:0] ? 4'hf : _GEN_7436; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7438 = 8'h91 == _T_368[7:0] ? 4'hf : _GEN_7437; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7439 = 8'h92 == _T_368[7:0] ? 4'hf : _GEN_7438; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7440 = 8'h93 == _T_368[7:0] ? 4'hf : _GEN_7439; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7441 = 8'h94 == _T_368[7:0] ? 4'hf : _GEN_7440; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7442 = 8'h95 == _T_368[7:0] ? 4'hf : _GEN_7441; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7443 = 8'h96 == _T_368[7:0] ? 4'hf : _GEN_7442; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7444 = 8'h97 == _T_368[7:0] ? 4'hf : _GEN_7443; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7445 = 8'h98 == _T_368[7:0] ? 4'hf : _GEN_7444; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7446 = 8'h99 == _T_368[7:0] ? 4'hf : _GEN_7445; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7447 = 8'h9a == _T_368[7:0] ? 4'hf : _GEN_7446; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7448 = 8'h9b == _T_368[7:0] ? 4'hf : _GEN_7447; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7449 = 8'h9c == _T_368[7:0] ? 4'hf : _GEN_7448; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7450 = 8'h9d == _T_368[7:0] ? 4'hf : _GEN_7449; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7451 = 8'h9e == _T_368[7:0] ? 4'hf : _GEN_7450; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7452 = 8'h9f == _T_368[7:0] ? 4'hf : _GEN_7451; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7453 = 8'ha0 == _T_368[7:0] ? 4'hf : _GEN_7452; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7454 = 8'ha1 == _T_368[7:0] ? 4'hf : _GEN_7453; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7455 = 8'ha2 == _T_368[7:0] ? 4'hf : _GEN_7454; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7456 = 8'ha3 == _T_368[7:0] ? 4'hf : _GEN_7455; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7457 = 8'ha4 == _T_368[7:0] ? 4'hf : _GEN_7456; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7458 = 8'ha5 == _T_368[7:0] ? 4'hf : _GEN_7457; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7459 = 8'ha6 == _T_368[7:0] ? 4'hf : _GEN_7458; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7460 = 8'ha7 == _T_368[7:0] ? 4'hf : _GEN_7459; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7461 = 8'ha8 == _T_368[7:0] ? 4'hf : _GEN_7460; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7462 = 8'ha9 == _T_368[7:0] ? 4'hf : _GEN_7461; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7463 = 8'haa == _T_368[7:0] ? 4'hf : _GEN_7462; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7464 = 8'hab == _T_368[7:0] ? 4'hf : _GEN_7463; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7465 = 8'hac == _T_368[7:0] ? 4'hf : _GEN_7464; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7466 = 8'had == _T_368[7:0] ? 4'hf : _GEN_7465; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7467 = 8'hae == _T_368[7:0] ? 4'hf : _GEN_7466; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7468 = 8'haf == _T_368[7:0] ? 4'hf : _GEN_7467; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7469 = 8'hb0 == _T_368[7:0] ? 4'hf : _GEN_7468; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7470 = 8'hb1 == _T_368[7:0] ? 4'hf : _GEN_7469; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7471 = 8'hb2 == _T_368[7:0] ? 4'hf : _GEN_7470; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7472 = 8'hb3 == _T_368[7:0] ? 4'hf : _GEN_7471; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7473 = 8'hb4 == _T_368[7:0] ? 4'hf : _GEN_7472; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7474 = 8'hb5 == _T_368[7:0] ? 4'hf : _GEN_7473; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7475 = 8'hb6 == _T_368[7:0] ? 4'hf : _GEN_7474; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7476 = 8'hb7 == _T_368[7:0] ? 4'hf : _GEN_7475; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7477 = 8'hb8 == _T_368[7:0] ? 4'hf : _GEN_7476; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7478 = 8'hb9 == _T_368[7:0] ? 4'hf : _GEN_7477; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7479 = 8'hba == _T_368[7:0] ? 4'hf : _GEN_7478; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7480 = 8'hbb == _T_368[7:0] ? 4'hf : _GEN_7479; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7481 = 8'hbc == _T_368[7:0] ? 4'hf : _GEN_7480; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7482 = 8'hbd == _T_368[7:0] ? 4'hf : _GEN_7481; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7483 = 8'hbe == _T_368[7:0] ? 4'hf : _GEN_7482; // @[Filter.scala 165:126]
  wire [3:0] _GEN_7484 = 8'hbf == _T_368[7:0] ? 4'hf : _GEN_7483; // @[Filter.scala 165:126]
  wire [6:0] _GEN_19066 = {{3'd0}, _GEN_7484}; // @[Filter.scala 165:126]
  wire [10:0] _T_375 = _GEN_19066 * 7'h46; // @[Filter.scala 165:126]
  wire [10:0] _GEN_19067 = {{2'd0}, _T_370}; // @[Filter.scala 165:93]
  wire [10:0] _T_377 = _GEN_19067 + _T_375; // @[Filter.scala 165:93]
  wire [3:0] _GEN_7493 = 8'h8 == _T_368[7:0] ? 4'hf : 4'h0; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7494 = 8'h9 == _T_368[7:0] ? 4'hf : _GEN_7493; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7495 = 8'ha == _T_368[7:0] ? 4'hf : _GEN_7494; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7496 = 8'hb == _T_368[7:0] ? 4'hf : _GEN_7495; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7497 = 8'hc == _T_368[7:0] ? 4'hf : _GEN_7496; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7498 = 8'hd == _T_368[7:0] ? 4'hf : _GEN_7497; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7499 = 8'he == _T_368[7:0] ? 4'hf : _GEN_7498; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7500 = 8'hf == _T_368[7:0] ? 4'hf : _GEN_7499; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7501 = 8'h10 == _T_368[7:0] ? 4'h0 : _GEN_7500; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7502 = 8'h11 == _T_368[7:0] ? 4'h0 : _GEN_7501; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7503 = 8'h12 == _T_368[7:0] ? 4'h0 : _GEN_7502; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7504 = 8'h13 == _T_368[7:0] ? 4'h0 : _GEN_7503; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7505 = 8'h14 == _T_368[7:0] ? 4'h0 : _GEN_7504; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7506 = 8'h15 == _T_368[7:0] ? 4'h0 : _GEN_7505; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7507 = 8'h16 == _T_368[7:0] ? 4'h0 : _GEN_7506; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7508 = 8'h17 == _T_368[7:0] ? 4'h0 : _GEN_7507; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7509 = 8'h18 == _T_368[7:0] ? 4'hf : _GEN_7508; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7510 = 8'h19 == _T_368[7:0] ? 4'hf : _GEN_7509; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7511 = 8'h1a == _T_368[7:0] ? 4'hf : _GEN_7510; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7512 = 8'h1b == _T_368[7:0] ? 4'hf : _GEN_7511; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7513 = 8'h1c == _T_368[7:0] ? 4'hf : _GEN_7512; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7514 = 8'h1d == _T_368[7:0] ? 4'hf : _GEN_7513; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7515 = 8'h1e == _T_368[7:0] ? 4'hf : _GEN_7514; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7516 = 8'h1f == _T_368[7:0] ? 4'hf : _GEN_7515; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7517 = 8'h20 == _T_368[7:0] ? 4'h0 : _GEN_7516; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7518 = 8'h21 == _T_368[7:0] ? 4'h0 : _GEN_7517; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7519 = 8'h22 == _T_368[7:0] ? 4'h0 : _GEN_7518; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7520 = 8'h23 == _T_368[7:0] ? 4'h0 : _GEN_7519; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7521 = 8'h24 == _T_368[7:0] ? 4'h0 : _GEN_7520; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7522 = 8'h25 == _T_368[7:0] ? 4'h0 : _GEN_7521; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7523 = 8'h26 == _T_368[7:0] ? 4'h0 : _GEN_7522; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7524 = 8'h27 == _T_368[7:0] ? 4'h0 : _GEN_7523; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7525 = 8'h28 == _T_368[7:0] ? 4'hf : _GEN_7524; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7526 = 8'h29 == _T_368[7:0] ? 4'hf : _GEN_7525; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7527 = 8'h2a == _T_368[7:0] ? 4'hf : _GEN_7526; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7528 = 8'h2b == _T_368[7:0] ? 4'hf : _GEN_7527; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7529 = 8'h2c == _T_368[7:0] ? 4'hf : _GEN_7528; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7530 = 8'h2d == _T_368[7:0] ? 4'hf : _GEN_7529; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7531 = 8'h2e == _T_368[7:0] ? 4'hf : _GEN_7530; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7532 = 8'h2f == _T_368[7:0] ? 4'hf : _GEN_7531; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7533 = 8'h30 == _T_368[7:0] ? 4'h0 : _GEN_7532; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7534 = 8'h31 == _T_368[7:0] ? 4'h0 : _GEN_7533; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7535 = 8'h32 == _T_368[7:0] ? 4'h0 : _GEN_7534; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7536 = 8'h33 == _T_368[7:0] ? 4'h0 : _GEN_7535; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7537 = 8'h34 == _T_368[7:0] ? 4'h0 : _GEN_7536; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7538 = 8'h35 == _T_368[7:0] ? 4'h0 : _GEN_7537; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7539 = 8'h36 == _T_368[7:0] ? 4'h0 : _GEN_7538; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7540 = 8'h37 == _T_368[7:0] ? 4'h0 : _GEN_7539; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7541 = 8'h38 == _T_368[7:0] ? 4'hf : _GEN_7540; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7542 = 8'h39 == _T_368[7:0] ? 4'hf : _GEN_7541; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7543 = 8'h3a == _T_368[7:0] ? 4'hf : _GEN_7542; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7544 = 8'h3b == _T_368[7:0] ? 4'hf : _GEN_7543; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7545 = 8'h3c == _T_368[7:0] ? 4'hf : _GEN_7544; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7546 = 8'h3d == _T_368[7:0] ? 4'hf : _GEN_7545; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7547 = 8'h3e == _T_368[7:0] ? 4'hf : _GEN_7546; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7548 = 8'h3f == _T_368[7:0] ? 4'hf : _GEN_7547; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7549 = 8'h40 == _T_368[7:0] ? 4'h0 : _GEN_7548; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7550 = 8'h41 == _T_368[7:0] ? 4'h0 : _GEN_7549; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7551 = 8'h42 == _T_368[7:0] ? 4'h0 : _GEN_7550; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7552 = 8'h43 == _T_368[7:0] ? 4'h0 : _GEN_7551; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7553 = 8'h44 == _T_368[7:0] ? 4'h0 : _GEN_7552; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7554 = 8'h45 == _T_368[7:0] ? 4'h0 : _GEN_7553; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7555 = 8'h46 == _T_368[7:0] ? 4'h0 : _GEN_7554; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7556 = 8'h47 == _T_368[7:0] ? 4'h0 : _GEN_7555; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7557 = 8'h48 == _T_368[7:0] ? 4'hf : _GEN_7556; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7558 = 8'h49 == _T_368[7:0] ? 4'hf : _GEN_7557; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7559 = 8'h4a == _T_368[7:0] ? 4'hf : _GEN_7558; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7560 = 8'h4b == _T_368[7:0] ? 4'hf : _GEN_7559; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7561 = 8'h4c == _T_368[7:0] ? 4'hf : _GEN_7560; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7562 = 8'h4d == _T_368[7:0] ? 4'hf : _GEN_7561; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7563 = 8'h4e == _T_368[7:0] ? 4'hf : _GEN_7562; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7564 = 8'h4f == _T_368[7:0] ? 4'hf : _GEN_7563; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7565 = 8'h50 == _T_368[7:0] ? 4'h0 : _GEN_7564; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7566 = 8'h51 == _T_368[7:0] ? 4'h0 : _GEN_7565; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7567 = 8'h52 == _T_368[7:0] ? 4'h0 : _GEN_7566; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7568 = 8'h53 == _T_368[7:0] ? 4'h0 : _GEN_7567; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7569 = 8'h54 == _T_368[7:0] ? 4'h0 : _GEN_7568; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7570 = 8'h55 == _T_368[7:0] ? 4'h0 : _GEN_7569; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7571 = 8'h56 == _T_368[7:0] ? 4'h0 : _GEN_7570; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7572 = 8'h57 == _T_368[7:0] ? 4'h0 : _GEN_7571; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7573 = 8'h58 == _T_368[7:0] ? 4'hf : _GEN_7572; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7574 = 8'h59 == _T_368[7:0] ? 4'hf : _GEN_7573; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7575 = 8'h5a == _T_368[7:0] ? 4'hf : _GEN_7574; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7576 = 8'h5b == _T_368[7:0] ? 4'hf : _GEN_7575; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7577 = 8'h5c == _T_368[7:0] ? 4'hf : _GEN_7576; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7578 = 8'h5d == _T_368[7:0] ? 4'hf : _GEN_7577; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7579 = 8'h5e == _T_368[7:0] ? 4'hf : _GEN_7578; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7580 = 8'h5f == _T_368[7:0] ? 4'hf : _GEN_7579; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7581 = 8'h60 == _T_368[7:0] ? 4'h0 : _GEN_7580; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7582 = 8'h61 == _T_368[7:0] ? 4'h0 : _GEN_7581; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7583 = 8'h62 == _T_368[7:0] ? 4'h0 : _GEN_7582; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7584 = 8'h63 == _T_368[7:0] ? 4'h0 : _GEN_7583; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7585 = 8'h64 == _T_368[7:0] ? 4'h0 : _GEN_7584; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7586 = 8'h65 == _T_368[7:0] ? 4'h0 : _GEN_7585; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7587 = 8'h66 == _T_368[7:0] ? 4'h0 : _GEN_7586; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7588 = 8'h67 == _T_368[7:0] ? 4'h0 : _GEN_7587; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7589 = 8'h68 == _T_368[7:0] ? 4'hf : _GEN_7588; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7590 = 8'h69 == _T_368[7:0] ? 4'hf : _GEN_7589; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7591 = 8'h6a == _T_368[7:0] ? 4'hf : _GEN_7590; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7592 = 8'h6b == _T_368[7:0] ? 4'hf : _GEN_7591; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7593 = 8'h6c == _T_368[7:0] ? 4'hf : _GEN_7592; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7594 = 8'h6d == _T_368[7:0] ? 4'hf : _GEN_7593; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7595 = 8'h6e == _T_368[7:0] ? 4'hf : _GEN_7594; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7596 = 8'h6f == _T_368[7:0] ? 4'hf : _GEN_7595; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7597 = 8'h70 == _T_368[7:0] ? 4'h0 : _GEN_7596; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7598 = 8'h71 == _T_368[7:0] ? 4'h0 : _GEN_7597; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7599 = 8'h72 == _T_368[7:0] ? 4'h0 : _GEN_7598; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7600 = 8'h73 == _T_368[7:0] ? 4'h0 : _GEN_7599; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7601 = 8'h74 == _T_368[7:0] ? 4'h0 : _GEN_7600; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7602 = 8'h75 == _T_368[7:0] ? 4'h0 : _GEN_7601; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7603 = 8'h76 == _T_368[7:0] ? 4'h0 : _GEN_7602; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7604 = 8'h77 == _T_368[7:0] ? 4'h0 : _GEN_7603; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7605 = 8'h78 == _T_368[7:0] ? 4'hf : _GEN_7604; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7606 = 8'h79 == _T_368[7:0] ? 4'hf : _GEN_7605; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7607 = 8'h7a == _T_368[7:0] ? 4'hf : _GEN_7606; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7608 = 8'h7b == _T_368[7:0] ? 4'hf : _GEN_7607; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7609 = 8'h7c == _T_368[7:0] ? 4'hf : _GEN_7608; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7610 = 8'h7d == _T_368[7:0] ? 4'hf : _GEN_7609; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7611 = 8'h7e == _T_368[7:0] ? 4'hf : _GEN_7610; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7612 = 8'h7f == _T_368[7:0] ? 4'hf : _GEN_7611; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7613 = 8'h80 == _T_368[7:0] ? 4'h0 : _GEN_7612; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7614 = 8'h81 == _T_368[7:0] ? 4'h0 : _GEN_7613; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7615 = 8'h82 == _T_368[7:0] ? 4'h0 : _GEN_7614; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7616 = 8'h83 == _T_368[7:0] ? 4'h0 : _GEN_7615; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7617 = 8'h84 == _T_368[7:0] ? 4'h0 : _GEN_7616; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7618 = 8'h85 == _T_368[7:0] ? 4'h0 : _GEN_7617; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7619 = 8'h86 == _T_368[7:0] ? 4'h0 : _GEN_7618; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7620 = 8'h87 == _T_368[7:0] ? 4'h0 : _GEN_7619; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7621 = 8'h88 == _T_368[7:0] ? 4'hf : _GEN_7620; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7622 = 8'h89 == _T_368[7:0] ? 4'hf : _GEN_7621; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7623 = 8'h8a == _T_368[7:0] ? 4'hf : _GEN_7622; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7624 = 8'h8b == _T_368[7:0] ? 4'hf : _GEN_7623; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7625 = 8'h8c == _T_368[7:0] ? 4'hf : _GEN_7624; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7626 = 8'h8d == _T_368[7:0] ? 4'hf : _GEN_7625; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7627 = 8'h8e == _T_368[7:0] ? 4'hf : _GEN_7626; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7628 = 8'h8f == _T_368[7:0] ? 4'hf : _GEN_7627; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7629 = 8'h90 == _T_368[7:0] ? 4'h0 : _GEN_7628; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7630 = 8'h91 == _T_368[7:0] ? 4'h0 : _GEN_7629; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7631 = 8'h92 == _T_368[7:0] ? 4'h0 : _GEN_7630; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7632 = 8'h93 == _T_368[7:0] ? 4'h0 : _GEN_7631; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7633 = 8'h94 == _T_368[7:0] ? 4'h0 : _GEN_7632; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7634 = 8'h95 == _T_368[7:0] ? 4'h0 : _GEN_7633; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7635 = 8'h96 == _T_368[7:0] ? 4'h0 : _GEN_7634; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7636 = 8'h97 == _T_368[7:0] ? 4'h0 : _GEN_7635; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7637 = 8'h98 == _T_368[7:0] ? 4'hf : _GEN_7636; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7638 = 8'h99 == _T_368[7:0] ? 4'hf : _GEN_7637; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7639 = 8'h9a == _T_368[7:0] ? 4'hf : _GEN_7638; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7640 = 8'h9b == _T_368[7:0] ? 4'hf : _GEN_7639; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7641 = 8'h9c == _T_368[7:0] ? 4'hf : _GEN_7640; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7642 = 8'h9d == _T_368[7:0] ? 4'hf : _GEN_7641; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7643 = 8'h9e == _T_368[7:0] ? 4'hf : _GEN_7642; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7644 = 8'h9f == _T_368[7:0] ? 4'hf : _GEN_7643; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7645 = 8'ha0 == _T_368[7:0] ? 4'h0 : _GEN_7644; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7646 = 8'ha1 == _T_368[7:0] ? 4'h0 : _GEN_7645; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7647 = 8'ha2 == _T_368[7:0] ? 4'h0 : _GEN_7646; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7648 = 8'ha3 == _T_368[7:0] ? 4'h0 : _GEN_7647; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7649 = 8'ha4 == _T_368[7:0] ? 4'h0 : _GEN_7648; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7650 = 8'ha5 == _T_368[7:0] ? 4'h0 : _GEN_7649; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7651 = 8'ha6 == _T_368[7:0] ? 4'h0 : _GEN_7650; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7652 = 8'ha7 == _T_368[7:0] ? 4'h0 : _GEN_7651; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7653 = 8'ha8 == _T_368[7:0] ? 4'hf : _GEN_7652; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7654 = 8'ha9 == _T_368[7:0] ? 4'hf : _GEN_7653; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7655 = 8'haa == _T_368[7:0] ? 4'hf : _GEN_7654; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7656 = 8'hab == _T_368[7:0] ? 4'hf : _GEN_7655; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7657 = 8'hac == _T_368[7:0] ? 4'hf : _GEN_7656; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7658 = 8'had == _T_368[7:0] ? 4'hf : _GEN_7657; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7659 = 8'hae == _T_368[7:0] ? 4'hf : _GEN_7658; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7660 = 8'haf == _T_368[7:0] ? 4'hf : _GEN_7659; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7661 = 8'hb0 == _T_368[7:0] ? 4'h0 : _GEN_7660; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7662 = 8'hb1 == _T_368[7:0] ? 4'h0 : _GEN_7661; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7663 = 8'hb2 == _T_368[7:0] ? 4'h0 : _GEN_7662; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7664 = 8'hb3 == _T_368[7:0] ? 4'h0 : _GEN_7663; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7665 = 8'hb4 == _T_368[7:0] ? 4'h0 : _GEN_7664; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7666 = 8'hb5 == _T_368[7:0] ? 4'h0 : _GEN_7665; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7667 = 8'hb6 == _T_368[7:0] ? 4'h0 : _GEN_7666; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7668 = 8'hb7 == _T_368[7:0] ? 4'h0 : _GEN_7667; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7669 = 8'hb8 == _T_368[7:0] ? 4'hf : _GEN_7668; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7670 = 8'hb9 == _T_368[7:0] ? 4'hf : _GEN_7669; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7671 = 8'hba == _T_368[7:0] ? 4'hf : _GEN_7670; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7672 = 8'hbb == _T_368[7:0] ? 4'hf : _GEN_7671; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7673 = 8'hbc == _T_368[7:0] ? 4'hf : _GEN_7672; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7674 = 8'hbd == _T_368[7:0] ? 4'hf : _GEN_7673; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7675 = 8'hbe == _T_368[7:0] ? 4'hf : _GEN_7674; // @[Filter.scala 165:166]
  wire [3:0] _GEN_7676 = 8'hbf == _T_368[7:0] ? 4'hf : _GEN_7675; // @[Filter.scala 165:166]
  wire [7:0] _T_382 = _GEN_7676 * 4'ha; // @[Filter.scala 165:166]
  wire [10:0] _GEN_19069 = {{3'd0}, _T_382}; // @[Filter.scala 165:133]
  wire [10:0] _T_384 = _T_377 + _GEN_19069; // @[Filter.scala 165:133]
  wire [10:0] _T_385 = _T_384 / 11'h64; // @[Filter.scala 165:174]
  wire [10:0] _GEN_7869 = io_SPI_distort ? _T_385 : {{7'd0}, _GEN_7292}; // @[Filter.scala 164:35]
  wire [10:0] _GEN_7870 = _T_365 ? 11'h0 : _GEN_7869; // @[Filter.scala 162:80]
  wire [10:0] _GEN_8639 = io_SPI_distort ? _T_385 : {{7'd0}, _GEN_7484}; // @[Filter.scala 164:35]
  wire [10:0] _GEN_8640 = _T_365 ? 11'h0 : _GEN_8639; // @[Filter.scala 162:80]
  wire [10:0] _GEN_9409 = io_SPI_distort ? _T_385 : {{7'd0}, _GEN_7676}; // @[Filter.scala 164:35]
  wire [10:0] _GEN_9410 = _T_365 ? 11'h0 : _GEN_9409; // @[Filter.scala 162:80]
  wire [31:0] _T_453 = pixelIndex + 32'h4; // @[Filter.scala 158:31]
  wire [31:0] _GEN_4 = _T_453 % 32'h10; // @[Filter.scala 158:38]
  wire [4:0] _T_454 = _GEN_4[4:0]; // @[Filter.scala 158:38]
  wire [4:0] _T_456 = _T_454 + _GEN_18983; // @[Filter.scala 158:53]
  wire [4:0] _T_458 = _T_456 - 5'h1; // @[Filter.scala 158:69]
  wire [31:0] _T_461 = _T_453 / 32'h10; // @[Filter.scala 159:38]
  wire [31:0] _T_463 = _T_461 + _GEN_18984; // @[Filter.scala 159:53]
  wire [31:0] _T_465 = _T_463 - 32'h1; // @[Filter.scala 159:69]
  wire  _T_467 = _T_458 >= 5'h10; // @[Filter.scala 162:31]
  wire  _T_471 = _T_465 >= 32'hc; // @[Filter.scala 162:63]
  wire  _T_472 = _T_467 | _T_471; // @[Filter.scala 162:58]
  wire [36:0] _T_473 = _T_465 * 32'h10; // @[Filter.scala 165:66]
  wire [36:0] _GEN_19089 = {{32'd0}, _T_458}; // @[Filter.scala 165:81]
  wire [36:0] _T_475 = _T_473 + _GEN_19089; // @[Filter.scala 165:81]
  wire [3:0] _GEN_9419 = 8'h8 == _T_475[7:0] ? 4'h0 : 4'hf; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9420 = 8'h9 == _T_475[7:0] ? 4'h0 : _GEN_9419; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9421 = 8'ha == _T_475[7:0] ? 4'h0 : _GEN_9420; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9422 = 8'hb == _T_475[7:0] ? 4'h0 : _GEN_9421; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9423 = 8'hc == _T_475[7:0] ? 4'h0 : _GEN_9422; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9424 = 8'hd == _T_475[7:0] ? 4'h0 : _GEN_9423; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9425 = 8'he == _T_475[7:0] ? 4'h0 : _GEN_9424; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9426 = 8'hf == _T_475[7:0] ? 4'h0 : _GEN_9425; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9427 = 8'h10 == _T_475[7:0] ? 4'hf : _GEN_9426; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9428 = 8'h11 == _T_475[7:0] ? 4'hf : _GEN_9427; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9429 = 8'h12 == _T_475[7:0] ? 4'hf : _GEN_9428; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9430 = 8'h13 == _T_475[7:0] ? 4'hf : _GEN_9429; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9431 = 8'h14 == _T_475[7:0] ? 4'hf : _GEN_9430; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9432 = 8'h15 == _T_475[7:0] ? 4'hf : _GEN_9431; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9433 = 8'h16 == _T_475[7:0] ? 4'hf : _GEN_9432; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9434 = 8'h17 == _T_475[7:0] ? 4'hf : _GEN_9433; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9435 = 8'h18 == _T_475[7:0] ? 4'h0 : _GEN_9434; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9436 = 8'h19 == _T_475[7:0] ? 4'h0 : _GEN_9435; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9437 = 8'h1a == _T_475[7:0] ? 4'h0 : _GEN_9436; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9438 = 8'h1b == _T_475[7:0] ? 4'h0 : _GEN_9437; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9439 = 8'h1c == _T_475[7:0] ? 4'h0 : _GEN_9438; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9440 = 8'h1d == _T_475[7:0] ? 4'h0 : _GEN_9439; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9441 = 8'h1e == _T_475[7:0] ? 4'h0 : _GEN_9440; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9442 = 8'h1f == _T_475[7:0] ? 4'h0 : _GEN_9441; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9443 = 8'h20 == _T_475[7:0] ? 4'hf : _GEN_9442; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9444 = 8'h21 == _T_475[7:0] ? 4'hf : _GEN_9443; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9445 = 8'h22 == _T_475[7:0] ? 4'hf : _GEN_9444; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9446 = 8'h23 == _T_475[7:0] ? 4'hf : _GEN_9445; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9447 = 8'h24 == _T_475[7:0] ? 4'hf : _GEN_9446; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9448 = 8'h25 == _T_475[7:0] ? 4'hf : _GEN_9447; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9449 = 8'h26 == _T_475[7:0] ? 4'hf : _GEN_9448; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9450 = 8'h27 == _T_475[7:0] ? 4'hf : _GEN_9449; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9451 = 8'h28 == _T_475[7:0] ? 4'h0 : _GEN_9450; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9452 = 8'h29 == _T_475[7:0] ? 4'h0 : _GEN_9451; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9453 = 8'h2a == _T_475[7:0] ? 4'h0 : _GEN_9452; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9454 = 8'h2b == _T_475[7:0] ? 4'h0 : _GEN_9453; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9455 = 8'h2c == _T_475[7:0] ? 4'h0 : _GEN_9454; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9456 = 8'h2d == _T_475[7:0] ? 4'h0 : _GEN_9455; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9457 = 8'h2e == _T_475[7:0] ? 4'h0 : _GEN_9456; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9458 = 8'h2f == _T_475[7:0] ? 4'h0 : _GEN_9457; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9459 = 8'h30 == _T_475[7:0] ? 4'hf : _GEN_9458; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9460 = 8'h31 == _T_475[7:0] ? 4'hf : _GEN_9459; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9461 = 8'h32 == _T_475[7:0] ? 4'hf : _GEN_9460; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9462 = 8'h33 == _T_475[7:0] ? 4'hf : _GEN_9461; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9463 = 8'h34 == _T_475[7:0] ? 4'hf : _GEN_9462; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9464 = 8'h35 == _T_475[7:0] ? 4'hf : _GEN_9463; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9465 = 8'h36 == _T_475[7:0] ? 4'hf : _GEN_9464; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9466 = 8'h37 == _T_475[7:0] ? 4'hf : _GEN_9465; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9467 = 8'h38 == _T_475[7:0] ? 4'h0 : _GEN_9466; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9468 = 8'h39 == _T_475[7:0] ? 4'h0 : _GEN_9467; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9469 = 8'h3a == _T_475[7:0] ? 4'h0 : _GEN_9468; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9470 = 8'h3b == _T_475[7:0] ? 4'h0 : _GEN_9469; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9471 = 8'h3c == _T_475[7:0] ? 4'h0 : _GEN_9470; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9472 = 8'h3d == _T_475[7:0] ? 4'h0 : _GEN_9471; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9473 = 8'h3e == _T_475[7:0] ? 4'h0 : _GEN_9472; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9474 = 8'h3f == _T_475[7:0] ? 4'h0 : _GEN_9473; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9475 = 8'h40 == _T_475[7:0] ? 4'hf : _GEN_9474; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9476 = 8'h41 == _T_475[7:0] ? 4'hf : _GEN_9475; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9477 = 8'h42 == _T_475[7:0] ? 4'hf : _GEN_9476; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9478 = 8'h43 == _T_475[7:0] ? 4'hf : _GEN_9477; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9479 = 8'h44 == _T_475[7:0] ? 4'hf : _GEN_9478; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9480 = 8'h45 == _T_475[7:0] ? 4'hf : _GEN_9479; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9481 = 8'h46 == _T_475[7:0] ? 4'hf : _GEN_9480; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9482 = 8'h47 == _T_475[7:0] ? 4'hf : _GEN_9481; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9483 = 8'h48 == _T_475[7:0] ? 4'h0 : _GEN_9482; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9484 = 8'h49 == _T_475[7:0] ? 4'h0 : _GEN_9483; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9485 = 8'h4a == _T_475[7:0] ? 4'h0 : _GEN_9484; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9486 = 8'h4b == _T_475[7:0] ? 4'h0 : _GEN_9485; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9487 = 8'h4c == _T_475[7:0] ? 4'h0 : _GEN_9486; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9488 = 8'h4d == _T_475[7:0] ? 4'h0 : _GEN_9487; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9489 = 8'h4e == _T_475[7:0] ? 4'h0 : _GEN_9488; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9490 = 8'h4f == _T_475[7:0] ? 4'h0 : _GEN_9489; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9491 = 8'h50 == _T_475[7:0] ? 4'hf : _GEN_9490; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9492 = 8'h51 == _T_475[7:0] ? 4'hf : _GEN_9491; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9493 = 8'h52 == _T_475[7:0] ? 4'hf : _GEN_9492; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9494 = 8'h53 == _T_475[7:0] ? 4'hf : _GEN_9493; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9495 = 8'h54 == _T_475[7:0] ? 4'hf : _GEN_9494; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9496 = 8'h55 == _T_475[7:0] ? 4'hf : _GEN_9495; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9497 = 8'h56 == _T_475[7:0] ? 4'hf : _GEN_9496; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9498 = 8'h57 == _T_475[7:0] ? 4'hf : _GEN_9497; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9499 = 8'h58 == _T_475[7:0] ? 4'h0 : _GEN_9498; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9500 = 8'h59 == _T_475[7:0] ? 4'h0 : _GEN_9499; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9501 = 8'h5a == _T_475[7:0] ? 4'h0 : _GEN_9500; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9502 = 8'h5b == _T_475[7:0] ? 4'h0 : _GEN_9501; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9503 = 8'h5c == _T_475[7:0] ? 4'h0 : _GEN_9502; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9504 = 8'h5d == _T_475[7:0] ? 4'h0 : _GEN_9503; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9505 = 8'h5e == _T_475[7:0] ? 4'h0 : _GEN_9504; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9506 = 8'h5f == _T_475[7:0] ? 4'h0 : _GEN_9505; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9507 = 8'h60 == _T_475[7:0] ? 4'h0 : _GEN_9506; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9508 = 8'h61 == _T_475[7:0] ? 4'h0 : _GEN_9507; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9509 = 8'h62 == _T_475[7:0] ? 4'h0 : _GEN_9508; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9510 = 8'h63 == _T_475[7:0] ? 4'h0 : _GEN_9509; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9511 = 8'h64 == _T_475[7:0] ? 4'h0 : _GEN_9510; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9512 = 8'h65 == _T_475[7:0] ? 4'h0 : _GEN_9511; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9513 = 8'h66 == _T_475[7:0] ? 4'h0 : _GEN_9512; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9514 = 8'h67 == _T_475[7:0] ? 4'h0 : _GEN_9513; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9515 = 8'h68 == _T_475[7:0] ? 4'hf : _GEN_9514; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9516 = 8'h69 == _T_475[7:0] ? 4'hf : _GEN_9515; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9517 = 8'h6a == _T_475[7:0] ? 4'hf : _GEN_9516; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9518 = 8'h6b == _T_475[7:0] ? 4'hf : _GEN_9517; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9519 = 8'h6c == _T_475[7:0] ? 4'hf : _GEN_9518; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9520 = 8'h6d == _T_475[7:0] ? 4'hf : _GEN_9519; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9521 = 8'h6e == _T_475[7:0] ? 4'hf : _GEN_9520; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9522 = 8'h6f == _T_475[7:0] ? 4'hf : _GEN_9521; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9523 = 8'h70 == _T_475[7:0] ? 4'h0 : _GEN_9522; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9524 = 8'h71 == _T_475[7:0] ? 4'h0 : _GEN_9523; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9525 = 8'h72 == _T_475[7:0] ? 4'h0 : _GEN_9524; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9526 = 8'h73 == _T_475[7:0] ? 4'h0 : _GEN_9525; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9527 = 8'h74 == _T_475[7:0] ? 4'h0 : _GEN_9526; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9528 = 8'h75 == _T_475[7:0] ? 4'h0 : _GEN_9527; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9529 = 8'h76 == _T_475[7:0] ? 4'h0 : _GEN_9528; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9530 = 8'h77 == _T_475[7:0] ? 4'h0 : _GEN_9529; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9531 = 8'h78 == _T_475[7:0] ? 4'hf : _GEN_9530; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9532 = 8'h79 == _T_475[7:0] ? 4'hf : _GEN_9531; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9533 = 8'h7a == _T_475[7:0] ? 4'hf : _GEN_9532; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9534 = 8'h7b == _T_475[7:0] ? 4'hf : _GEN_9533; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9535 = 8'h7c == _T_475[7:0] ? 4'hf : _GEN_9534; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9536 = 8'h7d == _T_475[7:0] ? 4'hf : _GEN_9535; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9537 = 8'h7e == _T_475[7:0] ? 4'hf : _GEN_9536; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9538 = 8'h7f == _T_475[7:0] ? 4'hf : _GEN_9537; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9539 = 8'h80 == _T_475[7:0] ? 4'h0 : _GEN_9538; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9540 = 8'h81 == _T_475[7:0] ? 4'h0 : _GEN_9539; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9541 = 8'h82 == _T_475[7:0] ? 4'h0 : _GEN_9540; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9542 = 8'h83 == _T_475[7:0] ? 4'h0 : _GEN_9541; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9543 = 8'h84 == _T_475[7:0] ? 4'h0 : _GEN_9542; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9544 = 8'h85 == _T_475[7:0] ? 4'h0 : _GEN_9543; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9545 = 8'h86 == _T_475[7:0] ? 4'h0 : _GEN_9544; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9546 = 8'h87 == _T_475[7:0] ? 4'h0 : _GEN_9545; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9547 = 8'h88 == _T_475[7:0] ? 4'hf : _GEN_9546; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9548 = 8'h89 == _T_475[7:0] ? 4'hf : _GEN_9547; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9549 = 8'h8a == _T_475[7:0] ? 4'hf : _GEN_9548; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9550 = 8'h8b == _T_475[7:0] ? 4'hf : _GEN_9549; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9551 = 8'h8c == _T_475[7:0] ? 4'hf : _GEN_9550; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9552 = 8'h8d == _T_475[7:0] ? 4'hf : _GEN_9551; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9553 = 8'h8e == _T_475[7:0] ? 4'hf : _GEN_9552; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9554 = 8'h8f == _T_475[7:0] ? 4'hf : _GEN_9553; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9555 = 8'h90 == _T_475[7:0] ? 4'h0 : _GEN_9554; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9556 = 8'h91 == _T_475[7:0] ? 4'h0 : _GEN_9555; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9557 = 8'h92 == _T_475[7:0] ? 4'h0 : _GEN_9556; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9558 = 8'h93 == _T_475[7:0] ? 4'h0 : _GEN_9557; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9559 = 8'h94 == _T_475[7:0] ? 4'h0 : _GEN_9558; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9560 = 8'h95 == _T_475[7:0] ? 4'h0 : _GEN_9559; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9561 = 8'h96 == _T_475[7:0] ? 4'h0 : _GEN_9560; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9562 = 8'h97 == _T_475[7:0] ? 4'h0 : _GEN_9561; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9563 = 8'h98 == _T_475[7:0] ? 4'hf : _GEN_9562; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9564 = 8'h99 == _T_475[7:0] ? 4'hf : _GEN_9563; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9565 = 8'h9a == _T_475[7:0] ? 4'hf : _GEN_9564; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9566 = 8'h9b == _T_475[7:0] ? 4'hf : _GEN_9565; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9567 = 8'h9c == _T_475[7:0] ? 4'hf : _GEN_9566; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9568 = 8'h9d == _T_475[7:0] ? 4'hf : _GEN_9567; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9569 = 8'h9e == _T_475[7:0] ? 4'hf : _GEN_9568; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9570 = 8'h9f == _T_475[7:0] ? 4'hf : _GEN_9569; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9571 = 8'ha0 == _T_475[7:0] ? 4'h0 : _GEN_9570; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9572 = 8'ha1 == _T_475[7:0] ? 4'h0 : _GEN_9571; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9573 = 8'ha2 == _T_475[7:0] ? 4'h0 : _GEN_9572; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9574 = 8'ha3 == _T_475[7:0] ? 4'h0 : _GEN_9573; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9575 = 8'ha4 == _T_475[7:0] ? 4'h0 : _GEN_9574; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9576 = 8'ha5 == _T_475[7:0] ? 4'h0 : _GEN_9575; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9577 = 8'ha6 == _T_475[7:0] ? 4'h0 : _GEN_9576; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9578 = 8'ha7 == _T_475[7:0] ? 4'h0 : _GEN_9577; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9579 = 8'ha8 == _T_475[7:0] ? 4'hf : _GEN_9578; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9580 = 8'ha9 == _T_475[7:0] ? 4'hf : _GEN_9579; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9581 = 8'haa == _T_475[7:0] ? 4'hf : _GEN_9580; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9582 = 8'hab == _T_475[7:0] ? 4'hf : _GEN_9581; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9583 = 8'hac == _T_475[7:0] ? 4'hf : _GEN_9582; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9584 = 8'had == _T_475[7:0] ? 4'hf : _GEN_9583; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9585 = 8'hae == _T_475[7:0] ? 4'hf : _GEN_9584; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9586 = 8'haf == _T_475[7:0] ? 4'hf : _GEN_9585; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9587 = 8'hb0 == _T_475[7:0] ? 4'h0 : _GEN_9586; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9588 = 8'hb1 == _T_475[7:0] ? 4'h0 : _GEN_9587; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9589 = 8'hb2 == _T_475[7:0] ? 4'h0 : _GEN_9588; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9590 = 8'hb3 == _T_475[7:0] ? 4'h0 : _GEN_9589; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9591 = 8'hb4 == _T_475[7:0] ? 4'h0 : _GEN_9590; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9592 = 8'hb5 == _T_475[7:0] ? 4'h0 : _GEN_9591; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9593 = 8'hb6 == _T_475[7:0] ? 4'h0 : _GEN_9592; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9594 = 8'hb7 == _T_475[7:0] ? 4'h0 : _GEN_9593; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9595 = 8'hb8 == _T_475[7:0] ? 4'hf : _GEN_9594; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9596 = 8'hb9 == _T_475[7:0] ? 4'hf : _GEN_9595; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9597 = 8'hba == _T_475[7:0] ? 4'hf : _GEN_9596; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9598 = 8'hbb == _T_475[7:0] ? 4'hf : _GEN_9597; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9599 = 8'hbc == _T_475[7:0] ? 4'hf : _GEN_9598; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9600 = 8'hbd == _T_475[7:0] ? 4'hf : _GEN_9599; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9601 = 8'hbe == _T_475[7:0] ? 4'hf : _GEN_9600; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9602 = 8'hbf == _T_475[7:0] ? 4'hf : _GEN_9601; // @[Filter.scala 165:86]
  wire [4:0] _GEN_19090 = {{1'd0}, _GEN_9602}; // @[Filter.scala 165:86]
  wire [8:0] _T_477 = _GEN_19090 * 5'h14; // @[Filter.scala 165:86]
  wire [3:0] _GEN_9699 = 8'h60 == _T_475[7:0] ? 4'hf : 4'h0; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9700 = 8'h61 == _T_475[7:0] ? 4'hf : _GEN_9699; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9701 = 8'h62 == _T_475[7:0] ? 4'hf : _GEN_9700; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9702 = 8'h63 == _T_475[7:0] ? 4'hf : _GEN_9701; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9703 = 8'h64 == _T_475[7:0] ? 4'hf : _GEN_9702; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9704 = 8'h65 == _T_475[7:0] ? 4'hf : _GEN_9703; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9705 = 8'h66 == _T_475[7:0] ? 4'hf : _GEN_9704; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9706 = 8'h67 == _T_475[7:0] ? 4'hf : _GEN_9705; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9707 = 8'h68 == _T_475[7:0] ? 4'hf : _GEN_9706; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9708 = 8'h69 == _T_475[7:0] ? 4'hf : _GEN_9707; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9709 = 8'h6a == _T_475[7:0] ? 4'hf : _GEN_9708; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9710 = 8'h6b == _T_475[7:0] ? 4'hf : _GEN_9709; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9711 = 8'h6c == _T_475[7:0] ? 4'hf : _GEN_9710; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9712 = 8'h6d == _T_475[7:0] ? 4'hf : _GEN_9711; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9713 = 8'h6e == _T_475[7:0] ? 4'hf : _GEN_9712; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9714 = 8'h6f == _T_475[7:0] ? 4'hf : _GEN_9713; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9715 = 8'h70 == _T_475[7:0] ? 4'hf : _GEN_9714; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9716 = 8'h71 == _T_475[7:0] ? 4'hf : _GEN_9715; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9717 = 8'h72 == _T_475[7:0] ? 4'hf : _GEN_9716; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9718 = 8'h73 == _T_475[7:0] ? 4'hf : _GEN_9717; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9719 = 8'h74 == _T_475[7:0] ? 4'hf : _GEN_9718; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9720 = 8'h75 == _T_475[7:0] ? 4'hf : _GEN_9719; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9721 = 8'h76 == _T_475[7:0] ? 4'hf : _GEN_9720; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9722 = 8'h77 == _T_475[7:0] ? 4'hf : _GEN_9721; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9723 = 8'h78 == _T_475[7:0] ? 4'hf : _GEN_9722; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9724 = 8'h79 == _T_475[7:0] ? 4'hf : _GEN_9723; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9725 = 8'h7a == _T_475[7:0] ? 4'hf : _GEN_9724; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9726 = 8'h7b == _T_475[7:0] ? 4'hf : _GEN_9725; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9727 = 8'h7c == _T_475[7:0] ? 4'hf : _GEN_9726; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9728 = 8'h7d == _T_475[7:0] ? 4'hf : _GEN_9727; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9729 = 8'h7e == _T_475[7:0] ? 4'hf : _GEN_9728; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9730 = 8'h7f == _T_475[7:0] ? 4'hf : _GEN_9729; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9731 = 8'h80 == _T_475[7:0] ? 4'hf : _GEN_9730; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9732 = 8'h81 == _T_475[7:0] ? 4'hf : _GEN_9731; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9733 = 8'h82 == _T_475[7:0] ? 4'hf : _GEN_9732; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9734 = 8'h83 == _T_475[7:0] ? 4'hf : _GEN_9733; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9735 = 8'h84 == _T_475[7:0] ? 4'hf : _GEN_9734; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9736 = 8'h85 == _T_475[7:0] ? 4'hf : _GEN_9735; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9737 = 8'h86 == _T_475[7:0] ? 4'hf : _GEN_9736; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9738 = 8'h87 == _T_475[7:0] ? 4'hf : _GEN_9737; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9739 = 8'h88 == _T_475[7:0] ? 4'hf : _GEN_9738; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9740 = 8'h89 == _T_475[7:0] ? 4'hf : _GEN_9739; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9741 = 8'h8a == _T_475[7:0] ? 4'hf : _GEN_9740; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9742 = 8'h8b == _T_475[7:0] ? 4'hf : _GEN_9741; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9743 = 8'h8c == _T_475[7:0] ? 4'hf : _GEN_9742; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9744 = 8'h8d == _T_475[7:0] ? 4'hf : _GEN_9743; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9745 = 8'h8e == _T_475[7:0] ? 4'hf : _GEN_9744; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9746 = 8'h8f == _T_475[7:0] ? 4'hf : _GEN_9745; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9747 = 8'h90 == _T_475[7:0] ? 4'hf : _GEN_9746; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9748 = 8'h91 == _T_475[7:0] ? 4'hf : _GEN_9747; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9749 = 8'h92 == _T_475[7:0] ? 4'hf : _GEN_9748; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9750 = 8'h93 == _T_475[7:0] ? 4'hf : _GEN_9749; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9751 = 8'h94 == _T_475[7:0] ? 4'hf : _GEN_9750; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9752 = 8'h95 == _T_475[7:0] ? 4'hf : _GEN_9751; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9753 = 8'h96 == _T_475[7:0] ? 4'hf : _GEN_9752; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9754 = 8'h97 == _T_475[7:0] ? 4'hf : _GEN_9753; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9755 = 8'h98 == _T_475[7:0] ? 4'hf : _GEN_9754; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9756 = 8'h99 == _T_475[7:0] ? 4'hf : _GEN_9755; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9757 = 8'h9a == _T_475[7:0] ? 4'hf : _GEN_9756; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9758 = 8'h9b == _T_475[7:0] ? 4'hf : _GEN_9757; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9759 = 8'h9c == _T_475[7:0] ? 4'hf : _GEN_9758; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9760 = 8'h9d == _T_475[7:0] ? 4'hf : _GEN_9759; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9761 = 8'h9e == _T_475[7:0] ? 4'hf : _GEN_9760; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9762 = 8'h9f == _T_475[7:0] ? 4'hf : _GEN_9761; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9763 = 8'ha0 == _T_475[7:0] ? 4'hf : _GEN_9762; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9764 = 8'ha1 == _T_475[7:0] ? 4'hf : _GEN_9763; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9765 = 8'ha2 == _T_475[7:0] ? 4'hf : _GEN_9764; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9766 = 8'ha3 == _T_475[7:0] ? 4'hf : _GEN_9765; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9767 = 8'ha4 == _T_475[7:0] ? 4'hf : _GEN_9766; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9768 = 8'ha5 == _T_475[7:0] ? 4'hf : _GEN_9767; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9769 = 8'ha6 == _T_475[7:0] ? 4'hf : _GEN_9768; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9770 = 8'ha7 == _T_475[7:0] ? 4'hf : _GEN_9769; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9771 = 8'ha8 == _T_475[7:0] ? 4'hf : _GEN_9770; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9772 = 8'ha9 == _T_475[7:0] ? 4'hf : _GEN_9771; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9773 = 8'haa == _T_475[7:0] ? 4'hf : _GEN_9772; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9774 = 8'hab == _T_475[7:0] ? 4'hf : _GEN_9773; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9775 = 8'hac == _T_475[7:0] ? 4'hf : _GEN_9774; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9776 = 8'had == _T_475[7:0] ? 4'hf : _GEN_9775; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9777 = 8'hae == _T_475[7:0] ? 4'hf : _GEN_9776; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9778 = 8'haf == _T_475[7:0] ? 4'hf : _GEN_9777; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9779 = 8'hb0 == _T_475[7:0] ? 4'hf : _GEN_9778; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9780 = 8'hb1 == _T_475[7:0] ? 4'hf : _GEN_9779; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9781 = 8'hb2 == _T_475[7:0] ? 4'hf : _GEN_9780; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9782 = 8'hb3 == _T_475[7:0] ? 4'hf : _GEN_9781; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9783 = 8'hb4 == _T_475[7:0] ? 4'hf : _GEN_9782; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9784 = 8'hb5 == _T_475[7:0] ? 4'hf : _GEN_9783; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9785 = 8'hb6 == _T_475[7:0] ? 4'hf : _GEN_9784; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9786 = 8'hb7 == _T_475[7:0] ? 4'hf : _GEN_9785; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9787 = 8'hb8 == _T_475[7:0] ? 4'hf : _GEN_9786; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9788 = 8'hb9 == _T_475[7:0] ? 4'hf : _GEN_9787; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9789 = 8'hba == _T_475[7:0] ? 4'hf : _GEN_9788; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9790 = 8'hbb == _T_475[7:0] ? 4'hf : _GEN_9789; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9791 = 8'hbc == _T_475[7:0] ? 4'hf : _GEN_9790; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9792 = 8'hbd == _T_475[7:0] ? 4'hf : _GEN_9791; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9793 = 8'hbe == _T_475[7:0] ? 4'hf : _GEN_9792; // @[Filter.scala 165:126]
  wire [3:0] _GEN_9794 = 8'hbf == _T_475[7:0] ? 4'hf : _GEN_9793; // @[Filter.scala 165:126]
  wire [6:0] _GEN_19092 = {{3'd0}, _GEN_9794}; // @[Filter.scala 165:126]
  wire [10:0] _T_482 = _GEN_19092 * 7'h46; // @[Filter.scala 165:126]
  wire [10:0] _GEN_19093 = {{2'd0}, _T_477}; // @[Filter.scala 165:93]
  wire [10:0] _T_484 = _GEN_19093 + _T_482; // @[Filter.scala 165:93]
  wire [3:0] _GEN_9803 = 8'h8 == _T_475[7:0] ? 4'hf : 4'h0; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9804 = 8'h9 == _T_475[7:0] ? 4'hf : _GEN_9803; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9805 = 8'ha == _T_475[7:0] ? 4'hf : _GEN_9804; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9806 = 8'hb == _T_475[7:0] ? 4'hf : _GEN_9805; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9807 = 8'hc == _T_475[7:0] ? 4'hf : _GEN_9806; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9808 = 8'hd == _T_475[7:0] ? 4'hf : _GEN_9807; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9809 = 8'he == _T_475[7:0] ? 4'hf : _GEN_9808; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9810 = 8'hf == _T_475[7:0] ? 4'hf : _GEN_9809; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9811 = 8'h10 == _T_475[7:0] ? 4'h0 : _GEN_9810; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9812 = 8'h11 == _T_475[7:0] ? 4'h0 : _GEN_9811; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9813 = 8'h12 == _T_475[7:0] ? 4'h0 : _GEN_9812; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9814 = 8'h13 == _T_475[7:0] ? 4'h0 : _GEN_9813; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9815 = 8'h14 == _T_475[7:0] ? 4'h0 : _GEN_9814; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9816 = 8'h15 == _T_475[7:0] ? 4'h0 : _GEN_9815; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9817 = 8'h16 == _T_475[7:0] ? 4'h0 : _GEN_9816; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9818 = 8'h17 == _T_475[7:0] ? 4'h0 : _GEN_9817; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9819 = 8'h18 == _T_475[7:0] ? 4'hf : _GEN_9818; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9820 = 8'h19 == _T_475[7:0] ? 4'hf : _GEN_9819; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9821 = 8'h1a == _T_475[7:0] ? 4'hf : _GEN_9820; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9822 = 8'h1b == _T_475[7:0] ? 4'hf : _GEN_9821; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9823 = 8'h1c == _T_475[7:0] ? 4'hf : _GEN_9822; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9824 = 8'h1d == _T_475[7:0] ? 4'hf : _GEN_9823; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9825 = 8'h1e == _T_475[7:0] ? 4'hf : _GEN_9824; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9826 = 8'h1f == _T_475[7:0] ? 4'hf : _GEN_9825; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9827 = 8'h20 == _T_475[7:0] ? 4'h0 : _GEN_9826; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9828 = 8'h21 == _T_475[7:0] ? 4'h0 : _GEN_9827; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9829 = 8'h22 == _T_475[7:0] ? 4'h0 : _GEN_9828; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9830 = 8'h23 == _T_475[7:0] ? 4'h0 : _GEN_9829; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9831 = 8'h24 == _T_475[7:0] ? 4'h0 : _GEN_9830; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9832 = 8'h25 == _T_475[7:0] ? 4'h0 : _GEN_9831; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9833 = 8'h26 == _T_475[7:0] ? 4'h0 : _GEN_9832; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9834 = 8'h27 == _T_475[7:0] ? 4'h0 : _GEN_9833; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9835 = 8'h28 == _T_475[7:0] ? 4'hf : _GEN_9834; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9836 = 8'h29 == _T_475[7:0] ? 4'hf : _GEN_9835; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9837 = 8'h2a == _T_475[7:0] ? 4'hf : _GEN_9836; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9838 = 8'h2b == _T_475[7:0] ? 4'hf : _GEN_9837; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9839 = 8'h2c == _T_475[7:0] ? 4'hf : _GEN_9838; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9840 = 8'h2d == _T_475[7:0] ? 4'hf : _GEN_9839; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9841 = 8'h2e == _T_475[7:0] ? 4'hf : _GEN_9840; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9842 = 8'h2f == _T_475[7:0] ? 4'hf : _GEN_9841; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9843 = 8'h30 == _T_475[7:0] ? 4'h0 : _GEN_9842; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9844 = 8'h31 == _T_475[7:0] ? 4'h0 : _GEN_9843; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9845 = 8'h32 == _T_475[7:0] ? 4'h0 : _GEN_9844; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9846 = 8'h33 == _T_475[7:0] ? 4'h0 : _GEN_9845; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9847 = 8'h34 == _T_475[7:0] ? 4'h0 : _GEN_9846; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9848 = 8'h35 == _T_475[7:0] ? 4'h0 : _GEN_9847; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9849 = 8'h36 == _T_475[7:0] ? 4'h0 : _GEN_9848; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9850 = 8'h37 == _T_475[7:0] ? 4'h0 : _GEN_9849; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9851 = 8'h38 == _T_475[7:0] ? 4'hf : _GEN_9850; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9852 = 8'h39 == _T_475[7:0] ? 4'hf : _GEN_9851; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9853 = 8'h3a == _T_475[7:0] ? 4'hf : _GEN_9852; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9854 = 8'h3b == _T_475[7:0] ? 4'hf : _GEN_9853; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9855 = 8'h3c == _T_475[7:0] ? 4'hf : _GEN_9854; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9856 = 8'h3d == _T_475[7:0] ? 4'hf : _GEN_9855; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9857 = 8'h3e == _T_475[7:0] ? 4'hf : _GEN_9856; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9858 = 8'h3f == _T_475[7:0] ? 4'hf : _GEN_9857; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9859 = 8'h40 == _T_475[7:0] ? 4'h0 : _GEN_9858; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9860 = 8'h41 == _T_475[7:0] ? 4'h0 : _GEN_9859; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9861 = 8'h42 == _T_475[7:0] ? 4'h0 : _GEN_9860; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9862 = 8'h43 == _T_475[7:0] ? 4'h0 : _GEN_9861; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9863 = 8'h44 == _T_475[7:0] ? 4'h0 : _GEN_9862; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9864 = 8'h45 == _T_475[7:0] ? 4'h0 : _GEN_9863; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9865 = 8'h46 == _T_475[7:0] ? 4'h0 : _GEN_9864; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9866 = 8'h47 == _T_475[7:0] ? 4'h0 : _GEN_9865; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9867 = 8'h48 == _T_475[7:0] ? 4'hf : _GEN_9866; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9868 = 8'h49 == _T_475[7:0] ? 4'hf : _GEN_9867; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9869 = 8'h4a == _T_475[7:0] ? 4'hf : _GEN_9868; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9870 = 8'h4b == _T_475[7:0] ? 4'hf : _GEN_9869; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9871 = 8'h4c == _T_475[7:0] ? 4'hf : _GEN_9870; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9872 = 8'h4d == _T_475[7:0] ? 4'hf : _GEN_9871; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9873 = 8'h4e == _T_475[7:0] ? 4'hf : _GEN_9872; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9874 = 8'h4f == _T_475[7:0] ? 4'hf : _GEN_9873; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9875 = 8'h50 == _T_475[7:0] ? 4'h0 : _GEN_9874; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9876 = 8'h51 == _T_475[7:0] ? 4'h0 : _GEN_9875; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9877 = 8'h52 == _T_475[7:0] ? 4'h0 : _GEN_9876; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9878 = 8'h53 == _T_475[7:0] ? 4'h0 : _GEN_9877; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9879 = 8'h54 == _T_475[7:0] ? 4'h0 : _GEN_9878; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9880 = 8'h55 == _T_475[7:0] ? 4'h0 : _GEN_9879; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9881 = 8'h56 == _T_475[7:0] ? 4'h0 : _GEN_9880; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9882 = 8'h57 == _T_475[7:0] ? 4'h0 : _GEN_9881; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9883 = 8'h58 == _T_475[7:0] ? 4'hf : _GEN_9882; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9884 = 8'h59 == _T_475[7:0] ? 4'hf : _GEN_9883; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9885 = 8'h5a == _T_475[7:0] ? 4'hf : _GEN_9884; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9886 = 8'h5b == _T_475[7:0] ? 4'hf : _GEN_9885; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9887 = 8'h5c == _T_475[7:0] ? 4'hf : _GEN_9886; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9888 = 8'h5d == _T_475[7:0] ? 4'hf : _GEN_9887; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9889 = 8'h5e == _T_475[7:0] ? 4'hf : _GEN_9888; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9890 = 8'h5f == _T_475[7:0] ? 4'hf : _GEN_9889; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9891 = 8'h60 == _T_475[7:0] ? 4'h0 : _GEN_9890; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9892 = 8'h61 == _T_475[7:0] ? 4'h0 : _GEN_9891; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9893 = 8'h62 == _T_475[7:0] ? 4'h0 : _GEN_9892; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9894 = 8'h63 == _T_475[7:0] ? 4'h0 : _GEN_9893; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9895 = 8'h64 == _T_475[7:0] ? 4'h0 : _GEN_9894; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9896 = 8'h65 == _T_475[7:0] ? 4'h0 : _GEN_9895; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9897 = 8'h66 == _T_475[7:0] ? 4'h0 : _GEN_9896; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9898 = 8'h67 == _T_475[7:0] ? 4'h0 : _GEN_9897; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9899 = 8'h68 == _T_475[7:0] ? 4'hf : _GEN_9898; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9900 = 8'h69 == _T_475[7:0] ? 4'hf : _GEN_9899; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9901 = 8'h6a == _T_475[7:0] ? 4'hf : _GEN_9900; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9902 = 8'h6b == _T_475[7:0] ? 4'hf : _GEN_9901; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9903 = 8'h6c == _T_475[7:0] ? 4'hf : _GEN_9902; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9904 = 8'h6d == _T_475[7:0] ? 4'hf : _GEN_9903; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9905 = 8'h6e == _T_475[7:0] ? 4'hf : _GEN_9904; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9906 = 8'h6f == _T_475[7:0] ? 4'hf : _GEN_9905; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9907 = 8'h70 == _T_475[7:0] ? 4'h0 : _GEN_9906; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9908 = 8'h71 == _T_475[7:0] ? 4'h0 : _GEN_9907; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9909 = 8'h72 == _T_475[7:0] ? 4'h0 : _GEN_9908; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9910 = 8'h73 == _T_475[7:0] ? 4'h0 : _GEN_9909; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9911 = 8'h74 == _T_475[7:0] ? 4'h0 : _GEN_9910; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9912 = 8'h75 == _T_475[7:0] ? 4'h0 : _GEN_9911; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9913 = 8'h76 == _T_475[7:0] ? 4'h0 : _GEN_9912; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9914 = 8'h77 == _T_475[7:0] ? 4'h0 : _GEN_9913; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9915 = 8'h78 == _T_475[7:0] ? 4'hf : _GEN_9914; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9916 = 8'h79 == _T_475[7:0] ? 4'hf : _GEN_9915; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9917 = 8'h7a == _T_475[7:0] ? 4'hf : _GEN_9916; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9918 = 8'h7b == _T_475[7:0] ? 4'hf : _GEN_9917; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9919 = 8'h7c == _T_475[7:0] ? 4'hf : _GEN_9918; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9920 = 8'h7d == _T_475[7:0] ? 4'hf : _GEN_9919; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9921 = 8'h7e == _T_475[7:0] ? 4'hf : _GEN_9920; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9922 = 8'h7f == _T_475[7:0] ? 4'hf : _GEN_9921; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9923 = 8'h80 == _T_475[7:0] ? 4'h0 : _GEN_9922; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9924 = 8'h81 == _T_475[7:0] ? 4'h0 : _GEN_9923; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9925 = 8'h82 == _T_475[7:0] ? 4'h0 : _GEN_9924; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9926 = 8'h83 == _T_475[7:0] ? 4'h0 : _GEN_9925; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9927 = 8'h84 == _T_475[7:0] ? 4'h0 : _GEN_9926; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9928 = 8'h85 == _T_475[7:0] ? 4'h0 : _GEN_9927; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9929 = 8'h86 == _T_475[7:0] ? 4'h0 : _GEN_9928; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9930 = 8'h87 == _T_475[7:0] ? 4'h0 : _GEN_9929; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9931 = 8'h88 == _T_475[7:0] ? 4'hf : _GEN_9930; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9932 = 8'h89 == _T_475[7:0] ? 4'hf : _GEN_9931; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9933 = 8'h8a == _T_475[7:0] ? 4'hf : _GEN_9932; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9934 = 8'h8b == _T_475[7:0] ? 4'hf : _GEN_9933; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9935 = 8'h8c == _T_475[7:0] ? 4'hf : _GEN_9934; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9936 = 8'h8d == _T_475[7:0] ? 4'hf : _GEN_9935; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9937 = 8'h8e == _T_475[7:0] ? 4'hf : _GEN_9936; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9938 = 8'h8f == _T_475[7:0] ? 4'hf : _GEN_9937; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9939 = 8'h90 == _T_475[7:0] ? 4'h0 : _GEN_9938; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9940 = 8'h91 == _T_475[7:0] ? 4'h0 : _GEN_9939; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9941 = 8'h92 == _T_475[7:0] ? 4'h0 : _GEN_9940; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9942 = 8'h93 == _T_475[7:0] ? 4'h0 : _GEN_9941; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9943 = 8'h94 == _T_475[7:0] ? 4'h0 : _GEN_9942; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9944 = 8'h95 == _T_475[7:0] ? 4'h0 : _GEN_9943; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9945 = 8'h96 == _T_475[7:0] ? 4'h0 : _GEN_9944; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9946 = 8'h97 == _T_475[7:0] ? 4'h0 : _GEN_9945; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9947 = 8'h98 == _T_475[7:0] ? 4'hf : _GEN_9946; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9948 = 8'h99 == _T_475[7:0] ? 4'hf : _GEN_9947; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9949 = 8'h9a == _T_475[7:0] ? 4'hf : _GEN_9948; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9950 = 8'h9b == _T_475[7:0] ? 4'hf : _GEN_9949; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9951 = 8'h9c == _T_475[7:0] ? 4'hf : _GEN_9950; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9952 = 8'h9d == _T_475[7:0] ? 4'hf : _GEN_9951; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9953 = 8'h9e == _T_475[7:0] ? 4'hf : _GEN_9952; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9954 = 8'h9f == _T_475[7:0] ? 4'hf : _GEN_9953; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9955 = 8'ha0 == _T_475[7:0] ? 4'h0 : _GEN_9954; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9956 = 8'ha1 == _T_475[7:0] ? 4'h0 : _GEN_9955; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9957 = 8'ha2 == _T_475[7:0] ? 4'h0 : _GEN_9956; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9958 = 8'ha3 == _T_475[7:0] ? 4'h0 : _GEN_9957; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9959 = 8'ha4 == _T_475[7:0] ? 4'h0 : _GEN_9958; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9960 = 8'ha5 == _T_475[7:0] ? 4'h0 : _GEN_9959; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9961 = 8'ha6 == _T_475[7:0] ? 4'h0 : _GEN_9960; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9962 = 8'ha7 == _T_475[7:0] ? 4'h0 : _GEN_9961; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9963 = 8'ha8 == _T_475[7:0] ? 4'hf : _GEN_9962; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9964 = 8'ha9 == _T_475[7:0] ? 4'hf : _GEN_9963; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9965 = 8'haa == _T_475[7:0] ? 4'hf : _GEN_9964; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9966 = 8'hab == _T_475[7:0] ? 4'hf : _GEN_9965; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9967 = 8'hac == _T_475[7:0] ? 4'hf : _GEN_9966; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9968 = 8'had == _T_475[7:0] ? 4'hf : _GEN_9967; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9969 = 8'hae == _T_475[7:0] ? 4'hf : _GEN_9968; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9970 = 8'haf == _T_475[7:0] ? 4'hf : _GEN_9969; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9971 = 8'hb0 == _T_475[7:0] ? 4'h0 : _GEN_9970; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9972 = 8'hb1 == _T_475[7:0] ? 4'h0 : _GEN_9971; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9973 = 8'hb2 == _T_475[7:0] ? 4'h0 : _GEN_9972; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9974 = 8'hb3 == _T_475[7:0] ? 4'h0 : _GEN_9973; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9975 = 8'hb4 == _T_475[7:0] ? 4'h0 : _GEN_9974; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9976 = 8'hb5 == _T_475[7:0] ? 4'h0 : _GEN_9975; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9977 = 8'hb6 == _T_475[7:0] ? 4'h0 : _GEN_9976; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9978 = 8'hb7 == _T_475[7:0] ? 4'h0 : _GEN_9977; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9979 = 8'hb8 == _T_475[7:0] ? 4'hf : _GEN_9978; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9980 = 8'hb9 == _T_475[7:0] ? 4'hf : _GEN_9979; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9981 = 8'hba == _T_475[7:0] ? 4'hf : _GEN_9980; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9982 = 8'hbb == _T_475[7:0] ? 4'hf : _GEN_9981; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9983 = 8'hbc == _T_475[7:0] ? 4'hf : _GEN_9982; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9984 = 8'hbd == _T_475[7:0] ? 4'hf : _GEN_9983; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9985 = 8'hbe == _T_475[7:0] ? 4'hf : _GEN_9984; // @[Filter.scala 165:166]
  wire [3:0] _GEN_9986 = 8'hbf == _T_475[7:0] ? 4'hf : _GEN_9985; // @[Filter.scala 165:166]
  wire [7:0] _T_489 = _GEN_9986 * 4'ha; // @[Filter.scala 165:166]
  wire [10:0] _GEN_19095 = {{3'd0}, _T_489}; // @[Filter.scala 165:133]
  wire [10:0] _T_491 = _T_484 + _GEN_19095; // @[Filter.scala 165:133]
  wire [10:0] _T_492 = _T_491 / 11'h64; // @[Filter.scala 165:174]
  wire [10:0] _GEN_10179 = io_SPI_distort ? _T_492 : {{7'd0}, _GEN_9602}; // @[Filter.scala 164:35]
  wire [10:0] _GEN_10180 = _T_472 ? 11'h0 : _GEN_10179; // @[Filter.scala 162:80]
  wire [10:0] _GEN_10949 = io_SPI_distort ? _T_492 : {{7'd0}, _GEN_9794}; // @[Filter.scala 164:35]
  wire [10:0] _GEN_10950 = _T_472 ? 11'h0 : _GEN_10949; // @[Filter.scala 162:80]
  wire [10:0] _GEN_11719 = io_SPI_distort ? _T_492 : {{7'd0}, _GEN_9986}; // @[Filter.scala 164:35]
  wire [10:0] _GEN_11720 = _T_472 ? 11'h0 : _GEN_11719; // @[Filter.scala 162:80]
  wire [31:0] _T_560 = pixelIndex + 32'h5; // @[Filter.scala 158:31]
  wire [31:0] _GEN_5 = _T_560 % 32'h10; // @[Filter.scala 158:38]
  wire [4:0] _T_561 = _GEN_5[4:0]; // @[Filter.scala 158:38]
  wire [4:0] _T_563 = _T_561 + _GEN_18983; // @[Filter.scala 158:53]
  wire [4:0] _T_565 = _T_563 - 5'h1; // @[Filter.scala 158:69]
  wire [31:0] _T_568 = _T_560 / 32'h10; // @[Filter.scala 159:38]
  wire [31:0] _T_570 = _T_568 + _GEN_18984; // @[Filter.scala 159:53]
  wire [31:0] _T_572 = _T_570 - 32'h1; // @[Filter.scala 159:69]
  wire  _T_574 = _T_565 >= 5'h10; // @[Filter.scala 162:31]
  wire  _T_578 = _T_572 >= 32'hc; // @[Filter.scala 162:63]
  wire  _T_579 = _T_574 | _T_578; // @[Filter.scala 162:58]
  wire [36:0] _T_580 = _T_572 * 32'h10; // @[Filter.scala 165:66]
  wire [36:0] _GEN_19115 = {{32'd0}, _T_565}; // @[Filter.scala 165:81]
  wire [36:0] _T_582 = _T_580 + _GEN_19115; // @[Filter.scala 165:81]
  wire [3:0] _GEN_11729 = 8'h8 == _T_582[7:0] ? 4'h0 : 4'hf; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11730 = 8'h9 == _T_582[7:0] ? 4'h0 : _GEN_11729; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11731 = 8'ha == _T_582[7:0] ? 4'h0 : _GEN_11730; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11732 = 8'hb == _T_582[7:0] ? 4'h0 : _GEN_11731; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11733 = 8'hc == _T_582[7:0] ? 4'h0 : _GEN_11732; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11734 = 8'hd == _T_582[7:0] ? 4'h0 : _GEN_11733; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11735 = 8'he == _T_582[7:0] ? 4'h0 : _GEN_11734; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11736 = 8'hf == _T_582[7:0] ? 4'h0 : _GEN_11735; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11737 = 8'h10 == _T_582[7:0] ? 4'hf : _GEN_11736; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11738 = 8'h11 == _T_582[7:0] ? 4'hf : _GEN_11737; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11739 = 8'h12 == _T_582[7:0] ? 4'hf : _GEN_11738; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11740 = 8'h13 == _T_582[7:0] ? 4'hf : _GEN_11739; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11741 = 8'h14 == _T_582[7:0] ? 4'hf : _GEN_11740; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11742 = 8'h15 == _T_582[7:0] ? 4'hf : _GEN_11741; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11743 = 8'h16 == _T_582[7:0] ? 4'hf : _GEN_11742; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11744 = 8'h17 == _T_582[7:0] ? 4'hf : _GEN_11743; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11745 = 8'h18 == _T_582[7:0] ? 4'h0 : _GEN_11744; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11746 = 8'h19 == _T_582[7:0] ? 4'h0 : _GEN_11745; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11747 = 8'h1a == _T_582[7:0] ? 4'h0 : _GEN_11746; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11748 = 8'h1b == _T_582[7:0] ? 4'h0 : _GEN_11747; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11749 = 8'h1c == _T_582[7:0] ? 4'h0 : _GEN_11748; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11750 = 8'h1d == _T_582[7:0] ? 4'h0 : _GEN_11749; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11751 = 8'h1e == _T_582[7:0] ? 4'h0 : _GEN_11750; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11752 = 8'h1f == _T_582[7:0] ? 4'h0 : _GEN_11751; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11753 = 8'h20 == _T_582[7:0] ? 4'hf : _GEN_11752; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11754 = 8'h21 == _T_582[7:0] ? 4'hf : _GEN_11753; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11755 = 8'h22 == _T_582[7:0] ? 4'hf : _GEN_11754; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11756 = 8'h23 == _T_582[7:0] ? 4'hf : _GEN_11755; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11757 = 8'h24 == _T_582[7:0] ? 4'hf : _GEN_11756; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11758 = 8'h25 == _T_582[7:0] ? 4'hf : _GEN_11757; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11759 = 8'h26 == _T_582[7:0] ? 4'hf : _GEN_11758; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11760 = 8'h27 == _T_582[7:0] ? 4'hf : _GEN_11759; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11761 = 8'h28 == _T_582[7:0] ? 4'h0 : _GEN_11760; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11762 = 8'h29 == _T_582[7:0] ? 4'h0 : _GEN_11761; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11763 = 8'h2a == _T_582[7:0] ? 4'h0 : _GEN_11762; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11764 = 8'h2b == _T_582[7:0] ? 4'h0 : _GEN_11763; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11765 = 8'h2c == _T_582[7:0] ? 4'h0 : _GEN_11764; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11766 = 8'h2d == _T_582[7:0] ? 4'h0 : _GEN_11765; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11767 = 8'h2e == _T_582[7:0] ? 4'h0 : _GEN_11766; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11768 = 8'h2f == _T_582[7:0] ? 4'h0 : _GEN_11767; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11769 = 8'h30 == _T_582[7:0] ? 4'hf : _GEN_11768; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11770 = 8'h31 == _T_582[7:0] ? 4'hf : _GEN_11769; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11771 = 8'h32 == _T_582[7:0] ? 4'hf : _GEN_11770; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11772 = 8'h33 == _T_582[7:0] ? 4'hf : _GEN_11771; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11773 = 8'h34 == _T_582[7:0] ? 4'hf : _GEN_11772; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11774 = 8'h35 == _T_582[7:0] ? 4'hf : _GEN_11773; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11775 = 8'h36 == _T_582[7:0] ? 4'hf : _GEN_11774; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11776 = 8'h37 == _T_582[7:0] ? 4'hf : _GEN_11775; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11777 = 8'h38 == _T_582[7:0] ? 4'h0 : _GEN_11776; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11778 = 8'h39 == _T_582[7:0] ? 4'h0 : _GEN_11777; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11779 = 8'h3a == _T_582[7:0] ? 4'h0 : _GEN_11778; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11780 = 8'h3b == _T_582[7:0] ? 4'h0 : _GEN_11779; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11781 = 8'h3c == _T_582[7:0] ? 4'h0 : _GEN_11780; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11782 = 8'h3d == _T_582[7:0] ? 4'h0 : _GEN_11781; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11783 = 8'h3e == _T_582[7:0] ? 4'h0 : _GEN_11782; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11784 = 8'h3f == _T_582[7:0] ? 4'h0 : _GEN_11783; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11785 = 8'h40 == _T_582[7:0] ? 4'hf : _GEN_11784; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11786 = 8'h41 == _T_582[7:0] ? 4'hf : _GEN_11785; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11787 = 8'h42 == _T_582[7:0] ? 4'hf : _GEN_11786; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11788 = 8'h43 == _T_582[7:0] ? 4'hf : _GEN_11787; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11789 = 8'h44 == _T_582[7:0] ? 4'hf : _GEN_11788; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11790 = 8'h45 == _T_582[7:0] ? 4'hf : _GEN_11789; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11791 = 8'h46 == _T_582[7:0] ? 4'hf : _GEN_11790; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11792 = 8'h47 == _T_582[7:0] ? 4'hf : _GEN_11791; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11793 = 8'h48 == _T_582[7:0] ? 4'h0 : _GEN_11792; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11794 = 8'h49 == _T_582[7:0] ? 4'h0 : _GEN_11793; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11795 = 8'h4a == _T_582[7:0] ? 4'h0 : _GEN_11794; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11796 = 8'h4b == _T_582[7:0] ? 4'h0 : _GEN_11795; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11797 = 8'h4c == _T_582[7:0] ? 4'h0 : _GEN_11796; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11798 = 8'h4d == _T_582[7:0] ? 4'h0 : _GEN_11797; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11799 = 8'h4e == _T_582[7:0] ? 4'h0 : _GEN_11798; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11800 = 8'h4f == _T_582[7:0] ? 4'h0 : _GEN_11799; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11801 = 8'h50 == _T_582[7:0] ? 4'hf : _GEN_11800; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11802 = 8'h51 == _T_582[7:0] ? 4'hf : _GEN_11801; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11803 = 8'h52 == _T_582[7:0] ? 4'hf : _GEN_11802; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11804 = 8'h53 == _T_582[7:0] ? 4'hf : _GEN_11803; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11805 = 8'h54 == _T_582[7:0] ? 4'hf : _GEN_11804; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11806 = 8'h55 == _T_582[7:0] ? 4'hf : _GEN_11805; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11807 = 8'h56 == _T_582[7:0] ? 4'hf : _GEN_11806; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11808 = 8'h57 == _T_582[7:0] ? 4'hf : _GEN_11807; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11809 = 8'h58 == _T_582[7:0] ? 4'h0 : _GEN_11808; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11810 = 8'h59 == _T_582[7:0] ? 4'h0 : _GEN_11809; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11811 = 8'h5a == _T_582[7:0] ? 4'h0 : _GEN_11810; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11812 = 8'h5b == _T_582[7:0] ? 4'h0 : _GEN_11811; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11813 = 8'h5c == _T_582[7:0] ? 4'h0 : _GEN_11812; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11814 = 8'h5d == _T_582[7:0] ? 4'h0 : _GEN_11813; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11815 = 8'h5e == _T_582[7:0] ? 4'h0 : _GEN_11814; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11816 = 8'h5f == _T_582[7:0] ? 4'h0 : _GEN_11815; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11817 = 8'h60 == _T_582[7:0] ? 4'h0 : _GEN_11816; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11818 = 8'h61 == _T_582[7:0] ? 4'h0 : _GEN_11817; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11819 = 8'h62 == _T_582[7:0] ? 4'h0 : _GEN_11818; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11820 = 8'h63 == _T_582[7:0] ? 4'h0 : _GEN_11819; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11821 = 8'h64 == _T_582[7:0] ? 4'h0 : _GEN_11820; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11822 = 8'h65 == _T_582[7:0] ? 4'h0 : _GEN_11821; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11823 = 8'h66 == _T_582[7:0] ? 4'h0 : _GEN_11822; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11824 = 8'h67 == _T_582[7:0] ? 4'h0 : _GEN_11823; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11825 = 8'h68 == _T_582[7:0] ? 4'hf : _GEN_11824; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11826 = 8'h69 == _T_582[7:0] ? 4'hf : _GEN_11825; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11827 = 8'h6a == _T_582[7:0] ? 4'hf : _GEN_11826; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11828 = 8'h6b == _T_582[7:0] ? 4'hf : _GEN_11827; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11829 = 8'h6c == _T_582[7:0] ? 4'hf : _GEN_11828; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11830 = 8'h6d == _T_582[7:0] ? 4'hf : _GEN_11829; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11831 = 8'h6e == _T_582[7:0] ? 4'hf : _GEN_11830; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11832 = 8'h6f == _T_582[7:0] ? 4'hf : _GEN_11831; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11833 = 8'h70 == _T_582[7:0] ? 4'h0 : _GEN_11832; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11834 = 8'h71 == _T_582[7:0] ? 4'h0 : _GEN_11833; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11835 = 8'h72 == _T_582[7:0] ? 4'h0 : _GEN_11834; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11836 = 8'h73 == _T_582[7:0] ? 4'h0 : _GEN_11835; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11837 = 8'h74 == _T_582[7:0] ? 4'h0 : _GEN_11836; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11838 = 8'h75 == _T_582[7:0] ? 4'h0 : _GEN_11837; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11839 = 8'h76 == _T_582[7:0] ? 4'h0 : _GEN_11838; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11840 = 8'h77 == _T_582[7:0] ? 4'h0 : _GEN_11839; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11841 = 8'h78 == _T_582[7:0] ? 4'hf : _GEN_11840; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11842 = 8'h79 == _T_582[7:0] ? 4'hf : _GEN_11841; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11843 = 8'h7a == _T_582[7:0] ? 4'hf : _GEN_11842; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11844 = 8'h7b == _T_582[7:0] ? 4'hf : _GEN_11843; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11845 = 8'h7c == _T_582[7:0] ? 4'hf : _GEN_11844; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11846 = 8'h7d == _T_582[7:0] ? 4'hf : _GEN_11845; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11847 = 8'h7e == _T_582[7:0] ? 4'hf : _GEN_11846; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11848 = 8'h7f == _T_582[7:0] ? 4'hf : _GEN_11847; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11849 = 8'h80 == _T_582[7:0] ? 4'h0 : _GEN_11848; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11850 = 8'h81 == _T_582[7:0] ? 4'h0 : _GEN_11849; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11851 = 8'h82 == _T_582[7:0] ? 4'h0 : _GEN_11850; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11852 = 8'h83 == _T_582[7:0] ? 4'h0 : _GEN_11851; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11853 = 8'h84 == _T_582[7:0] ? 4'h0 : _GEN_11852; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11854 = 8'h85 == _T_582[7:0] ? 4'h0 : _GEN_11853; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11855 = 8'h86 == _T_582[7:0] ? 4'h0 : _GEN_11854; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11856 = 8'h87 == _T_582[7:0] ? 4'h0 : _GEN_11855; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11857 = 8'h88 == _T_582[7:0] ? 4'hf : _GEN_11856; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11858 = 8'h89 == _T_582[7:0] ? 4'hf : _GEN_11857; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11859 = 8'h8a == _T_582[7:0] ? 4'hf : _GEN_11858; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11860 = 8'h8b == _T_582[7:0] ? 4'hf : _GEN_11859; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11861 = 8'h8c == _T_582[7:0] ? 4'hf : _GEN_11860; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11862 = 8'h8d == _T_582[7:0] ? 4'hf : _GEN_11861; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11863 = 8'h8e == _T_582[7:0] ? 4'hf : _GEN_11862; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11864 = 8'h8f == _T_582[7:0] ? 4'hf : _GEN_11863; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11865 = 8'h90 == _T_582[7:0] ? 4'h0 : _GEN_11864; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11866 = 8'h91 == _T_582[7:0] ? 4'h0 : _GEN_11865; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11867 = 8'h92 == _T_582[7:0] ? 4'h0 : _GEN_11866; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11868 = 8'h93 == _T_582[7:0] ? 4'h0 : _GEN_11867; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11869 = 8'h94 == _T_582[7:0] ? 4'h0 : _GEN_11868; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11870 = 8'h95 == _T_582[7:0] ? 4'h0 : _GEN_11869; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11871 = 8'h96 == _T_582[7:0] ? 4'h0 : _GEN_11870; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11872 = 8'h97 == _T_582[7:0] ? 4'h0 : _GEN_11871; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11873 = 8'h98 == _T_582[7:0] ? 4'hf : _GEN_11872; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11874 = 8'h99 == _T_582[7:0] ? 4'hf : _GEN_11873; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11875 = 8'h9a == _T_582[7:0] ? 4'hf : _GEN_11874; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11876 = 8'h9b == _T_582[7:0] ? 4'hf : _GEN_11875; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11877 = 8'h9c == _T_582[7:0] ? 4'hf : _GEN_11876; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11878 = 8'h9d == _T_582[7:0] ? 4'hf : _GEN_11877; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11879 = 8'h9e == _T_582[7:0] ? 4'hf : _GEN_11878; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11880 = 8'h9f == _T_582[7:0] ? 4'hf : _GEN_11879; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11881 = 8'ha0 == _T_582[7:0] ? 4'h0 : _GEN_11880; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11882 = 8'ha1 == _T_582[7:0] ? 4'h0 : _GEN_11881; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11883 = 8'ha2 == _T_582[7:0] ? 4'h0 : _GEN_11882; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11884 = 8'ha3 == _T_582[7:0] ? 4'h0 : _GEN_11883; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11885 = 8'ha4 == _T_582[7:0] ? 4'h0 : _GEN_11884; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11886 = 8'ha5 == _T_582[7:0] ? 4'h0 : _GEN_11885; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11887 = 8'ha6 == _T_582[7:0] ? 4'h0 : _GEN_11886; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11888 = 8'ha7 == _T_582[7:0] ? 4'h0 : _GEN_11887; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11889 = 8'ha8 == _T_582[7:0] ? 4'hf : _GEN_11888; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11890 = 8'ha9 == _T_582[7:0] ? 4'hf : _GEN_11889; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11891 = 8'haa == _T_582[7:0] ? 4'hf : _GEN_11890; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11892 = 8'hab == _T_582[7:0] ? 4'hf : _GEN_11891; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11893 = 8'hac == _T_582[7:0] ? 4'hf : _GEN_11892; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11894 = 8'had == _T_582[7:0] ? 4'hf : _GEN_11893; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11895 = 8'hae == _T_582[7:0] ? 4'hf : _GEN_11894; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11896 = 8'haf == _T_582[7:0] ? 4'hf : _GEN_11895; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11897 = 8'hb0 == _T_582[7:0] ? 4'h0 : _GEN_11896; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11898 = 8'hb1 == _T_582[7:0] ? 4'h0 : _GEN_11897; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11899 = 8'hb2 == _T_582[7:0] ? 4'h0 : _GEN_11898; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11900 = 8'hb3 == _T_582[7:0] ? 4'h0 : _GEN_11899; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11901 = 8'hb4 == _T_582[7:0] ? 4'h0 : _GEN_11900; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11902 = 8'hb5 == _T_582[7:0] ? 4'h0 : _GEN_11901; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11903 = 8'hb6 == _T_582[7:0] ? 4'h0 : _GEN_11902; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11904 = 8'hb7 == _T_582[7:0] ? 4'h0 : _GEN_11903; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11905 = 8'hb8 == _T_582[7:0] ? 4'hf : _GEN_11904; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11906 = 8'hb9 == _T_582[7:0] ? 4'hf : _GEN_11905; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11907 = 8'hba == _T_582[7:0] ? 4'hf : _GEN_11906; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11908 = 8'hbb == _T_582[7:0] ? 4'hf : _GEN_11907; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11909 = 8'hbc == _T_582[7:0] ? 4'hf : _GEN_11908; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11910 = 8'hbd == _T_582[7:0] ? 4'hf : _GEN_11909; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11911 = 8'hbe == _T_582[7:0] ? 4'hf : _GEN_11910; // @[Filter.scala 165:86]
  wire [3:0] _GEN_11912 = 8'hbf == _T_582[7:0] ? 4'hf : _GEN_11911; // @[Filter.scala 165:86]
  wire [4:0] _GEN_19116 = {{1'd0}, _GEN_11912}; // @[Filter.scala 165:86]
  wire [8:0] _T_584 = _GEN_19116 * 5'h14; // @[Filter.scala 165:86]
  wire [3:0] _GEN_12009 = 8'h60 == _T_582[7:0] ? 4'hf : 4'h0; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12010 = 8'h61 == _T_582[7:0] ? 4'hf : _GEN_12009; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12011 = 8'h62 == _T_582[7:0] ? 4'hf : _GEN_12010; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12012 = 8'h63 == _T_582[7:0] ? 4'hf : _GEN_12011; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12013 = 8'h64 == _T_582[7:0] ? 4'hf : _GEN_12012; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12014 = 8'h65 == _T_582[7:0] ? 4'hf : _GEN_12013; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12015 = 8'h66 == _T_582[7:0] ? 4'hf : _GEN_12014; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12016 = 8'h67 == _T_582[7:0] ? 4'hf : _GEN_12015; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12017 = 8'h68 == _T_582[7:0] ? 4'hf : _GEN_12016; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12018 = 8'h69 == _T_582[7:0] ? 4'hf : _GEN_12017; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12019 = 8'h6a == _T_582[7:0] ? 4'hf : _GEN_12018; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12020 = 8'h6b == _T_582[7:0] ? 4'hf : _GEN_12019; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12021 = 8'h6c == _T_582[7:0] ? 4'hf : _GEN_12020; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12022 = 8'h6d == _T_582[7:0] ? 4'hf : _GEN_12021; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12023 = 8'h6e == _T_582[7:0] ? 4'hf : _GEN_12022; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12024 = 8'h6f == _T_582[7:0] ? 4'hf : _GEN_12023; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12025 = 8'h70 == _T_582[7:0] ? 4'hf : _GEN_12024; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12026 = 8'h71 == _T_582[7:0] ? 4'hf : _GEN_12025; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12027 = 8'h72 == _T_582[7:0] ? 4'hf : _GEN_12026; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12028 = 8'h73 == _T_582[7:0] ? 4'hf : _GEN_12027; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12029 = 8'h74 == _T_582[7:0] ? 4'hf : _GEN_12028; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12030 = 8'h75 == _T_582[7:0] ? 4'hf : _GEN_12029; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12031 = 8'h76 == _T_582[7:0] ? 4'hf : _GEN_12030; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12032 = 8'h77 == _T_582[7:0] ? 4'hf : _GEN_12031; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12033 = 8'h78 == _T_582[7:0] ? 4'hf : _GEN_12032; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12034 = 8'h79 == _T_582[7:0] ? 4'hf : _GEN_12033; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12035 = 8'h7a == _T_582[7:0] ? 4'hf : _GEN_12034; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12036 = 8'h7b == _T_582[7:0] ? 4'hf : _GEN_12035; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12037 = 8'h7c == _T_582[7:0] ? 4'hf : _GEN_12036; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12038 = 8'h7d == _T_582[7:0] ? 4'hf : _GEN_12037; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12039 = 8'h7e == _T_582[7:0] ? 4'hf : _GEN_12038; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12040 = 8'h7f == _T_582[7:0] ? 4'hf : _GEN_12039; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12041 = 8'h80 == _T_582[7:0] ? 4'hf : _GEN_12040; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12042 = 8'h81 == _T_582[7:0] ? 4'hf : _GEN_12041; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12043 = 8'h82 == _T_582[7:0] ? 4'hf : _GEN_12042; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12044 = 8'h83 == _T_582[7:0] ? 4'hf : _GEN_12043; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12045 = 8'h84 == _T_582[7:0] ? 4'hf : _GEN_12044; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12046 = 8'h85 == _T_582[7:0] ? 4'hf : _GEN_12045; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12047 = 8'h86 == _T_582[7:0] ? 4'hf : _GEN_12046; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12048 = 8'h87 == _T_582[7:0] ? 4'hf : _GEN_12047; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12049 = 8'h88 == _T_582[7:0] ? 4'hf : _GEN_12048; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12050 = 8'h89 == _T_582[7:0] ? 4'hf : _GEN_12049; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12051 = 8'h8a == _T_582[7:0] ? 4'hf : _GEN_12050; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12052 = 8'h8b == _T_582[7:0] ? 4'hf : _GEN_12051; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12053 = 8'h8c == _T_582[7:0] ? 4'hf : _GEN_12052; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12054 = 8'h8d == _T_582[7:0] ? 4'hf : _GEN_12053; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12055 = 8'h8e == _T_582[7:0] ? 4'hf : _GEN_12054; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12056 = 8'h8f == _T_582[7:0] ? 4'hf : _GEN_12055; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12057 = 8'h90 == _T_582[7:0] ? 4'hf : _GEN_12056; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12058 = 8'h91 == _T_582[7:0] ? 4'hf : _GEN_12057; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12059 = 8'h92 == _T_582[7:0] ? 4'hf : _GEN_12058; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12060 = 8'h93 == _T_582[7:0] ? 4'hf : _GEN_12059; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12061 = 8'h94 == _T_582[7:0] ? 4'hf : _GEN_12060; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12062 = 8'h95 == _T_582[7:0] ? 4'hf : _GEN_12061; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12063 = 8'h96 == _T_582[7:0] ? 4'hf : _GEN_12062; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12064 = 8'h97 == _T_582[7:0] ? 4'hf : _GEN_12063; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12065 = 8'h98 == _T_582[7:0] ? 4'hf : _GEN_12064; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12066 = 8'h99 == _T_582[7:0] ? 4'hf : _GEN_12065; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12067 = 8'h9a == _T_582[7:0] ? 4'hf : _GEN_12066; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12068 = 8'h9b == _T_582[7:0] ? 4'hf : _GEN_12067; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12069 = 8'h9c == _T_582[7:0] ? 4'hf : _GEN_12068; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12070 = 8'h9d == _T_582[7:0] ? 4'hf : _GEN_12069; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12071 = 8'h9e == _T_582[7:0] ? 4'hf : _GEN_12070; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12072 = 8'h9f == _T_582[7:0] ? 4'hf : _GEN_12071; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12073 = 8'ha0 == _T_582[7:0] ? 4'hf : _GEN_12072; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12074 = 8'ha1 == _T_582[7:0] ? 4'hf : _GEN_12073; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12075 = 8'ha2 == _T_582[7:0] ? 4'hf : _GEN_12074; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12076 = 8'ha3 == _T_582[7:0] ? 4'hf : _GEN_12075; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12077 = 8'ha4 == _T_582[7:0] ? 4'hf : _GEN_12076; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12078 = 8'ha5 == _T_582[7:0] ? 4'hf : _GEN_12077; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12079 = 8'ha6 == _T_582[7:0] ? 4'hf : _GEN_12078; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12080 = 8'ha7 == _T_582[7:0] ? 4'hf : _GEN_12079; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12081 = 8'ha8 == _T_582[7:0] ? 4'hf : _GEN_12080; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12082 = 8'ha9 == _T_582[7:0] ? 4'hf : _GEN_12081; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12083 = 8'haa == _T_582[7:0] ? 4'hf : _GEN_12082; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12084 = 8'hab == _T_582[7:0] ? 4'hf : _GEN_12083; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12085 = 8'hac == _T_582[7:0] ? 4'hf : _GEN_12084; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12086 = 8'had == _T_582[7:0] ? 4'hf : _GEN_12085; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12087 = 8'hae == _T_582[7:0] ? 4'hf : _GEN_12086; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12088 = 8'haf == _T_582[7:0] ? 4'hf : _GEN_12087; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12089 = 8'hb0 == _T_582[7:0] ? 4'hf : _GEN_12088; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12090 = 8'hb1 == _T_582[7:0] ? 4'hf : _GEN_12089; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12091 = 8'hb2 == _T_582[7:0] ? 4'hf : _GEN_12090; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12092 = 8'hb3 == _T_582[7:0] ? 4'hf : _GEN_12091; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12093 = 8'hb4 == _T_582[7:0] ? 4'hf : _GEN_12092; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12094 = 8'hb5 == _T_582[7:0] ? 4'hf : _GEN_12093; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12095 = 8'hb6 == _T_582[7:0] ? 4'hf : _GEN_12094; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12096 = 8'hb7 == _T_582[7:0] ? 4'hf : _GEN_12095; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12097 = 8'hb8 == _T_582[7:0] ? 4'hf : _GEN_12096; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12098 = 8'hb9 == _T_582[7:0] ? 4'hf : _GEN_12097; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12099 = 8'hba == _T_582[7:0] ? 4'hf : _GEN_12098; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12100 = 8'hbb == _T_582[7:0] ? 4'hf : _GEN_12099; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12101 = 8'hbc == _T_582[7:0] ? 4'hf : _GEN_12100; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12102 = 8'hbd == _T_582[7:0] ? 4'hf : _GEN_12101; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12103 = 8'hbe == _T_582[7:0] ? 4'hf : _GEN_12102; // @[Filter.scala 165:126]
  wire [3:0] _GEN_12104 = 8'hbf == _T_582[7:0] ? 4'hf : _GEN_12103; // @[Filter.scala 165:126]
  wire [6:0] _GEN_19118 = {{3'd0}, _GEN_12104}; // @[Filter.scala 165:126]
  wire [10:0] _T_589 = _GEN_19118 * 7'h46; // @[Filter.scala 165:126]
  wire [10:0] _GEN_19119 = {{2'd0}, _T_584}; // @[Filter.scala 165:93]
  wire [10:0] _T_591 = _GEN_19119 + _T_589; // @[Filter.scala 165:93]
  wire [3:0] _GEN_12113 = 8'h8 == _T_582[7:0] ? 4'hf : 4'h0; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12114 = 8'h9 == _T_582[7:0] ? 4'hf : _GEN_12113; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12115 = 8'ha == _T_582[7:0] ? 4'hf : _GEN_12114; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12116 = 8'hb == _T_582[7:0] ? 4'hf : _GEN_12115; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12117 = 8'hc == _T_582[7:0] ? 4'hf : _GEN_12116; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12118 = 8'hd == _T_582[7:0] ? 4'hf : _GEN_12117; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12119 = 8'he == _T_582[7:0] ? 4'hf : _GEN_12118; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12120 = 8'hf == _T_582[7:0] ? 4'hf : _GEN_12119; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12121 = 8'h10 == _T_582[7:0] ? 4'h0 : _GEN_12120; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12122 = 8'h11 == _T_582[7:0] ? 4'h0 : _GEN_12121; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12123 = 8'h12 == _T_582[7:0] ? 4'h0 : _GEN_12122; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12124 = 8'h13 == _T_582[7:0] ? 4'h0 : _GEN_12123; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12125 = 8'h14 == _T_582[7:0] ? 4'h0 : _GEN_12124; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12126 = 8'h15 == _T_582[7:0] ? 4'h0 : _GEN_12125; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12127 = 8'h16 == _T_582[7:0] ? 4'h0 : _GEN_12126; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12128 = 8'h17 == _T_582[7:0] ? 4'h0 : _GEN_12127; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12129 = 8'h18 == _T_582[7:0] ? 4'hf : _GEN_12128; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12130 = 8'h19 == _T_582[7:0] ? 4'hf : _GEN_12129; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12131 = 8'h1a == _T_582[7:0] ? 4'hf : _GEN_12130; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12132 = 8'h1b == _T_582[7:0] ? 4'hf : _GEN_12131; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12133 = 8'h1c == _T_582[7:0] ? 4'hf : _GEN_12132; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12134 = 8'h1d == _T_582[7:0] ? 4'hf : _GEN_12133; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12135 = 8'h1e == _T_582[7:0] ? 4'hf : _GEN_12134; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12136 = 8'h1f == _T_582[7:0] ? 4'hf : _GEN_12135; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12137 = 8'h20 == _T_582[7:0] ? 4'h0 : _GEN_12136; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12138 = 8'h21 == _T_582[7:0] ? 4'h0 : _GEN_12137; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12139 = 8'h22 == _T_582[7:0] ? 4'h0 : _GEN_12138; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12140 = 8'h23 == _T_582[7:0] ? 4'h0 : _GEN_12139; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12141 = 8'h24 == _T_582[7:0] ? 4'h0 : _GEN_12140; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12142 = 8'h25 == _T_582[7:0] ? 4'h0 : _GEN_12141; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12143 = 8'h26 == _T_582[7:0] ? 4'h0 : _GEN_12142; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12144 = 8'h27 == _T_582[7:0] ? 4'h0 : _GEN_12143; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12145 = 8'h28 == _T_582[7:0] ? 4'hf : _GEN_12144; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12146 = 8'h29 == _T_582[7:0] ? 4'hf : _GEN_12145; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12147 = 8'h2a == _T_582[7:0] ? 4'hf : _GEN_12146; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12148 = 8'h2b == _T_582[7:0] ? 4'hf : _GEN_12147; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12149 = 8'h2c == _T_582[7:0] ? 4'hf : _GEN_12148; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12150 = 8'h2d == _T_582[7:0] ? 4'hf : _GEN_12149; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12151 = 8'h2e == _T_582[7:0] ? 4'hf : _GEN_12150; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12152 = 8'h2f == _T_582[7:0] ? 4'hf : _GEN_12151; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12153 = 8'h30 == _T_582[7:0] ? 4'h0 : _GEN_12152; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12154 = 8'h31 == _T_582[7:0] ? 4'h0 : _GEN_12153; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12155 = 8'h32 == _T_582[7:0] ? 4'h0 : _GEN_12154; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12156 = 8'h33 == _T_582[7:0] ? 4'h0 : _GEN_12155; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12157 = 8'h34 == _T_582[7:0] ? 4'h0 : _GEN_12156; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12158 = 8'h35 == _T_582[7:0] ? 4'h0 : _GEN_12157; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12159 = 8'h36 == _T_582[7:0] ? 4'h0 : _GEN_12158; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12160 = 8'h37 == _T_582[7:0] ? 4'h0 : _GEN_12159; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12161 = 8'h38 == _T_582[7:0] ? 4'hf : _GEN_12160; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12162 = 8'h39 == _T_582[7:0] ? 4'hf : _GEN_12161; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12163 = 8'h3a == _T_582[7:0] ? 4'hf : _GEN_12162; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12164 = 8'h3b == _T_582[7:0] ? 4'hf : _GEN_12163; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12165 = 8'h3c == _T_582[7:0] ? 4'hf : _GEN_12164; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12166 = 8'h3d == _T_582[7:0] ? 4'hf : _GEN_12165; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12167 = 8'h3e == _T_582[7:0] ? 4'hf : _GEN_12166; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12168 = 8'h3f == _T_582[7:0] ? 4'hf : _GEN_12167; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12169 = 8'h40 == _T_582[7:0] ? 4'h0 : _GEN_12168; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12170 = 8'h41 == _T_582[7:0] ? 4'h0 : _GEN_12169; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12171 = 8'h42 == _T_582[7:0] ? 4'h0 : _GEN_12170; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12172 = 8'h43 == _T_582[7:0] ? 4'h0 : _GEN_12171; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12173 = 8'h44 == _T_582[7:0] ? 4'h0 : _GEN_12172; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12174 = 8'h45 == _T_582[7:0] ? 4'h0 : _GEN_12173; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12175 = 8'h46 == _T_582[7:0] ? 4'h0 : _GEN_12174; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12176 = 8'h47 == _T_582[7:0] ? 4'h0 : _GEN_12175; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12177 = 8'h48 == _T_582[7:0] ? 4'hf : _GEN_12176; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12178 = 8'h49 == _T_582[7:0] ? 4'hf : _GEN_12177; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12179 = 8'h4a == _T_582[7:0] ? 4'hf : _GEN_12178; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12180 = 8'h4b == _T_582[7:0] ? 4'hf : _GEN_12179; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12181 = 8'h4c == _T_582[7:0] ? 4'hf : _GEN_12180; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12182 = 8'h4d == _T_582[7:0] ? 4'hf : _GEN_12181; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12183 = 8'h4e == _T_582[7:0] ? 4'hf : _GEN_12182; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12184 = 8'h4f == _T_582[7:0] ? 4'hf : _GEN_12183; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12185 = 8'h50 == _T_582[7:0] ? 4'h0 : _GEN_12184; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12186 = 8'h51 == _T_582[7:0] ? 4'h0 : _GEN_12185; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12187 = 8'h52 == _T_582[7:0] ? 4'h0 : _GEN_12186; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12188 = 8'h53 == _T_582[7:0] ? 4'h0 : _GEN_12187; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12189 = 8'h54 == _T_582[7:0] ? 4'h0 : _GEN_12188; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12190 = 8'h55 == _T_582[7:0] ? 4'h0 : _GEN_12189; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12191 = 8'h56 == _T_582[7:0] ? 4'h0 : _GEN_12190; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12192 = 8'h57 == _T_582[7:0] ? 4'h0 : _GEN_12191; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12193 = 8'h58 == _T_582[7:0] ? 4'hf : _GEN_12192; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12194 = 8'h59 == _T_582[7:0] ? 4'hf : _GEN_12193; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12195 = 8'h5a == _T_582[7:0] ? 4'hf : _GEN_12194; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12196 = 8'h5b == _T_582[7:0] ? 4'hf : _GEN_12195; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12197 = 8'h5c == _T_582[7:0] ? 4'hf : _GEN_12196; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12198 = 8'h5d == _T_582[7:0] ? 4'hf : _GEN_12197; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12199 = 8'h5e == _T_582[7:0] ? 4'hf : _GEN_12198; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12200 = 8'h5f == _T_582[7:0] ? 4'hf : _GEN_12199; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12201 = 8'h60 == _T_582[7:0] ? 4'h0 : _GEN_12200; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12202 = 8'h61 == _T_582[7:0] ? 4'h0 : _GEN_12201; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12203 = 8'h62 == _T_582[7:0] ? 4'h0 : _GEN_12202; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12204 = 8'h63 == _T_582[7:0] ? 4'h0 : _GEN_12203; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12205 = 8'h64 == _T_582[7:0] ? 4'h0 : _GEN_12204; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12206 = 8'h65 == _T_582[7:0] ? 4'h0 : _GEN_12205; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12207 = 8'h66 == _T_582[7:0] ? 4'h0 : _GEN_12206; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12208 = 8'h67 == _T_582[7:0] ? 4'h0 : _GEN_12207; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12209 = 8'h68 == _T_582[7:0] ? 4'hf : _GEN_12208; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12210 = 8'h69 == _T_582[7:0] ? 4'hf : _GEN_12209; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12211 = 8'h6a == _T_582[7:0] ? 4'hf : _GEN_12210; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12212 = 8'h6b == _T_582[7:0] ? 4'hf : _GEN_12211; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12213 = 8'h6c == _T_582[7:0] ? 4'hf : _GEN_12212; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12214 = 8'h6d == _T_582[7:0] ? 4'hf : _GEN_12213; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12215 = 8'h6e == _T_582[7:0] ? 4'hf : _GEN_12214; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12216 = 8'h6f == _T_582[7:0] ? 4'hf : _GEN_12215; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12217 = 8'h70 == _T_582[7:0] ? 4'h0 : _GEN_12216; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12218 = 8'h71 == _T_582[7:0] ? 4'h0 : _GEN_12217; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12219 = 8'h72 == _T_582[7:0] ? 4'h0 : _GEN_12218; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12220 = 8'h73 == _T_582[7:0] ? 4'h0 : _GEN_12219; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12221 = 8'h74 == _T_582[7:0] ? 4'h0 : _GEN_12220; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12222 = 8'h75 == _T_582[7:0] ? 4'h0 : _GEN_12221; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12223 = 8'h76 == _T_582[7:0] ? 4'h0 : _GEN_12222; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12224 = 8'h77 == _T_582[7:0] ? 4'h0 : _GEN_12223; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12225 = 8'h78 == _T_582[7:0] ? 4'hf : _GEN_12224; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12226 = 8'h79 == _T_582[7:0] ? 4'hf : _GEN_12225; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12227 = 8'h7a == _T_582[7:0] ? 4'hf : _GEN_12226; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12228 = 8'h7b == _T_582[7:0] ? 4'hf : _GEN_12227; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12229 = 8'h7c == _T_582[7:0] ? 4'hf : _GEN_12228; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12230 = 8'h7d == _T_582[7:0] ? 4'hf : _GEN_12229; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12231 = 8'h7e == _T_582[7:0] ? 4'hf : _GEN_12230; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12232 = 8'h7f == _T_582[7:0] ? 4'hf : _GEN_12231; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12233 = 8'h80 == _T_582[7:0] ? 4'h0 : _GEN_12232; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12234 = 8'h81 == _T_582[7:0] ? 4'h0 : _GEN_12233; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12235 = 8'h82 == _T_582[7:0] ? 4'h0 : _GEN_12234; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12236 = 8'h83 == _T_582[7:0] ? 4'h0 : _GEN_12235; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12237 = 8'h84 == _T_582[7:0] ? 4'h0 : _GEN_12236; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12238 = 8'h85 == _T_582[7:0] ? 4'h0 : _GEN_12237; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12239 = 8'h86 == _T_582[7:0] ? 4'h0 : _GEN_12238; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12240 = 8'h87 == _T_582[7:0] ? 4'h0 : _GEN_12239; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12241 = 8'h88 == _T_582[7:0] ? 4'hf : _GEN_12240; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12242 = 8'h89 == _T_582[7:0] ? 4'hf : _GEN_12241; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12243 = 8'h8a == _T_582[7:0] ? 4'hf : _GEN_12242; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12244 = 8'h8b == _T_582[7:0] ? 4'hf : _GEN_12243; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12245 = 8'h8c == _T_582[7:0] ? 4'hf : _GEN_12244; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12246 = 8'h8d == _T_582[7:0] ? 4'hf : _GEN_12245; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12247 = 8'h8e == _T_582[7:0] ? 4'hf : _GEN_12246; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12248 = 8'h8f == _T_582[7:0] ? 4'hf : _GEN_12247; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12249 = 8'h90 == _T_582[7:0] ? 4'h0 : _GEN_12248; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12250 = 8'h91 == _T_582[7:0] ? 4'h0 : _GEN_12249; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12251 = 8'h92 == _T_582[7:0] ? 4'h0 : _GEN_12250; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12252 = 8'h93 == _T_582[7:0] ? 4'h0 : _GEN_12251; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12253 = 8'h94 == _T_582[7:0] ? 4'h0 : _GEN_12252; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12254 = 8'h95 == _T_582[7:0] ? 4'h0 : _GEN_12253; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12255 = 8'h96 == _T_582[7:0] ? 4'h0 : _GEN_12254; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12256 = 8'h97 == _T_582[7:0] ? 4'h0 : _GEN_12255; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12257 = 8'h98 == _T_582[7:0] ? 4'hf : _GEN_12256; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12258 = 8'h99 == _T_582[7:0] ? 4'hf : _GEN_12257; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12259 = 8'h9a == _T_582[7:0] ? 4'hf : _GEN_12258; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12260 = 8'h9b == _T_582[7:0] ? 4'hf : _GEN_12259; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12261 = 8'h9c == _T_582[7:0] ? 4'hf : _GEN_12260; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12262 = 8'h9d == _T_582[7:0] ? 4'hf : _GEN_12261; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12263 = 8'h9e == _T_582[7:0] ? 4'hf : _GEN_12262; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12264 = 8'h9f == _T_582[7:0] ? 4'hf : _GEN_12263; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12265 = 8'ha0 == _T_582[7:0] ? 4'h0 : _GEN_12264; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12266 = 8'ha1 == _T_582[7:0] ? 4'h0 : _GEN_12265; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12267 = 8'ha2 == _T_582[7:0] ? 4'h0 : _GEN_12266; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12268 = 8'ha3 == _T_582[7:0] ? 4'h0 : _GEN_12267; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12269 = 8'ha4 == _T_582[7:0] ? 4'h0 : _GEN_12268; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12270 = 8'ha5 == _T_582[7:0] ? 4'h0 : _GEN_12269; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12271 = 8'ha6 == _T_582[7:0] ? 4'h0 : _GEN_12270; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12272 = 8'ha7 == _T_582[7:0] ? 4'h0 : _GEN_12271; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12273 = 8'ha8 == _T_582[7:0] ? 4'hf : _GEN_12272; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12274 = 8'ha9 == _T_582[7:0] ? 4'hf : _GEN_12273; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12275 = 8'haa == _T_582[7:0] ? 4'hf : _GEN_12274; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12276 = 8'hab == _T_582[7:0] ? 4'hf : _GEN_12275; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12277 = 8'hac == _T_582[7:0] ? 4'hf : _GEN_12276; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12278 = 8'had == _T_582[7:0] ? 4'hf : _GEN_12277; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12279 = 8'hae == _T_582[7:0] ? 4'hf : _GEN_12278; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12280 = 8'haf == _T_582[7:0] ? 4'hf : _GEN_12279; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12281 = 8'hb0 == _T_582[7:0] ? 4'h0 : _GEN_12280; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12282 = 8'hb1 == _T_582[7:0] ? 4'h0 : _GEN_12281; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12283 = 8'hb2 == _T_582[7:0] ? 4'h0 : _GEN_12282; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12284 = 8'hb3 == _T_582[7:0] ? 4'h0 : _GEN_12283; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12285 = 8'hb4 == _T_582[7:0] ? 4'h0 : _GEN_12284; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12286 = 8'hb5 == _T_582[7:0] ? 4'h0 : _GEN_12285; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12287 = 8'hb6 == _T_582[7:0] ? 4'h0 : _GEN_12286; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12288 = 8'hb7 == _T_582[7:0] ? 4'h0 : _GEN_12287; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12289 = 8'hb8 == _T_582[7:0] ? 4'hf : _GEN_12288; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12290 = 8'hb9 == _T_582[7:0] ? 4'hf : _GEN_12289; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12291 = 8'hba == _T_582[7:0] ? 4'hf : _GEN_12290; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12292 = 8'hbb == _T_582[7:0] ? 4'hf : _GEN_12291; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12293 = 8'hbc == _T_582[7:0] ? 4'hf : _GEN_12292; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12294 = 8'hbd == _T_582[7:0] ? 4'hf : _GEN_12293; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12295 = 8'hbe == _T_582[7:0] ? 4'hf : _GEN_12294; // @[Filter.scala 165:166]
  wire [3:0] _GEN_12296 = 8'hbf == _T_582[7:0] ? 4'hf : _GEN_12295; // @[Filter.scala 165:166]
  wire [7:0] _T_596 = _GEN_12296 * 4'ha; // @[Filter.scala 165:166]
  wire [10:0] _GEN_19121 = {{3'd0}, _T_596}; // @[Filter.scala 165:133]
  wire [10:0] _T_598 = _T_591 + _GEN_19121; // @[Filter.scala 165:133]
  wire [10:0] _T_599 = _T_598 / 11'h64; // @[Filter.scala 165:174]
  wire [10:0] _GEN_12489 = io_SPI_distort ? _T_599 : {{7'd0}, _GEN_11912}; // @[Filter.scala 164:35]
  wire [10:0] _GEN_12490 = _T_579 ? 11'h0 : _GEN_12489; // @[Filter.scala 162:80]
  wire [10:0] _GEN_13259 = io_SPI_distort ? _T_599 : {{7'd0}, _GEN_12104}; // @[Filter.scala 164:35]
  wire [10:0] _GEN_13260 = _T_579 ? 11'h0 : _GEN_13259; // @[Filter.scala 162:80]
  wire [10:0] _GEN_14029 = io_SPI_distort ? _T_599 : {{7'd0}, _GEN_12296}; // @[Filter.scala 164:35]
  wire [10:0] _GEN_14030 = _T_579 ? 11'h0 : _GEN_14029; // @[Filter.scala 162:80]
  wire [31:0] _T_667 = pixelIndex + 32'h6; // @[Filter.scala 158:31]
  wire [31:0] _GEN_6 = _T_667 % 32'h10; // @[Filter.scala 158:38]
  wire [4:0] _T_668 = _GEN_6[4:0]; // @[Filter.scala 158:38]
  wire [4:0] _T_670 = _T_668 + _GEN_18983; // @[Filter.scala 158:53]
  wire [4:0] _T_672 = _T_670 - 5'h1; // @[Filter.scala 158:69]
  wire [31:0] _T_675 = _T_667 / 32'h10; // @[Filter.scala 159:38]
  wire [31:0] _T_677 = _T_675 + _GEN_18984; // @[Filter.scala 159:53]
  wire [31:0] _T_679 = _T_677 - 32'h1; // @[Filter.scala 159:69]
  wire  _T_681 = _T_672 >= 5'h10; // @[Filter.scala 162:31]
  wire  _T_685 = _T_679 >= 32'hc; // @[Filter.scala 162:63]
  wire  _T_686 = _T_681 | _T_685; // @[Filter.scala 162:58]
  wire [36:0] _T_687 = _T_679 * 32'h10; // @[Filter.scala 165:66]
  wire [36:0] _GEN_19141 = {{32'd0}, _T_672}; // @[Filter.scala 165:81]
  wire [36:0] _T_689 = _T_687 + _GEN_19141; // @[Filter.scala 165:81]
  wire [3:0] _GEN_14039 = 8'h8 == _T_689[7:0] ? 4'h0 : 4'hf; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14040 = 8'h9 == _T_689[7:0] ? 4'h0 : _GEN_14039; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14041 = 8'ha == _T_689[7:0] ? 4'h0 : _GEN_14040; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14042 = 8'hb == _T_689[7:0] ? 4'h0 : _GEN_14041; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14043 = 8'hc == _T_689[7:0] ? 4'h0 : _GEN_14042; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14044 = 8'hd == _T_689[7:0] ? 4'h0 : _GEN_14043; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14045 = 8'he == _T_689[7:0] ? 4'h0 : _GEN_14044; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14046 = 8'hf == _T_689[7:0] ? 4'h0 : _GEN_14045; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14047 = 8'h10 == _T_689[7:0] ? 4'hf : _GEN_14046; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14048 = 8'h11 == _T_689[7:0] ? 4'hf : _GEN_14047; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14049 = 8'h12 == _T_689[7:0] ? 4'hf : _GEN_14048; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14050 = 8'h13 == _T_689[7:0] ? 4'hf : _GEN_14049; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14051 = 8'h14 == _T_689[7:0] ? 4'hf : _GEN_14050; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14052 = 8'h15 == _T_689[7:0] ? 4'hf : _GEN_14051; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14053 = 8'h16 == _T_689[7:0] ? 4'hf : _GEN_14052; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14054 = 8'h17 == _T_689[7:0] ? 4'hf : _GEN_14053; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14055 = 8'h18 == _T_689[7:0] ? 4'h0 : _GEN_14054; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14056 = 8'h19 == _T_689[7:0] ? 4'h0 : _GEN_14055; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14057 = 8'h1a == _T_689[7:0] ? 4'h0 : _GEN_14056; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14058 = 8'h1b == _T_689[7:0] ? 4'h0 : _GEN_14057; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14059 = 8'h1c == _T_689[7:0] ? 4'h0 : _GEN_14058; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14060 = 8'h1d == _T_689[7:0] ? 4'h0 : _GEN_14059; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14061 = 8'h1e == _T_689[7:0] ? 4'h0 : _GEN_14060; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14062 = 8'h1f == _T_689[7:0] ? 4'h0 : _GEN_14061; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14063 = 8'h20 == _T_689[7:0] ? 4'hf : _GEN_14062; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14064 = 8'h21 == _T_689[7:0] ? 4'hf : _GEN_14063; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14065 = 8'h22 == _T_689[7:0] ? 4'hf : _GEN_14064; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14066 = 8'h23 == _T_689[7:0] ? 4'hf : _GEN_14065; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14067 = 8'h24 == _T_689[7:0] ? 4'hf : _GEN_14066; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14068 = 8'h25 == _T_689[7:0] ? 4'hf : _GEN_14067; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14069 = 8'h26 == _T_689[7:0] ? 4'hf : _GEN_14068; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14070 = 8'h27 == _T_689[7:0] ? 4'hf : _GEN_14069; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14071 = 8'h28 == _T_689[7:0] ? 4'h0 : _GEN_14070; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14072 = 8'h29 == _T_689[7:0] ? 4'h0 : _GEN_14071; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14073 = 8'h2a == _T_689[7:0] ? 4'h0 : _GEN_14072; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14074 = 8'h2b == _T_689[7:0] ? 4'h0 : _GEN_14073; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14075 = 8'h2c == _T_689[7:0] ? 4'h0 : _GEN_14074; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14076 = 8'h2d == _T_689[7:0] ? 4'h0 : _GEN_14075; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14077 = 8'h2e == _T_689[7:0] ? 4'h0 : _GEN_14076; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14078 = 8'h2f == _T_689[7:0] ? 4'h0 : _GEN_14077; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14079 = 8'h30 == _T_689[7:0] ? 4'hf : _GEN_14078; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14080 = 8'h31 == _T_689[7:0] ? 4'hf : _GEN_14079; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14081 = 8'h32 == _T_689[7:0] ? 4'hf : _GEN_14080; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14082 = 8'h33 == _T_689[7:0] ? 4'hf : _GEN_14081; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14083 = 8'h34 == _T_689[7:0] ? 4'hf : _GEN_14082; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14084 = 8'h35 == _T_689[7:0] ? 4'hf : _GEN_14083; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14085 = 8'h36 == _T_689[7:0] ? 4'hf : _GEN_14084; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14086 = 8'h37 == _T_689[7:0] ? 4'hf : _GEN_14085; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14087 = 8'h38 == _T_689[7:0] ? 4'h0 : _GEN_14086; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14088 = 8'h39 == _T_689[7:0] ? 4'h0 : _GEN_14087; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14089 = 8'h3a == _T_689[7:0] ? 4'h0 : _GEN_14088; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14090 = 8'h3b == _T_689[7:0] ? 4'h0 : _GEN_14089; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14091 = 8'h3c == _T_689[7:0] ? 4'h0 : _GEN_14090; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14092 = 8'h3d == _T_689[7:0] ? 4'h0 : _GEN_14091; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14093 = 8'h3e == _T_689[7:0] ? 4'h0 : _GEN_14092; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14094 = 8'h3f == _T_689[7:0] ? 4'h0 : _GEN_14093; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14095 = 8'h40 == _T_689[7:0] ? 4'hf : _GEN_14094; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14096 = 8'h41 == _T_689[7:0] ? 4'hf : _GEN_14095; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14097 = 8'h42 == _T_689[7:0] ? 4'hf : _GEN_14096; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14098 = 8'h43 == _T_689[7:0] ? 4'hf : _GEN_14097; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14099 = 8'h44 == _T_689[7:0] ? 4'hf : _GEN_14098; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14100 = 8'h45 == _T_689[7:0] ? 4'hf : _GEN_14099; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14101 = 8'h46 == _T_689[7:0] ? 4'hf : _GEN_14100; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14102 = 8'h47 == _T_689[7:0] ? 4'hf : _GEN_14101; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14103 = 8'h48 == _T_689[7:0] ? 4'h0 : _GEN_14102; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14104 = 8'h49 == _T_689[7:0] ? 4'h0 : _GEN_14103; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14105 = 8'h4a == _T_689[7:0] ? 4'h0 : _GEN_14104; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14106 = 8'h4b == _T_689[7:0] ? 4'h0 : _GEN_14105; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14107 = 8'h4c == _T_689[7:0] ? 4'h0 : _GEN_14106; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14108 = 8'h4d == _T_689[7:0] ? 4'h0 : _GEN_14107; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14109 = 8'h4e == _T_689[7:0] ? 4'h0 : _GEN_14108; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14110 = 8'h4f == _T_689[7:0] ? 4'h0 : _GEN_14109; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14111 = 8'h50 == _T_689[7:0] ? 4'hf : _GEN_14110; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14112 = 8'h51 == _T_689[7:0] ? 4'hf : _GEN_14111; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14113 = 8'h52 == _T_689[7:0] ? 4'hf : _GEN_14112; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14114 = 8'h53 == _T_689[7:0] ? 4'hf : _GEN_14113; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14115 = 8'h54 == _T_689[7:0] ? 4'hf : _GEN_14114; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14116 = 8'h55 == _T_689[7:0] ? 4'hf : _GEN_14115; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14117 = 8'h56 == _T_689[7:0] ? 4'hf : _GEN_14116; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14118 = 8'h57 == _T_689[7:0] ? 4'hf : _GEN_14117; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14119 = 8'h58 == _T_689[7:0] ? 4'h0 : _GEN_14118; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14120 = 8'h59 == _T_689[7:0] ? 4'h0 : _GEN_14119; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14121 = 8'h5a == _T_689[7:0] ? 4'h0 : _GEN_14120; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14122 = 8'h5b == _T_689[7:0] ? 4'h0 : _GEN_14121; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14123 = 8'h5c == _T_689[7:0] ? 4'h0 : _GEN_14122; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14124 = 8'h5d == _T_689[7:0] ? 4'h0 : _GEN_14123; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14125 = 8'h5e == _T_689[7:0] ? 4'h0 : _GEN_14124; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14126 = 8'h5f == _T_689[7:0] ? 4'h0 : _GEN_14125; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14127 = 8'h60 == _T_689[7:0] ? 4'h0 : _GEN_14126; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14128 = 8'h61 == _T_689[7:0] ? 4'h0 : _GEN_14127; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14129 = 8'h62 == _T_689[7:0] ? 4'h0 : _GEN_14128; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14130 = 8'h63 == _T_689[7:0] ? 4'h0 : _GEN_14129; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14131 = 8'h64 == _T_689[7:0] ? 4'h0 : _GEN_14130; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14132 = 8'h65 == _T_689[7:0] ? 4'h0 : _GEN_14131; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14133 = 8'h66 == _T_689[7:0] ? 4'h0 : _GEN_14132; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14134 = 8'h67 == _T_689[7:0] ? 4'h0 : _GEN_14133; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14135 = 8'h68 == _T_689[7:0] ? 4'hf : _GEN_14134; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14136 = 8'h69 == _T_689[7:0] ? 4'hf : _GEN_14135; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14137 = 8'h6a == _T_689[7:0] ? 4'hf : _GEN_14136; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14138 = 8'h6b == _T_689[7:0] ? 4'hf : _GEN_14137; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14139 = 8'h6c == _T_689[7:0] ? 4'hf : _GEN_14138; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14140 = 8'h6d == _T_689[7:0] ? 4'hf : _GEN_14139; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14141 = 8'h6e == _T_689[7:0] ? 4'hf : _GEN_14140; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14142 = 8'h6f == _T_689[7:0] ? 4'hf : _GEN_14141; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14143 = 8'h70 == _T_689[7:0] ? 4'h0 : _GEN_14142; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14144 = 8'h71 == _T_689[7:0] ? 4'h0 : _GEN_14143; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14145 = 8'h72 == _T_689[7:0] ? 4'h0 : _GEN_14144; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14146 = 8'h73 == _T_689[7:0] ? 4'h0 : _GEN_14145; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14147 = 8'h74 == _T_689[7:0] ? 4'h0 : _GEN_14146; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14148 = 8'h75 == _T_689[7:0] ? 4'h0 : _GEN_14147; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14149 = 8'h76 == _T_689[7:0] ? 4'h0 : _GEN_14148; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14150 = 8'h77 == _T_689[7:0] ? 4'h0 : _GEN_14149; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14151 = 8'h78 == _T_689[7:0] ? 4'hf : _GEN_14150; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14152 = 8'h79 == _T_689[7:0] ? 4'hf : _GEN_14151; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14153 = 8'h7a == _T_689[7:0] ? 4'hf : _GEN_14152; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14154 = 8'h7b == _T_689[7:0] ? 4'hf : _GEN_14153; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14155 = 8'h7c == _T_689[7:0] ? 4'hf : _GEN_14154; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14156 = 8'h7d == _T_689[7:0] ? 4'hf : _GEN_14155; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14157 = 8'h7e == _T_689[7:0] ? 4'hf : _GEN_14156; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14158 = 8'h7f == _T_689[7:0] ? 4'hf : _GEN_14157; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14159 = 8'h80 == _T_689[7:0] ? 4'h0 : _GEN_14158; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14160 = 8'h81 == _T_689[7:0] ? 4'h0 : _GEN_14159; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14161 = 8'h82 == _T_689[7:0] ? 4'h0 : _GEN_14160; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14162 = 8'h83 == _T_689[7:0] ? 4'h0 : _GEN_14161; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14163 = 8'h84 == _T_689[7:0] ? 4'h0 : _GEN_14162; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14164 = 8'h85 == _T_689[7:0] ? 4'h0 : _GEN_14163; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14165 = 8'h86 == _T_689[7:0] ? 4'h0 : _GEN_14164; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14166 = 8'h87 == _T_689[7:0] ? 4'h0 : _GEN_14165; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14167 = 8'h88 == _T_689[7:0] ? 4'hf : _GEN_14166; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14168 = 8'h89 == _T_689[7:0] ? 4'hf : _GEN_14167; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14169 = 8'h8a == _T_689[7:0] ? 4'hf : _GEN_14168; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14170 = 8'h8b == _T_689[7:0] ? 4'hf : _GEN_14169; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14171 = 8'h8c == _T_689[7:0] ? 4'hf : _GEN_14170; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14172 = 8'h8d == _T_689[7:0] ? 4'hf : _GEN_14171; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14173 = 8'h8e == _T_689[7:0] ? 4'hf : _GEN_14172; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14174 = 8'h8f == _T_689[7:0] ? 4'hf : _GEN_14173; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14175 = 8'h90 == _T_689[7:0] ? 4'h0 : _GEN_14174; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14176 = 8'h91 == _T_689[7:0] ? 4'h0 : _GEN_14175; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14177 = 8'h92 == _T_689[7:0] ? 4'h0 : _GEN_14176; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14178 = 8'h93 == _T_689[7:0] ? 4'h0 : _GEN_14177; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14179 = 8'h94 == _T_689[7:0] ? 4'h0 : _GEN_14178; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14180 = 8'h95 == _T_689[7:0] ? 4'h0 : _GEN_14179; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14181 = 8'h96 == _T_689[7:0] ? 4'h0 : _GEN_14180; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14182 = 8'h97 == _T_689[7:0] ? 4'h0 : _GEN_14181; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14183 = 8'h98 == _T_689[7:0] ? 4'hf : _GEN_14182; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14184 = 8'h99 == _T_689[7:0] ? 4'hf : _GEN_14183; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14185 = 8'h9a == _T_689[7:0] ? 4'hf : _GEN_14184; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14186 = 8'h9b == _T_689[7:0] ? 4'hf : _GEN_14185; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14187 = 8'h9c == _T_689[7:0] ? 4'hf : _GEN_14186; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14188 = 8'h9d == _T_689[7:0] ? 4'hf : _GEN_14187; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14189 = 8'h9e == _T_689[7:0] ? 4'hf : _GEN_14188; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14190 = 8'h9f == _T_689[7:0] ? 4'hf : _GEN_14189; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14191 = 8'ha0 == _T_689[7:0] ? 4'h0 : _GEN_14190; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14192 = 8'ha1 == _T_689[7:0] ? 4'h0 : _GEN_14191; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14193 = 8'ha2 == _T_689[7:0] ? 4'h0 : _GEN_14192; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14194 = 8'ha3 == _T_689[7:0] ? 4'h0 : _GEN_14193; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14195 = 8'ha4 == _T_689[7:0] ? 4'h0 : _GEN_14194; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14196 = 8'ha5 == _T_689[7:0] ? 4'h0 : _GEN_14195; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14197 = 8'ha6 == _T_689[7:0] ? 4'h0 : _GEN_14196; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14198 = 8'ha7 == _T_689[7:0] ? 4'h0 : _GEN_14197; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14199 = 8'ha8 == _T_689[7:0] ? 4'hf : _GEN_14198; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14200 = 8'ha9 == _T_689[7:0] ? 4'hf : _GEN_14199; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14201 = 8'haa == _T_689[7:0] ? 4'hf : _GEN_14200; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14202 = 8'hab == _T_689[7:0] ? 4'hf : _GEN_14201; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14203 = 8'hac == _T_689[7:0] ? 4'hf : _GEN_14202; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14204 = 8'had == _T_689[7:0] ? 4'hf : _GEN_14203; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14205 = 8'hae == _T_689[7:0] ? 4'hf : _GEN_14204; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14206 = 8'haf == _T_689[7:0] ? 4'hf : _GEN_14205; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14207 = 8'hb0 == _T_689[7:0] ? 4'h0 : _GEN_14206; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14208 = 8'hb1 == _T_689[7:0] ? 4'h0 : _GEN_14207; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14209 = 8'hb2 == _T_689[7:0] ? 4'h0 : _GEN_14208; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14210 = 8'hb3 == _T_689[7:0] ? 4'h0 : _GEN_14209; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14211 = 8'hb4 == _T_689[7:0] ? 4'h0 : _GEN_14210; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14212 = 8'hb5 == _T_689[7:0] ? 4'h0 : _GEN_14211; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14213 = 8'hb6 == _T_689[7:0] ? 4'h0 : _GEN_14212; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14214 = 8'hb7 == _T_689[7:0] ? 4'h0 : _GEN_14213; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14215 = 8'hb8 == _T_689[7:0] ? 4'hf : _GEN_14214; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14216 = 8'hb9 == _T_689[7:0] ? 4'hf : _GEN_14215; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14217 = 8'hba == _T_689[7:0] ? 4'hf : _GEN_14216; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14218 = 8'hbb == _T_689[7:0] ? 4'hf : _GEN_14217; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14219 = 8'hbc == _T_689[7:0] ? 4'hf : _GEN_14218; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14220 = 8'hbd == _T_689[7:0] ? 4'hf : _GEN_14219; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14221 = 8'hbe == _T_689[7:0] ? 4'hf : _GEN_14220; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14222 = 8'hbf == _T_689[7:0] ? 4'hf : _GEN_14221; // @[Filter.scala 165:86]
  wire [4:0] _GEN_19142 = {{1'd0}, _GEN_14222}; // @[Filter.scala 165:86]
  wire [8:0] _T_691 = _GEN_19142 * 5'h14; // @[Filter.scala 165:86]
  wire [3:0] _GEN_14319 = 8'h60 == _T_689[7:0] ? 4'hf : 4'h0; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14320 = 8'h61 == _T_689[7:0] ? 4'hf : _GEN_14319; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14321 = 8'h62 == _T_689[7:0] ? 4'hf : _GEN_14320; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14322 = 8'h63 == _T_689[7:0] ? 4'hf : _GEN_14321; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14323 = 8'h64 == _T_689[7:0] ? 4'hf : _GEN_14322; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14324 = 8'h65 == _T_689[7:0] ? 4'hf : _GEN_14323; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14325 = 8'h66 == _T_689[7:0] ? 4'hf : _GEN_14324; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14326 = 8'h67 == _T_689[7:0] ? 4'hf : _GEN_14325; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14327 = 8'h68 == _T_689[7:0] ? 4'hf : _GEN_14326; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14328 = 8'h69 == _T_689[7:0] ? 4'hf : _GEN_14327; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14329 = 8'h6a == _T_689[7:0] ? 4'hf : _GEN_14328; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14330 = 8'h6b == _T_689[7:0] ? 4'hf : _GEN_14329; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14331 = 8'h6c == _T_689[7:0] ? 4'hf : _GEN_14330; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14332 = 8'h6d == _T_689[7:0] ? 4'hf : _GEN_14331; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14333 = 8'h6e == _T_689[7:0] ? 4'hf : _GEN_14332; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14334 = 8'h6f == _T_689[7:0] ? 4'hf : _GEN_14333; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14335 = 8'h70 == _T_689[7:0] ? 4'hf : _GEN_14334; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14336 = 8'h71 == _T_689[7:0] ? 4'hf : _GEN_14335; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14337 = 8'h72 == _T_689[7:0] ? 4'hf : _GEN_14336; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14338 = 8'h73 == _T_689[7:0] ? 4'hf : _GEN_14337; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14339 = 8'h74 == _T_689[7:0] ? 4'hf : _GEN_14338; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14340 = 8'h75 == _T_689[7:0] ? 4'hf : _GEN_14339; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14341 = 8'h76 == _T_689[7:0] ? 4'hf : _GEN_14340; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14342 = 8'h77 == _T_689[7:0] ? 4'hf : _GEN_14341; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14343 = 8'h78 == _T_689[7:0] ? 4'hf : _GEN_14342; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14344 = 8'h79 == _T_689[7:0] ? 4'hf : _GEN_14343; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14345 = 8'h7a == _T_689[7:0] ? 4'hf : _GEN_14344; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14346 = 8'h7b == _T_689[7:0] ? 4'hf : _GEN_14345; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14347 = 8'h7c == _T_689[7:0] ? 4'hf : _GEN_14346; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14348 = 8'h7d == _T_689[7:0] ? 4'hf : _GEN_14347; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14349 = 8'h7e == _T_689[7:0] ? 4'hf : _GEN_14348; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14350 = 8'h7f == _T_689[7:0] ? 4'hf : _GEN_14349; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14351 = 8'h80 == _T_689[7:0] ? 4'hf : _GEN_14350; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14352 = 8'h81 == _T_689[7:0] ? 4'hf : _GEN_14351; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14353 = 8'h82 == _T_689[7:0] ? 4'hf : _GEN_14352; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14354 = 8'h83 == _T_689[7:0] ? 4'hf : _GEN_14353; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14355 = 8'h84 == _T_689[7:0] ? 4'hf : _GEN_14354; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14356 = 8'h85 == _T_689[7:0] ? 4'hf : _GEN_14355; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14357 = 8'h86 == _T_689[7:0] ? 4'hf : _GEN_14356; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14358 = 8'h87 == _T_689[7:0] ? 4'hf : _GEN_14357; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14359 = 8'h88 == _T_689[7:0] ? 4'hf : _GEN_14358; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14360 = 8'h89 == _T_689[7:0] ? 4'hf : _GEN_14359; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14361 = 8'h8a == _T_689[7:0] ? 4'hf : _GEN_14360; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14362 = 8'h8b == _T_689[7:0] ? 4'hf : _GEN_14361; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14363 = 8'h8c == _T_689[7:0] ? 4'hf : _GEN_14362; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14364 = 8'h8d == _T_689[7:0] ? 4'hf : _GEN_14363; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14365 = 8'h8e == _T_689[7:0] ? 4'hf : _GEN_14364; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14366 = 8'h8f == _T_689[7:0] ? 4'hf : _GEN_14365; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14367 = 8'h90 == _T_689[7:0] ? 4'hf : _GEN_14366; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14368 = 8'h91 == _T_689[7:0] ? 4'hf : _GEN_14367; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14369 = 8'h92 == _T_689[7:0] ? 4'hf : _GEN_14368; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14370 = 8'h93 == _T_689[7:0] ? 4'hf : _GEN_14369; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14371 = 8'h94 == _T_689[7:0] ? 4'hf : _GEN_14370; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14372 = 8'h95 == _T_689[7:0] ? 4'hf : _GEN_14371; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14373 = 8'h96 == _T_689[7:0] ? 4'hf : _GEN_14372; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14374 = 8'h97 == _T_689[7:0] ? 4'hf : _GEN_14373; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14375 = 8'h98 == _T_689[7:0] ? 4'hf : _GEN_14374; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14376 = 8'h99 == _T_689[7:0] ? 4'hf : _GEN_14375; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14377 = 8'h9a == _T_689[7:0] ? 4'hf : _GEN_14376; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14378 = 8'h9b == _T_689[7:0] ? 4'hf : _GEN_14377; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14379 = 8'h9c == _T_689[7:0] ? 4'hf : _GEN_14378; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14380 = 8'h9d == _T_689[7:0] ? 4'hf : _GEN_14379; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14381 = 8'h9e == _T_689[7:0] ? 4'hf : _GEN_14380; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14382 = 8'h9f == _T_689[7:0] ? 4'hf : _GEN_14381; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14383 = 8'ha0 == _T_689[7:0] ? 4'hf : _GEN_14382; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14384 = 8'ha1 == _T_689[7:0] ? 4'hf : _GEN_14383; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14385 = 8'ha2 == _T_689[7:0] ? 4'hf : _GEN_14384; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14386 = 8'ha3 == _T_689[7:0] ? 4'hf : _GEN_14385; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14387 = 8'ha4 == _T_689[7:0] ? 4'hf : _GEN_14386; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14388 = 8'ha5 == _T_689[7:0] ? 4'hf : _GEN_14387; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14389 = 8'ha6 == _T_689[7:0] ? 4'hf : _GEN_14388; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14390 = 8'ha7 == _T_689[7:0] ? 4'hf : _GEN_14389; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14391 = 8'ha8 == _T_689[7:0] ? 4'hf : _GEN_14390; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14392 = 8'ha9 == _T_689[7:0] ? 4'hf : _GEN_14391; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14393 = 8'haa == _T_689[7:0] ? 4'hf : _GEN_14392; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14394 = 8'hab == _T_689[7:0] ? 4'hf : _GEN_14393; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14395 = 8'hac == _T_689[7:0] ? 4'hf : _GEN_14394; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14396 = 8'had == _T_689[7:0] ? 4'hf : _GEN_14395; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14397 = 8'hae == _T_689[7:0] ? 4'hf : _GEN_14396; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14398 = 8'haf == _T_689[7:0] ? 4'hf : _GEN_14397; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14399 = 8'hb0 == _T_689[7:0] ? 4'hf : _GEN_14398; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14400 = 8'hb1 == _T_689[7:0] ? 4'hf : _GEN_14399; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14401 = 8'hb2 == _T_689[7:0] ? 4'hf : _GEN_14400; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14402 = 8'hb3 == _T_689[7:0] ? 4'hf : _GEN_14401; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14403 = 8'hb4 == _T_689[7:0] ? 4'hf : _GEN_14402; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14404 = 8'hb5 == _T_689[7:0] ? 4'hf : _GEN_14403; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14405 = 8'hb6 == _T_689[7:0] ? 4'hf : _GEN_14404; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14406 = 8'hb7 == _T_689[7:0] ? 4'hf : _GEN_14405; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14407 = 8'hb8 == _T_689[7:0] ? 4'hf : _GEN_14406; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14408 = 8'hb9 == _T_689[7:0] ? 4'hf : _GEN_14407; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14409 = 8'hba == _T_689[7:0] ? 4'hf : _GEN_14408; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14410 = 8'hbb == _T_689[7:0] ? 4'hf : _GEN_14409; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14411 = 8'hbc == _T_689[7:0] ? 4'hf : _GEN_14410; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14412 = 8'hbd == _T_689[7:0] ? 4'hf : _GEN_14411; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14413 = 8'hbe == _T_689[7:0] ? 4'hf : _GEN_14412; // @[Filter.scala 165:126]
  wire [3:0] _GEN_14414 = 8'hbf == _T_689[7:0] ? 4'hf : _GEN_14413; // @[Filter.scala 165:126]
  wire [6:0] _GEN_19144 = {{3'd0}, _GEN_14414}; // @[Filter.scala 165:126]
  wire [10:0] _T_696 = _GEN_19144 * 7'h46; // @[Filter.scala 165:126]
  wire [10:0] _GEN_19145 = {{2'd0}, _T_691}; // @[Filter.scala 165:93]
  wire [10:0] _T_698 = _GEN_19145 + _T_696; // @[Filter.scala 165:93]
  wire [3:0] _GEN_14423 = 8'h8 == _T_689[7:0] ? 4'hf : 4'h0; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14424 = 8'h9 == _T_689[7:0] ? 4'hf : _GEN_14423; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14425 = 8'ha == _T_689[7:0] ? 4'hf : _GEN_14424; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14426 = 8'hb == _T_689[7:0] ? 4'hf : _GEN_14425; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14427 = 8'hc == _T_689[7:0] ? 4'hf : _GEN_14426; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14428 = 8'hd == _T_689[7:0] ? 4'hf : _GEN_14427; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14429 = 8'he == _T_689[7:0] ? 4'hf : _GEN_14428; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14430 = 8'hf == _T_689[7:0] ? 4'hf : _GEN_14429; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14431 = 8'h10 == _T_689[7:0] ? 4'h0 : _GEN_14430; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14432 = 8'h11 == _T_689[7:0] ? 4'h0 : _GEN_14431; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14433 = 8'h12 == _T_689[7:0] ? 4'h0 : _GEN_14432; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14434 = 8'h13 == _T_689[7:0] ? 4'h0 : _GEN_14433; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14435 = 8'h14 == _T_689[7:0] ? 4'h0 : _GEN_14434; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14436 = 8'h15 == _T_689[7:0] ? 4'h0 : _GEN_14435; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14437 = 8'h16 == _T_689[7:0] ? 4'h0 : _GEN_14436; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14438 = 8'h17 == _T_689[7:0] ? 4'h0 : _GEN_14437; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14439 = 8'h18 == _T_689[7:0] ? 4'hf : _GEN_14438; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14440 = 8'h19 == _T_689[7:0] ? 4'hf : _GEN_14439; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14441 = 8'h1a == _T_689[7:0] ? 4'hf : _GEN_14440; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14442 = 8'h1b == _T_689[7:0] ? 4'hf : _GEN_14441; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14443 = 8'h1c == _T_689[7:0] ? 4'hf : _GEN_14442; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14444 = 8'h1d == _T_689[7:0] ? 4'hf : _GEN_14443; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14445 = 8'h1e == _T_689[7:0] ? 4'hf : _GEN_14444; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14446 = 8'h1f == _T_689[7:0] ? 4'hf : _GEN_14445; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14447 = 8'h20 == _T_689[7:0] ? 4'h0 : _GEN_14446; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14448 = 8'h21 == _T_689[7:0] ? 4'h0 : _GEN_14447; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14449 = 8'h22 == _T_689[7:0] ? 4'h0 : _GEN_14448; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14450 = 8'h23 == _T_689[7:0] ? 4'h0 : _GEN_14449; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14451 = 8'h24 == _T_689[7:0] ? 4'h0 : _GEN_14450; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14452 = 8'h25 == _T_689[7:0] ? 4'h0 : _GEN_14451; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14453 = 8'h26 == _T_689[7:0] ? 4'h0 : _GEN_14452; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14454 = 8'h27 == _T_689[7:0] ? 4'h0 : _GEN_14453; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14455 = 8'h28 == _T_689[7:0] ? 4'hf : _GEN_14454; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14456 = 8'h29 == _T_689[7:0] ? 4'hf : _GEN_14455; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14457 = 8'h2a == _T_689[7:0] ? 4'hf : _GEN_14456; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14458 = 8'h2b == _T_689[7:0] ? 4'hf : _GEN_14457; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14459 = 8'h2c == _T_689[7:0] ? 4'hf : _GEN_14458; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14460 = 8'h2d == _T_689[7:0] ? 4'hf : _GEN_14459; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14461 = 8'h2e == _T_689[7:0] ? 4'hf : _GEN_14460; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14462 = 8'h2f == _T_689[7:0] ? 4'hf : _GEN_14461; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14463 = 8'h30 == _T_689[7:0] ? 4'h0 : _GEN_14462; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14464 = 8'h31 == _T_689[7:0] ? 4'h0 : _GEN_14463; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14465 = 8'h32 == _T_689[7:0] ? 4'h0 : _GEN_14464; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14466 = 8'h33 == _T_689[7:0] ? 4'h0 : _GEN_14465; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14467 = 8'h34 == _T_689[7:0] ? 4'h0 : _GEN_14466; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14468 = 8'h35 == _T_689[7:0] ? 4'h0 : _GEN_14467; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14469 = 8'h36 == _T_689[7:0] ? 4'h0 : _GEN_14468; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14470 = 8'h37 == _T_689[7:0] ? 4'h0 : _GEN_14469; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14471 = 8'h38 == _T_689[7:0] ? 4'hf : _GEN_14470; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14472 = 8'h39 == _T_689[7:0] ? 4'hf : _GEN_14471; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14473 = 8'h3a == _T_689[7:0] ? 4'hf : _GEN_14472; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14474 = 8'h3b == _T_689[7:0] ? 4'hf : _GEN_14473; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14475 = 8'h3c == _T_689[7:0] ? 4'hf : _GEN_14474; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14476 = 8'h3d == _T_689[7:0] ? 4'hf : _GEN_14475; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14477 = 8'h3e == _T_689[7:0] ? 4'hf : _GEN_14476; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14478 = 8'h3f == _T_689[7:0] ? 4'hf : _GEN_14477; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14479 = 8'h40 == _T_689[7:0] ? 4'h0 : _GEN_14478; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14480 = 8'h41 == _T_689[7:0] ? 4'h0 : _GEN_14479; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14481 = 8'h42 == _T_689[7:0] ? 4'h0 : _GEN_14480; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14482 = 8'h43 == _T_689[7:0] ? 4'h0 : _GEN_14481; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14483 = 8'h44 == _T_689[7:0] ? 4'h0 : _GEN_14482; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14484 = 8'h45 == _T_689[7:0] ? 4'h0 : _GEN_14483; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14485 = 8'h46 == _T_689[7:0] ? 4'h0 : _GEN_14484; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14486 = 8'h47 == _T_689[7:0] ? 4'h0 : _GEN_14485; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14487 = 8'h48 == _T_689[7:0] ? 4'hf : _GEN_14486; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14488 = 8'h49 == _T_689[7:0] ? 4'hf : _GEN_14487; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14489 = 8'h4a == _T_689[7:0] ? 4'hf : _GEN_14488; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14490 = 8'h4b == _T_689[7:0] ? 4'hf : _GEN_14489; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14491 = 8'h4c == _T_689[7:0] ? 4'hf : _GEN_14490; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14492 = 8'h4d == _T_689[7:0] ? 4'hf : _GEN_14491; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14493 = 8'h4e == _T_689[7:0] ? 4'hf : _GEN_14492; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14494 = 8'h4f == _T_689[7:0] ? 4'hf : _GEN_14493; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14495 = 8'h50 == _T_689[7:0] ? 4'h0 : _GEN_14494; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14496 = 8'h51 == _T_689[7:0] ? 4'h0 : _GEN_14495; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14497 = 8'h52 == _T_689[7:0] ? 4'h0 : _GEN_14496; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14498 = 8'h53 == _T_689[7:0] ? 4'h0 : _GEN_14497; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14499 = 8'h54 == _T_689[7:0] ? 4'h0 : _GEN_14498; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14500 = 8'h55 == _T_689[7:0] ? 4'h0 : _GEN_14499; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14501 = 8'h56 == _T_689[7:0] ? 4'h0 : _GEN_14500; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14502 = 8'h57 == _T_689[7:0] ? 4'h0 : _GEN_14501; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14503 = 8'h58 == _T_689[7:0] ? 4'hf : _GEN_14502; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14504 = 8'h59 == _T_689[7:0] ? 4'hf : _GEN_14503; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14505 = 8'h5a == _T_689[7:0] ? 4'hf : _GEN_14504; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14506 = 8'h5b == _T_689[7:0] ? 4'hf : _GEN_14505; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14507 = 8'h5c == _T_689[7:0] ? 4'hf : _GEN_14506; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14508 = 8'h5d == _T_689[7:0] ? 4'hf : _GEN_14507; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14509 = 8'h5e == _T_689[7:0] ? 4'hf : _GEN_14508; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14510 = 8'h5f == _T_689[7:0] ? 4'hf : _GEN_14509; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14511 = 8'h60 == _T_689[7:0] ? 4'h0 : _GEN_14510; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14512 = 8'h61 == _T_689[7:0] ? 4'h0 : _GEN_14511; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14513 = 8'h62 == _T_689[7:0] ? 4'h0 : _GEN_14512; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14514 = 8'h63 == _T_689[7:0] ? 4'h0 : _GEN_14513; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14515 = 8'h64 == _T_689[7:0] ? 4'h0 : _GEN_14514; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14516 = 8'h65 == _T_689[7:0] ? 4'h0 : _GEN_14515; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14517 = 8'h66 == _T_689[7:0] ? 4'h0 : _GEN_14516; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14518 = 8'h67 == _T_689[7:0] ? 4'h0 : _GEN_14517; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14519 = 8'h68 == _T_689[7:0] ? 4'hf : _GEN_14518; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14520 = 8'h69 == _T_689[7:0] ? 4'hf : _GEN_14519; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14521 = 8'h6a == _T_689[7:0] ? 4'hf : _GEN_14520; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14522 = 8'h6b == _T_689[7:0] ? 4'hf : _GEN_14521; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14523 = 8'h6c == _T_689[7:0] ? 4'hf : _GEN_14522; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14524 = 8'h6d == _T_689[7:0] ? 4'hf : _GEN_14523; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14525 = 8'h6e == _T_689[7:0] ? 4'hf : _GEN_14524; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14526 = 8'h6f == _T_689[7:0] ? 4'hf : _GEN_14525; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14527 = 8'h70 == _T_689[7:0] ? 4'h0 : _GEN_14526; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14528 = 8'h71 == _T_689[7:0] ? 4'h0 : _GEN_14527; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14529 = 8'h72 == _T_689[7:0] ? 4'h0 : _GEN_14528; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14530 = 8'h73 == _T_689[7:0] ? 4'h0 : _GEN_14529; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14531 = 8'h74 == _T_689[7:0] ? 4'h0 : _GEN_14530; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14532 = 8'h75 == _T_689[7:0] ? 4'h0 : _GEN_14531; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14533 = 8'h76 == _T_689[7:0] ? 4'h0 : _GEN_14532; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14534 = 8'h77 == _T_689[7:0] ? 4'h0 : _GEN_14533; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14535 = 8'h78 == _T_689[7:0] ? 4'hf : _GEN_14534; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14536 = 8'h79 == _T_689[7:0] ? 4'hf : _GEN_14535; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14537 = 8'h7a == _T_689[7:0] ? 4'hf : _GEN_14536; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14538 = 8'h7b == _T_689[7:0] ? 4'hf : _GEN_14537; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14539 = 8'h7c == _T_689[7:0] ? 4'hf : _GEN_14538; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14540 = 8'h7d == _T_689[7:0] ? 4'hf : _GEN_14539; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14541 = 8'h7e == _T_689[7:0] ? 4'hf : _GEN_14540; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14542 = 8'h7f == _T_689[7:0] ? 4'hf : _GEN_14541; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14543 = 8'h80 == _T_689[7:0] ? 4'h0 : _GEN_14542; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14544 = 8'h81 == _T_689[7:0] ? 4'h0 : _GEN_14543; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14545 = 8'h82 == _T_689[7:0] ? 4'h0 : _GEN_14544; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14546 = 8'h83 == _T_689[7:0] ? 4'h0 : _GEN_14545; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14547 = 8'h84 == _T_689[7:0] ? 4'h0 : _GEN_14546; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14548 = 8'h85 == _T_689[7:0] ? 4'h0 : _GEN_14547; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14549 = 8'h86 == _T_689[7:0] ? 4'h0 : _GEN_14548; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14550 = 8'h87 == _T_689[7:0] ? 4'h0 : _GEN_14549; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14551 = 8'h88 == _T_689[7:0] ? 4'hf : _GEN_14550; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14552 = 8'h89 == _T_689[7:0] ? 4'hf : _GEN_14551; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14553 = 8'h8a == _T_689[7:0] ? 4'hf : _GEN_14552; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14554 = 8'h8b == _T_689[7:0] ? 4'hf : _GEN_14553; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14555 = 8'h8c == _T_689[7:0] ? 4'hf : _GEN_14554; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14556 = 8'h8d == _T_689[7:0] ? 4'hf : _GEN_14555; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14557 = 8'h8e == _T_689[7:0] ? 4'hf : _GEN_14556; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14558 = 8'h8f == _T_689[7:0] ? 4'hf : _GEN_14557; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14559 = 8'h90 == _T_689[7:0] ? 4'h0 : _GEN_14558; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14560 = 8'h91 == _T_689[7:0] ? 4'h0 : _GEN_14559; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14561 = 8'h92 == _T_689[7:0] ? 4'h0 : _GEN_14560; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14562 = 8'h93 == _T_689[7:0] ? 4'h0 : _GEN_14561; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14563 = 8'h94 == _T_689[7:0] ? 4'h0 : _GEN_14562; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14564 = 8'h95 == _T_689[7:0] ? 4'h0 : _GEN_14563; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14565 = 8'h96 == _T_689[7:0] ? 4'h0 : _GEN_14564; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14566 = 8'h97 == _T_689[7:0] ? 4'h0 : _GEN_14565; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14567 = 8'h98 == _T_689[7:0] ? 4'hf : _GEN_14566; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14568 = 8'h99 == _T_689[7:0] ? 4'hf : _GEN_14567; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14569 = 8'h9a == _T_689[7:0] ? 4'hf : _GEN_14568; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14570 = 8'h9b == _T_689[7:0] ? 4'hf : _GEN_14569; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14571 = 8'h9c == _T_689[7:0] ? 4'hf : _GEN_14570; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14572 = 8'h9d == _T_689[7:0] ? 4'hf : _GEN_14571; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14573 = 8'h9e == _T_689[7:0] ? 4'hf : _GEN_14572; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14574 = 8'h9f == _T_689[7:0] ? 4'hf : _GEN_14573; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14575 = 8'ha0 == _T_689[7:0] ? 4'h0 : _GEN_14574; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14576 = 8'ha1 == _T_689[7:0] ? 4'h0 : _GEN_14575; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14577 = 8'ha2 == _T_689[7:0] ? 4'h0 : _GEN_14576; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14578 = 8'ha3 == _T_689[7:0] ? 4'h0 : _GEN_14577; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14579 = 8'ha4 == _T_689[7:0] ? 4'h0 : _GEN_14578; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14580 = 8'ha5 == _T_689[7:0] ? 4'h0 : _GEN_14579; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14581 = 8'ha6 == _T_689[7:0] ? 4'h0 : _GEN_14580; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14582 = 8'ha7 == _T_689[7:0] ? 4'h0 : _GEN_14581; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14583 = 8'ha8 == _T_689[7:0] ? 4'hf : _GEN_14582; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14584 = 8'ha9 == _T_689[7:0] ? 4'hf : _GEN_14583; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14585 = 8'haa == _T_689[7:0] ? 4'hf : _GEN_14584; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14586 = 8'hab == _T_689[7:0] ? 4'hf : _GEN_14585; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14587 = 8'hac == _T_689[7:0] ? 4'hf : _GEN_14586; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14588 = 8'had == _T_689[7:0] ? 4'hf : _GEN_14587; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14589 = 8'hae == _T_689[7:0] ? 4'hf : _GEN_14588; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14590 = 8'haf == _T_689[7:0] ? 4'hf : _GEN_14589; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14591 = 8'hb0 == _T_689[7:0] ? 4'h0 : _GEN_14590; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14592 = 8'hb1 == _T_689[7:0] ? 4'h0 : _GEN_14591; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14593 = 8'hb2 == _T_689[7:0] ? 4'h0 : _GEN_14592; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14594 = 8'hb3 == _T_689[7:0] ? 4'h0 : _GEN_14593; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14595 = 8'hb4 == _T_689[7:0] ? 4'h0 : _GEN_14594; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14596 = 8'hb5 == _T_689[7:0] ? 4'h0 : _GEN_14595; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14597 = 8'hb6 == _T_689[7:0] ? 4'h0 : _GEN_14596; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14598 = 8'hb7 == _T_689[7:0] ? 4'h0 : _GEN_14597; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14599 = 8'hb8 == _T_689[7:0] ? 4'hf : _GEN_14598; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14600 = 8'hb9 == _T_689[7:0] ? 4'hf : _GEN_14599; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14601 = 8'hba == _T_689[7:0] ? 4'hf : _GEN_14600; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14602 = 8'hbb == _T_689[7:0] ? 4'hf : _GEN_14601; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14603 = 8'hbc == _T_689[7:0] ? 4'hf : _GEN_14602; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14604 = 8'hbd == _T_689[7:0] ? 4'hf : _GEN_14603; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14605 = 8'hbe == _T_689[7:0] ? 4'hf : _GEN_14604; // @[Filter.scala 165:166]
  wire [3:0] _GEN_14606 = 8'hbf == _T_689[7:0] ? 4'hf : _GEN_14605; // @[Filter.scala 165:166]
  wire [7:0] _T_703 = _GEN_14606 * 4'ha; // @[Filter.scala 165:166]
  wire [10:0] _GEN_19147 = {{3'd0}, _T_703}; // @[Filter.scala 165:133]
  wire [10:0] _T_705 = _T_698 + _GEN_19147; // @[Filter.scala 165:133]
  wire [10:0] _T_706 = _T_705 / 11'h64; // @[Filter.scala 165:174]
  wire [10:0] _GEN_14799 = io_SPI_distort ? _T_706 : {{7'd0}, _GEN_14222}; // @[Filter.scala 164:35]
  wire [10:0] _GEN_14800 = _T_686 ? 11'h0 : _GEN_14799; // @[Filter.scala 162:80]
  wire [10:0] _GEN_15569 = io_SPI_distort ? _T_706 : {{7'd0}, _GEN_14414}; // @[Filter.scala 164:35]
  wire [10:0] _GEN_15570 = _T_686 ? 11'h0 : _GEN_15569; // @[Filter.scala 162:80]
  wire [10:0] _GEN_16339 = io_SPI_distort ? _T_706 : {{7'd0}, _GEN_14606}; // @[Filter.scala 164:35]
  wire [10:0] _GEN_16340 = _T_686 ? 11'h0 : _GEN_16339; // @[Filter.scala 162:80]
  wire [31:0] _T_774 = pixelIndex + 32'h7; // @[Filter.scala 158:31]
  wire [31:0] _GEN_56 = _T_774 % 32'h10; // @[Filter.scala 158:38]
  wire [4:0] _T_775 = _GEN_56[4:0]; // @[Filter.scala 158:38]
  wire [4:0] _T_777 = _T_775 + _GEN_18983; // @[Filter.scala 158:53]
  wire [4:0] _T_779 = _T_777 - 5'h1; // @[Filter.scala 158:69]
  wire [31:0] _T_782 = _T_774 / 32'h10; // @[Filter.scala 159:38]
  wire [31:0] _T_784 = _T_782 + _GEN_18984; // @[Filter.scala 159:53]
  wire [31:0] _T_786 = _T_784 - 32'h1; // @[Filter.scala 159:69]
  wire  _T_788 = _T_779 >= 5'h10; // @[Filter.scala 162:31]
  wire  _T_792 = _T_786 >= 32'hc; // @[Filter.scala 162:63]
  wire  _T_793 = _T_788 | _T_792; // @[Filter.scala 162:58]
  wire [36:0] _T_794 = _T_786 * 32'h10; // @[Filter.scala 165:66]
  wire [36:0] _GEN_19167 = {{32'd0}, _T_779}; // @[Filter.scala 165:81]
  wire [36:0] _T_796 = _T_794 + _GEN_19167; // @[Filter.scala 165:81]
  wire [3:0] _GEN_16349 = 8'h8 == _T_796[7:0] ? 4'h0 : 4'hf; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16350 = 8'h9 == _T_796[7:0] ? 4'h0 : _GEN_16349; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16351 = 8'ha == _T_796[7:0] ? 4'h0 : _GEN_16350; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16352 = 8'hb == _T_796[7:0] ? 4'h0 : _GEN_16351; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16353 = 8'hc == _T_796[7:0] ? 4'h0 : _GEN_16352; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16354 = 8'hd == _T_796[7:0] ? 4'h0 : _GEN_16353; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16355 = 8'he == _T_796[7:0] ? 4'h0 : _GEN_16354; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16356 = 8'hf == _T_796[7:0] ? 4'h0 : _GEN_16355; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16357 = 8'h10 == _T_796[7:0] ? 4'hf : _GEN_16356; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16358 = 8'h11 == _T_796[7:0] ? 4'hf : _GEN_16357; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16359 = 8'h12 == _T_796[7:0] ? 4'hf : _GEN_16358; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16360 = 8'h13 == _T_796[7:0] ? 4'hf : _GEN_16359; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16361 = 8'h14 == _T_796[7:0] ? 4'hf : _GEN_16360; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16362 = 8'h15 == _T_796[7:0] ? 4'hf : _GEN_16361; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16363 = 8'h16 == _T_796[7:0] ? 4'hf : _GEN_16362; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16364 = 8'h17 == _T_796[7:0] ? 4'hf : _GEN_16363; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16365 = 8'h18 == _T_796[7:0] ? 4'h0 : _GEN_16364; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16366 = 8'h19 == _T_796[7:0] ? 4'h0 : _GEN_16365; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16367 = 8'h1a == _T_796[7:0] ? 4'h0 : _GEN_16366; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16368 = 8'h1b == _T_796[7:0] ? 4'h0 : _GEN_16367; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16369 = 8'h1c == _T_796[7:0] ? 4'h0 : _GEN_16368; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16370 = 8'h1d == _T_796[7:0] ? 4'h0 : _GEN_16369; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16371 = 8'h1e == _T_796[7:0] ? 4'h0 : _GEN_16370; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16372 = 8'h1f == _T_796[7:0] ? 4'h0 : _GEN_16371; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16373 = 8'h20 == _T_796[7:0] ? 4'hf : _GEN_16372; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16374 = 8'h21 == _T_796[7:0] ? 4'hf : _GEN_16373; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16375 = 8'h22 == _T_796[7:0] ? 4'hf : _GEN_16374; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16376 = 8'h23 == _T_796[7:0] ? 4'hf : _GEN_16375; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16377 = 8'h24 == _T_796[7:0] ? 4'hf : _GEN_16376; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16378 = 8'h25 == _T_796[7:0] ? 4'hf : _GEN_16377; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16379 = 8'h26 == _T_796[7:0] ? 4'hf : _GEN_16378; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16380 = 8'h27 == _T_796[7:0] ? 4'hf : _GEN_16379; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16381 = 8'h28 == _T_796[7:0] ? 4'h0 : _GEN_16380; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16382 = 8'h29 == _T_796[7:0] ? 4'h0 : _GEN_16381; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16383 = 8'h2a == _T_796[7:0] ? 4'h0 : _GEN_16382; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16384 = 8'h2b == _T_796[7:0] ? 4'h0 : _GEN_16383; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16385 = 8'h2c == _T_796[7:0] ? 4'h0 : _GEN_16384; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16386 = 8'h2d == _T_796[7:0] ? 4'h0 : _GEN_16385; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16387 = 8'h2e == _T_796[7:0] ? 4'h0 : _GEN_16386; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16388 = 8'h2f == _T_796[7:0] ? 4'h0 : _GEN_16387; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16389 = 8'h30 == _T_796[7:0] ? 4'hf : _GEN_16388; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16390 = 8'h31 == _T_796[7:0] ? 4'hf : _GEN_16389; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16391 = 8'h32 == _T_796[7:0] ? 4'hf : _GEN_16390; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16392 = 8'h33 == _T_796[7:0] ? 4'hf : _GEN_16391; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16393 = 8'h34 == _T_796[7:0] ? 4'hf : _GEN_16392; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16394 = 8'h35 == _T_796[7:0] ? 4'hf : _GEN_16393; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16395 = 8'h36 == _T_796[7:0] ? 4'hf : _GEN_16394; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16396 = 8'h37 == _T_796[7:0] ? 4'hf : _GEN_16395; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16397 = 8'h38 == _T_796[7:0] ? 4'h0 : _GEN_16396; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16398 = 8'h39 == _T_796[7:0] ? 4'h0 : _GEN_16397; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16399 = 8'h3a == _T_796[7:0] ? 4'h0 : _GEN_16398; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16400 = 8'h3b == _T_796[7:0] ? 4'h0 : _GEN_16399; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16401 = 8'h3c == _T_796[7:0] ? 4'h0 : _GEN_16400; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16402 = 8'h3d == _T_796[7:0] ? 4'h0 : _GEN_16401; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16403 = 8'h3e == _T_796[7:0] ? 4'h0 : _GEN_16402; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16404 = 8'h3f == _T_796[7:0] ? 4'h0 : _GEN_16403; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16405 = 8'h40 == _T_796[7:0] ? 4'hf : _GEN_16404; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16406 = 8'h41 == _T_796[7:0] ? 4'hf : _GEN_16405; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16407 = 8'h42 == _T_796[7:0] ? 4'hf : _GEN_16406; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16408 = 8'h43 == _T_796[7:0] ? 4'hf : _GEN_16407; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16409 = 8'h44 == _T_796[7:0] ? 4'hf : _GEN_16408; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16410 = 8'h45 == _T_796[7:0] ? 4'hf : _GEN_16409; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16411 = 8'h46 == _T_796[7:0] ? 4'hf : _GEN_16410; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16412 = 8'h47 == _T_796[7:0] ? 4'hf : _GEN_16411; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16413 = 8'h48 == _T_796[7:0] ? 4'h0 : _GEN_16412; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16414 = 8'h49 == _T_796[7:0] ? 4'h0 : _GEN_16413; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16415 = 8'h4a == _T_796[7:0] ? 4'h0 : _GEN_16414; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16416 = 8'h4b == _T_796[7:0] ? 4'h0 : _GEN_16415; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16417 = 8'h4c == _T_796[7:0] ? 4'h0 : _GEN_16416; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16418 = 8'h4d == _T_796[7:0] ? 4'h0 : _GEN_16417; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16419 = 8'h4e == _T_796[7:0] ? 4'h0 : _GEN_16418; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16420 = 8'h4f == _T_796[7:0] ? 4'h0 : _GEN_16419; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16421 = 8'h50 == _T_796[7:0] ? 4'hf : _GEN_16420; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16422 = 8'h51 == _T_796[7:0] ? 4'hf : _GEN_16421; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16423 = 8'h52 == _T_796[7:0] ? 4'hf : _GEN_16422; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16424 = 8'h53 == _T_796[7:0] ? 4'hf : _GEN_16423; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16425 = 8'h54 == _T_796[7:0] ? 4'hf : _GEN_16424; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16426 = 8'h55 == _T_796[7:0] ? 4'hf : _GEN_16425; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16427 = 8'h56 == _T_796[7:0] ? 4'hf : _GEN_16426; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16428 = 8'h57 == _T_796[7:0] ? 4'hf : _GEN_16427; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16429 = 8'h58 == _T_796[7:0] ? 4'h0 : _GEN_16428; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16430 = 8'h59 == _T_796[7:0] ? 4'h0 : _GEN_16429; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16431 = 8'h5a == _T_796[7:0] ? 4'h0 : _GEN_16430; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16432 = 8'h5b == _T_796[7:0] ? 4'h0 : _GEN_16431; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16433 = 8'h5c == _T_796[7:0] ? 4'h0 : _GEN_16432; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16434 = 8'h5d == _T_796[7:0] ? 4'h0 : _GEN_16433; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16435 = 8'h5e == _T_796[7:0] ? 4'h0 : _GEN_16434; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16436 = 8'h5f == _T_796[7:0] ? 4'h0 : _GEN_16435; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16437 = 8'h60 == _T_796[7:0] ? 4'h0 : _GEN_16436; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16438 = 8'h61 == _T_796[7:0] ? 4'h0 : _GEN_16437; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16439 = 8'h62 == _T_796[7:0] ? 4'h0 : _GEN_16438; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16440 = 8'h63 == _T_796[7:0] ? 4'h0 : _GEN_16439; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16441 = 8'h64 == _T_796[7:0] ? 4'h0 : _GEN_16440; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16442 = 8'h65 == _T_796[7:0] ? 4'h0 : _GEN_16441; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16443 = 8'h66 == _T_796[7:0] ? 4'h0 : _GEN_16442; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16444 = 8'h67 == _T_796[7:0] ? 4'h0 : _GEN_16443; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16445 = 8'h68 == _T_796[7:0] ? 4'hf : _GEN_16444; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16446 = 8'h69 == _T_796[7:0] ? 4'hf : _GEN_16445; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16447 = 8'h6a == _T_796[7:0] ? 4'hf : _GEN_16446; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16448 = 8'h6b == _T_796[7:0] ? 4'hf : _GEN_16447; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16449 = 8'h6c == _T_796[7:0] ? 4'hf : _GEN_16448; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16450 = 8'h6d == _T_796[7:0] ? 4'hf : _GEN_16449; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16451 = 8'h6e == _T_796[7:0] ? 4'hf : _GEN_16450; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16452 = 8'h6f == _T_796[7:0] ? 4'hf : _GEN_16451; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16453 = 8'h70 == _T_796[7:0] ? 4'h0 : _GEN_16452; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16454 = 8'h71 == _T_796[7:0] ? 4'h0 : _GEN_16453; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16455 = 8'h72 == _T_796[7:0] ? 4'h0 : _GEN_16454; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16456 = 8'h73 == _T_796[7:0] ? 4'h0 : _GEN_16455; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16457 = 8'h74 == _T_796[7:0] ? 4'h0 : _GEN_16456; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16458 = 8'h75 == _T_796[7:0] ? 4'h0 : _GEN_16457; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16459 = 8'h76 == _T_796[7:0] ? 4'h0 : _GEN_16458; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16460 = 8'h77 == _T_796[7:0] ? 4'h0 : _GEN_16459; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16461 = 8'h78 == _T_796[7:0] ? 4'hf : _GEN_16460; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16462 = 8'h79 == _T_796[7:0] ? 4'hf : _GEN_16461; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16463 = 8'h7a == _T_796[7:0] ? 4'hf : _GEN_16462; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16464 = 8'h7b == _T_796[7:0] ? 4'hf : _GEN_16463; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16465 = 8'h7c == _T_796[7:0] ? 4'hf : _GEN_16464; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16466 = 8'h7d == _T_796[7:0] ? 4'hf : _GEN_16465; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16467 = 8'h7e == _T_796[7:0] ? 4'hf : _GEN_16466; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16468 = 8'h7f == _T_796[7:0] ? 4'hf : _GEN_16467; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16469 = 8'h80 == _T_796[7:0] ? 4'h0 : _GEN_16468; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16470 = 8'h81 == _T_796[7:0] ? 4'h0 : _GEN_16469; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16471 = 8'h82 == _T_796[7:0] ? 4'h0 : _GEN_16470; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16472 = 8'h83 == _T_796[7:0] ? 4'h0 : _GEN_16471; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16473 = 8'h84 == _T_796[7:0] ? 4'h0 : _GEN_16472; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16474 = 8'h85 == _T_796[7:0] ? 4'h0 : _GEN_16473; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16475 = 8'h86 == _T_796[7:0] ? 4'h0 : _GEN_16474; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16476 = 8'h87 == _T_796[7:0] ? 4'h0 : _GEN_16475; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16477 = 8'h88 == _T_796[7:0] ? 4'hf : _GEN_16476; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16478 = 8'h89 == _T_796[7:0] ? 4'hf : _GEN_16477; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16479 = 8'h8a == _T_796[7:0] ? 4'hf : _GEN_16478; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16480 = 8'h8b == _T_796[7:0] ? 4'hf : _GEN_16479; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16481 = 8'h8c == _T_796[7:0] ? 4'hf : _GEN_16480; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16482 = 8'h8d == _T_796[7:0] ? 4'hf : _GEN_16481; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16483 = 8'h8e == _T_796[7:0] ? 4'hf : _GEN_16482; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16484 = 8'h8f == _T_796[7:0] ? 4'hf : _GEN_16483; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16485 = 8'h90 == _T_796[7:0] ? 4'h0 : _GEN_16484; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16486 = 8'h91 == _T_796[7:0] ? 4'h0 : _GEN_16485; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16487 = 8'h92 == _T_796[7:0] ? 4'h0 : _GEN_16486; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16488 = 8'h93 == _T_796[7:0] ? 4'h0 : _GEN_16487; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16489 = 8'h94 == _T_796[7:0] ? 4'h0 : _GEN_16488; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16490 = 8'h95 == _T_796[7:0] ? 4'h0 : _GEN_16489; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16491 = 8'h96 == _T_796[7:0] ? 4'h0 : _GEN_16490; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16492 = 8'h97 == _T_796[7:0] ? 4'h0 : _GEN_16491; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16493 = 8'h98 == _T_796[7:0] ? 4'hf : _GEN_16492; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16494 = 8'h99 == _T_796[7:0] ? 4'hf : _GEN_16493; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16495 = 8'h9a == _T_796[7:0] ? 4'hf : _GEN_16494; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16496 = 8'h9b == _T_796[7:0] ? 4'hf : _GEN_16495; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16497 = 8'h9c == _T_796[7:0] ? 4'hf : _GEN_16496; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16498 = 8'h9d == _T_796[7:0] ? 4'hf : _GEN_16497; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16499 = 8'h9e == _T_796[7:0] ? 4'hf : _GEN_16498; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16500 = 8'h9f == _T_796[7:0] ? 4'hf : _GEN_16499; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16501 = 8'ha0 == _T_796[7:0] ? 4'h0 : _GEN_16500; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16502 = 8'ha1 == _T_796[7:0] ? 4'h0 : _GEN_16501; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16503 = 8'ha2 == _T_796[7:0] ? 4'h0 : _GEN_16502; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16504 = 8'ha3 == _T_796[7:0] ? 4'h0 : _GEN_16503; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16505 = 8'ha4 == _T_796[7:0] ? 4'h0 : _GEN_16504; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16506 = 8'ha5 == _T_796[7:0] ? 4'h0 : _GEN_16505; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16507 = 8'ha6 == _T_796[7:0] ? 4'h0 : _GEN_16506; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16508 = 8'ha7 == _T_796[7:0] ? 4'h0 : _GEN_16507; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16509 = 8'ha8 == _T_796[7:0] ? 4'hf : _GEN_16508; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16510 = 8'ha9 == _T_796[7:0] ? 4'hf : _GEN_16509; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16511 = 8'haa == _T_796[7:0] ? 4'hf : _GEN_16510; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16512 = 8'hab == _T_796[7:0] ? 4'hf : _GEN_16511; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16513 = 8'hac == _T_796[7:0] ? 4'hf : _GEN_16512; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16514 = 8'had == _T_796[7:0] ? 4'hf : _GEN_16513; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16515 = 8'hae == _T_796[7:0] ? 4'hf : _GEN_16514; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16516 = 8'haf == _T_796[7:0] ? 4'hf : _GEN_16515; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16517 = 8'hb0 == _T_796[7:0] ? 4'h0 : _GEN_16516; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16518 = 8'hb1 == _T_796[7:0] ? 4'h0 : _GEN_16517; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16519 = 8'hb2 == _T_796[7:0] ? 4'h0 : _GEN_16518; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16520 = 8'hb3 == _T_796[7:0] ? 4'h0 : _GEN_16519; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16521 = 8'hb4 == _T_796[7:0] ? 4'h0 : _GEN_16520; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16522 = 8'hb5 == _T_796[7:0] ? 4'h0 : _GEN_16521; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16523 = 8'hb6 == _T_796[7:0] ? 4'h0 : _GEN_16522; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16524 = 8'hb7 == _T_796[7:0] ? 4'h0 : _GEN_16523; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16525 = 8'hb8 == _T_796[7:0] ? 4'hf : _GEN_16524; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16526 = 8'hb9 == _T_796[7:0] ? 4'hf : _GEN_16525; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16527 = 8'hba == _T_796[7:0] ? 4'hf : _GEN_16526; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16528 = 8'hbb == _T_796[7:0] ? 4'hf : _GEN_16527; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16529 = 8'hbc == _T_796[7:0] ? 4'hf : _GEN_16528; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16530 = 8'hbd == _T_796[7:0] ? 4'hf : _GEN_16529; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16531 = 8'hbe == _T_796[7:0] ? 4'hf : _GEN_16530; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16532 = 8'hbf == _T_796[7:0] ? 4'hf : _GEN_16531; // @[Filter.scala 165:86]
  wire [4:0] _GEN_19168 = {{1'd0}, _GEN_16532}; // @[Filter.scala 165:86]
  wire [8:0] _T_798 = _GEN_19168 * 5'h14; // @[Filter.scala 165:86]
  wire [3:0] _GEN_16629 = 8'h60 == _T_796[7:0] ? 4'hf : 4'h0; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16630 = 8'h61 == _T_796[7:0] ? 4'hf : _GEN_16629; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16631 = 8'h62 == _T_796[7:0] ? 4'hf : _GEN_16630; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16632 = 8'h63 == _T_796[7:0] ? 4'hf : _GEN_16631; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16633 = 8'h64 == _T_796[7:0] ? 4'hf : _GEN_16632; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16634 = 8'h65 == _T_796[7:0] ? 4'hf : _GEN_16633; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16635 = 8'h66 == _T_796[7:0] ? 4'hf : _GEN_16634; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16636 = 8'h67 == _T_796[7:0] ? 4'hf : _GEN_16635; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16637 = 8'h68 == _T_796[7:0] ? 4'hf : _GEN_16636; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16638 = 8'h69 == _T_796[7:0] ? 4'hf : _GEN_16637; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16639 = 8'h6a == _T_796[7:0] ? 4'hf : _GEN_16638; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16640 = 8'h6b == _T_796[7:0] ? 4'hf : _GEN_16639; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16641 = 8'h6c == _T_796[7:0] ? 4'hf : _GEN_16640; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16642 = 8'h6d == _T_796[7:0] ? 4'hf : _GEN_16641; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16643 = 8'h6e == _T_796[7:0] ? 4'hf : _GEN_16642; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16644 = 8'h6f == _T_796[7:0] ? 4'hf : _GEN_16643; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16645 = 8'h70 == _T_796[7:0] ? 4'hf : _GEN_16644; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16646 = 8'h71 == _T_796[7:0] ? 4'hf : _GEN_16645; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16647 = 8'h72 == _T_796[7:0] ? 4'hf : _GEN_16646; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16648 = 8'h73 == _T_796[7:0] ? 4'hf : _GEN_16647; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16649 = 8'h74 == _T_796[7:0] ? 4'hf : _GEN_16648; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16650 = 8'h75 == _T_796[7:0] ? 4'hf : _GEN_16649; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16651 = 8'h76 == _T_796[7:0] ? 4'hf : _GEN_16650; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16652 = 8'h77 == _T_796[7:0] ? 4'hf : _GEN_16651; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16653 = 8'h78 == _T_796[7:0] ? 4'hf : _GEN_16652; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16654 = 8'h79 == _T_796[7:0] ? 4'hf : _GEN_16653; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16655 = 8'h7a == _T_796[7:0] ? 4'hf : _GEN_16654; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16656 = 8'h7b == _T_796[7:0] ? 4'hf : _GEN_16655; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16657 = 8'h7c == _T_796[7:0] ? 4'hf : _GEN_16656; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16658 = 8'h7d == _T_796[7:0] ? 4'hf : _GEN_16657; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16659 = 8'h7e == _T_796[7:0] ? 4'hf : _GEN_16658; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16660 = 8'h7f == _T_796[7:0] ? 4'hf : _GEN_16659; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16661 = 8'h80 == _T_796[7:0] ? 4'hf : _GEN_16660; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16662 = 8'h81 == _T_796[7:0] ? 4'hf : _GEN_16661; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16663 = 8'h82 == _T_796[7:0] ? 4'hf : _GEN_16662; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16664 = 8'h83 == _T_796[7:0] ? 4'hf : _GEN_16663; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16665 = 8'h84 == _T_796[7:0] ? 4'hf : _GEN_16664; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16666 = 8'h85 == _T_796[7:0] ? 4'hf : _GEN_16665; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16667 = 8'h86 == _T_796[7:0] ? 4'hf : _GEN_16666; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16668 = 8'h87 == _T_796[7:0] ? 4'hf : _GEN_16667; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16669 = 8'h88 == _T_796[7:0] ? 4'hf : _GEN_16668; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16670 = 8'h89 == _T_796[7:0] ? 4'hf : _GEN_16669; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16671 = 8'h8a == _T_796[7:0] ? 4'hf : _GEN_16670; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16672 = 8'h8b == _T_796[7:0] ? 4'hf : _GEN_16671; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16673 = 8'h8c == _T_796[7:0] ? 4'hf : _GEN_16672; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16674 = 8'h8d == _T_796[7:0] ? 4'hf : _GEN_16673; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16675 = 8'h8e == _T_796[7:0] ? 4'hf : _GEN_16674; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16676 = 8'h8f == _T_796[7:0] ? 4'hf : _GEN_16675; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16677 = 8'h90 == _T_796[7:0] ? 4'hf : _GEN_16676; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16678 = 8'h91 == _T_796[7:0] ? 4'hf : _GEN_16677; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16679 = 8'h92 == _T_796[7:0] ? 4'hf : _GEN_16678; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16680 = 8'h93 == _T_796[7:0] ? 4'hf : _GEN_16679; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16681 = 8'h94 == _T_796[7:0] ? 4'hf : _GEN_16680; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16682 = 8'h95 == _T_796[7:0] ? 4'hf : _GEN_16681; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16683 = 8'h96 == _T_796[7:0] ? 4'hf : _GEN_16682; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16684 = 8'h97 == _T_796[7:0] ? 4'hf : _GEN_16683; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16685 = 8'h98 == _T_796[7:0] ? 4'hf : _GEN_16684; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16686 = 8'h99 == _T_796[7:0] ? 4'hf : _GEN_16685; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16687 = 8'h9a == _T_796[7:0] ? 4'hf : _GEN_16686; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16688 = 8'h9b == _T_796[7:0] ? 4'hf : _GEN_16687; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16689 = 8'h9c == _T_796[7:0] ? 4'hf : _GEN_16688; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16690 = 8'h9d == _T_796[7:0] ? 4'hf : _GEN_16689; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16691 = 8'h9e == _T_796[7:0] ? 4'hf : _GEN_16690; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16692 = 8'h9f == _T_796[7:0] ? 4'hf : _GEN_16691; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16693 = 8'ha0 == _T_796[7:0] ? 4'hf : _GEN_16692; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16694 = 8'ha1 == _T_796[7:0] ? 4'hf : _GEN_16693; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16695 = 8'ha2 == _T_796[7:0] ? 4'hf : _GEN_16694; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16696 = 8'ha3 == _T_796[7:0] ? 4'hf : _GEN_16695; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16697 = 8'ha4 == _T_796[7:0] ? 4'hf : _GEN_16696; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16698 = 8'ha5 == _T_796[7:0] ? 4'hf : _GEN_16697; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16699 = 8'ha6 == _T_796[7:0] ? 4'hf : _GEN_16698; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16700 = 8'ha7 == _T_796[7:0] ? 4'hf : _GEN_16699; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16701 = 8'ha8 == _T_796[7:0] ? 4'hf : _GEN_16700; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16702 = 8'ha9 == _T_796[7:0] ? 4'hf : _GEN_16701; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16703 = 8'haa == _T_796[7:0] ? 4'hf : _GEN_16702; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16704 = 8'hab == _T_796[7:0] ? 4'hf : _GEN_16703; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16705 = 8'hac == _T_796[7:0] ? 4'hf : _GEN_16704; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16706 = 8'had == _T_796[7:0] ? 4'hf : _GEN_16705; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16707 = 8'hae == _T_796[7:0] ? 4'hf : _GEN_16706; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16708 = 8'haf == _T_796[7:0] ? 4'hf : _GEN_16707; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16709 = 8'hb0 == _T_796[7:0] ? 4'hf : _GEN_16708; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16710 = 8'hb1 == _T_796[7:0] ? 4'hf : _GEN_16709; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16711 = 8'hb2 == _T_796[7:0] ? 4'hf : _GEN_16710; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16712 = 8'hb3 == _T_796[7:0] ? 4'hf : _GEN_16711; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16713 = 8'hb4 == _T_796[7:0] ? 4'hf : _GEN_16712; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16714 = 8'hb5 == _T_796[7:0] ? 4'hf : _GEN_16713; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16715 = 8'hb6 == _T_796[7:0] ? 4'hf : _GEN_16714; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16716 = 8'hb7 == _T_796[7:0] ? 4'hf : _GEN_16715; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16717 = 8'hb8 == _T_796[7:0] ? 4'hf : _GEN_16716; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16718 = 8'hb9 == _T_796[7:0] ? 4'hf : _GEN_16717; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16719 = 8'hba == _T_796[7:0] ? 4'hf : _GEN_16718; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16720 = 8'hbb == _T_796[7:0] ? 4'hf : _GEN_16719; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16721 = 8'hbc == _T_796[7:0] ? 4'hf : _GEN_16720; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16722 = 8'hbd == _T_796[7:0] ? 4'hf : _GEN_16721; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16723 = 8'hbe == _T_796[7:0] ? 4'hf : _GEN_16722; // @[Filter.scala 165:126]
  wire [3:0] _GEN_16724 = 8'hbf == _T_796[7:0] ? 4'hf : _GEN_16723; // @[Filter.scala 165:126]
  wire [6:0] _GEN_19170 = {{3'd0}, _GEN_16724}; // @[Filter.scala 165:126]
  wire [10:0] _T_803 = _GEN_19170 * 7'h46; // @[Filter.scala 165:126]
  wire [10:0] _GEN_19171 = {{2'd0}, _T_798}; // @[Filter.scala 165:93]
  wire [10:0] _T_805 = _GEN_19171 + _T_803; // @[Filter.scala 165:93]
  wire [3:0] _GEN_16733 = 8'h8 == _T_796[7:0] ? 4'hf : 4'h0; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16734 = 8'h9 == _T_796[7:0] ? 4'hf : _GEN_16733; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16735 = 8'ha == _T_796[7:0] ? 4'hf : _GEN_16734; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16736 = 8'hb == _T_796[7:0] ? 4'hf : _GEN_16735; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16737 = 8'hc == _T_796[7:0] ? 4'hf : _GEN_16736; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16738 = 8'hd == _T_796[7:0] ? 4'hf : _GEN_16737; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16739 = 8'he == _T_796[7:0] ? 4'hf : _GEN_16738; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16740 = 8'hf == _T_796[7:0] ? 4'hf : _GEN_16739; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16741 = 8'h10 == _T_796[7:0] ? 4'h0 : _GEN_16740; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16742 = 8'h11 == _T_796[7:0] ? 4'h0 : _GEN_16741; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16743 = 8'h12 == _T_796[7:0] ? 4'h0 : _GEN_16742; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16744 = 8'h13 == _T_796[7:0] ? 4'h0 : _GEN_16743; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16745 = 8'h14 == _T_796[7:0] ? 4'h0 : _GEN_16744; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16746 = 8'h15 == _T_796[7:0] ? 4'h0 : _GEN_16745; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16747 = 8'h16 == _T_796[7:0] ? 4'h0 : _GEN_16746; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16748 = 8'h17 == _T_796[7:0] ? 4'h0 : _GEN_16747; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16749 = 8'h18 == _T_796[7:0] ? 4'hf : _GEN_16748; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16750 = 8'h19 == _T_796[7:0] ? 4'hf : _GEN_16749; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16751 = 8'h1a == _T_796[7:0] ? 4'hf : _GEN_16750; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16752 = 8'h1b == _T_796[7:0] ? 4'hf : _GEN_16751; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16753 = 8'h1c == _T_796[7:0] ? 4'hf : _GEN_16752; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16754 = 8'h1d == _T_796[7:0] ? 4'hf : _GEN_16753; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16755 = 8'h1e == _T_796[7:0] ? 4'hf : _GEN_16754; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16756 = 8'h1f == _T_796[7:0] ? 4'hf : _GEN_16755; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16757 = 8'h20 == _T_796[7:0] ? 4'h0 : _GEN_16756; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16758 = 8'h21 == _T_796[7:0] ? 4'h0 : _GEN_16757; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16759 = 8'h22 == _T_796[7:0] ? 4'h0 : _GEN_16758; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16760 = 8'h23 == _T_796[7:0] ? 4'h0 : _GEN_16759; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16761 = 8'h24 == _T_796[7:0] ? 4'h0 : _GEN_16760; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16762 = 8'h25 == _T_796[7:0] ? 4'h0 : _GEN_16761; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16763 = 8'h26 == _T_796[7:0] ? 4'h0 : _GEN_16762; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16764 = 8'h27 == _T_796[7:0] ? 4'h0 : _GEN_16763; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16765 = 8'h28 == _T_796[7:0] ? 4'hf : _GEN_16764; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16766 = 8'h29 == _T_796[7:0] ? 4'hf : _GEN_16765; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16767 = 8'h2a == _T_796[7:0] ? 4'hf : _GEN_16766; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16768 = 8'h2b == _T_796[7:0] ? 4'hf : _GEN_16767; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16769 = 8'h2c == _T_796[7:0] ? 4'hf : _GEN_16768; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16770 = 8'h2d == _T_796[7:0] ? 4'hf : _GEN_16769; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16771 = 8'h2e == _T_796[7:0] ? 4'hf : _GEN_16770; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16772 = 8'h2f == _T_796[7:0] ? 4'hf : _GEN_16771; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16773 = 8'h30 == _T_796[7:0] ? 4'h0 : _GEN_16772; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16774 = 8'h31 == _T_796[7:0] ? 4'h0 : _GEN_16773; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16775 = 8'h32 == _T_796[7:0] ? 4'h0 : _GEN_16774; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16776 = 8'h33 == _T_796[7:0] ? 4'h0 : _GEN_16775; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16777 = 8'h34 == _T_796[7:0] ? 4'h0 : _GEN_16776; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16778 = 8'h35 == _T_796[7:0] ? 4'h0 : _GEN_16777; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16779 = 8'h36 == _T_796[7:0] ? 4'h0 : _GEN_16778; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16780 = 8'h37 == _T_796[7:0] ? 4'h0 : _GEN_16779; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16781 = 8'h38 == _T_796[7:0] ? 4'hf : _GEN_16780; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16782 = 8'h39 == _T_796[7:0] ? 4'hf : _GEN_16781; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16783 = 8'h3a == _T_796[7:0] ? 4'hf : _GEN_16782; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16784 = 8'h3b == _T_796[7:0] ? 4'hf : _GEN_16783; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16785 = 8'h3c == _T_796[7:0] ? 4'hf : _GEN_16784; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16786 = 8'h3d == _T_796[7:0] ? 4'hf : _GEN_16785; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16787 = 8'h3e == _T_796[7:0] ? 4'hf : _GEN_16786; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16788 = 8'h3f == _T_796[7:0] ? 4'hf : _GEN_16787; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16789 = 8'h40 == _T_796[7:0] ? 4'h0 : _GEN_16788; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16790 = 8'h41 == _T_796[7:0] ? 4'h0 : _GEN_16789; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16791 = 8'h42 == _T_796[7:0] ? 4'h0 : _GEN_16790; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16792 = 8'h43 == _T_796[7:0] ? 4'h0 : _GEN_16791; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16793 = 8'h44 == _T_796[7:0] ? 4'h0 : _GEN_16792; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16794 = 8'h45 == _T_796[7:0] ? 4'h0 : _GEN_16793; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16795 = 8'h46 == _T_796[7:0] ? 4'h0 : _GEN_16794; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16796 = 8'h47 == _T_796[7:0] ? 4'h0 : _GEN_16795; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16797 = 8'h48 == _T_796[7:0] ? 4'hf : _GEN_16796; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16798 = 8'h49 == _T_796[7:0] ? 4'hf : _GEN_16797; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16799 = 8'h4a == _T_796[7:0] ? 4'hf : _GEN_16798; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16800 = 8'h4b == _T_796[7:0] ? 4'hf : _GEN_16799; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16801 = 8'h4c == _T_796[7:0] ? 4'hf : _GEN_16800; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16802 = 8'h4d == _T_796[7:0] ? 4'hf : _GEN_16801; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16803 = 8'h4e == _T_796[7:0] ? 4'hf : _GEN_16802; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16804 = 8'h4f == _T_796[7:0] ? 4'hf : _GEN_16803; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16805 = 8'h50 == _T_796[7:0] ? 4'h0 : _GEN_16804; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16806 = 8'h51 == _T_796[7:0] ? 4'h0 : _GEN_16805; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16807 = 8'h52 == _T_796[7:0] ? 4'h0 : _GEN_16806; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16808 = 8'h53 == _T_796[7:0] ? 4'h0 : _GEN_16807; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16809 = 8'h54 == _T_796[7:0] ? 4'h0 : _GEN_16808; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16810 = 8'h55 == _T_796[7:0] ? 4'h0 : _GEN_16809; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16811 = 8'h56 == _T_796[7:0] ? 4'h0 : _GEN_16810; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16812 = 8'h57 == _T_796[7:0] ? 4'h0 : _GEN_16811; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16813 = 8'h58 == _T_796[7:0] ? 4'hf : _GEN_16812; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16814 = 8'h59 == _T_796[7:0] ? 4'hf : _GEN_16813; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16815 = 8'h5a == _T_796[7:0] ? 4'hf : _GEN_16814; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16816 = 8'h5b == _T_796[7:0] ? 4'hf : _GEN_16815; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16817 = 8'h5c == _T_796[7:0] ? 4'hf : _GEN_16816; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16818 = 8'h5d == _T_796[7:0] ? 4'hf : _GEN_16817; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16819 = 8'h5e == _T_796[7:0] ? 4'hf : _GEN_16818; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16820 = 8'h5f == _T_796[7:0] ? 4'hf : _GEN_16819; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16821 = 8'h60 == _T_796[7:0] ? 4'h0 : _GEN_16820; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16822 = 8'h61 == _T_796[7:0] ? 4'h0 : _GEN_16821; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16823 = 8'h62 == _T_796[7:0] ? 4'h0 : _GEN_16822; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16824 = 8'h63 == _T_796[7:0] ? 4'h0 : _GEN_16823; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16825 = 8'h64 == _T_796[7:0] ? 4'h0 : _GEN_16824; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16826 = 8'h65 == _T_796[7:0] ? 4'h0 : _GEN_16825; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16827 = 8'h66 == _T_796[7:0] ? 4'h0 : _GEN_16826; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16828 = 8'h67 == _T_796[7:0] ? 4'h0 : _GEN_16827; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16829 = 8'h68 == _T_796[7:0] ? 4'hf : _GEN_16828; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16830 = 8'h69 == _T_796[7:0] ? 4'hf : _GEN_16829; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16831 = 8'h6a == _T_796[7:0] ? 4'hf : _GEN_16830; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16832 = 8'h6b == _T_796[7:0] ? 4'hf : _GEN_16831; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16833 = 8'h6c == _T_796[7:0] ? 4'hf : _GEN_16832; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16834 = 8'h6d == _T_796[7:0] ? 4'hf : _GEN_16833; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16835 = 8'h6e == _T_796[7:0] ? 4'hf : _GEN_16834; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16836 = 8'h6f == _T_796[7:0] ? 4'hf : _GEN_16835; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16837 = 8'h70 == _T_796[7:0] ? 4'h0 : _GEN_16836; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16838 = 8'h71 == _T_796[7:0] ? 4'h0 : _GEN_16837; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16839 = 8'h72 == _T_796[7:0] ? 4'h0 : _GEN_16838; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16840 = 8'h73 == _T_796[7:0] ? 4'h0 : _GEN_16839; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16841 = 8'h74 == _T_796[7:0] ? 4'h0 : _GEN_16840; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16842 = 8'h75 == _T_796[7:0] ? 4'h0 : _GEN_16841; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16843 = 8'h76 == _T_796[7:0] ? 4'h0 : _GEN_16842; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16844 = 8'h77 == _T_796[7:0] ? 4'h0 : _GEN_16843; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16845 = 8'h78 == _T_796[7:0] ? 4'hf : _GEN_16844; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16846 = 8'h79 == _T_796[7:0] ? 4'hf : _GEN_16845; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16847 = 8'h7a == _T_796[7:0] ? 4'hf : _GEN_16846; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16848 = 8'h7b == _T_796[7:0] ? 4'hf : _GEN_16847; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16849 = 8'h7c == _T_796[7:0] ? 4'hf : _GEN_16848; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16850 = 8'h7d == _T_796[7:0] ? 4'hf : _GEN_16849; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16851 = 8'h7e == _T_796[7:0] ? 4'hf : _GEN_16850; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16852 = 8'h7f == _T_796[7:0] ? 4'hf : _GEN_16851; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16853 = 8'h80 == _T_796[7:0] ? 4'h0 : _GEN_16852; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16854 = 8'h81 == _T_796[7:0] ? 4'h0 : _GEN_16853; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16855 = 8'h82 == _T_796[7:0] ? 4'h0 : _GEN_16854; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16856 = 8'h83 == _T_796[7:0] ? 4'h0 : _GEN_16855; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16857 = 8'h84 == _T_796[7:0] ? 4'h0 : _GEN_16856; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16858 = 8'h85 == _T_796[7:0] ? 4'h0 : _GEN_16857; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16859 = 8'h86 == _T_796[7:0] ? 4'h0 : _GEN_16858; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16860 = 8'h87 == _T_796[7:0] ? 4'h0 : _GEN_16859; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16861 = 8'h88 == _T_796[7:0] ? 4'hf : _GEN_16860; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16862 = 8'h89 == _T_796[7:0] ? 4'hf : _GEN_16861; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16863 = 8'h8a == _T_796[7:0] ? 4'hf : _GEN_16862; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16864 = 8'h8b == _T_796[7:0] ? 4'hf : _GEN_16863; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16865 = 8'h8c == _T_796[7:0] ? 4'hf : _GEN_16864; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16866 = 8'h8d == _T_796[7:0] ? 4'hf : _GEN_16865; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16867 = 8'h8e == _T_796[7:0] ? 4'hf : _GEN_16866; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16868 = 8'h8f == _T_796[7:0] ? 4'hf : _GEN_16867; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16869 = 8'h90 == _T_796[7:0] ? 4'h0 : _GEN_16868; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16870 = 8'h91 == _T_796[7:0] ? 4'h0 : _GEN_16869; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16871 = 8'h92 == _T_796[7:0] ? 4'h0 : _GEN_16870; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16872 = 8'h93 == _T_796[7:0] ? 4'h0 : _GEN_16871; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16873 = 8'h94 == _T_796[7:0] ? 4'h0 : _GEN_16872; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16874 = 8'h95 == _T_796[7:0] ? 4'h0 : _GEN_16873; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16875 = 8'h96 == _T_796[7:0] ? 4'h0 : _GEN_16874; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16876 = 8'h97 == _T_796[7:0] ? 4'h0 : _GEN_16875; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16877 = 8'h98 == _T_796[7:0] ? 4'hf : _GEN_16876; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16878 = 8'h99 == _T_796[7:0] ? 4'hf : _GEN_16877; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16879 = 8'h9a == _T_796[7:0] ? 4'hf : _GEN_16878; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16880 = 8'h9b == _T_796[7:0] ? 4'hf : _GEN_16879; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16881 = 8'h9c == _T_796[7:0] ? 4'hf : _GEN_16880; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16882 = 8'h9d == _T_796[7:0] ? 4'hf : _GEN_16881; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16883 = 8'h9e == _T_796[7:0] ? 4'hf : _GEN_16882; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16884 = 8'h9f == _T_796[7:0] ? 4'hf : _GEN_16883; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16885 = 8'ha0 == _T_796[7:0] ? 4'h0 : _GEN_16884; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16886 = 8'ha1 == _T_796[7:0] ? 4'h0 : _GEN_16885; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16887 = 8'ha2 == _T_796[7:0] ? 4'h0 : _GEN_16886; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16888 = 8'ha3 == _T_796[7:0] ? 4'h0 : _GEN_16887; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16889 = 8'ha4 == _T_796[7:0] ? 4'h0 : _GEN_16888; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16890 = 8'ha5 == _T_796[7:0] ? 4'h0 : _GEN_16889; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16891 = 8'ha6 == _T_796[7:0] ? 4'h0 : _GEN_16890; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16892 = 8'ha7 == _T_796[7:0] ? 4'h0 : _GEN_16891; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16893 = 8'ha8 == _T_796[7:0] ? 4'hf : _GEN_16892; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16894 = 8'ha9 == _T_796[7:0] ? 4'hf : _GEN_16893; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16895 = 8'haa == _T_796[7:0] ? 4'hf : _GEN_16894; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16896 = 8'hab == _T_796[7:0] ? 4'hf : _GEN_16895; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16897 = 8'hac == _T_796[7:0] ? 4'hf : _GEN_16896; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16898 = 8'had == _T_796[7:0] ? 4'hf : _GEN_16897; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16899 = 8'hae == _T_796[7:0] ? 4'hf : _GEN_16898; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16900 = 8'haf == _T_796[7:0] ? 4'hf : _GEN_16899; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16901 = 8'hb0 == _T_796[7:0] ? 4'h0 : _GEN_16900; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16902 = 8'hb1 == _T_796[7:0] ? 4'h0 : _GEN_16901; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16903 = 8'hb2 == _T_796[7:0] ? 4'h0 : _GEN_16902; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16904 = 8'hb3 == _T_796[7:0] ? 4'h0 : _GEN_16903; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16905 = 8'hb4 == _T_796[7:0] ? 4'h0 : _GEN_16904; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16906 = 8'hb5 == _T_796[7:0] ? 4'h0 : _GEN_16905; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16907 = 8'hb6 == _T_796[7:0] ? 4'h0 : _GEN_16906; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16908 = 8'hb7 == _T_796[7:0] ? 4'h0 : _GEN_16907; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16909 = 8'hb8 == _T_796[7:0] ? 4'hf : _GEN_16908; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16910 = 8'hb9 == _T_796[7:0] ? 4'hf : _GEN_16909; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16911 = 8'hba == _T_796[7:0] ? 4'hf : _GEN_16910; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16912 = 8'hbb == _T_796[7:0] ? 4'hf : _GEN_16911; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16913 = 8'hbc == _T_796[7:0] ? 4'hf : _GEN_16912; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16914 = 8'hbd == _T_796[7:0] ? 4'hf : _GEN_16913; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16915 = 8'hbe == _T_796[7:0] ? 4'hf : _GEN_16914; // @[Filter.scala 165:166]
  wire [3:0] _GEN_16916 = 8'hbf == _T_796[7:0] ? 4'hf : _GEN_16915; // @[Filter.scala 165:166]
  wire [7:0] _T_810 = _GEN_16916 * 4'ha; // @[Filter.scala 165:166]
  wire [10:0] _GEN_19173 = {{3'd0}, _T_810}; // @[Filter.scala 165:133]
  wire [10:0] _T_812 = _T_805 + _GEN_19173; // @[Filter.scala 165:133]
  wire [10:0] _T_813 = _T_812 / 11'h64; // @[Filter.scala 165:174]
  wire [10:0] _GEN_17109 = io_SPI_distort ? _T_813 : {{7'd0}, _GEN_16532}; // @[Filter.scala 164:35]
  wire [10:0] _GEN_17110 = _T_793 ? 11'h0 : _GEN_17109; // @[Filter.scala 162:80]
  wire [10:0] _GEN_17879 = io_SPI_distort ? _T_813 : {{7'd0}, _GEN_16724}; // @[Filter.scala 164:35]
  wire [10:0] _GEN_17880 = _T_793 ? 11'h0 : _GEN_17879; // @[Filter.scala 162:80]
  wire [10:0] _GEN_18649 = io_SPI_distort ? _T_813 : {{7'd0}, _GEN_16916}; // @[Filter.scala 164:35]
  wire [10:0] _GEN_18650 = _T_793 ? 11'h0 : _GEN_18649; // @[Filter.scala 162:80]
  wire [7:0] _GEN_18652 = 3'h1 == io_SPI_filterIndex[2:0] ? $signed(8'sh9) : $signed(8'sh1); // @[Filter.scala 185:33]
  wire [7:0] _GEN_18653 = 3'h2 == io_SPI_filterIndex[2:0] ? $signed(8'sh10) : $signed(_GEN_18652); // @[Filter.scala 185:33]
  wire [7:0] _GEN_18654 = 3'h3 == io_SPI_filterIndex[2:0] ? $signed(8'sh1) : $signed(_GEN_18653); // @[Filter.scala 185:33]
  wire [7:0] _GEN_18655 = 3'h4 == io_SPI_filterIndex[2:0] ? $signed(8'sh1) : $signed(_GEN_18654); // @[Filter.scala 185:33]
  wire [7:0] _GEN_18656 = 3'h5 == io_SPI_filterIndex[2:0] ? $signed(8'sh1) : $signed(_GEN_18655); // @[Filter.scala 185:33]
  wire [8:0] _GEN_19191 = {{1{_GEN_18656[7]}},_GEN_18656}; // @[Filter.scala 185:33]
  wire [9:0] _T_884 = $signed(KernelConvolution_io_pixelVal_out_0) / $signed(_GEN_19191); // @[Filter.scala 185:44]
  wire [9:0] _T_890 = $signed(KernelConvolution_io_pixelVal_out_1) / $signed(_GEN_19191); // @[Filter.scala 185:44]
  wire [9:0] _T_896 = $signed(KernelConvolution_io_pixelVal_out_2) / $signed(_GEN_19191); // @[Filter.scala 185:44]
  wire [9:0] _T_902 = $signed(KernelConvolution_io_pixelVal_out_3) / $signed(_GEN_19191); // @[Filter.scala 185:44]
  wire [9:0] _T_908 = $signed(KernelConvolution_io_pixelVal_out_4) / $signed(_GEN_19191); // @[Filter.scala 185:44]
  wire [9:0] _T_914 = $signed(KernelConvolution_io_pixelVal_out_5) / $signed(_GEN_19191); // @[Filter.scala 185:44]
  wire [9:0] _T_920 = $signed(KernelConvolution_io_pixelVal_out_6) / $signed(_GEN_19191); // @[Filter.scala 185:44]
  wire [9:0] _T_926 = $signed(KernelConvolution_io_pixelVal_out_7) / $signed(_GEN_19191); // @[Filter.scala 185:44]
  wire [9:0] _T_932 = $signed(KernelConvolution_1_io_pixelVal_out_0) / $signed(_GEN_19191); // @[Filter.scala 185:44]
  wire [9:0] _T_938 = $signed(KernelConvolution_1_io_pixelVal_out_1) / $signed(_GEN_19191); // @[Filter.scala 185:44]
  wire [9:0] _T_944 = $signed(KernelConvolution_1_io_pixelVal_out_2) / $signed(_GEN_19191); // @[Filter.scala 185:44]
  wire [9:0] _T_950 = $signed(KernelConvolution_1_io_pixelVal_out_3) / $signed(_GEN_19191); // @[Filter.scala 185:44]
  wire [9:0] _T_956 = $signed(KernelConvolution_1_io_pixelVal_out_4) / $signed(_GEN_19191); // @[Filter.scala 185:44]
  wire [9:0] _T_962 = $signed(KernelConvolution_1_io_pixelVal_out_5) / $signed(_GEN_19191); // @[Filter.scala 185:44]
  wire [9:0] _T_968 = $signed(KernelConvolution_1_io_pixelVal_out_6) / $signed(_GEN_19191); // @[Filter.scala 185:44]
  wire [9:0] _T_974 = $signed(KernelConvolution_1_io_pixelVal_out_7) / $signed(_GEN_19191); // @[Filter.scala 185:44]
  wire [9:0] _T_980 = $signed(KernelConvolution_2_io_pixelVal_out_0) / $signed(_GEN_19191); // @[Filter.scala 185:44]
  wire [9:0] _T_986 = $signed(KernelConvolution_2_io_pixelVal_out_1) / $signed(_GEN_19191); // @[Filter.scala 185:44]
  wire [9:0] _T_992 = $signed(KernelConvolution_2_io_pixelVal_out_2) / $signed(_GEN_19191); // @[Filter.scala 185:44]
  wire [9:0] _T_998 = $signed(KernelConvolution_2_io_pixelVal_out_3) / $signed(_GEN_19191); // @[Filter.scala 185:44]
  wire [9:0] _T_1004 = $signed(KernelConvolution_2_io_pixelVal_out_4) / $signed(_GEN_19191); // @[Filter.scala 185:44]
  wire [9:0] _T_1010 = $signed(KernelConvolution_2_io_pixelVal_out_5) / $signed(_GEN_19191); // @[Filter.scala 185:44]
  wire [9:0] _T_1016 = $signed(KernelConvolution_2_io_pixelVal_out_6) / $signed(_GEN_19191); // @[Filter.scala 185:44]
  wire [9:0] _T_1022 = $signed(KernelConvolution_2_io_pixelVal_out_7) / $signed(_GEN_19191); // @[Filter.scala 185:44]
  wire [31:0] _T_1026 = pixelIndex + 32'h8; // @[Filter.scala 199:34]
  wire [8:0] _T_1027 = 5'h10 * 5'hc; // @[Filter.scala 200:42]
  wire [31:0] _GEN_19215 = {{23'd0}, _T_1027}; // @[Filter.scala 200:25]
  wire  _T_1028 = pixelIndex == _GEN_19215; // @[Filter.scala 200:25]
  KernelConvolution KernelConvolution ( // @[Filter.scala 142:36]
    .clock(KernelConvolution_clock),
    .reset(KernelConvolution_reset),
    .io_kernelVal_in(KernelConvolution_io_kernelVal_in),
    .io_pixelVal_in_0(KernelConvolution_io_pixelVal_in_0),
    .io_pixelVal_in_1(KernelConvolution_io_pixelVal_in_1),
    .io_pixelVal_in_2(KernelConvolution_io_pixelVal_in_2),
    .io_pixelVal_in_3(KernelConvolution_io_pixelVal_in_3),
    .io_pixelVal_in_4(KernelConvolution_io_pixelVal_in_4),
    .io_pixelVal_in_5(KernelConvolution_io_pixelVal_in_5),
    .io_pixelVal_in_6(KernelConvolution_io_pixelVal_in_6),
    .io_pixelVal_in_7(KernelConvolution_io_pixelVal_in_7),
    .io_pixelVal_out_0(KernelConvolution_io_pixelVal_out_0),
    .io_pixelVal_out_1(KernelConvolution_io_pixelVal_out_1),
    .io_pixelVal_out_2(KernelConvolution_io_pixelVal_out_2),
    .io_pixelVal_out_3(KernelConvolution_io_pixelVal_out_3),
    .io_pixelVal_out_4(KernelConvolution_io_pixelVal_out_4),
    .io_pixelVal_out_5(KernelConvolution_io_pixelVal_out_5),
    .io_pixelVal_out_6(KernelConvolution_io_pixelVal_out_6),
    .io_pixelVal_out_7(KernelConvolution_io_pixelVal_out_7),
    .io_valid_out(KernelConvolution_io_valid_out)
  );
  KernelConvolution KernelConvolution_1 ( // @[Filter.scala 143:36]
    .clock(KernelConvolution_1_clock),
    .reset(KernelConvolution_1_reset),
    .io_kernelVal_in(KernelConvolution_1_io_kernelVal_in),
    .io_pixelVal_in_0(KernelConvolution_1_io_pixelVal_in_0),
    .io_pixelVal_in_1(KernelConvolution_1_io_pixelVal_in_1),
    .io_pixelVal_in_2(KernelConvolution_1_io_pixelVal_in_2),
    .io_pixelVal_in_3(KernelConvolution_1_io_pixelVal_in_3),
    .io_pixelVal_in_4(KernelConvolution_1_io_pixelVal_in_4),
    .io_pixelVal_in_5(KernelConvolution_1_io_pixelVal_in_5),
    .io_pixelVal_in_6(KernelConvolution_1_io_pixelVal_in_6),
    .io_pixelVal_in_7(KernelConvolution_1_io_pixelVal_in_7),
    .io_pixelVal_out_0(KernelConvolution_1_io_pixelVal_out_0),
    .io_pixelVal_out_1(KernelConvolution_1_io_pixelVal_out_1),
    .io_pixelVal_out_2(KernelConvolution_1_io_pixelVal_out_2),
    .io_pixelVal_out_3(KernelConvolution_1_io_pixelVal_out_3),
    .io_pixelVal_out_4(KernelConvolution_1_io_pixelVal_out_4),
    .io_pixelVal_out_5(KernelConvolution_1_io_pixelVal_out_5),
    .io_pixelVal_out_6(KernelConvolution_1_io_pixelVal_out_6),
    .io_pixelVal_out_7(KernelConvolution_1_io_pixelVal_out_7),
    .io_valid_out(KernelConvolution_1_io_valid_out)
  );
  KernelConvolution KernelConvolution_2 ( // @[Filter.scala 144:36]
    .clock(KernelConvolution_2_clock),
    .reset(KernelConvolution_2_reset),
    .io_kernelVal_in(KernelConvolution_2_io_kernelVal_in),
    .io_pixelVal_in_0(KernelConvolution_2_io_pixelVal_in_0),
    .io_pixelVal_in_1(KernelConvolution_2_io_pixelVal_in_1),
    .io_pixelVal_in_2(KernelConvolution_2_io_pixelVal_in_2),
    .io_pixelVal_in_3(KernelConvolution_2_io_pixelVal_in_3),
    .io_pixelVal_in_4(KernelConvolution_2_io_pixelVal_in_4),
    .io_pixelVal_in_5(KernelConvolution_2_io_pixelVal_in_5),
    .io_pixelVal_in_6(KernelConvolution_2_io_pixelVal_in_6),
    .io_pixelVal_in_7(KernelConvolution_2_io_pixelVal_in_7),
    .io_pixelVal_out_0(KernelConvolution_2_io_pixelVal_out_0),
    .io_pixelVal_out_1(KernelConvolution_2_io_pixelVal_out_1),
    .io_pixelVal_out_2(KernelConvolution_2_io_pixelVal_out_2),
    .io_pixelVal_out_3(KernelConvolution_2_io_pixelVal_out_3),
    .io_pixelVal_out_4(KernelConvolution_2_io_pixelVal_out_4),
    .io_pixelVal_out_5(KernelConvolution_2_io_pixelVal_out_5),
    .io_pixelVal_out_6(KernelConvolution_2_io_pixelVal_out_6),
    .io_pixelVal_out_7(KernelConvolution_2_io_pixelVal_out_7),
    .io_valid_out(KernelConvolution_2_io_valid_out)
  );
  assign io_pixelVal_out_0_0 = _T_884[3:0]; // @[Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_0_1 = _T_890[3:0]; // @[Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_0_2 = _T_896[3:0]; // @[Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_0_3 = _T_902[3:0]; // @[Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_0_4 = _T_908[3:0]; // @[Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_0_5 = _T_914[3:0]; // @[Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_0_6 = _T_920[3:0]; // @[Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_0_7 = _T_926[3:0]; // @[Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_1_0 = _T_932[3:0]; // @[Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_1_1 = _T_938[3:0]; // @[Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_1_2 = _T_944[3:0]; // @[Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_1_3 = _T_950[3:0]; // @[Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_1_4 = _T_956[3:0]; // @[Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_1_5 = _T_962[3:0]; // @[Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_1_6 = _T_968[3:0]; // @[Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_1_7 = _T_974[3:0]; // @[Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_2_0 = _T_980[3:0]; // @[Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_2_1 = _T_986[3:0]; // @[Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_2_2 = _T_992[3:0]; // @[Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_2_3 = _T_998[3:0]; // @[Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_2_4 = _T_1004[3:0]; // @[Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_2_5 = _T_1010[3:0]; // @[Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_2_6 = _T_1016[3:0]; // @[Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_2_7 = _T_1022[3:0]; // @[Filter.scala 189:35 Filter.scala 191:35]
  assign io_valid_out = KernelConvolution_io_valid_out; // @[Filter.scala 196:18]
  assign KernelConvolution_clock = clock;
  assign KernelConvolution_reset = reset;
  assign KernelConvolution_io_kernelVal_in = _GEN_18765 & _GEN_18692 ? $signed(5'sh0) : $signed(_GEN_55); // @[Filter.scala 150:41]
  assign KernelConvolution_io_pixelVal_in_0 = _GEN_940[3:0]; // @[Filter.scala 163:53 Filter.scala 165:51 Filter.scala 167:51]
  assign KernelConvolution_io_pixelVal_in_1 = _GEN_3250[3:0]; // @[Filter.scala 163:53 Filter.scala 165:51 Filter.scala 167:51]
  assign KernelConvolution_io_pixelVal_in_2 = _GEN_5560[3:0]; // @[Filter.scala 163:53 Filter.scala 165:51 Filter.scala 167:51]
  assign KernelConvolution_io_pixelVal_in_3 = _GEN_7870[3:0]; // @[Filter.scala 163:53 Filter.scala 165:51 Filter.scala 167:51]
  assign KernelConvolution_io_pixelVal_in_4 = _GEN_10180[3:0]; // @[Filter.scala 163:53 Filter.scala 165:51 Filter.scala 167:51]
  assign KernelConvolution_io_pixelVal_in_5 = _GEN_12490[3:0]; // @[Filter.scala 163:53 Filter.scala 165:51 Filter.scala 167:51]
  assign KernelConvolution_io_pixelVal_in_6 = _GEN_14800[3:0]; // @[Filter.scala 163:53 Filter.scala 165:51 Filter.scala 167:51]
  assign KernelConvolution_io_pixelVal_in_7 = _GEN_17110[3:0]; // @[Filter.scala 163:53 Filter.scala 165:51 Filter.scala 167:51]
  assign KernelConvolution_1_clock = clock;
  assign KernelConvolution_1_reset = reset;
  assign KernelConvolution_1_io_kernelVal_in = _GEN_18765 & _GEN_18692 ? $signed(5'sh0) : $signed(_GEN_55); // @[Filter.scala 150:41]
  assign KernelConvolution_1_io_pixelVal_in_0 = _GEN_1710[3:0]; // @[Filter.scala 163:53 Filter.scala 165:51 Filter.scala 167:51]
  assign KernelConvolution_1_io_pixelVal_in_1 = _GEN_4020[3:0]; // @[Filter.scala 163:53 Filter.scala 165:51 Filter.scala 167:51]
  assign KernelConvolution_1_io_pixelVal_in_2 = _GEN_6330[3:0]; // @[Filter.scala 163:53 Filter.scala 165:51 Filter.scala 167:51]
  assign KernelConvolution_1_io_pixelVal_in_3 = _GEN_8640[3:0]; // @[Filter.scala 163:53 Filter.scala 165:51 Filter.scala 167:51]
  assign KernelConvolution_1_io_pixelVal_in_4 = _GEN_10950[3:0]; // @[Filter.scala 163:53 Filter.scala 165:51 Filter.scala 167:51]
  assign KernelConvolution_1_io_pixelVal_in_5 = _GEN_13260[3:0]; // @[Filter.scala 163:53 Filter.scala 165:51 Filter.scala 167:51]
  assign KernelConvolution_1_io_pixelVal_in_6 = _GEN_15570[3:0]; // @[Filter.scala 163:53 Filter.scala 165:51 Filter.scala 167:51]
  assign KernelConvolution_1_io_pixelVal_in_7 = _GEN_17880[3:0]; // @[Filter.scala 163:53 Filter.scala 165:51 Filter.scala 167:51]
  assign KernelConvolution_2_clock = clock;
  assign KernelConvolution_2_reset = reset;
  assign KernelConvolution_2_io_kernelVal_in = _GEN_18765 & _GEN_18692 ? $signed(5'sh0) : $signed(_GEN_55); // @[Filter.scala 150:41]
  assign KernelConvolution_2_io_pixelVal_in_0 = _GEN_2480[3:0]; // @[Filter.scala 163:53 Filter.scala 165:51 Filter.scala 167:51]
  assign KernelConvolution_2_io_pixelVal_in_1 = _GEN_4790[3:0]; // @[Filter.scala 163:53 Filter.scala 165:51 Filter.scala 167:51]
  assign KernelConvolution_2_io_pixelVal_in_2 = _GEN_7100[3:0]; // @[Filter.scala 163:53 Filter.scala 165:51 Filter.scala 167:51]
  assign KernelConvolution_2_io_pixelVal_in_3 = _GEN_9410[3:0]; // @[Filter.scala 163:53 Filter.scala 165:51 Filter.scala 167:51]
  assign KernelConvolution_2_io_pixelVal_in_4 = _GEN_11720[3:0]; // @[Filter.scala 163:53 Filter.scala 165:51 Filter.scala 167:51]
  assign KernelConvolution_2_io_pixelVal_in_5 = _GEN_14030[3:0]; // @[Filter.scala 163:53 Filter.scala 165:51 Filter.scala 167:51]
  assign KernelConvolution_2_io_pixelVal_in_6 = _GEN_16340[3:0]; // @[Filter.scala 163:53 Filter.scala 165:51 Filter.scala 167:51]
  assign KernelConvolution_2_io_pixelVal_in_7 = _GEN_18650[3:0]; // @[Filter.scala 163:53 Filter.scala 165:51 Filter.scala 167:51]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  kernelCounter = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  imageCounterX = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  imageCounterY = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  pixelIndex = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      kernelCounter <= 4'h0;
    end else if (kernelCountReset) begin
      kernelCounter <= 4'h0;
    end else begin
      kernelCounter <= _T_14;
    end
    if (reset) begin
      imageCounterX <= 2'h0;
    end else if (imageCounterXReset) begin
      imageCounterX <= 2'h0;
    end else begin
      imageCounterX <= _T_20;
    end
    if (reset) begin
      imageCounterY <= 2'h0;
    end else if (imageCounterXReset) begin
      if (_T_21) begin
        imageCounterY <= 2'h0;
      end else begin
        imageCounterY <= _T_23;
      end
    end
    if (reset) begin
      pixelIndex <= 32'h0;
    end else if (kernelCountReset) begin
      if (_T_1028) begin
        pixelIndex <= 32'h0;
      end else begin
        pixelIndex <= _T_1026;
      end
    end
  end
endmodule
module VideoBuffer(
  input         clock,
  input         reset,
  input  [3:0]  io_pixelVal_in_0_0,
  input  [3:0]  io_pixelVal_in_0_1,
  input  [3:0]  io_pixelVal_in_0_2,
  input  [3:0]  io_pixelVal_in_0_3,
  input  [3:0]  io_pixelVal_in_0_4,
  input  [3:0]  io_pixelVal_in_0_5,
  input  [3:0]  io_pixelVal_in_0_6,
  input  [3:0]  io_pixelVal_in_0_7,
  input  [3:0]  io_pixelVal_in_1_0,
  input  [3:0]  io_pixelVal_in_1_1,
  input  [3:0]  io_pixelVal_in_1_2,
  input  [3:0]  io_pixelVal_in_1_3,
  input  [3:0]  io_pixelVal_in_1_4,
  input  [3:0]  io_pixelVal_in_1_5,
  input  [3:0]  io_pixelVal_in_1_6,
  input  [3:0]  io_pixelVal_in_1_7,
  input  [3:0]  io_pixelVal_in_2_0,
  input  [3:0]  io_pixelVal_in_2_1,
  input  [3:0]  io_pixelVal_in_2_2,
  input  [3:0]  io_pixelVal_in_2_3,
  input  [3:0]  io_pixelVal_in_2_4,
  input  [3:0]  io_pixelVal_in_2_5,
  input  [3:0]  io_pixelVal_in_2_6,
  input  [3:0]  io_pixelVal_in_2_7,
  input         io_valid_in,
  input  [10:0] io_rowIndex,
  input  [10:0] io_colIndex,
  output [3:0]  io_pixelVal_out_0,
  output [3:0]  io_pixelVal_out_1,
  output [3:0]  io_pixelVal_out_2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] image_0_0; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_1; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_2; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_3; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_4; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_5; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_6; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_7; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_8; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_9; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_10; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_11; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_12; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_13; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_14; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_15; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_16; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_17; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_18; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_19; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_20; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_21; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_22; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_23; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_24; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_25; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_26; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_27; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_28; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_29; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_30; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_31; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_32; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_33; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_34; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_35; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_36; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_37; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_38; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_39; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_40; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_41; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_42; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_43; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_44; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_45; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_46; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_47; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_48; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_49; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_50; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_51; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_52; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_53; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_54; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_55; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_56; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_57; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_58; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_59; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_60; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_61; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_62; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_63; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_64; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_65; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_66; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_67; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_68; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_69; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_70; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_71; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_72; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_73; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_74; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_75; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_76; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_77; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_78; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_79; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_80; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_81; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_82; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_83; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_84; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_85; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_86; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_87; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_88; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_89; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_90; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_91; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_92; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_93; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_94; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_95; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_96; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_97; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_98; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_99; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_100; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_101; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_102; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_103; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_104; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_105; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_106; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_107; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_108; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_109; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_110; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_111; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_112; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_113; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_114; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_115; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_116; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_117; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_118; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_119; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_120; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_121; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_122; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_123; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_124; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_125; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_126; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_127; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_128; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_129; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_130; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_131; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_132; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_133; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_134; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_135; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_136; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_137; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_138; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_139; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_140; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_141; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_142; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_143; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_144; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_145; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_146; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_147; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_148; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_149; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_150; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_151; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_152; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_153; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_154; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_155; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_156; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_157; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_158; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_159; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_160; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_161; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_162; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_163; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_164; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_165; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_166; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_167; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_168; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_169; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_170; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_171; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_172; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_173; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_174; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_175; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_176; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_177; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_178; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_179; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_180; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_181; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_182; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_183; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_184; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_185; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_186; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_187; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_188; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_189; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_190; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_191; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_1_0; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_1; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_2; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_3; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_4; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_5; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_6; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_7; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_8; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_9; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_10; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_11; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_12; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_13; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_14; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_15; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_16; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_17; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_18; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_19; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_20; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_21; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_22; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_23; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_24; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_25; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_26; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_27; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_28; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_29; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_30; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_31; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_32; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_33; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_34; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_35; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_36; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_37; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_38; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_39; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_40; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_41; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_42; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_43; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_44; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_45; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_46; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_47; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_48; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_49; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_50; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_51; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_52; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_53; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_54; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_55; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_56; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_57; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_58; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_59; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_60; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_61; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_62; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_63; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_64; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_65; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_66; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_67; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_68; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_69; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_70; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_71; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_72; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_73; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_74; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_75; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_76; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_77; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_78; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_79; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_80; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_81; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_82; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_83; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_84; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_85; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_86; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_87; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_88; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_89; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_90; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_91; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_92; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_93; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_94; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_95; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_96; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_97; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_98; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_99; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_100; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_101; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_102; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_103; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_104; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_105; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_106; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_107; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_108; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_109; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_110; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_111; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_112; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_113; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_114; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_115; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_116; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_117; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_118; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_119; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_120; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_121; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_122; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_123; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_124; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_125; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_126; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_127; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_128; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_129; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_130; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_131; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_132; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_133; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_134; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_135; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_136; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_137; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_138; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_139; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_140; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_141; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_142; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_143; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_144; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_145; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_146; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_147; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_148; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_149; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_150; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_151; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_152; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_153; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_154; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_155; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_156; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_157; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_158; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_159; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_160; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_161; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_162; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_163; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_164; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_165; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_166; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_167; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_168; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_169; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_170; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_171; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_172; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_173; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_174; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_175; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_176; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_177; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_178; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_179; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_180; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_181; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_182; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_183; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_184; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_185; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_186; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_187; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_188; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_189; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_190; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_191; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_2_0; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_1; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_2; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_3; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_4; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_5; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_6; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_7; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_8; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_9; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_10; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_11; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_12; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_13; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_14; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_15; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_16; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_17; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_18; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_19; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_20; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_21; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_22; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_23; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_24; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_25; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_26; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_27; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_28; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_29; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_30; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_31; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_32; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_33; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_34; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_35; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_36; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_37; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_38; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_39; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_40; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_41; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_42; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_43; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_44; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_45; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_46; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_47; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_48; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_49; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_50; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_51; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_52; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_53; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_54; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_55; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_56; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_57; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_58; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_59; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_60; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_61; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_62; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_63; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_64; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_65; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_66; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_67; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_68; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_69; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_70; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_71; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_72; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_73; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_74; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_75; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_76; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_77; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_78; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_79; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_80; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_81; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_82; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_83; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_84; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_85; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_86; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_87; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_88; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_89; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_90; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_91; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_92; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_93; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_94; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_95; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_96; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_97; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_98; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_99; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_100; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_101; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_102; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_103; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_104; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_105; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_106; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_107; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_108; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_109; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_110; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_111; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_112; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_113; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_114; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_115; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_116; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_117; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_118; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_119; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_120; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_121; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_122; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_123; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_124; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_125; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_126; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_127; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_128; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_129; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_130; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_131; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_132; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_133; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_134; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_135; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_136; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_137; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_138; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_139; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_140; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_141; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_142; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_143; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_144; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_145; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_146; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_147; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_148; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_149; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_150; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_151; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_152; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_153; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_154; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_155; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_156; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_157; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_158; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_159; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_160; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_161; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_162; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_163; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_164; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_165; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_166; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_167; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_168; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_169; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_170; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_171; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_172; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_173; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_174; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_175; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_176; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_177; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_178; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_179; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_180; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_181; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_182; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_183; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_184; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_185; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_186; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_187; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_188; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_189; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_190; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_191; // @[VideoBuffer.scala 21:25]
  reg [31:0] pixelIndex; // @[VideoBuffer.scala 24:33]
  wire [15:0] _T_3 = io_rowIndex * 11'h10; // @[VideoBuffer.scala 27:54]
  wire [15:0] _GEN_5761 = {{5'd0}, io_colIndex}; // @[VideoBuffer.scala 27:69]
  wire [15:0] _T_5 = _T_3 + _GEN_5761; // @[VideoBuffer.scala 27:69]
  wire [3:0] _GEN_1 = 8'h1 == _T_5[7:0] ? image_0_1 : image_0_0; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2 = 8'h2 == _T_5[7:0] ? image_0_2 : _GEN_1; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3 = 8'h3 == _T_5[7:0] ? image_0_3 : _GEN_2; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4 = 8'h4 == _T_5[7:0] ? image_0_4 : _GEN_3; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_5 = 8'h5 == _T_5[7:0] ? image_0_5 : _GEN_4; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_6 = 8'h6 == _T_5[7:0] ? image_0_6 : _GEN_5; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_7 = 8'h7 == _T_5[7:0] ? image_0_7 : _GEN_6; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_8 = 8'h8 == _T_5[7:0] ? image_0_8 : _GEN_7; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_9 = 8'h9 == _T_5[7:0] ? image_0_9 : _GEN_8; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_10 = 8'ha == _T_5[7:0] ? image_0_10 : _GEN_9; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_11 = 8'hb == _T_5[7:0] ? image_0_11 : _GEN_10; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_12 = 8'hc == _T_5[7:0] ? image_0_12 : _GEN_11; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_13 = 8'hd == _T_5[7:0] ? image_0_13 : _GEN_12; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_14 = 8'he == _T_5[7:0] ? image_0_14 : _GEN_13; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_15 = 8'hf == _T_5[7:0] ? image_0_15 : _GEN_14; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_16 = 8'h10 == _T_5[7:0] ? image_0_16 : _GEN_15; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_17 = 8'h11 == _T_5[7:0] ? image_0_17 : _GEN_16; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_18 = 8'h12 == _T_5[7:0] ? image_0_18 : _GEN_17; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_19 = 8'h13 == _T_5[7:0] ? image_0_19 : _GEN_18; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_20 = 8'h14 == _T_5[7:0] ? image_0_20 : _GEN_19; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_21 = 8'h15 == _T_5[7:0] ? image_0_21 : _GEN_20; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_22 = 8'h16 == _T_5[7:0] ? image_0_22 : _GEN_21; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_23 = 8'h17 == _T_5[7:0] ? image_0_23 : _GEN_22; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_24 = 8'h18 == _T_5[7:0] ? image_0_24 : _GEN_23; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_25 = 8'h19 == _T_5[7:0] ? image_0_25 : _GEN_24; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_26 = 8'h1a == _T_5[7:0] ? image_0_26 : _GEN_25; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_27 = 8'h1b == _T_5[7:0] ? image_0_27 : _GEN_26; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_28 = 8'h1c == _T_5[7:0] ? image_0_28 : _GEN_27; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_29 = 8'h1d == _T_5[7:0] ? image_0_29 : _GEN_28; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_30 = 8'h1e == _T_5[7:0] ? image_0_30 : _GEN_29; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_31 = 8'h1f == _T_5[7:0] ? image_0_31 : _GEN_30; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_32 = 8'h20 == _T_5[7:0] ? image_0_32 : _GEN_31; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_33 = 8'h21 == _T_5[7:0] ? image_0_33 : _GEN_32; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_34 = 8'h22 == _T_5[7:0] ? image_0_34 : _GEN_33; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_35 = 8'h23 == _T_5[7:0] ? image_0_35 : _GEN_34; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_36 = 8'h24 == _T_5[7:0] ? image_0_36 : _GEN_35; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_37 = 8'h25 == _T_5[7:0] ? image_0_37 : _GEN_36; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_38 = 8'h26 == _T_5[7:0] ? image_0_38 : _GEN_37; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_39 = 8'h27 == _T_5[7:0] ? image_0_39 : _GEN_38; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_40 = 8'h28 == _T_5[7:0] ? image_0_40 : _GEN_39; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_41 = 8'h29 == _T_5[7:0] ? image_0_41 : _GEN_40; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_42 = 8'h2a == _T_5[7:0] ? image_0_42 : _GEN_41; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_43 = 8'h2b == _T_5[7:0] ? image_0_43 : _GEN_42; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_44 = 8'h2c == _T_5[7:0] ? image_0_44 : _GEN_43; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_45 = 8'h2d == _T_5[7:0] ? image_0_45 : _GEN_44; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_46 = 8'h2e == _T_5[7:0] ? image_0_46 : _GEN_45; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_47 = 8'h2f == _T_5[7:0] ? image_0_47 : _GEN_46; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_48 = 8'h30 == _T_5[7:0] ? image_0_48 : _GEN_47; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_49 = 8'h31 == _T_5[7:0] ? image_0_49 : _GEN_48; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_50 = 8'h32 == _T_5[7:0] ? image_0_50 : _GEN_49; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_51 = 8'h33 == _T_5[7:0] ? image_0_51 : _GEN_50; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_52 = 8'h34 == _T_5[7:0] ? image_0_52 : _GEN_51; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_53 = 8'h35 == _T_5[7:0] ? image_0_53 : _GEN_52; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_54 = 8'h36 == _T_5[7:0] ? image_0_54 : _GEN_53; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_55 = 8'h37 == _T_5[7:0] ? image_0_55 : _GEN_54; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_56 = 8'h38 == _T_5[7:0] ? image_0_56 : _GEN_55; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_57 = 8'h39 == _T_5[7:0] ? image_0_57 : _GEN_56; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_58 = 8'h3a == _T_5[7:0] ? image_0_58 : _GEN_57; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_59 = 8'h3b == _T_5[7:0] ? image_0_59 : _GEN_58; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_60 = 8'h3c == _T_5[7:0] ? image_0_60 : _GEN_59; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_61 = 8'h3d == _T_5[7:0] ? image_0_61 : _GEN_60; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_62 = 8'h3e == _T_5[7:0] ? image_0_62 : _GEN_61; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_63 = 8'h3f == _T_5[7:0] ? image_0_63 : _GEN_62; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_64 = 8'h40 == _T_5[7:0] ? image_0_64 : _GEN_63; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_65 = 8'h41 == _T_5[7:0] ? image_0_65 : _GEN_64; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_66 = 8'h42 == _T_5[7:0] ? image_0_66 : _GEN_65; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_67 = 8'h43 == _T_5[7:0] ? image_0_67 : _GEN_66; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_68 = 8'h44 == _T_5[7:0] ? image_0_68 : _GEN_67; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_69 = 8'h45 == _T_5[7:0] ? image_0_69 : _GEN_68; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_70 = 8'h46 == _T_5[7:0] ? image_0_70 : _GEN_69; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_71 = 8'h47 == _T_5[7:0] ? image_0_71 : _GEN_70; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_72 = 8'h48 == _T_5[7:0] ? image_0_72 : _GEN_71; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_73 = 8'h49 == _T_5[7:0] ? image_0_73 : _GEN_72; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_74 = 8'h4a == _T_5[7:0] ? image_0_74 : _GEN_73; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_75 = 8'h4b == _T_5[7:0] ? image_0_75 : _GEN_74; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_76 = 8'h4c == _T_5[7:0] ? image_0_76 : _GEN_75; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_77 = 8'h4d == _T_5[7:0] ? image_0_77 : _GEN_76; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_78 = 8'h4e == _T_5[7:0] ? image_0_78 : _GEN_77; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_79 = 8'h4f == _T_5[7:0] ? image_0_79 : _GEN_78; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_80 = 8'h50 == _T_5[7:0] ? image_0_80 : _GEN_79; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_81 = 8'h51 == _T_5[7:0] ? image_0_81 : _GEN_80; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_82 = 8'h52 == _T_5[7:0] ? image_0_82 : _GEN_81; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_83 = 8'h53 == _T_5[7:0] ? image_0_83 : _GEN_82; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_84 = 8'h54 == _T_5[7:0] ? image_0_84 : _GEN_83; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_85 = 8'h55 == _T_5[7:0] ? image_0_85 : _GEN_84; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_86 = 8'h56 == _T_5[7:0] ? image_0_86 : _GEN_85; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_87 = 8'h57 == _T_5[7:0] ? image_0_87 : _GEN_86; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_88 = 8'h58 == _T_5[7:0] ? image_0_88 : _GEN_87; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_89 = 8'h59 == _T_5[7:0] ? image_0_89 : _GEN_88; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_90 = 8'h5a == _T_5[7:0] ? image_0_90 : _GEN_89; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_91 = 8'h5b == _T_5[7:0] ? image_0_91 : _GEN_90; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_92 = 8'h5c == _T_5[7:0] ? image_0_92 : _GEN_91; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_93 = 8'h5d == _T_5[7:0] ? image_0_93 : _GEN_92; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_94 = 8'h5e == _T_5[7:0] ? image_0_94 : _GEN_93; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_95 = 8'h5f == _T_5[7:0] ? image_0_95 : _GEN_94; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_96 = 8'h60 == _T_5[7:0] ? image_0_96 : _GEN_95; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_97 = 8'h61 == _T_5[7:0] ? image_0_97 : _GEN_96; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_98 = 8'h62 == _T_5[7:0] ? image_0_98 : _GEN_97; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_99 = 8'h63 == _T_5[7:0] ? image_0_99 : _GEN_98; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_100 = 8'h64 == _T_5[7:0] ? image_0_100 : _GEN_99; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_101 = 8'h65 == _T_5[7:0] ? image_0_101 : _GEN_100; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_102 = 8'h66 == _T_5[7:0] ? image_0_102 : _GEN_101; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_103 = 8'h67 == _T_5[7:0] ? image_0_103 : _GEN_102; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_104 = 8'h68 == _T_5[7:0] ? image_0_104 : _GEN_103; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_105 = 8'h69 == _T_5[7:0] ? image_0_105 : _GEN_104; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_106 = 8'h6a == _T_5[7:0] ? image_0_106 : _GEN_105; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_107 = 8'h6b == _T_5[7:0] ? image_0_107 : _GEN_106; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_108 = 8'h6c == _T_5[7:0] ? image_0_108 : _GEN_107; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_109 = 8'h6d == _T_5[7:0] ? image_0_109 : _GEN_108; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_110 = 8'h6e == _T_5[7:0] ? image_0_110 : _GEN_109; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_111 = 8'h6f == _T_5[7:0] ? image_0_111 : _GEN_110; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_112 = 8'h70 == _T_5[7:0] ? image_0_112 : _GEN_111; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_113 = 8'h71 == _T_5[7:0] ? image_0_113 : _GEN_112; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_114 = 8'h72 == _T_5[7:0] ? image_0_114 : _GEN_113; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_115 = 8'h73 == _T_5[7:0] ? image_0_115 : _GEN_114; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_116 = 8'h74 == _T_5[7:0] ? image_0_116 : _GEN_115; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_117 = 8'h75 == _T_5[7:0] ? image_0_117 : _GEN_116; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_118 = 8'h76 == _T_5[7:0] ? image_0_118 : _GEN_117; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_119 = 8'h77 == _T_5[7:0] ? image_0_119 : _GEN_118; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_120 = 8'h78 == _T_5[7:0] ? image_0_120 : _GEN_119; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_121 = 8'h79 == _T_5[7:0] ? image_0_121 : _GEN_120; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_122 = 8'h7a == _T_5[7:0] ? image_0_122 : _GEN_121; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_123 = 8'h7b == _T_5[7:0] ? image_0_123 : _GEN_122; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_124 = 8'h7c == _T_5[7:0] ? image_0_124 : _GEN_123; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_125 = 8'h7d == _T_5[7:0] ? image_0_125 : _GEN_124; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_126 = 8'h7e == _T_5[7:0] ? image_0_126 : _GEN_125; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_127 = 8'h7f == _T_5[7:0] ? image_0_127 : _GEN_126; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_128 = 8'h80 == _T_5[7:0] ? image_0_128 : _GEN_127; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_129 = 8'h81 == _T_5[7:0] ? image_0_129 : _GEN_128; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_130 = 8'h82 == _T_5[7:0] ? image_0_130 : _GEN_129; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_131 = 8'h83 == _T_5[7:0] ? image_0_131 : _GEN_130; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_132 = 8'h84 == _T_5[7:0] ? image_0_132 : _GEN_131; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_133 = 8'h85 == _T_5[7:0] ? image_0_133 : _GEN_132; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_134 = 8'h86 == _T_5[7:0] ? image_0_134 : _GEN_133; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_135 = 8'h87 == _T_5[7:0] ? image_0_135 : _GEN_134; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_136 = 8'h88 == _T_5[7:0] ? image_0_136 : _GEN_135; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_137 = 8'h89 == _T_5[7:0] ? image_0_137 : _GEN_136; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_138 = 8'h8a == _T_5[7:0] ? image_0_138 : _GEN_137; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_139 = 8'h8b == _T_5[7:0] ? image_0_139 : _GEN_138; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_140 = 8'h8c == _T_5[7:0] ? image_0_140 : _GEN_139; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_141 = 8'h8d == _T_5[7:0] ? image_0_141 : _GEN_140; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_142 = 8'h8e == _T_5[7:0] ? image_0_142 : _GEN_141; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_143 = 8'h8f == _T_5[7:0] ? image_0_143 : _GEN_142; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_144 = 8'h90 == _T_5[7:0] ? image_0_144 : _GEN_143; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_145 = 8'h91 == _T_5[7:0] ? image_0_145 : _GEN_144; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_146 = 8'h92 == _T_5[7:0] ? image_0_146 : _GEN_145; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_147 = 8'h93 == _T_5[7:0] ? image_0_147 : _GEN_146; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_148 = 8'h94 == _T_5[7:0] ? image_0_148 : _GEN_147; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_149 = 8'h95 == _T_5[7:0] ? image_0_149 : _GEN_148; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_150 = 8'h96 == _T_5[7:0] ? image_0_150 : _GEN_149; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_151 = 8'h97 == _T_5[7:0] ? image_0_151 : _GEN_150; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_152 = 8'h98 == _T_5[7:0] ? image_0_152 : _GEN_151; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_153 = 8'h99 == _T_5[7:0] ? image_0_153 : _GEN_152; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_154 = 8'h9a == _T_5[7:0] ? image_0_154 : _GEN_153; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_155 = 8'h9b == _T_5[7:0] ? image_0_155 : _GEN_154; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_156 = 8'h9c == _T_5[7:0] ? image_0_156 : _GEN_155; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_157 = 8'h9d == _T_5[7:0] ? image_0_157 : _GEN_156; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_158 = 8'h9e == _T_5[7:0] ? image_0_158 : _GEN_157; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_159 = 8'h9f == _T_5[7:0] ? image_0_159 : _GEN_158; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_160 = 8'ha0 == _T_5[7:0] ? image_0_160 : _GEN_159; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_161 = 8'ha1 == _T_5[7:0] ? image_0_161 : _GEN_160; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_162 = 8'ha2 == _T_5[7:0] ? image_0_162 : _GEN_161; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_163 = 8'ha3 == _T_5[7:0] ? image_0_163 : _GEN_162; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_164 = 8'ha4 == _T_5[7:0] ? image_0_164 : _GEN_163; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_165 = 8'ha5 == _T_5[7:0] ? image_0_165 : _GEN_164; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_166 = 8'ha6 == _T_5[7:0] ? image_0_166 : _GEN_165; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_167 = 8'ha7 == _T_5[7:0] ? image_0_167 : _GEN_166; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_168 = 8'ha8 == _T_5[7:0] ? image_0_168 : _GEN_167; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_169 = 8'ha9 == _T_5[7:0] ? image_0_169 : _GEN_168; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_170 = 8'haa == _T_5[7:0] ? image_0_170 : _GEN_169; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_171 = 8'hab == _T_5[7:0] ? image_0_171 : _GEN_170; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_172 = 8'hac == _T_5[7:0] ? image_0_172 : _GEN_171; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_173 = 8'had == _T_5[7:0] ? image_0_173 : _GEN_172; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_174 = 8'hae == _T_5[7:0] ? image_0_174 : _GEN_173; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_175 = 8'haf == _T_5[7:0] ? image_0_175 : _GEN_174; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_176 = 8'hb0 == _T_5[7:0] ? image_0_176 : _GEN_175; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_177 = 8'hb1 == _T_5[7:0] ? image_0_177 : _GEN_176; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_178 = 8'hb2 == _T_5[7:0] ? image_0_178 : _GEN_177; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_179 = 8'hb3 == _T_5[7:0] ? image_0_179 : _GEN_178; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_180 = 8'hb4 == _T_5[7:0] ? image_0_180 : _GEN_179; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_181 = 8'hb5 == _T_5[7:0] ? image_0_181 : _GEN_180; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_182 = 8'hb6 == _T_5[7:0] ? image_0_182 : _GEN_181; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_183 = 8'hb7 == _T_5[7:0] ? image_0_183 : _GEN_182; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_184 = 8'hb8 == _T_5[7:0] ? image_0_184 : _GEN_183; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_185 = 8'hb9 == _T_5[7:0] ? image_0_185 : _GEN_184; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_186 = 8'hba == _T_5[7:0] ? image_0_186 : _GEN_185; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_187 = 8'hbb == _T_5[7:0] ? image_0_187 : _GEN_186; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_188 = 8'hbc == _T_5[7:0] ? image_0_188 : _GEN_187; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_189 = 8'hbd == _T_5[7:0] ? image_0_189 : _GEN_188; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_190 = 8'hbe == _T_5[7:0] ? image_0_190 : _GEN_189; // @[VideoBuffer.scala 27:30]
  wire [32:0] _T_7 = {{1'd0}, pixelIndex}; // @[VideoBuffer.scala 31:35]
  wire [31:0] _T_11 = pixelIndex + 32'h1; // @[VideoBuffer.scala 31:35]
  wire [31:0] _T_14 = pixelIndex + 32'h2; // @[VideoBuffer.scala 31:35]
  wire [31:0] _T_17 = pixelIndex + 32'h3; // @[VideoBuffer.scala 31:35]
  wire [31:0] _T_20 = pixelIndex + 32'h4; // @[VideoBuffer.scala 31:35]
  wire [31:0] _T_23 = pixelIndex + 32'h5; // @[VideoBuffer.scala 31:35]
  wire [31:0] _T_26 = pixelIndex + 32'h6; // @[VideoBuffer.scala 31:35]
  wire [31:0] _T_29 = pixelIndex + 32'h7; // @[VideoBuffer.scala 31:35]
  wire [3:0] _GEN_1921 = 8'h1 == _T_5[7:0] ? image_1_1 : image_1_0; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1922 = 8'h2 == _T_5[7:0] ? image_1_2 : _GEN_1921; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1923 = 8'h3 == _T_5[7:0] ? image_1_3 : _GEN_1922; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1924 = 8'h4 == _T_5[7:0] ? image_1_4 : _GEN_1923; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1925 = 8'h5 == _T_5[7:0] ? image_1_5 : _GEN_1924; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1926 = 8'h6 == _T_5[7:0] ? image_1_6 : _GEN_1925; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1927 = 8'h7 == _T_5[7:0] ? image_1_7 : _GEN_1926; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1928 = 8'h8 == _T_5[7:0] ? image_1_8 : _GEN_1927; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1929 = 8'h9 == _T_5[7:0] ? image_1_9 : _GEN_1928; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1930 = 8'ha == _T_5[7:0] ? image_1_10 : _GEN_1929; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1931 = 8'hb == _T_5[7:0] ? image_1_11 : _GEN_1930; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1932 = 8'hc == _T_5[7:0] ? image_1_12 : _GEN_1931; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1933 = 8'hd == _T_5[7:0] ? image_1_13 : _GEN_1932; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1934 = 8'he == _T_5[7:0] ? image_1_14 : _GEN_1933; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1935 = 8'hf == _T_5[7:0] ? image_1_15 : _GEN_1934; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1936 = 8'h10 == _T_5[7:0] ? image_1_16 : _GEN_1935; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1937 = 8'h11 == _T_5[7:0] ? image_1_17 : _GEN_1936; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1938 = 8'h12 == _T_5[7:0] ? image_1_18 : _GEN_1937; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1939 = 8'h13 == _T_5[7:0] ? image_1_19 : _GEN_1938; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1940 = 8'h14 == _T_5[7:0] ? image_1_20 : _GEN_1939; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1941 = 8'h15 == _T_5[7:0] ? image_1_21 : _GEN_1940; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1942 = 8'h16 == _T_5[7:0] ? image_1_22 : _GEN_1941; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1943 = 8'h17 == _T_5[7:0] ? image_1_23 : _GEN_1942; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1944 = 8'h18 == _T_5[7:0] ? image_1_24 : _GEN_1943; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1945 = 8'h19 == _T_5[7:0] ? image_1_25 : _GEN_1944; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1946 = 8'h1a == _T_5[7:0] ? image_1_26 : _GEN_1945; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1947 = 8'h1b == _T_5[7:0] ? image_1_27 : _GEN_1946; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1948 = 8'h1c == _T_5[7:0] ? image_1_28 : _GEN_1947; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1949 = 8'h1d == _T_5[7:0] ? image_1_29 : _GEN_1948; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1950 = 8'h1e == _T_5[7:0] ? image_1_30 : _GEN_1949; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1951 = 8'h1f == _T_5[7:0] ? image_1_31 : _GEN_1950; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1952 = 8'h20 == _T_5[7:0] ? image_1_32 : _GEN_1951; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1953 = 8'h21 == _T_5[7:0] ? image_1_33 : _GEN_1952; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1954 = 8'h22 == _T_5[7:0] ? image_1_34 : _GEN_1953; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1955 = 8'h23 == _T_5[7:0] ? image_1_35 : _GEN_1954; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1956 = 8'h24 == _T_5[7:0] ? image_1_36 : _GEN_1955; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1957 = 8'h25 == _T_5[7:0] ? image_1_37 : _GEN_1956; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1958 = 8'h26 == _T_5[7:0] ? image_1_38 : _GEN_1957; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1959 = 8'h27 == _T_5[7:0] ? image_1_39 : _GEN_1958; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1960 = 8'h28 == _T_5[7:0] ? image_1_40 : _GEN_1959; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1961 = 8'h29 == _T_5[7:0] ? image_1_41 : _GEN_1960; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1962 = 8'h2a == _T_5[7:0] ? image_1_42 : _GEN_1961; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1963 = 8'h2b == _T_5[7:0] ? image_1_43 : _GEN_1962; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1964 = 8'h2c == _T_5[7:0] ? image_1_44 : _GEN_1963; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1965 = 8'h2d == _T_5[7:0] ? image_1_45 : _GEN_1964; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1966 = 8'h2e == _T_5[7:0] ? image_1_46 : _GEN_1965; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1967 = 8'h2f == _T_5[7:0] ? image_1_47 : _GEN_1966; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1968 = 8'h30 == _T_5[7:0] ? image_1_48 : _GEN_1967; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1969 = 8'h31 == _T_5[7:0] ? image_1_49 : _GEN_1968; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1970 = 8'h32 == _T_5[7:0] ? image_1_50 : _GEN_1969; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1971 = 8'h33 == _T_5[7:0] ? image_1_51 : _GEN_1970; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1972 = 8'h34 == _T_5[7:0] ? image_1_52 : _GEN_1971; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1973 = 8'h35 == _T_5[7:0] ? image_1_53 : _GEN_1972; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1974 = 8'h36 == _T_5[7:0] ? image_1_54 : _GEN_1973; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1975 = 8'h37 == _T_5[7:0] ? image_1_55 : _GEN_1974; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1976 = 8'h38 == _T_5[7:0] ? image_1_56 : _GEN_1975; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1977 = 8'h39 == _T_5[7:0] ? image_1_57 : _GEN_1976; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1978 = 8'h3a == _T_5[7:0] ? image_1_58 : _GEN_1977; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1979 = 8'h3b == _T_5[7:0] ? image_1_59 : _GEN_1978; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1980 = 8'h3c == _T_5[7:0] ? image_1_60 : _GEN_1979; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1981 = 8'h3d == _T_5[7:0] ? image_1_61 : _GEN_1980; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1982 = 8'h3e == _T_5[7:0] ? image_1_62 : _GEN_1981; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1983 = 8'h3f == _T_5[7:0] ? image_1_63 : _GEN_1982; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1984 = 8'h40 == _T_5[7:0] ? image_1_64 : _GEN_1983; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1985 = 8'h41 == _T_5[7:0] ? image_1_65 : _GEN_1984; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1986 = 8'h42 == _T_5[7:0] ? image_1_66 : _GEN_1985; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1987 = 8'h43 == _T_5[7:0] ? image_1_67 : _GEN_1986; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1988 = 8'h44 == _T_5[7:0] ? image_1_68 : _GEN_1987; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1989 = 8'h45 == _T_5[7:0] ? image_1_69 : _GEN_1988; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1990 = 8'h46 == _T_5[7:0] ? image_1_70 : _GEN_1989; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1991 = 8'h47 == _T_5[7:0] ? image_1_71 : _GEN_1990; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1992 = 8'h48 == _T_5[7:0] ? image_1_72 : _GEN_1991; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1993 = 8'h49 == _T_5[7:0] ? image_1_73 : _GEN_1992; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1994 = 8'h4a == _T_5[7:0] ? image_1_74 : _GEN_1993; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1995 = 8'h4b == _T_5[7:0] ? image_1_75 : _GEN_1994; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1996 = 8'h4c == _T_5[7:0] ? image_1_76 : _GEN_1995; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1997 = 8'h4d == _T_5[7:0] ? image_1_77 : _GEN_1996; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1998 = 8'h4e == _T_5[7:0] ? image_1_78 : _GEN_1997; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1999 = 8'h4f == _T_5[7:0] ? image_1_79 : _GEN_1998; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2000 = 8'h50 == _T_5[7:0] ? image_1_80 : _GEN_1999; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2001 = 8'h51 == _T_5[7:0] ? image_1_81 : _GEN_2000; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2002 = 8'h52 == _T_5[7:0] ? image_1_82 : _GEN_2001; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2003 = 8'h53 == _T_5[7:0] ? image_1_83 : _GEN_2002; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2004 = 8'h54 == _T_5[7:0] ? image_1_84 : _GEN_2003; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2005 = 8'h55 == _T_5[7:0] ? image_1_85 : _GEN_2004; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2006 = 8'h56 == _T_5[7:0] ? image_1_86 : _GEN_2005; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2007 = 8'h57 == _T_5[7:0] ? image_1_87 : _GEN_2006; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2008 = 8'h58 == _T_5[7:0] ? image_1_88 : _GEN_2007; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2009 = 8'h59 == _T_5[7:0] ? image_1_89 : _GEN_2008; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2010 = 8'h5a == _T_5[7:0] ? image_1_90 : _GEN_2009; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2011 = 8'h5b == _T_5[7:0] ? image_1_91 : _GEN_2010; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2012 = 8'h5c == _T_5[7:0] ? image_1_92 : _GEN_2011; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2013 = 8'h5d == _T_5[7:0] ? image_1_93 : _GEN_2012; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2014 = 8'h5e == _T_5[7:0] ? image_1_94 : _GEN_2013; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2015 = 8'h5f == _T_5[7:0] ? image_1_95 : _GEN_2014; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2016 = 8'h60 == _T_5[7:0] ? image_1_96 : _GEN_2015; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2017 = 8'h61 == _T_5[7:0] ? image_1_97 : _GEN_2016; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2018 = 8'h62 == _T_5[7:0] ? image_1_98 : _GEN_2017; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2019 = 8'h63 == _T_5[7:0] ? image_1_99 : _GEN_2018; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2020 = 8'h64 == _T_5[7:0] ? image_1_100 : _GEN_2019; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2021 = 8'h65 == _T_5[7:0] ? image_1_101 : _GEN_2020; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2022 = 8'h66 == _T_5[7:0] ? image_1_102 : _GEN_2021; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2023 = 8'h67 == _T_5[7:0] ? image_1_103 : _GEN_2022; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2024 = 8'h68 == _T_5[7:0] ? image_1_104 : _GEN_2023; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2025 = 8'h69 == _T_5[7:0] ? image_1_105 : _GEN_2024; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2026 = 8'h6a == _T_5[7:0] ? image_1_106 : _GEN_2025; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2027 = 8'h6b == _T_5[7:0] ? image_1_107 : _GEN_2026; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2028 = 8'h6c == _T_5[7:0] ? image_1_108 : _GEN_2027; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2029 = 8'h6d == _T_5[7:0] ? image_1_109 : _GEN_2028; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2030 = 8'h6e == _T_5[7:0] ? image_1_110 : _GEN_2029; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2031 = 8'h6f == _T_5[7:0] ? image_1_111 : _GEN_2030; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2032 = 8'h70 == _T_5[7:0] ? image_1_112 : _GEN_2031; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2033 = 8'h71 == _T_5[7:0] ? image_1_113 : _GEN_2032; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2034 = 8'h72 == _T_5[7:0] ? image_1_114 : _GEN_2033; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2035 = 8'h73 == _T_5[7:0] ? image_1_115 : _GEN_2034; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2036 = 8'h74 == _T_5[7:0] ? image_1_116 : _GEN_2035; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2037 = 8'h75 == _T_5[7:0] ? image_1_117 : _GEN_2036; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2038 = 8'h76 == _T_5[7:0] ? image_1_118 : _GEN_2037; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2039 = 8'h77 == _T_5[7:0] ? image_1_119 : _GEN_2038; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2040 = 8'h78 == _T_5[7:0] ? image_1_120 : _GEN_2039; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2041 = 8'h79 == _T_5[7:0] ? image_1_121 : _GEN_2040; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2042 = 8'h7a == _T_5[7:0] ? image_1_122 : _GEN_2041; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2043 = 8'h7b == _T_5[7:0] ? image_1_123 : _GEN_2042; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2044 = 8'h7c == _T_5[7:0] ? image_1_124 : _GEN_2043; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2045 = 8'h7d == _T_5[7:0] ? image_1_125 : _GEN_2044; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2046 = 8'h7e == _T_5[7:0] ? image_1_126 : _GEN_2045; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2047 = 8'h7f == _T_5[7:0] ? image_1_127 : _GEN_2046; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2048 = 8'h80 == _T_5[7:0] ? image_1_128 : _GEN_2047; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2049 = 8'h81 == _T_5[7:0] ? image_1_129 : _GEN_2048; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2050 = 8'h82 == _T_5[7:0] ? image_1_130 : _GEN_2049; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2051 = 8'h83 == _T_5[7:0] ? image_1_131 : _GEN_2050; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2052 = 8'h84 == _T_5[7:0] ? image_1_132 : _GEN_2051; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2053 = 8'h85 == _T_5[7:0] ? image_1_133 : _GEN_2052; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2054 = 8'h86 == _T_5[7:0] ? image_1_134 : _GEN_2053; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2055 = 8'h87 == _T_5[7:0] ? image_1_135 : _GEN_2054; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2056 = 8'h88 == _T_5[7:0] ? image_1_136 : _GEN_2055; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2057 = 8'h89 == _T_5[7:0] ? image_1_137 : _GEN_2056; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2058 = 8'h8a == _T_5[7:0] ? image_1_138 : _GEN_2057; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2059 = 8'h8b == _T_5[7:0] ? image_1_139 : _GEN_2058; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2060 = 8'h8c == _T_5[7:0] ? image_1_140 : _GEN_2059; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2061 = 8'h8d == _T_5[7:0] ? image_1_141 : _GEN_2060; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2062 = 8'h8e == _T_5[7:0] ? image_1_142 : _GEN_2061; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2063 = 8'h8f == _T_5[7:0] ? image_1_143 : _GEN_2062; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2064 = 8'h90 == _T_5[7:0] ? image_1_144 : _GEN_2063; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2065 = 8'h91 == _T_5[7:0] ? image_1_145 : _GEN_2064; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2066 = 8'h92 == _T_5[7:0] ? image_1_146 : _GEN_2065; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2067 = 8'h93 == _T_5[7:0] ? image_1_147 : _GEN_2066; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2068 = 8'h94 == _T_5[7:0] ? image_1_148 : _GEN_2067; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2069 = 8'h95 == _T_5[7:0] ? image_1_149 : _GEN_2068; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2070 = 8'h96 == _T_5[7:0] ? image_1_150 : _GEN_2069; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2071 = 8'h97 == _T_5[7:0] ? image_1_151 : _GEN_2070; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2072 = 8'h98 == _T_5[7:0] ? image_1_152 : _GEN_2071; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2073 = 8'h99 == _T_5[7:0] ? image_1_153 : _GEN_2072; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2074 = 8'h9a == _T_5[7:0] ? image_1_154 : _GEN_2073; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2075 = 8'h9b == _T_5[7:0] ? image_1_155 : _GEN_2074; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2076 = 8'h9c == _T_5[7:0] ? image_1_156 : _GEN_2075; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2077 = 8'h9d == _T_5[7:0] ? image_1_157 : _GEN_2076; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2078 = 8'h9e == _T_5[7:0] ? image_1_158 : _GEN_2077; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2079 = 8'h9f == _T_5[7:0] ? image_1_159 : _GEN_2078; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2080 = 8'ha0 == _T_5[7:0] ? image_1_160 : _GEN_2079; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2081 = 8'ha1 == _T_5[7:0] ? image_1_161 : _GEN_2080; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2082 = 8'ha2 == _T_5[7:0] ? image_1_162 : _GEN_2081; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2083 = 8'ha3 == _T_5[7:0] ? image_1_163 : _GEN_2082; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2084 = 8'ha4 == _T_5[7:0] ? image_1_164 : _GEN_2083; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2085 = 8'ha5 == _T_5[7:0] ? image_1_165 : _GEN_2084; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2086 = 8'ha6 == _T_5[7:0] ? image_1_166 : _GEN_2085; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2087 = 8'ha7 == _T_5[7:0] ? image_1_167 : _GEN_2086; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2088 = 8'ha8 == _T_5[7:0] ? image_1_168 : _GEN_2087; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2089 = 8'ha9 == _T_5[7:0] ? image_1_169 : _GEN_2088; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2090 = 8'haa == _T_5[7:0] ? image_1_170 : _GEN_2089; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2091 = 8'hab == _T_5[7:0] ? image_1_171 : _GEN_2090; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2092 = 8'hac == _T_5[7:0] ? image_1_172 : _GEN_2091; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2093 = 8'had == _T_5[7:0] ? image_1_173 : _GEN_2092; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2094 = 8'hae == _T_5[7:0] ? image_1_174 : _GEN_2093; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2095 = 8'haf == _T_5[7:0] ? image_1_175 : _GEN_2094; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2096 = 8'hb0 == _T_5[7:0] ? image_1_176 : _GEN_2095; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2097 = 8'hb1 == _T_5[7:0] ? image_1_177 : _GEN_2096; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2098 = 8'hb2 == _T_5[7:0] ? image_1_178 : _GEN_2097; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2099 = 8'hb3 == _T_5[7:0] ? image_1_179 : _GEN_2098; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2100 = 8'hb4 == _T_5[7:0] ? image_1_180 : _GEN_2099; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2101 = 8'hb5 == _T_5[7:0] ? image_1_181 : _GEN_2100; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2102 = 8'hb6 == _T_5[7:0] ? image_1_182 : _GEN_2101; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2103 = 8'hb7 == _T_5[7:0] ? image_1_183 : _GEN_2102; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2104 = 8'hb8 == _T_5[7:0] ? image_1_184 : _GEN_2103; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2105 = 8'hb9 == _T_5[7:0] ? image_1_185 : _GEN_2104; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2106 = 8'hba == _T_5[7:0] ? image_1_186 : _GEN_2105; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2107 = 8'hbb == _T_5[7:0] ? image_1_187 : _GEN_2106; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2108 = 8'hbc == _T_5[7:0] ? image_1_188 : _GEN_2107; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2109 = 8'hbd == _T_5[7:0] ? image_1_189 : _GEN_2108; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2110 = 8'hbe == _T_5[7:0] ? image_1_190 : _GEN_2109; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3841 = 8'h1 == _T_5[7:0] ? image_2_1 : image_2_0; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3842 = 8'h2 == _T_5[7:0] ? image_2_2 : _GEN_3841; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3843 = 8'h3 == _T_5[7:0] ? image_2_3 : _GEN_3842; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3844 = 8'h4 == _T_5[7:0] ? image_2_4 : _GEN_3843; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3845 = 8'h5 == _T_5[7:0] ? image_2_5 : _GEN_3844; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3846 = 8'h6 == _T_5[7:0] ? image_2_6 : _GEN_3845; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3847 = 8'h7 == _T_5[7:0] ? image_2_7 : _GEN_3846; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3848 = 8'h8 == _T_5[7:0] ? image_2_8 : _GEN_3847; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3849 = 8'h9 == _T_5[7:0] ? image_2_9 : _GEN_3848; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3850 = 8'ha == _T_5[7:0] ? image_2_10 : _GEN_3849; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3851 = 8'hb == _T_5[7:0] ? image_2_11 : _GEN_3850; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3852 = 8'hc == _T_5[7:0] ? image_2_12 : _GEN_3851; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3853 = 8'hd == _T_5[7:0] ? image_2_13 : _GEN_3852; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3854 = 8'he == _T_5[7:0] ? image_2_14 : _GEN_3853; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3855 = 8'hf == _T_5[7:0] ? image_2_15 : _GEN_3854; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3856 = 8'h10 == _T_5[7:0] ? image_2_16 : _GEN_3855; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3857 = 8'h11 == _T_5[7:0] ? image_2_17 : _GEN_3856; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3858 = 8'h12 == _T_5[7:0] ? image_2_18 : _GEN_3857; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3859 = 8'h13 == _T_5[7:0] ? image_2_19 : _GEN_3858; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3860 = 8'h14 == _T_5[7:0] ? image_2_20 : _GEN_3859; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3861 = 8'h15 == _T_5[7:0] ? image_2_21 : _GEN_3860; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3862 = 8'h16 == _T_5[7:0] ? image_2_22 : _GEN_3861; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3863 = 8'h17 == _T_5[7:0] ? image_2_23 : _GEN_3862; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3864 = 8'h18 == _T_5[7:0] ? image_2_24 : _GEN_3863; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3865 = 8'h19 == _T_5[7:0] ? image_2_25 : _GEN_3864; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3866 = 8'h1a == _T_5[7:0] ? image_2_26 : _GEN_3865; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3867 = 8'h1b == _T_5[7:0] ? image_2_27 : _GEN_3866; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3868 = 8'h1c == _T_5[7:0] ? image_2_28 : _GEN_3867; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3869 = 8'h1d == _T_5[7:0] ? image_2_29 : _GEN_3868; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3870 = 8'h1e == _T_5[7:0] ? image_2_30 : _GEN_3869; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3871 = 8'h1f == _T_5[7:0] ? image_2_31 : _GEN_3870; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3872 = 8'h20 == _T_5[7:0] ? image_2_32 : _GEN_3871; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3873 = 8'h21 == _T_5[7:0] ? image_2_33 : _GEN_3872; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3874 = 8'h22 == _T_5[7:0] ? image_2_34 : _GEN_3873; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3875 = 8'h23 == _T_5[7:0] ? image_2_35 : _GEN_3874; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3876 = 8'h24 == _T_5[7:0] ? image_2_36 : _GEN_3875; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3877 = 8'h25 == _T_5[7:0] ? image_2_37 : _GEN_3876; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3878 = 8'h26 == _T_5[7:0] ? image_2_38 : _GEN_3877; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3879 = 8'h27 == _T_5[7:0] ? image_2_39 : _GEN_3878; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3880 = 8'h28 == _T_5[7:0] ? image_2_40 : _GEN_3879; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3881 = 8'h29 == _T_5[7:0] ? image_2_41 : _GEN_3880; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3882 = 8'h2a == _T_5[7:0] ? image_2_42 : _GEN_3881; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3883 = 8'h2b == _T_5[7:0] ? image_2_43 : _GEN_3882; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3884 = 8'h2c == _T_5[7:0] ? image_2_44 : _GEN_3883; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3885 = 8'h2d == _T_5[7:0] ? image_2_45 : _GEN_3884; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3886 = 8'h2e == _T_5[7:0] ? image_2_46 : _GEN_3885; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3887 = 8'h2f == _T_5[7:0] ? image_2_47 : _GEN_3886; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3888 = 8'h30 == _T_5[7:0] ? image_2_48 : _GEN_3887; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3889 = 8'h31 == _T_5[7:0] ? image_2_49 : _GEN_3888; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3890 = 8'h32 == _T_5[7:0] ? image_2_50 : _GEN_3889; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3891 = 8'h33 == _T_5[7:0] ? image_2_51 : _GEN_3890; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3892 = 8'h34 == _T_5[7:0] ? image_2_52 : _GEN_3891; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3893 = 8'h35 == _T_5[7:0] ? image_2_53 : _GEN_3892; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3894 = 8'h36 == _T_5[7:0] ? image_2_54 : _GEN_3893; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3895 = 8'h37 == _T_5[7:0] ? image_2_55 : _GEN_3894; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3896 = 8'h38 == _T_5[7:0] ? image_2_56 : _GEN_3895; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3897 = 8'h39 == _T_5[7:0] ? image_2_57 : _GEN_3896; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3898 = 8'h3a == _T_5[7:0] ? image_2_58 : _GEN_3897; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3899 = 8'h3b == _T_5[7:0] ? image_2_59 : _GEN_3898; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3900 = 8'h3c == _T_5[7:0] ? image_2_60 : _GEN_3899; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3901 = 8'h3d == _T_5[7:0] ? image_2_61 : _GEN_3900; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3902 = 8'h3e == _T_5[7:0] ? image_2_62 : _GEN_3901; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3903 = 8'h3f == _T_5[7:0] ? image_2_63 : _GEN_3902; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3904 = 8'h40 == _T_5[7:0] ? image_2_64 : _GEN_3903; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3905 = 8'h41 == _T_5[7:0] ? image_2_65 : _GEN_3904; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3906 = 8'h42 == _T_5[7:0] ? image_2_66 : _GEN_3905; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3907 = 8'h43 == _T_5[7:0] ? image_2_67 : _GEN_3906; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3908 = 8'h44 == _T_5[7:0] ? image_2_68 : _GEN_3907; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3909 = 8'h45 == _T_5[7:0] ? image_2_69 : _GEN_3908; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3910 = 8'h46 == _T_5[7:0] ? image_2_70 : _GEN_3909; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3911 = 8'h47 == _T_5[7:0] ? image_2_71 : _GEN_3910; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3912 = 8'h48 == _T_5[7:0] ? image_2_72 : _GEN_3911; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3913 = 8'h49 == _T_5[7:0] ? image_2_73 : _GEN_3912; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3914 = 8'h4a == _T_5[7:0] ? image_2_74 : _GEN_3913; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3915 = 8'h4b == _T_5[7:0] ? image_2_75 : _GEN_3914; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3916 = 8'h4c == _T_5[7:0] ? image_2_76 : _GEN_3915; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3917 = 8'h4d == _T_5[7:0] ? image_2_77 : _GEN_3916; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3918 = 8'h4e == _T_5[7:0] ? image_2_78 : _GEN_3917; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3919 = 8'h4f == _T_5[7:0] ? image_2_79 : _GEN_3918; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3920 = 8'h50 == _T_5[7:0] ? image_2_80 : _GEN_3919; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3921 = 8'h51 == _T_5[7:0] ? image_2_81 : _GEN_3920; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3922 = 8'h52 == _T_5[7:0] ? image_2_82 : _GEN_3921; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3923 = 8'h53 == _T_5[7:0] ? image_2_83 : _GEN_3922; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3924 = 8'h54 == _T_5[7:0] ? image_2_84 : _GEN_3923; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3925 = 8'h55 == _T_5[7:0] ? image_2_85 : _GEN_3924; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3926 = 8'h56 == _T_5[7:0] ? image_2_86 : _GEN_3925; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3927 = 8'h57 == _T_5[7:0] ? image_2_87 : _GEN_3926; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3928 = 8'h58 == _T_5[7:0] ? image_2_88 : _GEN_3927; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3929 = 8'h59 == _T_5[7:0] ? image_2_89 : _GEN_3928; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3930 = 8'h5a == _T_5[7:0] ? image_2_90 : _GEN_3929; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3931 = 8'h5b == _T_5[7:0] ? image_2_91 : _GEN_3930; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3932 = 8'h5c == _T_5[7:0] ? image_2_92 : _GEN_3931; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3933 = 8'h5d == _T_5[7:0] ? image_2_93 : _GEN_3932; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3934 = 8'h5e == _T_5[7:0] ? image_2_94 : _GEN_3933; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3935 = 8'h5f == _T_5[7:0] ? image_2_95 : _GEN_3934; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3936 = 8'h60 == _T_5[7:0] ? image_2_96 : _GEN_3935; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3937 = 8'h61 == _T_5[7:0] ? image_2_97 : _GEN_3936; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3938 = 8'h62 == _T_5[7:0] ? image_2_98 : _GEN_3937; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3939 = 8'h63 == _T_5[7:0] ? image_2_99 : _GEN_3938; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3940 = 8'h64 == _T_5[7:0] ? image_2_100 : _GEN_3939; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3941 = 8'h65 == _T_5[7:0] ? image_2_101 : _GEN_3940; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3942 = 8'h66 == _T_5[7:0] ? image_2_102 : _GEN_3941; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3943 = 8'h67 == _T_5[7:0] ? image_2_103 : _GEN_3942; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3944 = 8'h68 == _T_5[7:0] ? image_2_104 : _GEN_3943; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3945 = 8'h69 == _T_5[7:0] ? image_2_105 : _GEN_3944; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3946 = 8'h6a == _T_5[7:0] ? image_2_106 : _GEN_3945; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3947 = 8'h6b == _T_5[7:0] ? image_2_107 : _GEN_3946; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3948 = 8'h6c == _T_5[7:0] ? image_2_108 : _GEN_3947; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3949 = 8'h6d == _T_5[7:0] ? image_2_109 : _GEN_3948; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3950 = 8'h6e == _T_5[7:0] ? image_2_110 : _GEN_3949; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3951 = 8'h6f == _T_5[7:0] ? image_2_111 : _GEN_3950; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3952 = 8'h70 == _T_5[7:0] ? image_2_112 : _GEN_3951; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3953 = 8'h71 == _T_5[7:0] ? image_2_113 : _GEN_3952; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3954 = 8'h72 == _T_5[7:0] ? image_2_114 : _GEN_3953; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3955 = 8'h73 == _T_5[7:0] ? image_2_115 : _GEN_3954; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3956 = 8'h74 == _T_5[7:0] ? image_2_116 : _GEN_3955; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3957 = 8'h75 == _T_5[7:0] ? image_2_117 : _GEN_3956; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3958 = 8'h76 == _T_5[7:0] ? image_2_118 : _GEN_3957; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3959 = 8'h77 == _T_5[7:0] ? image_2_119 : _GEN_3958; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3960 = 8'h78 == _T_5[7:0] ? image_2_120 : _GEN_3959; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3961 = 8'h79 == _T_5[7:0] ? image_2_121 : _GEN_3960; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3962 = 8'h7a == _T_5[7:0] ? image_2_122 : _GEN_3961; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3963 = 8'h7b == _T_5[7:0] ? image_2_123 : _GEN_3962; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3964 = 8'h7c == _T_5[7:0] ? image_2_124 : _GEN_3963; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3965 = 8'h7d == _T_5[7:0] ? image_2_125 : _GEN_3964; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3966 = 8'h7e == _T_5[7:0] ? image_2_126 : _GEN_3965; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3967 = 8'h7f == _T_5[7:0] ? image_2_127 : _GEN_3966; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3968 = 8'h80 == _T_5[7:0] ? image_2_128 : _GEN_3967; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3969 = 8'h81 == _T_5[7:0] ? image_2_129 : _GEN_3968; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3970 = 8'h82 == _T_5[7:0] ? image_2_130 : _GEN_3969; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3971 = 8'h83 == _T_5[7:0] ? image_2_131 : _GEN_3970; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3972 = 8'h84 == _T_5[7:0] ? image_2_132 : _GEN_3971; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3973 = 8'h85 == _T_5[7:0] ? image_2_133 : _GEN_3972; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3974 = 8'h86 == _T_5[7:0] ? image_2_134 : _GEN_3973; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3975 = 8'h87 == _T_5[7:0] ? image_2_135 : _GEN_3974; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3976 = 8'h88 == _T_5[7:0] ? image_2_136 : _GEN_3975; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3977 = 8'h89 == _T_5[7:0] ? image_2_137 : _GEN_3976; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3978 = 8'h8a == _T_5[7:0] ? image_2_138 : _GEN_3977; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3979 = 8'h8b == _T_5[7:0] ? image_2_139 : _GEN_3978; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3980 = 8'h8c == _T_5[7:0] ? image_2_140 : _GEN_3979; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3981 = 8'h8d == _T_5[7:0] ? image_2_141 : _GEN_3980; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3982 = 8'h8e == _T_5[7:0] ? image_2_142 : _GEN_3981; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3983 = 8'h8f == _T_5[7:0] ? image_2_143 : _GEN_3982; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3984 = 8'h90 == _T_5[7:0] ? image_2_144 : _GEN_3983; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3985 = 8'h91 == _T_5[7:0] ? image_2_145 : _GEN_3984; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3986 = 8'h92 == _T_5[7:0] ? image_2_146 : _GEN_3985; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3987 = 8'h93 == _T_5[7:0] ? image_2_147 : _GEN_3986; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3988 = 8'h94 == _T_5[7:0] ? image_2_148 : _GEN_3987; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3989 = 8'h95 == _T_5[7:0] ? image_2_149 : _GEN_3988; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3990 = 8'h96 == _T_5[7:0] ? image_2_150 : _GEN_3989; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3991 = 8'h97 == _T_5[7:0] ? image_2_151 : _GEN_3990; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3992 = 8'h98 == _T_5[7:0] ? image_2_152 : _GEN_3991; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3993 = 8'h99 == _T_5[7:0] ? image_2_153 : _GEN_3992; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3994 = 8'h9a == _T_5[7:0] ? image_2_154 : _GEN_3993; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3995 = 8'h9b == _T_5[7:0] ? image_2_155 : _GEN_3994; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3996 = 8'h9c == _T_5[7:0] ? image_2_156 : _GEN_3995; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3997 = 8'h9d == _T_5[7:0] ? image_2_157 : _GEN_3996; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3998 = 8'h9e == _T_5[7:0] ? image_2_158 : _GEN_3997; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3999 = 8'h9f == _T_5[7:0] ? image_2_159 : _GEN_3998; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4000 = 8'ha0 == _T_5[7:0] ? image_2_160 : _GEN_3999; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4001 = 8'ha1 == _T_5[7:0] ? image_2_161 : _GEN_4000; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4002 = 8'ha2 == _T_5[7:0] ? image_2_162 : _GEN_4001; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4003 = 8'ha3 == _T_5[7:0] ? image_2_163 : _GEN_4002; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4004 = 8'ha4 == _T_5[7:0] ? image_2_164 : _GEN_4003; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4005 = 8'ha5 == _T_5[7:0] ? image_2_165 : _GEN_4004; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4006 = 8'ha6 == _T_5[7:0] ? image_2_166 : _GEN_4005; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4007 = 8'ha7 == _T_5[7:0] ? image_2_167 : _GEN_4006; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4008 = 8'ha8 == _T_5[7:0] ? image_2_168 : _GEN_4007; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4009 = 8'ha9 == _T_5[7:0] ? image_2_169 : _GEN_4008; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4010 = 8'haa == _T_5[7:0] ? image_2_170 : _GEN_4009; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4011 = 8'hab == _T_5[7:0] ? image_2_171 : _GEN_4010; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4012 = 8'hac == _T_5[7:0] ? image_2_172 : _GEN_4011; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4013 = 8'had == _T_5[7:0] ? image_2_173 : _GEN_4012; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4014 = 8'hae == _T_5[7:0] ? image_2_174 : _GEN_4013; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4015 = 8'haf == _T_5[7:0] ? image_2_175 : _GEN_4014; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4016 = 8'hb0 == _T_5[7:0] ? image_2_176 : _GEN_4015; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4017 = 8'hb1 == _T_5[7:0] ? image_2_177 : _GEN_4016; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4018 = 8'hb2 == _T_5[7:0] ? image_2_178 : _GEN_4017; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4019 = 8'hb3 == _T_5[7:0] ? image_2_179 : _GEN_4018; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4020 = 8'hb4 == _T_5[7:0] ? image_2_180 : _GEN_4019; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4021 = 8'hb5 == _T_5[7:0] ? image_2_181 : _GEN_4020; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4022 = 8'hb6 == _T_5[7:0] ? image_2_182 : _GEN_4021; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4023 = 8'hb7 == _T_5[7:0] ? image_2_183 : _GEN_4022; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4024 = 8'hb8 == _T_5[7:0] ? image_2_184 : _GEN_4023; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4025 = 8'hb9 == _T_5[7:0] ? image_2_185 : _GEN_4024; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4026 = 8'hba == _T_5[7:0] ? image_2_186 : _GEN_4025; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4027 = 8'hbb == _T_5[7:0] ? image_2_187 : _GEN_4026; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4028 = 8'hbc == _T_5[7:0] ? image_2_188 : _GEN_4027; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4029 = 8'hbd == _T_5[7:0] ? image_2_189 : _GEN_4028; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4030 = 8'hbe == _T_5[7:0] ? image_2_190 : _GEN_4029; // @[VideoBuffer.scala 27:30]
  wire [31:0] _T_88 = pixelIndex + 32'h8; // @[VideoBuffer.scala 35:30]
  wire [8:0] _T_89 = 5'h10 * 5'hc; // @[VideoBuffer.scala 36:38]
  wire [31:0] _GEN_5764 = {{23'd0}, _T_89}; // @[VideoBuffer.scala 36:21]
  wire  _T_90 = pixelIndex == _GEN_5764; // @[VideoBuffer.scala 36:21]
  assign io_pixelVal_out_0 = 8'hbf == _T_5[7:0] ? image_0_191 : _GEN_190; // @[VideoBuffer.scala 27:30]
  assign io_pixelVal_out_1 = 8'hbf == _T_5[7:0] ? image_1_191 : _GEN_2110; // @[VideoBuffer.scala 27:30]
  assign io_pixelVal_out_2 = 8'hbf == _T_5[7:0] ? image_2_191 : _GEN_4030; // @[VideoBuffer.scala 27:30]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  image_0_0 = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  image_0_1 = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  image_0_2 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  image_0_3 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  image_0_4 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  image_0_5 = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  image_0_6 = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  image_0_7 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  image_0_8 = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  image_0_9 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  image_0_10 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  image_0_11 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  image_0_12 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  image_0_13 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  image_0_14 = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  image_0_15 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  image_0_16 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  image_0_17 = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  image_0_18 = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  image_0_19 = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  image_0_20 = _RAND_20[3:0];
  _RAND_21 = {1{`RANDOM}};
  image_0_21 = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  image_0_22 = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  image_0_23 = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  image_0_24 = _RAND_24[3:0];
  _RAND_25 = {1{`RANDOM}};
  image_0_25 = _RAND_25[3:0];
  _RAND_26 = {1{`RANDOM}};
  image_0_26 = _RAND_26[3:0];
  _RAND_27 = {1{`RANDOM}};
  image_0_27 = _RAND_27[3:0];
  _RAND_28 = {1{`RANDOM}};
  image_0_28 = _RAND_28[3:0];
  _RAND_29 = {1{`RANDOM}};
  image_0_29 = _RAND_29[3:0];
  _RAND_30 = {1{`RANDOM}};
  image_0_30 = _RAND_30[3:0];
  _RAND_31 = {1{`RANDOM}};
  image_0_31 = _RAND_31[3:0];
  _RAND_32 = {1{`RANDOM}};
  image_0_32 = _RAND_32[3:0];
  _RAND_33 = {1{`RANDOM}};
  image_0_33 = _RAND_33[3:0];
  _RAND_34 = {1{`RANDOM}};
  image_0_34 = _RAND_34[3:0];
  _RAND_35 = {1{`RANDOM}};
  image_0_35 = _RAND_35[3:0];
  _RAND_36 = {1{`RANDOM}};
  image_0_36 = _RAND_36[3:0];
  _RAND_37 = {1{`RANDOM}};
  image_0_37 = _RAND_37[3:0];
  _RAND_38 = {1{`RANDOM}};
  image_0_38 = _RAND_38[3:0];
  _RAND_39 = {1{`RANDOM}};
  image_0_39 = _RAND_39[3:0];
  _RAND_40 = {1{`RANDOM}};
  image_0_40 = _RAND_40[3:0];
  _RAND_41 = {1{`RANDOM}};
  image_0_41 = _RAND_41[3:0];
  _RAND_42 = {1{`RANDOM}};
  image_0_42 = _RAND_42[3:0];
  _RAND_43 = {1{`RANDOM}};
  image_0_43 = _RAND_43[3:0];
  _RAND_44 = {1{`RANDOM}};
  image_0_44 = _RAND_44[3:0];
  _RAND_45 = {1{`RANDOM}};
  image_0_45 = _RAND_45[3:0];
  _RAND_46 = {1{`RANDOM}};
  image_0_46 = _RAND_46[3:0];
  _RAND_47 = {1{`RANDOM}};
  image_0_47 = _RAND_47[3:0];
  _RAND_48 = {1{`RANDOM}};
  image_0_48 = _RAND_48[3:0];
  _RAND_49 = {1{`RANDOM}};
  image_0_49 = _RAND_49[3:0];
  _RAND_50 = {1{`RANDOM}};
  image_0_50 = _RAND_50[3:0];
  _RAND_51 = {1{`RANDOM}};
  image_0_51 = _RAND_51[3:0];
  _RAND_52 = {1{`RANDOM}};
  image_0_52 = _RAND_52[3:0];
  _RAND_53 = {1{`RANDOM}};
  image_0_53 = _RAND_53[3:0];
  _RAND_54 = {1{`RANDOM}};
  image_0_54 = _RAND_54[3:0];
  _RAND_55 = {1{`RANDOM}};
  image_0_55 = _RAND_55[3:0];
  _RAND_56 = {1{`RANDOM}};
  image_0_56 = _RAND_56[3:0];
  _RAND_57 = {1{`RANDOM}};
  image_0_57 = _RAND_57[3:0];
  _RAND_58 = {1{`RANDOM}};
  image_0_58 = _RAND_58[3:0];
  _RAND_59 = {1{`RANDOM}};
  image_0_59 = _RAND_59[3:0];
  _RAND_60 = {1{`RANDOM}};
  image_0_60 = _RAND_60[3:0];
  _RAND_61 = {1{`RANDOM}};
  image_0_61 = _RAND_61[3:0];
  _RAND_62 = {1{`RANDOM}};
  image_0_62 = _RAND_62[3:0];
  _RAND_63 = {1{`RANDOM}};
  image_0_63 = _RAND_63[3:0];
  _RAND_64 = {1{`RANDOM}};
  image_0_64 = _RAND_64[3:0];
  _RAND_65 = {1{`RANDOM}};
  image_0_65 = _RAND_65[3:0];
  _RAND_66 = {1{`RANDOM}};
  image_0_66 = _RAND_66[3:0];
  _RAND_67 = {1{`RANDOM}};
  image_0_67 = _RAND_67[3:0];
  _RAND_68 = {1{`RANDOM}};
  image_0_68 = _RAND_68[3:0];
  _RAND_69 = {1{`RANDOM}};
  image_0_69 = _RAND_69[3:0];
  _RAND_70 = {1{`RANDOM}};
  image_0_70 = _RAND_70[3:0];
  _RAND_71 = {1{`RANDOM}};
  image_0_71 = _RAND_71[3:0];
  _RAND_72 = {1{`RANDOM}};
  image_0_72 = _RAND_72[3:0];
  _RAND_73 = {1{`RANDOM}};
  image_0_73 = _RAND_73[3:0];
  _RAND_74 = {1{`RANDOM}};
  image_0_74 = _RAND_74[3:0];
  _RAND_75 = {1{`RANDOM}};
  image_0_75 = _RAND_75[3:0];
  _RAND_76 = {1{`RANDOM}};
  image_0_76 = _RAND_76[3:0];
  _RAND_77 = {1{`RANDOM}};
  image_0_77 = _RAND_77[3:0];
  _RAND_78 = {1{`RANDOM}};
  image_0_78 = _RAND_78[3:0];
  _RAND_79 = {1{`RANDOM}};
  image_0_79 = _RAND_79[3:0];
  _RAND_80 = {1{`RANDOM}};
  image_0_80 = _RAND_80[3:0];
  _RAND_81 = {1{`RANDOM}};
  image_0_81 = _RAND_81[3:0];
  _RAND_82 = {1{`RANDOM}};
  image_0_82 = _RAND_82[3:0];
  _RAND_83 = {1{`RANDOM}};
  image_0_83 = _RAND_83[3:0];
  _RAND_84 = {1{`RANDOM}};
  image_0_84 = _RAND_84[3:0];
  _RAND_85 = {1{`RANDOM}};
  image_0_85 = _RAND_85[3:0];
  _RAND_86 = {1{`RANDOM}};
  image_0_86 = _RAND_86[3:0];
  _RAND_87 = {1{`RANDOM}};
  image_0_87 = _RAND_87[3:0];
  _RAND_88 = {1{`RANDOM}};
  image_0_88 = _RAND_88[3:0];
  _RAND_89 = {1{`RANDOM}};
  image_0_89 = _RAND_89[3:0];
  _RAND_90 = {1{`RANDOM}};
  image_0_90 = _RAND_90[3:0];
  _RAND_91 = {1{`RANDOM}};
  image_0_91 = _RAND_91[3:0];
  _RAND_92 = {1{`RANDOM}};
  image_0_92 = _RAND_92[3:0];
  _RAND_93 = {1{`RANDOM}};
  image_0_93 = _RAND_93[3:0];
  _RAND_94 = {1{`RANDOM}};
  image_0_94 = _RAND_94[3:0];
  _RAND_95 = {1{`RANDOM}};
  image_0_95 = _RAND_95[3:0];
  _RAND_96 = {1{`RANDOM}};
  image_0_96 = _RAND_96[3:0];
  _RAND_97 = {1{`RANDOM}};
  image_0_97 = _RAND_97[3:0];
  _RAND_98 = {1{`RANDOM}};
  image_0_98 = _RAND_98[3:0];
  _RAND_99 = {1{`RANDOM}};
  image_0_99 = _RAND_99[3:0];
  _RAND_100 = {1{`RANDOM}};
  image_0_100 = _RAND_100[3:0];
  _RAND_101 = {1{`RANDOM}};
  image_0_101 = _RAND_101[3:0];
  _RAND_102 = {1{`RANDOM}};
  image_0_102 = _RAND_102[3:0];
  _RAND_103 = {1{`RANDOM}};
  image_0_103 = _RAND_103[3:0];
  _RAND_104 = {1{`RANDOM}};
  image_0_104 = _RAND_104[3:0];
  _RAND_105 = {1{`RANDOM}};
  image_0_105 = _RAND_105[3:0];
  _RAND_106 = {1{`RANDOM}};
  image_0_106 = _RAND_106[3:0];
  _RAND_107 = {1{`RANDOM}};
  image_0_107 = _RAND_107[3:0];
  _RAND_108 = {1{`RANDOM}};
  image_0_108 = _RAND_108[3:0];
  _RAND_109 = {1{`RANDOM}};
  image_0_109 = _RAND_109[3:0];
  _RAND_110 = {1{`RANDOM}};
  image_0_110 = _RAND_110[3:0];
  _RAND_111 = {1{`RANDOM}};
  image_0_111 = _RAND_111[3:0];
  _RAND_112 = {1{`RANDOM}};
  image_0_112 = _RAND_112[3:0];
  _RAND_113 = {1{`RANDOM}};
  image_0_113 = _RAND_113[3:0];
  _RAND_114 = {1{`RANDOM}};
  image_0_114 = _RAND_114[3:0];
  _RAND_115 = {1{`RANDOM}};
  image_0_115 = _RAND_115[3:0];
  _RAND_116 = {1{`RANDOM}};
  image_0_116 = _RAND_116[3:0];
  _RAND_117 = {1{`RANDOM}};
  image_0_117 = _RAND_117[3:0];
  _RAND_118 = {1{`RANDOM}};
  image_0_118 = _RAND_118[3:0];
  _RAND_119 = {1{`RANDOM}};
  image_0_119 = _RAND_119[3:0];
  _RAND_120 = {1{`RANDOM}};
  image_0_120 = _RAND_120[3:0];
  _RAND_121 = {1{`RANDOM}};
  image_0_121 = _RAND_121[3:0];
  _RAND_122 = {1{`RANDOM}};
  image_0_122 = _RAND_122[3:0];
  _RAND_123 = {1{`RANDOM}};
  image_0_123 = _RAND_123[3:0];
  _RAND_124 = {1{`RANDOM}};
  image_0_124 = _RAND_124[3:0];
  _RAND_125 = {1{`RANDOM}};
  image_0_125 = _RAND_125[3:0];
  _RAND_126 = {1{`RANDOM}};
  image_0_126 = _RAND_126[3:0];
  _RAND_127 = {1{`RANDOM}};
  image_0_127 = _RAND_127[3:0];
  _RAND_128 = {1{`RANDOM}};
  image_0_128 = _RAND_128[3:0];
  _RAND_129 = {1{`RANDOM}};
  image_0_129 = _RAND_129[3:0];
  _RAND_130 = {1{`RANDOM}};
  image_0_130 = _RAND_130[3:0];
  _RAND_131 = {1{`RANDOM}};
  image_0_131 = _RAND_131[3:0];
  _RAND_132 = {1{`RANDOM}};
  image_0_132 = _RAND_132[3:0];
  _RAND_133 = {1{`RANDOM}};
  image_0_133 = _RAND_133[3:0];
  _RAND_134 = {1{`RANDOM}};
  image_0_134 = _RAND_134[3:0];
  _RAND_135 = {1{`RANDOM}};
  image_0_135 = _RAND_135[3:0];
  _RAND_136 = {1{`RANDOM}};
  image_0_136 = _RAND_136[3:0];
  _RAND_137 = {1{`RANDOM}};
  image_0_137 = _RAND_137[3:0];
  _RAND_138 = {1{`RANDOM}};
  image_0_138 = _RAND_138[3:0];
  _RAND_139 = {1{`RANDOM}};
  image_0_139 = _RAND_139[3:0];
  _RAND_140 = {1{`RANDOM}};
  image_0_140 = _RAND_140[3:0];
  _RAND_141 = {1{`RANDOM}};
  image_0_141 = _RAND_141[3:0];
  _RAND_142 = {1{`RANDOM}};
  image_0_142 = _RAND_142[3:0];
  _RAND_143 = {1{`RANDOM}};
  image_0_143 = _RAND_143[3:0];
  _RAND_144 = {1{`RANDOM}};
  image_0_144 = _RAND_144[3:0];
  _RAND_145 = {1{`RANDOM}};
  image_0_145 = _RAND_145[3:0];
  _RAND_146 = {1{`RANDOM}};
  image_0_146 = _RAND_146[3:0];
  _RAND_147 = {1{`RANDOM}};
  image_0_147 = _RAND_147[3:0];
  _RAND_148 = {1{`RANDOM}};
  image_0_148 = _RAND_148[3:0];
  _RAND_149 = {1{`RANDOM}};
  image_0_149 = _RAND_149[3:0];
  _RAND_150 = {1{`RANDOM}};
  image_0_150 = _RAND_150[3:0];
  _RAND_151 = {1{`RANDOM}};
  image_0_151 = _RAND_151[3:0];
  _RAND_152 = {1{`RANDOM}};
  image_0_152 = _RAND_152[3:0];
  _RAND_153 = {1{`RANDOM}};
  image_0_153 = _RAND_153[3:0];
  _RAND_154 = {1{`RANDOM}};
  image_0_154 = _RAND_154[3:0];
  _RAND_155 = {1{`RANDOM}};
  image_0_155 = _RAND_155[3:0];
  _RAND_156 = {1{`RANDOM}};
  image_0_156 = _RAND_156[3:0];
  _RAND_157 = {1{`RANDOM}};
  image_0_157 = _RAND_157[3:0];
  _RAND_158 = {1{`RANDOM}};
  image_0_158 = _RAND_158[3:0];
  _RAND_159 = {1{`RANDOM}};
  image_0_159 = _RAND_159[3:0];
  _RAND_160 = {1{`RANDOM}};
  image_0_160 = _RAND_160[3:0];
  _RAND_161 = {1{`RANDOM}};
  image_0_161 = _RAND_161[3:0];
  _RAND_162 = {1{`RANDOM}};
  image_0_162 = _RAND_162[3:0];
  _RAND_163 = {1{`RANDOM}};
  image_0_163 = _RAND_163[3:0];
  _RAND_164 = {1{`RANDOM}};
  image_0_164 = _RAND_164[3:0];
  _RAND_165 = {1{`RANDOM}};
  image_0_165 = _RAND_165[3:0];
  _RAND_166 = {1{`RANDOM}};
  image_0_166 = _RAND_166[3:0];
  _RAND_167 = {1{`RANDOM}};
  image_0_167 = _RAND_167[3:0];
  _RAND_168 = {1{`RANDOM}};
  image_0_168 = _RAND_168[3:0];
  _RAND_169 = {1{`RANDOM}};
  image_0_169 = _RAND_169[3:0];
  _RAND_170 = {1{`RANDOM}};
  image_0_170 = _RAND_170[3:0];
  _RAND_171 = {1{`RANDOM}};
  image_0_171 = _RAND_171[3:0];
  _RAND_172 = {1{`RANDOM}};
  image_0_172 = _RAND_172[3:0];
  _RAND_173 = {1{`RANDOM}};
  image_0_173 = _RAND_173[3:0];
  _RAND_174 = {1{`RANDOM}};
  image_0_174 = _RAND_174[3:0];
  _RAND_175 = {1{`RANDOM}};
  image_0_175 = _RAND_175[3:0];
  _RAND_176 = {1{`RANDOM}};
  image_0_176 = _RAND_176[3:0];
  _RAND_177 = {1{`RANDOM}};
  image_0_177 = _RAND_177[3:0];
  _RAND_178 = {1{`RANDOM}};
  image_0_178 = _RAND_178[3:0];
  _RAND_179 = {1{`RANDOM}};
  image_0_179 = _RAND_179[3:0];
  _RAND_180 = {1{`RANDOM}};
  image_0_180 = _RAND_180[3:0];
  _RAND_181 = {1{`RANDOM}};
  image_0_181 = _RAND_181[3:0];
  _RAND_182 = {1{`RANDOM}};
  image_0_182 = _RAND_182[3:0];
  _RAND_183 = {1{`RANDOM}};
  image_0_183 = _RAND_183[3:0];
  _RAND_184 = {1{`RANDOM}};
  image_0_184 = _RAND_184[3:0];
  _RAND_185 = {1{`RANDOM}};
  image_0_185 = _RAND_185[3:0];
  _RAND_186 = {1{`RANDOM}};
  image_0_186 = _RAND_186[3:0];
  _RAND_187 = {1{`RANDOM}};
  image_0_187 = _RAND_187[3:0];
  _RAND_188 = {1{`RANDOM}};
  image_0_188 = _RAND_188[3:0];
  _RAND_189 = {1{`RANDOM}};
  image_0_189 = _RAND_189[3:0];
  _RAND_190 = {1{`RANDOM}};
  image_0_190 = _RAND_190[3:0];
  _RAND_191 = {1{`RANDOM}};
  image_0_191 = _RAND_191[3:0];
  _RAND_192 = {1{`RANDOM}};
  image_1_0 = _RAND_192[3:0];
  _RAND_193 = {1{`RANDOM}};
  image_1_1 = _RAND_193[3:0];
  _RAND_194 = {1{`RANDOM}};
  image_1_2 = _RAND_194[3:0];
  _RAND_195 = {1{`RANDOM}};
  image_1_3 = _RAND_195[3:0];
  _RAND_196 = {1{`RANDOM}};
  image_1_4 = _RAND_196[3:0];
  _RAND_197 = {1{`RANDOM}};
  image_1_5 = _RAND_197[3:0];
  _RAND_198 = {1{`RANDOM}};
  image_1_6 = _RAND_198[3:0];
  _RAND_199 = {1{`RANDOM}};
  image_1_7 = _RAND_199[3:0];
  _RAND_200 = {1{`RANDOM}};
  image_1_8 = _RAND_200[3:0];
  _RAND_201 = {1{`RANDOM}};
  image_1_9 = _RAND_201[3:0];
  _RAND_202 = {1{`RANDOM}};
  image_1_10 = _RAND_202[3:0];
  _RAND_203 = {1{`RANDOM}};
  image_1_11 = _RAND_203[3:0];
  _RAND_204 = {1{`RANDOM}};
  image_1_12 = _RAND_204[3:0];
  _RAND_205 = {1{`RANDOM}};
  image_1_13 = _RAND_205[3:0];
  _RAND_206 = {1{`RANDOM}};
  image_1_14 = _RAND_206[3:0];
  _RAND_207 = {1{`RANDOM}};
  image_1_15 = _RAND_207[3:0];
  _RAND_208 = {1{`RANDOM}};
  image_1_16 = _RAND_208[3:0];
  _RAND_209 = {1{`RANDOM}};
  image_1_17 = _RAND_209[3:0];
  _RAND_210 = {1{`RANDOM}};
  image_1_18 = _RAND_210[3:0];
  _RAND_211 = {1{`RANDOM}};
  image_1_19 = _RAND_211[3:0];
  _RAND_212 = {1{`RANDOM}};
  image_1_20 = _RAND_212[3:0];
  _RAND_213 = {1{`RANDOM}};
  image_1_21 = _RAND_213[3:0];
  _RAND_214 = {1{`RANDOM}};
  image_1_22 = _RAND_214[3:0];
  _RAND_215 = {1{`RANDOM}};
  image_1_23 = _RAND_215[3:0];
  _RAND_216 = {1{`RANDOM}};
  image_1_24 = _RAND_216[3:0];
  _RAND_217 = {1{`RANDOM}};
  image_1_25 = _RAND_217[3:0];
  _RAND_218 = {1{`RANDOM}};
  image_1_26 = _RAND_218[3:0];
  _RAND_219 = {1{`RANDOM}};
  image_1_27 = _RAND_219[3:0];
  _RAND_220 = {1{`RANDOM}};
  image_1_28 = _RAND_220[3:0];
  _RAND_221 = {1{`RANDOM}};
  image_1_29 = _RAND_221[3:0];
  _RAND_222 = {1{`RANDOM}};
  image_1_30 = _RAND_222[3:0];
  _RAND_223 = {1{`RANDOM}};
  image_1_31 = _RAND_223[3:0];
  _RAND_224 = {1{`RANDOM}};
  image_1_32 = _RAND_224[3:0];
  _RAND_225 = {1{`RANDOM}};
  image_1_33 = _RAND_225[3:0];
  _RAND_226 = {1{`RANDOM}};
  image_1_34 = _RAND_226[3:0];
  _RAND_227 = {1{`RANDOM}};
  image_1_35 = _RAND_227[3:0];
  _RAND_228 = {1{`RANDOM}};
  image_1_36 = _RAND_228[3:0];
  _RAND_229 = {1{`RANDOM}};
  image_1_37 = _RAND_229[3:0];
  _RAND_230 = {1{`RANDOM}};
  image_1_38 = _RAND_230[3:0];
  _RAND_231 = {1{`RANDOM}};
  image_1_39 = _RAND_231[3:0];
  _RAND_232 = {1{`RANDOM}};
  image_1_40 = _RAND_232[3:0];
  _RAND_233 = {1{`RANDOM}};
  image_1_41 = _RAND_233[3:0];
  _RAND_234 = {1{`RANDOM}};
  image_1_42 = _RAND_234[3:0];
  _RAND_235 = {1{`RANDOM}};
  image_1_43 = _RAND_235[3:0];
  _RAND_236 = {1{`RANDOM}};
  image_1_44 = _RAND_236[3:0];
  _RAND_237 = {1{`RANDOM}};
  image_1_45 = _RAND_237[3:0];
  _RAND_238 = {1{`RANDOM}};
  image_1_46 = _RAND_238[3:0];
  _RAND_239 = {1{`RANDOM}};
  image_1_47 = _RAND_239[3:0];
  _RAND_240 = {1{`RANDOM}};
  image_1_48 = _RAND_240[3:0];
  _RAND_241 = {1{`RANDOM}};
  image_1_49 = _RAND_241[3:0];
  _RAND_242 = {1{`RANDOM}};
  image_1_50 = _RAND_242[3:0];
  _RAND_243 = {1{`RANDOM}};
  image_1_51 = _RAND_243[3:0];
  _RAND_244 = {1{`RANDOM}};
  image_1_52 = _RAND_244[3:0];
  _RAND_245 = {1{`RANDOM}};
  image_1_53 = _RAND_245[3:0];
  _RAND_246 = {1{`RANDOM}};
  image_1_54 = _RAND_246[3:0];
  _RAND_247 = {1{`RANDOM}};
  image_1_55 = _RAND_247[3:0];
  _RAND_248 = {1{`RANDOM}};
  image_1_56 = _RAND_248[3:0];
  _RAND_249 = {1{`RANDOM}};
  image_1_57 = _RAND_249[3:0];
  _RAND_250 = {1{`RANDOM}};
  image_1_58 = _RAND_250[3:0];
  _RAND_251 = {1{`RANDOM}};
  image_1_59 = _RAND_251[3:0];
  _RAND_252 = {1{`RANDOM}};
  image_1_60 = _RAND_252[3:0];
  _RAND_253 = {1{`RANDOM}};
  image_1_61 = _RAND_253[3:0];
  _RAND_254 = {1{`RANDOM}};
  image_1_62 = _RAND_254[3:0];
  _RAND_255 = {1{`RANDOM}};
  image_1_63 = _RAND_255[3:0];
  _RAND_256 = {1{`RANDOM}};
  image_1_64 = _RAND_256[3:0];
  _RAND_257 = {1{`RANDOM}};
  image_1_65 = _RAND_257[3:0];
  _RAND_258 = {1{`RANDOM}};
  image_1_66 = _RAND_258[3:0];
  _RAND_259 = {1{`RANDOM}};
  image_1_67 = _RAND_259[3:0];
  _RAND_260 = {1{`RANDOM}};
  image_1_68 = _RAND_260[3:0];
  _RAND_261 = {1{`RANDOM}};
  image_1_69 = _RAND_261[3:0];
  _RAND_262 = {1{`RANDOM}};
  image_1_70 = _RAND_262[3:0];
  _RAND_263 = {1{`RANDOM}};
  image_1_71 = _RAND_263[3:0];
  _RAND_264 = {1{`RANDOM}};
  image_1_72 = _RAND_264[3:0];
  _RAND_265 = {1{`RANDOM}};
  image_1_73 = _RAND_265[3:0];
  _RAND_266 = {1{`RANDOM}};
  image_1_74 = _RAND_266[3:0];
  _RAND_267 = {1{`RANDOM}};
  image_1_75 = _RAND_267[3:0];
  _RAND_268 = {1{`RANDOM}};
  image_1_76 = _RAND_268[3:0];
  _RAND_269 = {1{`RANDOM}};
  image_1_77 = _RAND_269[3:0];
  _RAND_270 = {1{`RANDOM}};
  image_1_78 = _RAND_270[3:0];
  _RAND_271 = {1{`RANDOM}};
  image_1_79 = _RAND_271[3:0];
  _RAND_272 = {1{`RANDOM}};
  image_1_80 = _RAND_272[3:0];
  _RAND_273 = {1{`RANDOM}};
  image_1_81 = _RAND_273[3:0];
  _RAND_274 = {1{`RANDOM}};
  image_1_82 = _RAND_274[3:0];
  _RAND_275 = {1{`RANDOM}};
  image_1_83 = _RAND_275[3:0];
  _RAND_276 = {1{`RANDOM}};
  image_1_84 = _RAND_276[3:0];
  _RAND_277 = {1{`RANDOM}};
  image_1_85 = _RAND_277[3:0];
  _RAND_278 = {1{`RANDOM}};
  image_1_86 = _RAND_278[3:0];
  _RAND_279 = {1{`RANDOM}};
  image_1_87 = _RAND_279[3:0];
  _RAND_280 = {1{`RANDOM}};
  image_1_88 = _RAND_280[3:0];
  _RAND_281 = {1{`RANDOM}};
  image_1_89 = _RAND_281[3:0];
  _RAND_282 = {1{`RANDOM}};
  image_1_90 = _RAND_282[3:0];
  _RAND_283 = {1{`RANDOM}};
  image_1_91 = _RAND_283[3:0];
  _RAND_284 = {1{`RANDOM}};
  image_1_92 = _RAND_284[3:0];
  _RAND_285 = {1{`RANDOM}};
  image_1_93 = _RAND_285[3:0];
  _RAND_286 = {1{`RANDOM}};
  image_1_94 = _RAND_286[3:0];
  _RAND_287 = {1{`RANDOM}};
  image_1_95 = _RAND_287[3:0];
  _RAND_288 = {1{`RANDOM}};
  image_1_96 = _RAND_288[3:0];
  _RAND_289 = {1{`RANDOM}};
  image_1_97 = _RAND_289[3:0];
  _RAND_290 = {1{`RANDOM}};
  image_1_98 = _RAND_290[3:0];
  _RAND_291 = {1{`RANDOM}};
  image_1_99 = _RAND_291[3:0];
  _RAND_292 = {1{`RANDOM}};
  image_1_100 = _RAND_292[3:0];
  _RAND_293 = {1{`RANDOM}};
  image_1_101 = _RAND_293[3:0];
  _RAND_294 = {1{`RANDOM}};
  image_1_102 = _RAND_294[3:0];
  _RAND_295 = {1{`RANDOM}};
  image_1_103 = _RAND_295[3:0];
  _RAND_296 = {1{`RANDOM}};
  image_1_104 = _RAND_296[3:0];
  _RAND_297 = {1{`RANDOM}};
  image_1_105 = _RAND_297[3:0];
  _RAND_298 = {1{`RANDOM}};
  image_1_106 = _RAND_298[3:0];
  _RAND_299 = {1{`RANDOM}};
  image_1_107 = _RAND_299[3:0];
  _RAND_300 = {1{`RANDOM}};
  image_1_108 = _RAND_300[3:0];
  _RAND_301 = {1{`RANDOM}};
  image_1_109 = _RAND_301[3:0];
  _RAND_302 = {1{`RANDOM}};
  image_1_110 = _RAND_302[3:0];
  _RAND_303 = {1{`RANDOM}};
  image_1_111 = _RAND_303[3:0];
  _RAND_304 = {1{`RANDOM}};
  image_1_112 = _RAND_304[3:0];
  _RAND_305 = {1{`RANDOM}};
  image_1_113 = _RAND_305[3:0];
  _RAND_306 = {1{`RANDOM}};
  image_1_114 = _RAND_306[3:0];
  _RAND_307 = {1{`RANDOM}};
  image_1_115 = _RAND_307[3:0];
  _RAND_308 = {1{`RANDOM}};
  image_1_116 = _RAND_308[3:0];
  _RAND_309 = {1{`RANDOM}};
  image_1_117 = _RAND_309[3:0];
  _RAND_310 = {1{`RANDOM}};
  image_1_118 = _RAND_310[3:0];
  _RAND_311 = {1{`RANDOM}};
  image_1_119 = _RAND_311[3:0];
  _RAND_312 = {1{`RANDOM}};
  image_1_120 = _RAND_312[3:0];
  _RAND_313 = {1{`RANDOM}};
  image_1_121 = _RAND_313[3:0];
  _RAND_314 = {1{`RANDOM}};
  image_1_122 = _RAND_314[3:0];
  _RAND_315 = {1{`RANDOM}};
  image_1_123 = _RAND_315[3:0];
  _RAND_316 = {1{`RANDOM}};
  image_1_124 = _RAND_316[3:0];
  _RAND_317 = {1{`RANDOM}};
  image_1_125 = _RAND_317[3:0];
  _RAND_318 = {1{`RANDOM}};
  image_1_126 = _RAND_318[3:0];
  _RAND_319 = {1{`RANDOM}};
  image_1_127 = _RAND_319[3:0];
  _RAND_320 = {1{`RANDOM}};
  image_1_128 = _RAND_320[3:0];
  _RAND_321 = {1{`RANDOM}};
  image_1_129 = _RAND_321[3:0];
  _RAND_322 = {1{`RANDOM}};
  image_1_130 = _RAND_322[3:0];
  _RAND_323 = {1{`RANDOM}};
  image_1_131 = _RAND_323[3:0];
  _RAND_324 = {1{`RANDOM}};
  image_1_132 = _RAND_324[3:0];
  _RAND_325 = {1{`RANDOM}};
  image_1_133 = _RAND_325[3:0];
  _RAND_326 = {1{`RANDOM}};
  image_1_134 = _RAND_326[3:0];
  _RAND_327 = {1{`RANDOM}};
  image_1_135 = _RAND_327[3:0];
  _RAND_328 = {1{`RANDOM}};
  image_1_136 = _RAND_328[3:0];
  _RAND_329 = {1{`RANDOM}};
  image_1_137 = _RAND_329[3:0];
  _RAND_330 = {1{`RANDOM}};
  image_1_138 = _RAND_330[3:0];
  _RAND_331 = {1{`RANDOM}};
  image_1_139 = _RAND_331[3:0];
  _RAND_332 = {1{`RANDOM}};
  image_1_140 = _RAND_332[3:0];
  _RAND_333 = {1{`RANDOM}};
  image_1_141 = _RAND_333[3:0];
  _RAND_334 = {1{`RANDOM}};
  image_1_142 = _RAND_334[3:0];
  _RAND_335 = {1{`RANDOM}};
  image_1_143 = _RAND_335[3:0];
  _RAND_336 = {1{`RANDOM}};
  image_1_144 = _RAND_336[3:0];
  _RAND_337 = {1{`RANDOM}};
  image_1_145 = _RAND_337[3:0];
  _RAND_338 = {1{`RANDOM}};
  image_1_146 = _RAND_338[3:0];
  _RAND_339 = {1{`RANDOM}};
  image_1_147 = _RAND_339[3:0];
  _RAND_340 = {1{`RANDOM}};
  image_1_148 = _RAND_340[3:0];
  _RAND_341 = {1{`RANDOM}};
  image_1_149 = _RAND_341[3:0];
  _RAND_342 = {1{`RANDOM}};
  image_1_150 = _RAND_342[3:0];
  _RAND_343 = {1{`RANDOM}};
  image_1_151 = _RAND_343[3:0];
  _RAND_344 = {1{`RANDOM}};
  image_1_152 = _RAND_344[3:0];
  _RAND_345 = {1{`RANDOM}};
  image_1_153 = _RAND_345[3:0];
  _RAND_346 = {1{`RANDOM}};
  image_1_154 = _RAND_346[3:0];
  _RAND_347 = {1{`RANDOM}};
  image_1_155 = _RAND_347[3:0];
  _RAND_348 = {1{`RANDOM}};
  image_1_156 = _RAND_348[3:0];
  _RAND_349 = {1{`RANDOM}};
  image_1_157 = _RAND_349[3:0];
  _RAND_350 = {1{`RANDOM}};
  image_1_158 = _RAND_350[3:0];
  _RAND_351 = {1{`RANDOM}};
  image_1_159 = _RAND_351[3:0];
  _RAND_352 = {1{`RANDOM}};
  image_1_160 = _RAND_352[3:0];
  _RAND_353 = {1{`RANDOM}};
  image_1_161 = _RAND_353[3:0];
  _RAND_354 = {1{`RANDOM}};
  image_1_162 = _RAND_354[3:0];
  _RAND_355 = {1{`RANDOM}};
  image_1_163 = _RAND_355[3:0];
  _RAND_356 = {1{`RANDOM}};
  image_1_164 = _RAND_356[3:0];
  _RAND_357 = {1{`RANDOM}};
  image_1_165 = _RAND_357[3:0];
  _RAND_358 = {1{`RANDOM}};
  image_1_166 = _RAND_358[3:0];
  _RAND_359 = {1{`RANDOM}};
  image_1_167 = _RAND_359[3:0];
  _RAND_360 = {1{`RANDOM}};
  image_1_168 = _RAND_360[3:0];
  _RAND_361 = {1{`RANDOM}};
  image_1_169 = _RAND_361[3:0];
  _RAND_362 = {1{`RANDOM}};
  image_1_170 = _RAND_362[3:0];
  _RAND_363 = {1{`RANDOM}};
  image_1_171 = _RAND_363[3:0];
  _RAND_364 = {1{`RANDOM}};
  image_1_172 = _RAND_364[3:0];
  _RAND_365 = {1{`RANDOM}};
  image_1_173 = _RAND_365[3:0];
  _RAND_366 = {1{`RANDOM}};
  image_1_174 = _RAND_366[3:0];
  _RAND_367 = {1{`RANDOM}};
  image_1_175 = _RAND_367[3:0];
  _RAND_368 = {1{`RANDOM}};
  image_1_176 = _RAND_368[3:0];
  _RAND_369 = {1{`RANDOM}};
  image_1_177 = _RAND_369[3:0];
  _RAND_370 = {1{`RANDOM}};
  image_1_178 = _RAND_370[3:0];
  _RAND_371 = {1{`RANDOM}};
  image_1_179 = _RAND_371[3:0];
  _RAND_372 = {1{`RANDOM}};
  image_1_180 = _RAND_372[3:0];
  _RAND_373 = {1{`RANDOM}};
  image_1_181 = _RAND_373[3:0];
  _RAND_374 = {1{`RANDOM}};
  image_1_182 = _RAND_374[3:0];
  _RAND_375 = {1{`RANDOM}};
  image_1_183 = _RAND_375[3:0];
  _RAND_376 = {1{`RANDOM}};
  image_1_184 = _RAND_376[3:0];
  _RAND_377 = {1{`RANDOM}};
  image_1_185 = _RAND_377[3:0];
  _RAND_378 = {1{`RANDOM}};
  image_1_186 = _RAND_378[3:0];
  _RAND_379 = {1{`RANDOM}};
  image_1_187 = _RAND_379[3:0];
  _RAND_380 = {1{`RANDOM}};
  image_1_188 = _RAND_380[3:0];
  _RAND_381 = {1{`RANDOM}};
  image_1_189 = _RAND_381[3:0];
  _RAND_382 = {1{`RANDOM}};
  image_1_190 = _RAND_382[3:0];
  _RAND_383 = {1{`RANDOM}};
  image_1_191 = _RAND_383[3:0];
  _RAND_384 = {1{`RANDOM}};
  image_2_0 = _RAND_384[3:0];
  _RAND_385 = {1{`RANDOM}};
  image_2_1 = _RAND_385[3:0];
  _RAND_386 = {1{`RANDOM}};
  image_2_2 = _RAND_386[3:0];
  _RAND_387 = {1{`RANDOM}};
  image_2_3 = _RAND_387[3:0];
  _RAND_388 = {1{`RANDOM}};
  image_2_4 = _RAND_388[3:0];
  _RAND_389 = {1{`RANDOM}};
  image_2_5 = _RAND_389[3:0];
  _RAND_390 = {1{`RANDOM}};
  image_2_6 = _RAND_390[3:0];
  _RAND_391 = {1{`RANDOM}};
  image_2_7 = _RAND_391[3:0];
  _RAND_392 = {1{`RANDOM}};
  image_2_8 = _RAND_392[3:0];
  _RAND_393 = {1{`RANDOM}};
  image_2_9 = _RAND_393[3:0];
  _RAND_394 = {1{`RANDOM}};
  image_2_10 = _RAND_394[3:0];
  _RAND_395 = {1{`RANDOM}};
  image_2_11 = _RAND_395[3:0];
  _RAND_396 = {1{`RANDOM}};
  image_2_12 = _RAND_396[3:0];
  _RAND_397 = {1{`RANDOM}};
  image_2_13 = _RAND_397[3:0];
  _RAND_398 = {1{`RANDOM}};
  image_2_14 = _RAND_398[3:0];
  _RAND_399 = {1{`RANDOM}};
  image_2_15 = _RAND_399[3:0];
  _RAND_400 = {1{`RANDOM}};
  image_2_16 = _RAND_400[3:0];
  _RAND_401 = {1{`RANDOM}};
  image_2_17 = _RAND_401[3:0];
  _RAND_402 = {1{`RANDOM}};
  image_2_18 = _RAND_402[3:0];
  _RAND_403 = {1{`RANDOM}};
  image_2_19 = _RAND_403[3:0];
  _RAND_404 = {1{`RANDOM}};
  image_2_20 = _RAND_404[3:0];
  _RAND_405 = {1{`RANDOM}};
  image_2_21 = _RAND_405[3:0];
  _RAND_406 = {1{`RANDOM}};
  image_2_22 = _RAND_406[3:0];
  _RAND_407 = {1{`RANDOM}};
  image_2_23 = _RAND_407[3:0];
  _RAND_408 = {1{`RANDOM}};
  image_2_24 = _RAND_408[3:0];
  _RAND_409 = {1{`RANDOM}};
  image_2_25 = _RAND_409[3:0];
  _RAND_410 = {1{`RANDOM}};
  image_2_26 = _RAND_410[3:0];
  _RAND_411 = {1{`RANDOM}};
  image_2_27 = _RAND_411[3:0];
  _RAND_412 = {1{`RANDOM}};
  image_2_28 = _RAND_412[3:0];
  _RAND_413 = {1{`RANDOM}};
  image_2_29 = _RAND_413[3:0];
  _RAND_414 = {1{`RANDOM}};
  image_2_30 = _RAND_414[3:0];
  _RAND_415 = {1{`RANDOM}};
  image_2_31 = _RAND_415[3:0];
  _RAND_416 = {1{`RANDOM}};
  image_2_32 = _RAND_416[3:0];
  _RAND_417 = {1{`RANDOM}};
  image_2_33 = _RAND_417[3:0];
  _RAND_418 = {1{`RANDOM}};
  image_2_34 = _RAND_418[3:0];
  _RAND_419 = {1{`RANDOM}};
  image_2_35 = _RAND_419[3:0];
  _RAND_420 = {1{`RANDOM}};
  image_2_36 = _RAND_420[3:0];
  _RAND_421 = {1{`RANDOM}};
  image_2_37 = _RAND_421[3:0];
  _RAND_422 = {1{`RANDOM}};
  image_2_38 = _RAND_422[3:0];
  _RAND_423 = {1{`RANDOM}};
  image_2_39 = _RAND_423[3:0];
  _RAND_424 = {1{`RANDOM}};
  image_2_40 = _RAND_424[3:0];
  _RAND_425 = {1{`RANDOM}};
  image_2_41 = _RAND_425[3:0];
  _RAND_426 = {1{`RANDOM}};
  image_2_42 = _RAND_426[3:0];
  _RAND_427 = {1{`RANDOM}};
  image_2_43 = _RAND_427[3:0];
  _RAND_428 = {1{`RANDOM}};
  image_2_44 = _RAND_428[3:0];
  _RAND_429 = {1{`RANDOM}};
  image_2_45 = _RAND_429[3:0];
  _RAND_430 = {1{`RANDOM}};
  image_2_46 = _RAND_430[3:0];
  _RAND_431 = {1{`RANDOM}};
  image_2_47 = _RAND_431[3:0];
  _RAND_432 = {1{`RANDOM}};
  image_2_48 = _RAND_432[3:0];
  _RAND_433 = {1{`RANDOM}};
  image_2_49 = _RAND_433[3:0];
  _RAND_434 = {1{`RANDOM}};
  image_2_50 = _RAND_434[3:0];
  _RAND_435 = {1{`RANDOM}};
  image_2_51 = _RAND_435[3:0];
  _RAND_436 = {1{`RANDOM}};
  image_2_52 = _RAND_436[3:0];
  _RAND_437 = {1{`RANDOM}};
  image_2_53 = _RAND_437[3:0];
  _RAND_438 = {1{`RANDOM}};
  image_2_54 = _RAND_438[3:0];
  _RAND_439 = {1{`RANDOM}};
  image_2_55 = _RAND_439[3:0];
  _RAND_440 = {1{`RANDOM}};
  image_2_56 = _RAND_440[3:0];
  _RAND_441 = {1{`RANDOM}};
  image_2_57 = _RAND_441[3:0];
  _RAND_442 = {1{`RANDOM}};
  image_2_58 = _RAND_442[3:0];
  _RAND_443 = {1{`RANDOM}};
  image_2_59 = _RAND_443[3:0];
  _RAND_444 = {1{`RANDOM}};
  image_2_60 = _RAND_444[3:0];
  _RAND_445 = {1{`RANDOM}};
  image_2_61 = _RAND_445[3:0];
  _RAND_446 = {1{`RANDOM}};
  image_2_62 = _RAND_446[3:0];
  _RAND_447 = {1{`RANDOM}};
  image_2_63 = _RAND_447[3:0];
  _RAND_448 = {1{`RANDOM}};
  image_2_64 = _RAND_448[3:0];
  _RAND_449 = {1{`RANDOM}};
  image_2_65 = _RAND_449[3:0];
  _RAND_450 = {1{`RANDOM}};
  image_2_66 = _RAND_450[3:0];
  _RAND_451 = {1{`RANDOM}};
  image_2_67 = _RAND_451[3:0];
  _RAND_452 = {1{`RANDOM}};
  image_2_68 = _RAND_452[3:0];
  _RAND_453 = {1{`RANDOM}};
  image_2_69 = _RAND_453[3:0];
  _RAND_454 = {1{`RANDOM}};
  image_2_70 = _RAND_454[3:0];
  _RAND_455 = {1{`RANDOM}};
  image_2_71 = _RAND_455[3:0];
  _RAND_456 = {1{`RANDOM}};
  image_2_72 = _RAND_456[3:0];
  _RAND_457 = {1{`RANDOM}};
  image_2_73 = _RAND_457[3:0];
  _RAND_458 = {1{`RANDOM}};
  image_2_74 = _RAND_458[3:0];
  _RAND_459 = {1{`RANDOM}};
  image_2_75 = _RAND_459[3:0];
  _RAND_460 = {1{`RANDOM}};
  image_2_76 = _RAND_460[3:0];
  _RAND_461 = {1{`RANDOM}};
  image_2_77 = _RAND_461[3:0];
  _RAND_462 = {1{`RANDOM}};
  image_2_78 = _RAND_462[3:0];
  _RAND_463 = {1{`RANDOM}};
  image_2_79 = _RAND_463[3:0];
  _RAND_464 = {1{`RANDOM}};
  image_2_80 = _RAND_464[3:0];
  _RAND_465 = {1{`RANDOM}};
  image_2_81 = _RAND_465[3:0];
  _RAND_466 = {1{`RANDOM}};
  image_2_82 = _RAND_466[3:0];
  _RAND_467 = {1{`RANDOM}};
  image_2_83 = _RAND_467[3:0];
  _RAND_468 = {1{`RANDOM}};
  image_2_84 = _RAND_468[3:0];
  _RAND_469 = {1{`RANDOM}};
  image_2_85 = _RAND_469[3:0];
  _RAND_470 = {1{`RANDOM}};
  image_2_86 = _RAND_470[3:0];
  _RAND_471 = {1{`RANDOM}};
  image_2_87 = _RAND_471[3:0];
  _RAND_472 = {1{`RANDOM}};
  image_2_88 = _RAND_472[3:0];
  _RAND_473 = {1{`RANDOM}};
  image_2_89 = _RAND_473[3:0];
  _RAND_474 = {1{`RANDOM}};
  image_2_90 = _RAND_474[3:0];
  _RAND_475 = {1{`RANDOM}};
  image_2_91 = _RAND_475[3:0];
  _RAND_476 = {1{`RANDOM}};
  image_2_92 = _RAND_476[3:0];
  _RAND_477 = {1{`RANDOM}};
  image_2_93 = _RAND_477[3:0];
  _RAND_478 = {1{`RANDOM}};
  image_2_94 = _RAND_478[3:0];
  _RAND_479 = {1{`RANDOM}};
  image_2_95 = _RAND_479[3:0];
  _RAND_480 = {1{`RANDOM}};
  image_2_96 = _RAND_480[3:0];
  _RAND_481 = {1{`RANDOM}};
  image_2_97 = _RAND_481[3:0];
  _RAND_482 = {1{`RANDOM}};
  image_2_98 = _RAND_482[3:0];
  _RAND_483 = {1{`RANDOM}};
  image_2_99 = _RAND_483[3:0];
  _RAND_484 = {1{`RANDOM}};
  image_2_100 = _RAND_484[3:0];
  _RAND_485 = {1{`RANDOM}};
  image_2_101 = _RAND_485[3:0];
  _RAND_486 = {1{`RANDOM}};
  image_2_102 = _RAND_486[3:0];
  _RAND_487 = {1{`RANDOM}};
  image_2_103 = _RAND_487[3:0];
  _RAND_488 = {1{`RANDOM}};
  image_2_104 = _RAND_488[3:0];
  _RAND_489 = {1{`RANDOM}};
  image_2_105 = _RAND_489[3:0];
  _RAND_490 = {1{`RANDOM}};
  image_2_106 = _RAND_490[3:0];
  _RAND_491 = {1{`RANDOM}};
  image_2_107 = _RAND_491[3:0];
  _RAND_492 = {1{`RANDOM}};
  image_2_108 = _RAND_492[3:0];
  _RAND_493 = {1{`RANDOM}};
  image_2_109 = _RAND_493[3:0];
  _RAND_494 = {1{`RANDOM}};
  image_2_110 = _RAND_494[3:0];
  _RAND_495 = {1{`RANDOM}};
  image_2_111 = _RAND_495[3:0];
  _RAND_496 = {1{`RANDOM}};
  image_2_112 = _RAND_496[3:0];
  _RAND_497 = {1{`RANDOM}};
  image_2_113 = _RAND_497[3:0];
  _RAND_498 = {1{`RANDOM}};
  image_2_114 = _RAND_498[3:0];
  _RAND_499 = {1{`RANDOM}};
  image_2_115 = _RAND_499[3:0];
  _RAND_500 = {1{`RANDOM}};
  image_2_116 = _RAND_500[3:0];
  _RAND_501 = {1{`RANDOM}};
  image_2_117 = _RAND_501[3:0];
  _RAND_502 = {1{`RANDOM}};
  image_2_118 = _RAND_502[3:0];
  _RAND_503 = {1{`RANDOM}};
  image_2_119 = _RAND_503[3:0];
  _RAND_504 = {1{`RANDOM}};
  image_2_120 = _RAND_504[3:0];
  _RAND_505 = {1{`RANDOM}};
  image_2_121 = _RAND_505[3:0];
  _RAND_506 = {1{`RANDOM}};
  image_2_122 = _RAND_506[3:0];
  _RAND_507 = {1{`RANDOM}};
  image_2_123 = _RAND_507[3:0];
  _RAND_508 = {1{`RANDOM}};
  image_2_124 = _RAND_508[3:0];
  _RAND_509 = {1{`RANDOM}};
  image_2_125 = _RAND_509[3:0];
  _RAND_510 = {1{`RANDOM}};
  image_2_126 = _RAND_510[3:0];
  _RAND_511 = {1{`RANDOM}};
  image_2_127 = _RAND_511[3:0];
  _RAND_512 = {1{`RANDOM}};
  image_2_128 = _RAND_512[3:0];
  _RAND_513 = {1{`RANDOM}};
  image_2_129 = _RAND_513[3:0];
  _RAND_514 = {1{`RANDOM}};
  image_2_130 = _RAND_514[3:0];
  _RAND_515 = {1{`RANDOM}};
  image_2_131 = _RAND_515[3:0];
  _RAND_516 = {1{`RANDOM}};
  image_2_132 = _RAND_516[3:0];
  _RAND_517 = {1{`RANDOM}};
  image_2_133 = _RAND_517[3:0];
  _RAND_518 = {1{`RANDOM}};
  image_2_134 = _RAND_518[3:0];
  _RAND_519 = {1{`RANDOM}};
  image_2_135 = _RAND_519[3:0];
  _RAND_520 = {1{`RANDOM}};
  image_2_136 = _RAND_520[3:0];
  _RAND_521 = {1{`RANDOM}};
  image_2_137 = _RAND_521[3:0];
  _RAND_522 = {1{`RANDOM}};
  image_2_138 = _RAND_522[3:0];
  _RAND_523 = {1{`RANDOM}};
  image_2_139 = _RAND_523[3:0];
  _RAND_524 = {1{`RANDOM}};
  image_2_140 = _RAND_524[3:0];
  _RAND_525 = {1{`RANDOM}};
  image_2_141 = _RAND_525[3:0];
  _RAND_526 = {1{`RANDOM}};
  image_2_142 = _RAND_526[3:0];
  _RAND_527 = {1{`RANDOM}};
  image_2_143 = _RAND_527[3:0];
  _RAND_528 = {1{`RANDOM}};
  image_2_144 = _RAND_528[3:0];
  _RAND_529 = {1{`RANDOM}};
  image_2_145 = _RAND_529[3:0];
  _RAND_530 = {1{`RANDOM}};
  image_2_146 = _RAND_530[3:0];
  _RAND_531 = {1{`RANDOM}};
  image_2_147 = _RAND_531[3:0];
  _RAND_532 = {1{`RANDOM}};
  image_2_148 = _RAND_532[3:0];
  _RAND_533 = {1{`RANDOM}};
  image_2_149 = _RAND_533[3:0];
  _RAND_534 = {1{`RANDOM}};
  image_2_150 = _RAND_534[3:0];
  _RAND_535 = {1{`RANDOM}};
  image_2_151 = _RAND_535[3:0];
  _RAND_536 = {1{`RANDOM}};
  image_2_152 = _RAND_536[3:0];
  _RAND_537 = {1{`RANDOM}};
  image_2_153 = _RAND_537[3:0];
  _RAND_538 = {1{`RANDOM}};
  image_2_154 = _RAND_538[3:0];
  _RAND_539 = {1{`RANDOM}};
  image_2_155 = _RAND_539[3:0];
  _RAND_540 = {1{`RANDOM}};
  image_2_156 = _RAND_540[3:0];
  _RAND_541 = {1{`RANDOM}};
  image_2_157 = _RAND_541[3:0];
  _RAND_542 = {1{`RANDOM}};
  image_2_158 = _RAND_542[3:0];
  _RAND_543 = {1{`RANDOM}};
  image_2_159 = _RAND_543[3:0];
  _RAND_544 = {1{`RANDOM}};
  image_2_160 = _RAND_544[3:0];
  _RAND_545 = {1{`RANDOM}};
  image_2_161 = _RAND_545[3:0];
  _RAND_546 = {1{`RANDOM}};
  image_2_162 = _RAND_546[3:0];
  _RAND_547 = {1{`RANDOM}};
  image_2_163 = _RAND_547[3:0];
  _RAND_548 = {1{`RANDOM}};
  image_2_164 = _RAND_548[3:0];
  _RAND_549 = {1{`RANDOM}};
  image_2_165 = _RAND_549[3:0];
  _RAND_550 = {1{`RANDOM}};
  image_2_166 = _RAND_550[3:0];
  _RAND_551 = {1{`RANDOM}};
  image_2_167 = _RAND_551[3:0];
  _RAND_552 = {1{`RANDOM}};
  image_2_168 = _RAND_552[3:0];
  _RAND_553 = {1{`RANDOM}};
  image_2_169 = _RAND_553[3:0];
  _RAND_554 = {1{`RANDOM}};
  image_2_170 = _RAND_554[3:0];
  _RAND_555 = {1{`RANDOM}};
  image_2_171 = _RAND_555[3:0];
  _RAND_556 = {1{`RANDOM}};
  image_2_172 = _RAND_556[3:0];
  _RAND_557 = {1{`RANDOM}};
  image_2_173 = _RAND_557[3:0];
  _RAND_558 = {1{`RANDOM}};
  image_2_174 = _RAND_558[3:0];
  _RAND_559 = {1{`RANDOM}};
  image_2_175 = _RAND_559[3:0];
  _RAND_560 = {1{`RANDOM}};
  image_2_176 = _RAND_560[3:0];
  _RAND_561 = {1{`RANDOM}};
  image_2_177 = _RAND_561[3:0];
  _RAND_562 = {1{`RANDOM}};
  image_2_178 = _RAND_562[3:0];
  _RAND_563 = {1{`RANDOM}};
  image_2_179 = _RAND_563[3:0];
  _RAND_564 = {1{`RANDOM}};
  image_2_180 = _RAND_564[3:0];
  _RAND_565 = {1{`RANDOM}};
  image_2_181 = _RAND_565[3:0];
  _RAND_566 = {1{`RANDOM}};
  image_2_182 = _RAND_566[3:0];
  _RAND_567 = {1{`RANDOM}};
  image_2_183 = _RAND_567[3:0];
  _RAND_568 = {1{`RANDOM}};
  image_2_184 = _RAND_568[3:0];
  _RAND_569 = {1{`RANDOM}};
  image_2_185 = _RAND_569[3:0];
  _RAND_570 = {1{`RANDOM}};
  image_2_186 = _RAND_570[3:0];
  _RAND_571 = {1{`RANDOM}};
  image_2_187 = _RAND_571[3:0];
  _RAND_572 = {1{`RANDOM}};
  image_2_188 = _RAND_572[3:0];
  _RAND_573 = {1{`RANDOM}};
  image_2_189 = _RAND_573[3:0];
  _RAND_574 = {1{`RANDOM}};
  image_2_190 = _RAND_574[3:0];
  _RAND_575 = {1{`RANDOM}};
  image_2_191 = _RAND_575[3:0];
  _RAND_576 = {1{`RANDOM}};
  pixelIndex = _RAND_576[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      image_0_0 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h0 == _T_29[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_7;
      end else if (8'h0 == _T_26[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_6;
      end else if (8'h0 == _T_23[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_5;
      end else if (8'h0 == _T_20[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_4;
      end else if (8'h0 == _T_17[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_3;
      end else if (8'h0 == _T_14[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_2;
      end else if (8'h0 == _T_11[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_1;
      end else if (8'h0 == _T_7[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_1 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1 == _T_29[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_7;
      end else if (8'h1 == _T_26[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_6;
      end else if (8'h1 == _T_23[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_5;
      end else if (8'h1 == _T_20[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_4;
      end else if (8'h1 == _T_17[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_3;
      end else if (8'h1 == _T_14[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_2;
      end else if (8'h1 == _T_11[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_1;
      end else if (8'h1 == _T_7[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_2 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2 == _T_29[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_7;
      end else if (8'h2 == _T_26[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_6;
      end else if (8'h2 == _T_23[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_5;
      end else if (8'h2 == _T_20[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_4;
      end else if (8'h2 == _T_17[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_3;
      end else if (8'h2 == _T_14[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_2;
      end else if (8'h2 == _T_11[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_1;
      end else if (8'h2 == _T_7[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_3 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3 == _T_29[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_7;
      end else if (8'h3 == _T_26[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_6;
      end else if (8'h3 == _T_23[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_5;
      end else if (8'h3 == _T_20[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_4;
      end else if (8'h3 == _T_17[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_3;
      end else if (8'h3 == _T_14[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_2;
      end else if (8'h3 == _T_11[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_1;
      end else if (8'h3 == _T_7[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_4 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4 == _T_29[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_7;
      end else if (8'h4 == _T_26[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_6;
      end else if (8'h4 == _T_23[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_5;
      end else if (8'h4 == _T_20[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_4;
      end else if (8'h4 == _T_17[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_3;
      end else if (8'h4 == _T_14[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_2;
      end else if (8'h4 == _T_11[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_1;
      end else if (8'h4 == _T_7[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_5 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5 == _T_29[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_7;
      end else if (8'h5 == _T_26[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_6;
      end else if (8'h5 == _T_23[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_5;
      end else if (8'h5 == _T_20[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_4;
      end else if (8'h5 == _T_17[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_3;
      end else if (8'h5 == _T_14[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_2;
      end else if (8'h5 == _T_11[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_1;
      end else if (8'h5 == _T_7[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_6 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6 == _T_29[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_7;
      end else if (8'h6 == _T_26[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_6;
      end else if (8'h6 == _T_23[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_5;
      end else if (8'h6 == _T_20[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_4;
      end else if (8'h6 == _T_17[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_3;
      end else if (8'h6 == _T_14[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_2;
      end else if (8'h6 == _T_11[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_1;
      end else if (8'h6 == _T_7[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_7 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7 == _T_29[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_7;
      end else if (8'h7 == _T_26[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_6;
      end else if (8'h7 == _T_23[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_5;
      end else if (8'h7 == _T_20[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_4;
      end else if (8'h7 == _T_17[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_3;
      end else if (8'h7 == _T_14[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_2;
      end else if (8'h7 == _T_11[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_1;
      end else if (8'h7 == _T_7[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_8 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8 == _T_29[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_7;
      end else if (8'h8 == _T_26[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_6;
      end else if (8'h8 == _T_23[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_5;
      end else if (8'h8 == _T_20[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_4;
      end else if (8'h8 == _T_17[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_3;
      end else if (8'h8 == _T_14[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_2;
      end else if (8'h8 == _T_11[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_1;
      end else if (8'h8 == _T_7[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_9 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h9 == _T_29[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_7;
      end else if (8'h9 == _T_26[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_6;
      end else if (8'h9 == _T_23[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_5;
      end else if (8'h9 == _T_20[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_4;
      end else if (8'h9 == _T_17[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_3;
      end else if (8'h9 == _T_14[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_2;
      end else if (8'h9 == _T_11[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_1;
      end else if (8'h9 == _T_7[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_10 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha == _T_29[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_7;
      end else if (8'ha == _T_26[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_6;
      end else if (8'ha == _T_23[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_5;
      end else if (8'ha == _T_20[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_4;
      end else if (8'ha == _T_17[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_3;
      end else if (8'ha == _T_14[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_2;
      end else if (8'ha == _T_11[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_1;
      end else if (8'ha == _T_7[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_11 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb == _T_29[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_7;
      end else if (8'hb == _T_26[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_6;
      end else if (8'hb == _T_23[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_5;
      end else if (8'hb == _T_20[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_4;
      end else if (8'hb == _T_17[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_3;
      end else if (8'hb == _T_14[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_2;
      end else if (8'hb == _T_11[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_1;
      end else if (8'hb == _T_7[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_12 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hc == _T_29[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_7;
      end else if (8'hc == _T_26[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_6;
      end else if (8'hc == _T_23[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_5;
      end else if (8'hc == _T_20[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_4;
      end else if (8'hc == _T_17[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_3;
      end else if (8'hc == _T_14[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_2;
      end else if (8'hc == _T_11[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_1;
      end else if (8'hc == _T_7[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_13 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hd == _T_29[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_7;
      end else if (8'hd == _T_26[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_6;
      end else if (8'hd == _T_23[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_5;
      end else if (8'hd == _T_20[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_4;
      end else if (8'hd == _T_17[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_3;
      end else if (8'hd == _T_14[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_2;
      end else if (8'hd == _T_11[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_1;
      end else if (8'hd == _T_7[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_14 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'he == _T_29[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_7;
      end else if (8'he == _T_26[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_6;
      end else if (8'he == _T_23[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_5;
      end else if (8'he == _T_20[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_4;
      end else if (8'he == _T_17[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_3;
      end else if (8'he == _T_14[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_2;
      end else if (8'he == _T_11[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_1;
      end else if (8'he == _T_7[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_15 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hf == _T_29[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_7;
      end else if (8'hf == _T_26[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_6;
      end else if (8'hf == _T_23[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_5;
      end else if (8'hf == _T_20[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_4;
      end else if (8'hf == _T_17[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_3;
      end else if (8'hf == _T_14[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_2;
      end else if (8'hf == _T_11[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_1;
      end else if (8'hf == _T_7[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_16 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h10 == _T_29[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_7;
      end else if (8'h10 == _T_26[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_6;
      end else if (8'h10 == _T_23[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_5;
      end else if (8'h10 == _T_20[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_4;
      end else if (8'h10 == _T_17[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_3;
      end else if (8'h10 == _T_14[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_2;
      end else if (8'h10 == _T_11[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_1;
      end else if (8'h10 == _T_7[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_17 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h11 == _T_29[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_7;
      end else if (8'h11 == _T_26[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_6;
      end else if (8'h11 == _T_23[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_5;
      end else if (8'h11 == _T_20[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_4;
      end else if (8'h11 == _T_17[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_3;
      end else if (8'h11 == _T_14[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_2;
      end else if (8'h11 == _T_11[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_1;
      end else if (8'h11 == _T_7[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_18 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h12 == _T_29[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_7;
      end else if (8'h12 == _T_26[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_6;
      end else if (8'h12 == _T_23[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_5;
      end else if (8'h12 == _T_20[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_4;
      end else if (8'h12 == _T_17[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_3;
      end else if (8'h12 == _T_14[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_2;
      end else if (8'h12 == _T_11[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_1;
      end else if (8'h12 == _T_7[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_19 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h13 == _T_29[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_7;
      end else if (8'h13 == _T_26[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_6;
      end else if (8'h13 == _T_23[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_5;
      end else if (8'h13 == _T_20[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_4;
      end else if (8'h13 == _T_17[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_3;
      end else if (8'h13 == _T_14[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_2;
      end else if (8'h13 == _T_11[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_1;
      end else if (8'h13 == _T_7[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_20 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h14 == _T_29[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_7;
      end else if (8'h14 == _T_26[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_6;
      end else if (8'h14 == _T_23[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_5;
      end else if (8'h14 == _T_20[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_4;
      end else if (8'h14 == _T_17[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_3;
      end else if (8'h14 == _T_14[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_2;
      end else if (8'h14 == _T_11[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_1;
      end else if (8'h14 == _T_7[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_21 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h15 == _T_29[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_7;
      end else if (8'h15 == _T_26[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_6;
      end else if (8'h15 == _T_23[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_5;
      end else if (8'h15 == _T_20[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_4;
      end else if (8'h15 == _T_17[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_3;
      end else if (8'h15 == _T_14[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_2;
      end else if (8'h15 == _T_11[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_1;
      end else if (8'h15 == _T_7[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_22 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h16 == _T_29[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_7;
      end else if (8'h16 == _T_26[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_6;
      end else if (8'h16 == _T_23[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_5;
      end else if (8'h16 == _T_20[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_4;
      end else if (8'h16 == _T_17[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_3;
      end else if (8'h16 == _T_14[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_2;
      end else if (8'h16 == _T_11[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_1;
      end else if (8'h16 == _T_7[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_23 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h17 == _T_29[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_7;
      end else if (8'h17 == _T_26[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_6;
      end else if (8'h17 == _T_23[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_5;
      end else if (8'h17 == _T_20[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_4;
      end else if (8'h17 == _T_17[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_3;
      end else if (8'h17 == _T_14[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_2;
      end else if (8'h17 == _T_11[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_1;
      end else if (8'h17 == _T_7[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_24 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h18 == _T_29[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_7;
      end else if (8'h18 == _T_26[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_6;
      end else if (8'h18 == _T_23[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_5;
      end else if (8'h18 == _T_20[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_4;
      end else if (8'h18 == _T_17[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_3;
      end else if (8'h18 == _T_14[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_2;
      end else if (8'h18 == _T_11[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_1;
      end else if (8'h18 == _T_7[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_25 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h19 == _T_29[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_7;
      end else if (8'h19 == _T_26[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_6;
      end else if (8'h19 == _T_23[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_5;
      end else if (8'h19 == _T_20[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_4;
      end else if (8'h19 == _T_17[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_3;
      end else if (8'h19 == _T_14[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_2;
      end else if (8'h19 == _T_11[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_1;
      end else if (8'h19 == _T_7[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_26 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1a == _T_29[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_7;
      end else if (8'h1a == _T_26[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_6;
      end else if (8'h1a == _T_23[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_5;
      end else if (8'h1a == _T_20[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_4;
      end else if (8'h1a == _T_17[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_3;
      end else if (8'h1a == _T_14[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_2;
      end else if (8'h1a == _T_11[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_1;
      end else if (8'h1a == _T_7[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_27 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1b == _T_29[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_7;
      end else if (8'h1b == _T_26[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_6;
      end else if (8'h1b == _T_23[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_5;
      end else if (8'h1b == _T_20[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_4;
      end else if (8'h1b == _T_17[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_3;
      end else if (8'h1b == _T_14[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_2;
      end else if (8'h1b == _T_11[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_1;
      end else if (8'h1b == _T_7[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_28 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1c == _T_29[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_7;
      end else if (8'h1c == _T_26[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_6;
      end else if (8'h1c == _T_23[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_5;
      end else if (8'h1c == _T_20[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_4;
      end else if (8'h1c == _T_17[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_3;
      end else if (8'h1c == _T_14[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_2;
      end else if (8'h1c == _T_11[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_1;
      end else if (8'h1c == _T_7[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_29 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1d == _T_29[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_7;
      end else if (8'h1d == _T_26[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_6;
      end else if (8'h1d == _T_23[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_5;
      end else if (8'h1d == _T_20[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_4;
      end else if (8'h1d == _T_17[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_3;
      end else if (8'h1d == _T_14[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_2;
      end else if (8'h1d == _T_11[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_1;
      end else if (8'h1d == _T_7[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_30 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1e == _T_29[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_7;
      end else if (8'h1e == _T_26[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_6;
      end else if (8'h1e == _T_23[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_5;
      end else if (8'h1e == _T_20[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_4;
      end else if (8'h1e == _T_17[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_3;
      end else if (8'h1e == _T_14[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_2;
      end else if (8'h1e == _T_11[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_1;
      end else if (8'h1e == _T_7[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_31 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1f == _T_29[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_7;
      end else if (8'h1f == _T_26[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_6;
      end else if (8'h1f == _T_23[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_5;
      end else if (8'h1f == _T_20[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_4;
      end else if (8'h1f == _T_17[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_3;
      end else if (8'h1f == _T_14[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_2;
      end else if (8'h1f == _T_11[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_1;
      end else if (8'h1f == _T_7[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_32 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h20 == _T_29[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_7;
      end else if (8'h20 == _T_26[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_6;
      end else if (8'h20 == _T_23[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_5;
      end else if (8'h20 == _T_20[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_4;
      end else if (8'h20 == _T_17[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_3;
      end else if (8'h20 == _T_14[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_2;
      end else if (8'h20 == _T_11[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_1;
      end else if (8'h20 == _T_7[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_33 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h21 == _T_29[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_7;
      end else if (8'h21 == _T_26[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_6;
      end else if (8'h21 == _T_23[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_5;
      end else if (8'h21 == _T_20[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_4;
      end else if (8'h21 == _T_17[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_3;
      end else if (8'h21 == _T_14[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_2;
      end else if (8'h21 == _T_11[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_1;
      end else if (8'h21 == _T_7[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_34 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h22 == _T_29[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_7;
      end else if (8'h22 == _T_26[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_6;
      end else if (8'h22 == _T_23[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_5;
      end else if (8'h22 == _T_20[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_4;
      end else if (8'h22 == _T_17[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_3;
      end else if (8'h22 == _T_14[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_2;
      end else if (8'h22 == _T_11[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_1;
      end else if (8'h22 == _T_7[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_35 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h23 == _T_29[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_7;
      end else if (8'h23 == _T_26[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_6;
      end else if (8'h23 == _T_23[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_5;
      end else if (8'h23 == _T_20[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_4;
      end else if (8'h23 == _T_17[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_3;
      end else if (8'h23 == _T_14[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_2;
      end else if (8'h23 == _T_11[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_1;
      end else if (8'h23 == _T_7[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_36 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h24 == _T_29[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_7;
      end else if (8'h24 == _T_26[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_6;
      end else if (8'h24 == _T_23[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_5;
      end else if (8'h24 == _T_20[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_4;
      end else if (8'h24 == _T_17[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_3;
      end else if (8'h24 == _T_14[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_2;
      end else if (8'h24 == _T_11[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_1;
      end else if (8'h24 == _T_7[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_37 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h25 == _T_29[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_7;
      end else if (8'h25 == _T_26[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_6;
      end else if (8'h25 == _T_23[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_5;
      end else if (8'h25 == _T_20[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_4;
      end else if (8'h25 == _T_17[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_3;
      end else if (8'h25 == _T_14[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_2;
      end else if (8'h25 == _T_11[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_1;
      end else if (8'h25 == _T_7[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_38 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h26 == _T_29[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_7;
      end else if (8'h26 == _T_26[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_6;
      end else if (8'h26 == _T_23[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_5;
      end else if (8'h26 == _T_20[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_4;
      end else if (8'h26 == _T_17[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_3;
      end else if (8'h26 == _T_14[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_2;
      end else if (8'h26 == _T_11[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_1;
      end else if (8'h26 == _T_7[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_39 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h27 == _T_29[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_7;
      end else if (8'h27 == _T_26[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_6;
      end else if (8'h27 == _T_23[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_5;
      end else if (8'h27 == _T_20[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_4;
      end else if (8'h27 == _T_17[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_3;
      end else if (8'h27 == _T_14[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_2;
      end else if (8'h27 == _T_11[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_1;
      end else if (8'h27 == _T_7[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_40 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h28 == _T_29[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_7;
      end else if (8'h28 == _T_26[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_6;
      end else if (8'h28 == _T_23[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_5;
      end else if (8'h28 == _T_20[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_4;
      end else if (8'h28 == _T_17[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_3;
      end else if (8'h28 == _T_14[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_2;
      end else if (8'h28 == _T_11[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_1;
      end else if (8'h28 == _T_7[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_41 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h29 == _T_29[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_7;
      end else if (8'h29 == _T_26[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_6;
      end else if (8'h29 == _T_23[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_5;
      end else if (8'h29 == _T_20[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_4;
      end else if (8'h29 == _T_17[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_3;
      end else if (8'h29 == _T_14[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_2;
      end else if (8'h29 == _T_11[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_1;
      end else if (8'h29 == _T_7[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_42 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2a == _T_29[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_7;
      end else if (8'h2a == _T_26[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_6;
      end else if (8'h2a == _T_23[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_5;
      end else if (8'h2a == _T_20[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_4;
      end else if (8'h2a == _T_17[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_3;
      end else if (8'h2a == _T_14[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_2;
      end else if (8'h2a == _T_11[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_1;
      end else if (8'h2a == _T_7[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_43 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2b == _T_29[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_7;
      end else if (8'h2b == _T_26[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_6;
      end else if (8'h2b == _T_23[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_5;
      end else if (8'h2b == _T_20[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_4;
      end else if (8'h2b == _T_17[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_3;
      end else if (8'h2b == _T_14[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_2;
      end else if (8'h2b == _T_11[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_1;
      end else if (8'h2b == _T_7[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_44 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2c == _T_29[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_7;
      end else if (8'h2c == _T_26[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_6;
      end else if (8'h2c == _T_23[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_5;
      end else if (8'h2c == _T_20[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_4;
      end else if (8'h2c == _T_17[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_3;
      end else if (8'h2c == _T_14[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_2;
      end else if (8'h2c == _T_11[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_1;
      end else if (8'h2c == _T_7[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_45 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2d == _T_29[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_7;
      end else if (8'h2d == _T_26[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_6;
      end else if (8'h2d == _T_23[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_5;
      end else if (8'h2d == _T_20[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_4;
      end else if (8'h2d == _T_17[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_3;
      end else if (8'h2d == _T_14[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_2;
      end else if (8'h2d == _T_11[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_1;
      end else if (8'h2d == _T_7[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_46 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2e == _T_29[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_7;
      end else if (8'h2e == _T_26[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_6;
      end else if (8'h2e == _T_23[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_5;
      end else if (8'h2e == _T_20[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_4;
      end else if (8'h2e == _T_17[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_3;
      end else if (8'h2e == _T_14[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_2;
      end else if (8'h2e == _T_11[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_1;
      end else if (8'h2e == _T_7[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_47 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2f == _T_29[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_7;
      end else if (8'h2f == _T_26[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_6;
      end else if (8'h2f == _T_23[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_5;
      end else if (8'h2f == _T_20[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_4;
      end else if (8'h2f == _T_17[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_3;
      end else if (8'h2f == _T_14[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_2;
      end else if (8'h2f == _T_11[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_1;
      end else if (8'h2f == _T_7[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_48 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h30 == _T_29[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_7;
      end else if (8'h30 == _T_26[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_6;
      end else if (8'h30 == _T_23[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_5;
      end else if (8'h30 == _T_20[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_4;
      end else if (8'h30 == _T_17[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_3;
      end else if (8'h30 == _T_14[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_2;
      end else if (8'h30 == _T_11[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_1;
      end else if (8'h30 == _T_7[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_49 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h31 == _T_29[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_7;
      end else if (8'h31 == _T_26[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_6;
      end else if (8'h31 == _T_23[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_5;
      end else if (8'h31 == _T_20[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_4;
      end else if (8'h31 == _T_17[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_3;
      end else if (8'h31 == _T_14[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_2;
      end else if (8'h31 == _T_11[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_1;
      end else if (8'h31 == _T_7[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_50 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h32 == _T_29[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_7;
      end else if (8'h32 == _T_26[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_6;
      end else if (8'h32 == _T_23[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_5;
      end else if (8'h32 == _T_20[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_4;
      end else if (8'h32 == _T_17[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_3;
      end else if (8'h32 == _T_14[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_2;
      end else if (8'h32 == _T_11[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_1;
      end else if (8'h32 == _T_7[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_51 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h33 == _T_29[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_7;
      end else if (8'h33 == _T_26[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_6;
      end else if (8'h33 == _T_23[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_5;
      end else if (8'h33 == _T_20[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_4;
      end else if (8'h33 == _T_17[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_3;
      end else if (8'h33 == _T_14[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_2;
      end else if (8'h33 == _T_11[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_1;
      end else if (8'h33 == _T_7[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_52 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h34 == _T_29[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_7;
      end else if (8'h34 == _T_26[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_6;
      end else if (8'h34 == _T_23[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_5;
      end else if (8'h34 == _T_20[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_4;
      end else if (8'h34 == _T_17[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_3;
      end else if (8'h34 == _T_14[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_2;
      end else if (8'h34 == _T_11[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_1;
      end else if (8'h34 == _T_7[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_53 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h35 == _T_29[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_7;
      end else if (8'h35 == _T_26[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_6;
      end else if (8'h35 == _T_23[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_5;
      end else if (8'h35 == _T_20[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_4;
      end else if (8'h35 == _T_17[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_3;
      end else if (8'h35 == _T_14[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_2;
      end else if (8'h35 == _T_11[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_1;
      end else if (8'h35 == _T_7[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_54 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h36 == _T_29[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_7;
      end else if (8'h36 == _T_26[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_6;
      end else if (8'h36 == _T_23[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_5;
      end else if (8'h36 == _T_20[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_4;
      end else if (8'h36 == _T_17[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_3;
      end else if (8'h36 == _T_14[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_2;
      end else if (8'h36 == _T_11[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_1;
      end else if (8'h36 == _T_7[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_55 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h37 == _T_29[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_7;
      end else if (8'h37 == _T_26[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_6;
      end else if (8'h37 == _T_23[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_5;
      end else if (8'h37 == _T_20[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_4;
      end else if (8'h37 == _T_17[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_3;
      end else if (8'h37 == _T_14[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_2;
      end else if (8'h37 == _T_11[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_1;
      end else if (8'h37 == _T_7[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_56 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h38 == _T_29[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_7;
      end else if (8'h38 == _T_26[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_6;
      end else if (8'h38 == _T_23[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_5;
      end else if (8'h38 == _T_20[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_4;
      end else if (8'h38 == _T_17[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_3;
      end else if (8'h38 == _T_14[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_2;
      end else if (8'h38 == _T_11[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_1;
      end else if (8'h38 == _T_7[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_57 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h39 == _T_29[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_7;
      end else if (8'h39 == _T_26[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_6;
      end else if (8'h39 == _T_23[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_5;
      end else if (8'h39 == _T_20[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_4;
      end else if (8'h39 == _T_17[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_3;
      end else if (8'h39 == _T_14[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_2;
      end else if (8'h39 == _T_11[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_1;
      end else if (8'h39 == _T_7[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_58 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3a == _T_29[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_7;
      end else if (8'h3a == _T_26[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_6;
      end else if (8'h3a == _T_23[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_5;
      end else if (8'h3a == _T_20[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_4;
      end else if (8'h3a == _T_17[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_3;
      end else if (8'h3a == _T_14[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_2;
      end else if (8'h3a == _T_11[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_1;
      end else if (8'h3a == _T_7[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_59 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3b == _T_29[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_7;
      end else if (8'h3b == _T_26[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_6;
      end else if (8'h3b == _T_23[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_5;
      end else if (8'h3b == _T_20[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_4;
      end else if (8'h3b == _T_17[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_3;
      end else if (8'h3b == _T_14[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_2;
      end else if (8'h3b == _T_11[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_1;
      end else if (8'h3b == _T_7[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_60 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3c == _T_29[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_7;
      end else if (8'h3c == _T_26[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_6;
      end else if (8'h3c == _T_23[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_5;
      end else if (8'h3c == _T_20[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_4;
      end else if (8'h3c == _T_17[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_3;
      end else if (8'h3c == _T_14[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_2;
      end else if (8'h3c == _T_11[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_1;
      end else if (8'h3c == _T_7[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_61 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3d == _T_29[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_7;
      end else if (8'h3d == _T_26[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_6;
      end else if (8'h3d == _T_23[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_5;
      end else if (8'h3d == _T_20[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_4;
      end else if (8'h3d == _T_17[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_3;
      end else if (8'h3d == _T_14[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_2;
      end else if (8'h3d == _T_11[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_1;
      end else if (8'h3d == _T_7[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_62 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3e == _T_29[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_7;
      end else if (8'h3e == _T_26[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_6;
      end else if (8'h3e == _T_23[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_5;
      end else if (8'h3e == _T_20[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_4;
      end else if (8'h3e == _T_17[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_3;
      end else if (8'h3e == _T_14[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_2;
      end else if (8'h3e == _T_11[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_1;
      end else if (8'h3e == _T_7[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_63 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3f == _T_29[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_7;
      end else if (8'h3f == _T_26[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_6;
      end else if (8'h3f == _T_23[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_5;
      end else if (8'h3f == _T_20[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_4;
      end else if (8'h3f == _T_17[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_3;
      end else if (8'h3f == _T_14[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_2;
      end else if (8'h3f == _T_11[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_1;
      end else if (8'h3f == _T_7[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_64 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h40 == _T_29[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_7;
      end else if (8'h40 == _T_26[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_6;
      end else if (8'h40 == _T_23[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_5;
      end else if (8'h40 == _T_20[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_4;
      end else if (8'h40 == _T_17[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_3;
      end else if (8'h40 == _T_14[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_2;
      end else if (8'h40 == _T_11[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_1;
      end else if (8'h40 == _T_7[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_65 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h41 == _T_29[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_7;
      end else if (8'h41 == _T_26[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_6;
      end else if (8'h41 == _T_23[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_5;
      end else if (8'h41 == _T_20[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_4;
      end else if (8'h41 == _T_17[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_3;
      end else if (8'h41 == _T_14[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_2;
      end else if (8'h41 == _T_11[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_1;
      end else if (8'h41 == _T_7[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_66 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h42 == _T_29[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_7;
      end else if (8'h42 == _T_26[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_6;
      end else if (8'h42 == _T_23[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_5;
      end else if (8'h42 == _T_20[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_4;
      end else if (8'h42 == _T_17[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_3;
      end else if (8'h42 == _T_14[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_2;
      end else if (8'h42 == _T_11[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_1;
      end else if (8'h42 == _T_7[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_67 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h43 == _T_29[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_7;
      end else if (8'h43 == _T_26[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_6;
      end else if (8'h43 == _T_23[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_5;
      end else if (8'h43 == _T_20[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_4;
      end else if (8'h43 == _T_17[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_3;
      end else if (8'h43 == _T_14[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_2;
      end else if (8'h43 == _T_11[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_1;
      end else if (8'h43 == _T_7[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_68 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h44 == _T_29[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_7;
      end else if (8'h44 == _T_26[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_6;
      end else if (8'h44 == _T_23[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_5;
      end else if (8'h44 == _T_20[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_4;
      end else if (8'h44 == _T_17[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_3;
      end else if (8'h44 == _T_14[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_2;
      end else if (8'h44 == _T_11[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_1;
      end else if (8'h44 == _T_7[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_69 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h45 == _T_29[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_7;
      end else if (8'h45 == _T_26[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_6;
      end else if (8'h45 == _T_23[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_5;
      end else if (8'h45 == _T_20[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_4;
      end else if (8'h45 == _T_17[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_3;
      end else if (8'h45 == _T_14[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_2;
      end else if (8'h45 == _T_11[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_1;
      end else if (8'h45 == _T_7[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_70 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h46 == _T_29[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_7;
      end else if (8'h46 == _T_26[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_6;
      end else if (8'h46 == _T_23[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_5;
      end else if (8'h46 == _T_20[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_4;
      end else if (8'h46 == _T_17[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_3;
      end else if (8'h46 == _T_14[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_2;
      end else if (8'h46 == _T_11[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_1;
      end else if (8'h46 == _T_7[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_71 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h47 == _T_29[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_7;
      end else if (8'h47 == _T_26[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_6;
      end else if (8'h47 == _T_23[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_5;
      end else if (8'h47 == _T_20[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_4;
      end else if (8'h47 == _T_17[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_3;
      end else if (8'h47 == _T_14[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_2;
      end else if (8'h47 == _T_11[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_1;
      end else if (8'h47 == _T_7[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_72 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h48 == _T_29[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_7;
      end else if (8'h48 == _T_26[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_6;
      end else if (8'h48 == _T_23[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_5;
      end else if (8'h48 == _T_20[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_4;
      end else if (8'h48 == _T_17[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_3;
      end else if (8'h48 == _T_14[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_2;
      end else if (8'h48 == _T_11[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_1;
      end else if (8'h48 == _T_7[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_73 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h49 == _T_29[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_7;
      end else if (8'h49 == _T_26[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_6;
      end else if (8'h49 == _T_23[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_5;
      end else if (8'h49 == _T_20[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_4;
      end else if (8'h49 == _T_17[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_3;
      end else if (8'h49 == _T_14[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_2;
      end else if (8'h49 == _T_11[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_1;
      end else if (8'h49 == _T_7[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_74 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4a == _T_29[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_7;
      end else if (8'h4a == _T_26[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_6;
      end else if (8'h4a == _T_23[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_5;
      end else if (8'h4a == _T_20[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_4;
      end else if (8'h4a == _T_17[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_3;
      end else if (8'h4a == _T_14[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_2;
      end else if (8'h4a == _T_11[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_1;
      end else if (8'h4a == _T_7[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_75 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4b == _T_29[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_7;
      end else if (8'h4b == _T_26[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_6;
      end else if (8'h4b == _T_23[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_5;
      end else if (8'h4b == _T_20[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_4;
      end else if (8'h4b == _T_17[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_3;
      end else if (8'h4b == _T_14[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_2;
      end else if (8'h4b == _T_11[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_1;
      end else if (8'h4b == _T_7[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_76 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4c == _T_29[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_7;
      end else if (8'h4c == _T_26[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_6;
      end else if (8'h4c == _T_23[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_5;
      end else if (8'h4c == _T_20[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_4;
      end else if (8'h4c == _T_17[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_3;
      end else if (8'h4c == _T_14[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_2;
      end else if (8'h4c == _T_11[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_1;
      end else if (8'h4c == _T_7[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_77 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4d == _T_29[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_7;
      end else if (8'h4d == _T_26[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_6;
      end else if (8'h4d == _T_23[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_5;
      end else if (8'h4d == _T_20[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_4;
      end else if (8'h4d == _T_17[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_3;
      end else if (8'h4d == _T_14[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_2;
      end else if (8'h4d == _T_11[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_1;
      end else if (8'h4d == _T_7[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_78 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4e == _T_29[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_7;
      end else if (8'h4e == _T_26[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_6;
      end else if (8'h4e == _T_23[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_5;
      end else if (8'h4e == _T_20[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_4;
      end else if (8'h4e == _T_17[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_3;
      end else if (8'h4e == _T_14[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_2;
      end else if (8'h4e == _T_11[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_1;
      end else if (8'h4e == _T_7[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_79 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4f == _T_29[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_7;
      end else if (8'h4f == _T_26[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_6;
      end else if (8'h4f == _T_23[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_5;
      end else if (8'h4f == _T_20[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_4;
      end else if (8'h4f == _T_17[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_3;
      end else if (8'h4f == _T_14[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_2;
      end else if (8'h4f == _T_11[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_1;
      end else if (8'h4f == _T_7[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_80 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h50 == _T_29[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_7;
      end else if (8'h50 == _T_26[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_6;
      end else if (8'h50 == _T_23[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_5;
      end else if (8'h50 == _T_20[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_4;
      end else if (8'h50 == _T_17[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_3;
      end else if (8'h50 == _T_14[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_2;
      end else if (8'h50 == _T_11[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_1;
      end else if (8'h50 == _T_7[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_81 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h51 == _T_29[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_7;
      end else if (8'h51 == _T_26[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_6;
      end else if (8'h51 == _T_23[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_5;
      end else if (8'h51 == _T_20[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_4;
      end else if (8'h51 == _T_17[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_3;
      end else if (8'h51 == _T_14[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_2;
      end else if (8'h51 == _T_11[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_1;
      end else if (8'h51 == _T_7[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_82 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h52 == _T_29[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_7;
      end else if (8'h52 == _T_26[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_6;
      end else if (8'h52 == _T_23[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_5;
      end else if (8'h52 == _T_20[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_4;
      end else if (8'h52 == _T_17[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_3;
      end else if (8'h52 == _T_14[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_2;
      end else if (8'h52 == _T_11[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_1;
      end else if (8'h52 == _T_7[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_83 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h53 == _T_29[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_7;
      end else if (8'h53 == _T_26[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_6;
      end else if (8'h53 == _T_23[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_5;
      end else if (8'h53 == _T_20[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_4;
      end else if (8'h53 == _T_17[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_3;
      end else if (8'h53 == _T_14[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_2;
      end else if (8'h53 == _T_11[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_1;
      end else if (8'h53 == _T_7[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_84 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h54 == _T_29[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_7;
      end else if (8'h54 == _T_26[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_6;
      end else if (8'h54 == _T_23[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_5;
      end else if (8'h54 == _T_20[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_4;
      end else if (8'h54 == _T_17[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_3;
      end else if (8'h54 == _T_14[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_2;
      end else if (8'h54 == _T_11[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_1;
      end else if (8'h54 == _T_7[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_85 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h55 == _T_29[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_7;
      end else if (8'h55 == _T_26[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_6;
      end else if (8'h55 == _T_23[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_5;
      end else if (8'h55 == _T_20[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_4;
      end else if (8'h55 == _T_17[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_3;
      end else if (8'h55 == _T_14[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_2;
      end else if (8'h55 == _T_11[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_1;
      end else if (8'h55 == _T_7[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_86 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h56 == _T_29[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_7;
      end else if (8'h56 == _T_26[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_6;
      end else if (8'h56 == _T_23[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_5;
      end else if (8'h56 == _T_20[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_4;
      end else if (8'h56 == _T_17[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_3;
      end else if (8'h56 == _T_14[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_2;
      end else if (8'h56 == _T_11[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_1;
      end else if (8'h56 == _T_7[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_87 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h57 == _T_29[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_7;
      end else if (8'h57 == _T_26[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_6;
      end else if (8'h57 == _T_23[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_5;
      end else if (8'h57 == _T_20[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_4;
      end else if (8'h57 == _T_17[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_3;
      end else if (8'h57 == _T_14[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_2;
      end else if (8'h57 == _T_11[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_1;
      end else if (8'h57 == _T_7[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_88 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h58 == _T_29[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_7;
      end else if (8'h58 == _T_26[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_6;
      end else if (8'h58 == _T_23[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_5;
      end else if (8'h58 == _T_20[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_4;
      end else if (8'h58 == _T_17[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_3;
      end else if (8'h58 == _T_14[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_2;
      end else if (8'h58 == _T_11[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_1;
      end else if (8'h58 == _T_7[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_89 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h59 == _T_29[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_7;
      end else if (8'h59 == _T_26[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_6;
      end else if (8'h59 == _T_23[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_5;
      end else if (8'h59 == _T_20[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_4;
      end else if (8'h59 == _T_17[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_3;
      end else if (8'h59 == _T_14[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_2;
      end else if (8'h59 == _T_11[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_1;
      end else if (8'h59 == _T_7[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_90 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5a == _T_29[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_7;
      end else if (8'h5a == _T_26[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_6;
      end else if (8'h5a == _T_23[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_5;
      end else if (8'h5a == _T_20[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_4;
      end else if (8'h5a == _T_17[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_3;
      end else if (8'h5a == _T_14[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_2;
      end else if (8'h5a == _T_11[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_1;
      end else if (8'h5a == _T_7[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_91 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5b == _T_29[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_7;
      end else if (8'h5b == _T_26[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_6;
      end else if (8'h5b == _T_23[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_5;
      end else if (8'h5b == _T_20[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_4;
      end else if (8'h5b == _T_17[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_3;
      end else if (8'h5b == _T_14[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_2;
      end else if (8'h5b == _T_11[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_1;
      end else if (8'h5b == _T_7[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_92 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5c == _T_29[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_7;
      end else if (8'h5c == _T_26[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_6;
      end else if (8'h5c == _T_23[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_5;
      end else if (8'h5c == _T_20[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_4;
      end else if (8'h5c == _T_17[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_3;
      end else if (8'h5c == _T_14[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_2;
      end else if (8'h5c == _T_11[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_1;
      end else if (8'h5c == _T_7[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_93 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5d == _T_29[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_7;
      end else if (8'h5d == _T_26[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_6;
      end else if (8'h5d == _T_23[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_5;
      end else if (8'h5d == _T_20[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_4;
      end else if (8'h5d == _T_17[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_3;
      end else if (8'h5d == _T_14[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_2;
      end else if (8'h5d == _T_11[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_1;
      end else if (8'h5d == _T_7[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_94 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5e == _T_29[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_7;
      end else if (8'h5e == _T_26[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_6;
      end else if (8'h5e == _T_23[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_5;
      end else if (8'h5e == _T_20[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_4;
      end else if (8'h5e == _T_17[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_3;
      end else if (8'h5e == _T_14[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_2;
      end else if (8'h5e == _T_11[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_1;
      end else if (8'h5e == _T_7[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_95 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5f == _T_29[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_7;
      end else if (8'h5f == _T_26[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_6;
      end else if (8'h5f == _T_23[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_5;
      end else if (8'h5f == _T_20[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_4;
      end else if (8'h5f == _T_17[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_3;
      end else if (8'h5f == _T_14[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_2;
      end else if (8'h5f == _T_11[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_1;
      end else if (8'h5f == _T_7[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_96 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h60 == _T_29[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_7;
      end else if (8'h60 == _T_26[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_6;
      end else if (8'h60 == _T_23[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_5;
      end else if (8'h60 == _T_20[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_4;
      end else if (8'h60 == _T_17[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_3;
      end else if (8'h60 == _T_14[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_2;
      end else if (8'h60 == _T_11[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_1;
      end else if (8'h60 == _T_7[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_97 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h61 == _T_29[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_7;
      end else if (8'h61 == _T_26[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_6;
      end else if (8'h61 == _T_23[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_5;
      end else if (8'h61 == _T_20[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_4;
      end else if (8'h61 == _T_17[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_3;
      end else if (8'h61 == _T_14[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_2;
      end else if (8'h61 == _T_11[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_1;
      end else if (8'h61 == _T_7[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_98 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h62 == _T_29[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_7;
      end else if (8'h62 == _T_26[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_6;
      end else if (8'h62 == _T_23[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_5;
      end else if (8'h62 == _T_20[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_4;
      end else if (8'h62 == _T_17[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_3;
      end else if (8'h62 == _T_14[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_2;
      end else if (8'h62 == _T_11[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_1;
      end else if (8'h62 == _T_7[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_99 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h63 == _T_29[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_7;
      end else if (8'h63 == _T_26[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_6;
      end else if (8'h63 == _T_23[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_5;
      end else if (8'h63 == _T_20[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_4;
      end else if (8'h63 == _T_17[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_3;
      end else if (8'h63 == _T_14[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_2;
      end else if (8'h63 == _T_11[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_1;
      end else if (8'h63 == _T_7[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_100 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h64 == _T_29[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_7;
      end else if (8'h64 == _T_26[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_6;
      end else if (8'h64 == _T_23[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_5;
      end else if (8'h64 == _T_20[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_4;
      end else if (8'h64 == _T_17[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_3;
      end else if (8'h64 == _T_14[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_2;
      end else if (8'h64 == _T_11[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_1;
      end else if (8'h64 == _T_7[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_101 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h65 == _T_29[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_7;
      end else if (8'h65 == _T_26[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_6;
      end else if (8'h65 == _T_23[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_5;
      end else if (8'h65 == _T_20[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_4;
      end else if (8'h65 == _T_17[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_3;
      end else if (8'h65 == _T_14[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_2;
      end else if (8'h65 == _T_11[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_1;
      end else if (8'h65 == _T_7[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_102 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h66 == _T_29[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_7;
      end else if (8'h66 == _T_26[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_6;
      end else if (8'h66 == _T_23[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_5;
      end else if (8'h66 == _T_20[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_4;
      end else if (8'h66 == _T_17[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_3;
      end else if (8'h66 == _T_14[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_2;
      end else if (8'h66 == _T_11[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_1;
      end else if (8'h66 == _T_7[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_103 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h67 == _T_29[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_7;
      end else if (8'h67 == _T_26[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_6;
      end else if (8'h67 == _T_23[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_5;
      end else if (8'h67 == _T_20[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_4;
      end else if (8'h67 == _T_17[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_3;
      end else if (8'h67 == _T_14[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_2;
      end else if (8'h67 == _T_11[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_1;
      end else if (8'h67 == _T_7[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_104 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h68 == _T_29[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_7;
      end else if (8'h68 == _T_26[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_6;
      end else if (8'h68 == _T_23[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_5;
      end else if (8'h68 == _T_20[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_4;
      end else if (8'h68 == _T_17[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_3;
      end else if (8'h68 == _T_14[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_2;
      end else if (8'h68 == _T_11[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_1;
      end else if (8'h68 == _T_7[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_105 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h69 == _T_29[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_7;
      end else if (8'h69 == _T_26[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_6;
      end else if (8'h69 == _T_23[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_5;
      end else if (8'h69 == _T_20[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_4;
      end else if (8'h69 == _T_17[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_3;
      end else if (8'h69 == _T_14[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_2;
      end else if (8'h69 == _T_11[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_1;
      end else if (8'h69 == _T_7[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_106 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6a == _T_29[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_7;
      end else if (8'h6a == _T_26[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_6;
      end else if (8'h6a == _T_23[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_5;
      end else if (8'h6a == _T_20[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_4;
      end else if (8'h6a == _T_17[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_3;
      end else if (8'h6a == _T_14[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_2;
      end else if (8'h6a == _T_11[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_1;
      end else if (8'h6a == _T_7[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_107 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6b == _T_29[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_7;
      end else if (8'h6b == _T_26[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_6;
      end else if (8'h6b == _T_23[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_5;
      end else if (8'h6b == _T_20[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_4;
      end else if (8'h6b == _T_17[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_3;
      end else if (8'h6b == _T_14[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_2;
      end else if (8'h6b == _T_11[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_1;
      end else if (8'h6b == _T_7[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_108 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6c == _T_29[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_7;
      end else if (8'h6c == _T_26[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_6;
      end else if (8'h6c == _T_23[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_5;
      end else if (8'h6c == _T_20[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_4;
      end else if (8'h6c == _T_17[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_3;
      end else if (8'h6c == _T_14[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_2;
      end else if (8'h6c == _T_11[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_1;
      end else if (8'h6c == _T_7[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_109 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6d == _T_29[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_7;
      end else if (8'h6d == _T_26[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_6;
      end else if (8'h6d == _T_23[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_5;
      end else if (8'h6d == _T_20[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_4;
      end else if (8'h6d == _T_17[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_3;
      end else if (8'h6d == _T_14[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_2;
      end else if (8'h6d == _T_11[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_1;
      end else if (8'h6d == _T_7[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_110 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6e == _T_29[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_7;
      end else if (8'h6e == _T_26[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_6;
      end else if (8'h6e == _T_23[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_5;
      end else if (8'h6e == _T_20[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_4;
      end else if (8'h6e == _T_17[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_3;
      end else if (8'h6e == _T_14[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_2;
      end else if (8'h6e == _T_11[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_1;
      end else if (8'h6e == _T_7[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_111 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6f == _T_29[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_7;
      end else if (8'h6f == _T_26[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_6;
      end else if (8'h6f == _T_23[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_5;
      end else if (8'h6f == _T_20[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_4;
      end else if (8'h6f == _T_17[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_3;
      end else if (8'h6f == _T_14[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_2;
      end else if (8'h6f == _T_11[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_1;
      end else if (8'h6f == _T_7[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_112 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h70 == _T_29[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_7;
      end else if (8'h70 == _T_26[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_6;
      end else if (8'h70 == _T_23[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_5;
      end else if (8'h70 == _T_20[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_4;
      end else if (8'h70 == _T_17[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_3;
      end else if (8'h70 == _T_14[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_2;
      end else if (8'h70 == _T_11[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_1;
      end else if (8'h70 == _T_7[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_113 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h71 == _T_29[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_7;
      end else if (8'h71 == _T_26[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_6;
      end else if (8'h71 == _T_23[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_5;
      end else if (8'h71 == _T_20[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_4;
      end else if (8'h71 == _T_17[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_3;
      end else if (8'h71 == _T_14[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_2;
      end else if (8'h71 == _T_11[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_1;
      end else if (8'h71 == _T_7[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_114 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h72 == _T_29[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_7;
      end else if (8'h72 == _T_26[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_6;
      end else if (8'h72 == _T_23[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_5;
      end else if (8'h72 == _T_20[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_4;
      end else if (8'h72 == _T_17[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_3;
      end else if (8'h72 == _T_14[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_2;
      end else if (8'h72 == _T_11[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_1;
      end else if (8'h72 == _T_7[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_115 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h73 == _T_29[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_7;
      end else if (8'h73 == _T_26[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_6;
      end else if (8'h73 == _T_23[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_5;
      end else if (8'h73 == _T_20[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_4;
      end else if (8'h73 == _T_17[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_3;
      end else if (8'h73 == _T_14[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_2;
      end else if (8'h73 == _T_11[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_1;
      end else if (8'h73 == _T_7[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_116 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h74 == _T_29[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_7;
      end else if (8'h74 == _T_26[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_6;
      end else if (8'h74 == _T_23[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_5;
      end else if (8'h74 == _T_20[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_4;
      end else if (8'h74 == _T_17[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_3;
      end else if (8'h74 == _T_14[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_2;
      end else if (8'h74 == _T_11[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_1;
      end else if (8'h74 == _T_7[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_117 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h75 == _T_29[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_7;
      end else if (8'h75 == _T_26[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_6;
      end else if (8'h75 == _T_23[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_5;
      end else if (8'h75 == _T_20[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_4;
      end else if (8'h75 == _T_17[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_3;
      end else if (8'h75 == _T_14[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_2;
      end else if (8'h75 == _T_11[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_1;
      end else if (8'h75 == _T_7[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_118 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h76 == _T_29[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_7;
      end else if (8'h76 == _T_26[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_6;
      end else if (8'h76 == _T_23[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_5;
      end else if (8'h76 == _T_20[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_4;
      end else if (8'h76 == _T_17[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_3;
      end else if (8'h76 == _T_14[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_2;
      end else if (8'h76 == _T_11[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_1;
      end else if (8'h76 == _T_7[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_119 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h77 == _T_29[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_7;
      end else if (8'h77 == _T_26[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_6;
      end else if (8'h77 == _T_23[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_5;
      end else if (8'h77 == _T_20[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_4;
      end else if (8'h77 == _T_17[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_3;
      end else if (8'h77 == _T_14[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_2;
      end else if (8'h77 == _T_11[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_1;
      end else if (8'h77 == _T_7[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_120 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h78 == _T_29[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_7;
      end else if (8'h78 == _T_26[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_6;
      end else if (8'h78 == _T_23[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_5;
      end else if (8'h78 == _T_20[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_4;
      end else if (8'h78 == _T_17[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_3;
      end else if (8'h78 == _T_14[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_2;
      end else if (8'h78 == _T_11[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_1;
      end else if (8'h78 == _T_7[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_121 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h79 == _T_29[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_7;
      end else if (8'h79 == _T_26[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_6;
      end else if (8'h79 == _T_23[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_5;
      end else if (8'h79 == _T_20[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_4;
      end else if (8'h79 == _T_17[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_3;
      end else if (8'h79 == _T_14[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_2;
      end else if (8'h79 == _T_11[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_1;
      end else if (8'h79 == _T_7[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_122 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7a == _T_29[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_7;
      end else if (8'h7a == _T_26[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_6;
      end else if (8'h7a == _T_23[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_5;
      end else if (8'h7a == _T_20[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_4;
      end else if (8'h7a == _T_17[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_3;
      end else if (8'h7a == _T_14[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_2;
      end else if (8'h7a == _T_11[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_1;
      end else if (8'h7a == _T_7[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_123 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7b == _T_29[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_7;
      end else if (8'h7b == _T_26[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_6;
      end else if (8'h7b == _T_23[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_5;
      end else if (8'h7b == _T_20[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_4;
      end else if (8'h7b == _T_17[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_3;
      end else if (8'h7b == _T_14[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_2;
      end else if (8'h7b == _T_11[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_1;
      end else if (8'h7b == _T_7[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_124 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7c == _T_29[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_7;
      end else if (8'h7c == _T_26[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_6;
      end else if (8'h7c == _T_23[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_5;
      end else if (8'h7c == _T_20[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_4;
      end else if (8'h7c == _T_17[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_3;
      end else if (8'h7c == _T_14[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_2;
      end else if (8'h7c == _T_11[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_1;
      end else if (8'h7c == _T_7[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_125 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7d == _T_29[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_7;
      end else if (8'h7d == _T_26[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_6;
      end else if (8'h7d == _T_23[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_5;
      end else if (8'h7d == _T_20[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_4;
      end else if (8'h7d == _T_17[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_3;
      end else if (8'h7d == _T_14[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_2;
      end else if (8'h7d == _T_11[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_1;
      end else if (8'h7d == _T_7[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_126 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7e == _T_29[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_7;
      end else if (8'h7e == _T_26[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_6;
      end else if (8'h7e == _T_23[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_5;
      end else if (8'h7e == _T_20[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_4;
      end else if (8'h7e == _T_17[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_3;
      end else if (8'h7e == _T_14[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_2;
      end else if (8'h7e == _T_11[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_1;
      end else if (8'h7e == _T_7[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_127 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7f == _T_29[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_7;
      end else if (8'h7f == _T_26[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_6;
      end else if (8'h7f == _T_23[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_5;
      end else if (8'h7f == _T_20[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_4;
      end else if (8'h7f == _T_17[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_3;
      end else if (8'h7f == _T_14[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_2;
      end else if (8'h7f == _T_11[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_1;
      end else if (8'h7f == _T_7[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_128 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h80 == _T_29[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_7;
      end else if (8'h80 == _T_26[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_6;
      end else if (8'h80 == _T_23[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_5;
      end else if (8'h80 == _T_20[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_4;
      end else if (8'h80 == _T_17[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_3;
      end else if (8'h80 == _T_14[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_2;
      end else if (8'h80 == _T_11[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_1;
      end else if (8'h80 == _T_7[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_129 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h81 == _T_29[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_7;
      end else if (8'h81 == _T_26[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_6;
      end else if (8'h81 == _T_23[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_5;
      end else if (8'h81 == _T_20[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_4;
      end else if (8'h81 == _T_17[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_3;
      end else if (8'h81 == _T_14[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_2;
      end else if (8'h81 == _T_11[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_1;
      end else if (8'h81 == _T_7[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_130 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h82 == _T_29[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_7;
      end else if (8'h82 == _T_26[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_6;
      end else if (8'h82 == _T_23[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_5;
      end else if (8'h82 == _T_20[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_4;
      end else if (8'h82 == _T_17[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_3;
      end else if (8'h82 == _T_14[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_2;
      end else if (8'h82 == _T_11[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_1;
      end else if (8'h82 == _T_7[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_131 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h83 == _T_29[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_7;
      end else if (8'h83 == _T_26[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_6;
      end else if (8'h83 == _T_23[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_5;
      end else if (8'h83 == _T_20[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_4;
      end else if (8'h83 == _T_17[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_3;
      end else if (8'h83 == _T_14[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_2;
      end else if (8'h83 == _T_11[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_1;
      end else if (8'h83 == _T_7[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_132 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h84 == _T_29[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_7;
      end else if (8'h84 == _T_26[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_6;
      end else if (8'h84 == _T_23[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_5;
      end else if (8'h84 == _T_20[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_4;
      end else if (8'h84 == _T_17[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_3;
      end else if (8'h84 == _T_14[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_2;
      end else if (8'h84 == _T_11[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_1;
      end else if (8'h84 == _T_7[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_133 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h85 == _T_29[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_7;
      end else if (8'h85 == _T_26[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_6;
      end else if (8'h85 == _T_23[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_5;
      end else if (8'h85 == _T_20[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_4;
      end else if (8'h85 == _T_17[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_3;
      end else if (8'h85 == _T_14[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_2;
      end else if (8'h85 == _T_11[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_1;
      end else if (8'h85 == _T_7[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_134 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h86 == _T_29[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_7;
      end else if (8'h86 == _T_26[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_6;
      end else if (8'h86 == _T_23[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_5;
      end else if (8'h86 == _T_20[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_4;
      end else if (8'h86 == _T_17[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_3;
      end else if (8'h86 == _T_14[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_2;
      end else if (8'h86 == _T_11[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_1;
      end else if (8'h86 == _T_7[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_135 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h87 == _T_29[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_7;
      end else if (8'h87 == _T_26[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_6;
      end else if (8'h87 == _T_23[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_5;
      end else if (8'h87 == _T_20[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_4;
      end else if (8'h87 == _T_17[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_3;
      end else if (8'h87 == _T_14[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_2;
      end else if (8'h87 == _T_11[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_1;
      end else if (8'h87 == _T_7[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_136 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h88 == _T_29[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_7;
      end else if (8'h88 == _T_26[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_6;
      end else if (8'h88 == _T_23[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_5;
      end else if (8'h88 == _T_20[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_4;
      end else if (8'h88 == _T_17[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_3;
      end else if (8'h88 == _T_14[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_2;
      end else if (8'h88 == _T_11[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_1;
      end else if (8'h88 == _T_7[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_137 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h89 == _T_29[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_7;
      end else if (8'h89 == _T_26[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_6;
      end else if (8'h89 == _T_23[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_5;
      end else if (8'h89 == _T_20[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_4;
      end else if (8'h89 == _T_17[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_3;
      end else if (8'h89 == _T_14[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_2;
      end else if (8'h89 == _T_11[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_1;
      end else if (8'h89 == _T_7[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_138 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8a == _T_29[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_7;
      end else if (8'h8a == _T_26[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_6;
      end else if (8'h8a == _T_23[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_5;
      end else if (8'h8a == _T_20[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_4;
      end else if (8'h8a == _T_17[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_3;
      end else if (8'h8a == _T_14[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_2;
      end else if (8'h8a == _T_11[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_1;
      end else if (8'h8a == _T_7[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_139 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8b == _T_29[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_7;
      end else if (8'h8b == _T_26[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_6;
      end else if (8'h8b == _T_23[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_5;
      end else if (8'h8b == _T_20[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_4;
      end else if (8'h8b == _T_17[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_3;
      end else if (8'h8b == _T_14[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_2;
      end else if (8'h8b == _T_11[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_1;
      end else if (8'h8b == _T_7[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_140 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8c == _T_29[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_7;
      end else if (8'h8c == _T_26[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_6;
      end else if (8'h8c == _T_23[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_5;
      end else if (8'h8c == _T_20[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_4;
      end else if (8'h8c == _T_17[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_3;
      end else if (8'h8c == _T_14[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_2;
      end else if (8'h8c == _T_11[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_1;
      end else if (8'h8c == _T_7[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_141 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8d == _T_29[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_7;
      end else if (8'h8d == _T_26[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_6;
      end else if (8'h8d == _T_23[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_5;
      end else if (8'h8d == _T_20[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_4;
      end else if (8'h8d == _T_17[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_3;
      end else if (8'h8d == _T_14[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_2;
      end else if (8'h8d == _T_11[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_1;
      end else if (8'h8d == _T_7[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_142 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8e == _T_29[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_7;
      end else if (8'h8e == _T_26[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_6;
      end else if (8'h8e == _T_23[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_5;
      end else if (8'h8e == _T_20[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_4;
      end else if (8'h8e == _T_17[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_3;
      end else if (8'h8e == _T_14[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_2;
      end else if (8'h8e == _T_11[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_1;
      end else if (8'h8e == _T_7[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_143 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8f == _T_29[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_7;
      end else if (8'h8f == _T_26[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_6;
      end else if (8'h8f == _T_23[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_5;
      end else if (8'h8f == _T_20[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_4;
      end else if (8'h8f == _T_17[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_3;
      end else if (8'h8f == _T_14[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_2;
      end else if (8'h8f == _T_11[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_1;
      end else if (8'h8f == _T_7[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_144 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h90 == _T_29[7:0]) begin
        image_0_144 <= io_pixelVal_in_0_7;
      end else if (8'h90 == _T_26[7:0]) begin
        image_0_144 <= io_pixelVal_in_0_6;
      end else if (8'h90 == _T_23[7:0]) begin
        image_0_144 <= io_pixelVal_in_0_5;
      end else if (8'h90 == _T_20[7:0]) begin
        image_0_144 <= io_pixelVal_in_0_4;
      end else if (8'h90 == _T_17[7:0]) begin
        image_0_144 <= io_pixelVal_in_0_3;
      end else if (8'h90 == _T_14[7:0]) begin
        image_0_144 <= io_pixelVal_in_0_2;
      end else if (8'h90 == _T_11[7:0]) begin
        image_0_144 <= io_pixelVal_in_0_1;
      end else if (8'h90 == _T_7[7:0]) begin
        image_0_144 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_145 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h91 == _T_29[7:0]) begin
        image_0_145 <= io_pixelVal_in_0_7;
      end else if (8'h91 == _T_26[7:0]) begin
        image_0_145 <= io_pixelVal_in_0_6;
      end else if (8'h91 == _T_23[7:0]) begin
        image_0_145 <= io_pixelVal_in_0_5;
      end else if (8'h91 == _T_20[7:0]) begin
        image_0_145 <= io_pixelVal_in_0_4;
      end else if (8'h91 == _T_17[7:0]) begin
        image_0_145 <= io_pixelVal_in_0_3;
      end else if (8'h91 == _T_14[7:0]) begin
        image_0_145 <= io_pixelVal_in_0_2;
      end else if (8'h91 == _T_11[7:0]) begin
        image_0_145 <= io_pixelVal_in_0_1;
      end else if (8'h91 == _T_7[7:0]) begin
        image_0_145 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_146 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h92 == _T_29[7:0]) begin
        image_0_146 <= io_pixelVal_in_0_7;
      end else if (8'h92 == _T_26[7:0]) begin
        image_0_146 <= io_pixelVal_in_0_6;
      end else if (8'h92 == _T_23[7:0]) begin
        image_0_146 <= io_pixelVal_in_0_5;
      end else if (8'h92 == _T_20[7:0]) begin
        image_0_146 <= io_pixelVal_in_0_4;
      end else if (8'h92 == _T_17[7:0]) begin
        image_0_146 <= io_pixelVal_in_0_3;
      end else if (8'h92 == _T_14[7:0]) begin
        image_0_146 <= io_pixelVal_in_0_2;
      end else if (8'h92 == _T_11[7:0]) begin
        image_0_146 <= io_pixelVal_in_0_1;
      end else if (8'h92 == _T_7[7:0]) begin
        image_0_146 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_147 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h93 == _T_29[7:0]) begin
        image_0_147 <= io_pixelVal_in_0_7;
      end else if (8'h93 == _T_26[7:0]) begin
        image_0_147 <= io_pixelVal_in_0_6;
      end else if (8'h93 == _T_23[7:0]) begin
        image_0_147 <= io_pixelVal_in_0_5;
      end else if (8'h93 == _T_20[7:0]) begin
        image_0_147 <= io_pixelVal_in_0_4;
      end else if (8'h93 == _T_17[7:0]) begin
        image_0_147 <= io_pixelVal_in_0_3;
      end else if (8'h93 == _T_14[7:0]) begin
        image_0_147 <= io_pixelVal_in_0_2;
      end else if (8'h93 == _T_11[7:0]) begin
        image_0_147 <= io_pixelVal_in_0_1;
      end else if (8'h93 == _T_7[7:0]) begin
        image_0_147 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_148 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h94 == _T_29[7:0]) begin
        image_0_148 <= io_pixelVal_in_0_7;
      end else if (8'h94 == _T_26[7:0]) begin
        image_0_148 <= io_pixelVal_in_0_6;
      end else if (8'h94 == _T_23[7:0]) begin
        image_0_148 <= io_pixelVal_in_0_5;
      end else if (8'h94 == _T_20[7:0]) begin
        image_0_148 <= io_pixelVal_in_0_4;
      end else if (8'h94 == _T_17[7:0]) begin
        image_0_148 <= io_pixelVal_in_0_3;
      end else if (8'h94 == _T_14[7:0]) begin
        image_0_148 <= io_pixelVal_in_0_2;
      end else if (8'h94 == _T_11[7:0]) begin
        image_0_148 <= io_pixelVal_in_0_1;
      end else if (8'h94 == _T_7[7:0]) begin
        image_0_148 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_149 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h95 == _T_29[7:0]) begin
        image_0_149 <= io_pixelVal_in_0_7;
      end else if (8'h95 == _T_26[7:0]) begin
        image_0_149 <= io_pixelVal_in_0_6;
      end else if (8'h95 == _T_23[7:0]) begin
        image_0_149 <= io_pixelVal_in_0_5;
      end else if (8'h95 == _T_20[7:0]) begin
        image_0_149 <= io_pixelVal_in_0_4;
      end else if (8'h95 == _T_17[7:0]) begin
        image_0_149 <= io_pixelVal_in_0_3;
      end else if (8'h95 == _T_14[7:0]) begin
        image_0_149 <= io_pixelVal_in_0_2;
      end else if (8'h95 == _T_11[7:0]) begin
        image_0_149 <= io_pixelVal_in_0_1;
      end else if (8'h95 == _T_7[7:0]) begin
        image_0_149 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_150 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h96 == _T_29[7:0]) begin
        image_0_150 <= io_pixelVal_in_0_7;
      end else if (8'h96 == _T_26[7:0]) begin
        image_0_150 <= io_pixelVal_in_0_6;
      end else if (8'h96 == _T_23[7:0]) begin
        image_0_150 <= io_pixelVal_in_0_5;
      end else if (8'h96 == _T_20[7:0]) begin
        image_0_150 <= io_pixelVal_in_0_4;
      end else if (8'h96 == _T_17[7:0]) begin
        image_0_150 <= io_pixelVal_in_0_3;
      end else if (8'h96 == _T_14[7:0]) begin
        image_0_150 <= io_pixelVal_in_0_2;
      end else if (8'h96 == _T_11[7:0]) begin
        image_0_150 <= io_pixelVal_in_0_1;
      end else if (8'h96 == _T_7[7:0]) begin
        image_0_150 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_151 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h97 == _T_29[7:0]) begin
        image_0_151 <= io_pixelVal_in_0_7;
      end else if (8'h97 == _T_26[7:0]) begin
        image_0_151 <= io_pixelVal_in_0_6;
      end else if (8'h97 == _T_23[7:0]) begin
        image_0_151 <= io_pixelVal_in_0_5;
      end else if (8'h97 == _T_20[7:0]) begin
        image_0_151 <= io_pixelVal_in_0_4;
      end else if (8'h97 == _T_17[7:0]) begin
        image_0_151 <= io_pixelVal_in_0_3;
      end else if (8'h97 == _T_14[7:0]) begin
        image_0_151 <= io_pixelVal_in_0_2;
      end else if (8'h97 == _T_11[7:0]) begin
        image_0_151 <= io_pixelVal_in_0_1;
      end else if (8'h97 == _T_7[7:0]) begin
        image_0_151 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_152 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h98 == _T_29[7:0]) begin
        image_0_152 <= io_pixelVal_in_0_7;
      end else if (8'h98 == _T_26[7:0]) begin
        image_0_152 <= io_pixelVal_in_0_6;
      end else if (8'h98 == _T_23[7:0]) begin
        image_0_152 <= io_pixelVal_in_0_5;
      end else if (8'h98 == _T_20[7:0]) begin
        image_0_152 <= io_pixelVal_in_0_4;
      end else if (8'h98 == _T_17[7:0]) begin
        image_0_152 <= io_pixelVal_in_0_3;
      end else if (8'h98 == _T_14[7:0]) begin
        image_0_152 <= io_pixelVal_in_0_2;
      end else if (8'h98 == _T_11[7:0]) begin
        image_0_152 <= io_pixelVal_in_0_1;
      end else if (8'h98 == _T_7[7:0]) begin
        image_0_152 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_153 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h99 == _T_29[7:0]) begin
        image_0_153 <= io_pixelVal_in_0_7;
      end else if (8'h99 == _T_26[7:0]) begin
        image_0_153 <= io_pixelVal_in_0_6;
      end else if (8'h99 == _T_23[7:0]) begin
        image_0_153 <= io_pixelVal_in_0_5;
      end else if (8'h99 == _T_20[7:0]) begin
        image_0_153 <= io_pixelVal_in_0_4;
      end else if (8'h99 == _T_17[7:0]) begin
        image_0_153 <= io_pixelVal_in_0_3;
      end else if (8'h99 == _T_14[7:0]) begin
        image_0_153 <= io_pixelVal_in_0_2;
      end else if (8'h99 == _T_11[7:0]) begin
        image_0_153 <= io_pixelVal_in_0_1;
      end else if (8'h99 == _T_7[7:0]) begin
        image_0_153 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_154 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h9a == _T_29[7:0]) begin
        image_0_154 <= io_pixelVal_in_0_7;
      end else if (8'h9a == _T_26[7:0]) begin
        image_0_154 <= io_pixelVal_in_0_6;
      end else if (8'h9a == _T_23[7:0]) begin
        image_0_154 <= io_pixelVal_in_0_5;
      end else if (8'h9a == _T_20[7:0]) begin
        image_0_154 <= io_pixelVal_in_0_4;
      end else if (8'h9a == _T_17[7:0]) begin
        image_0_154 <= io_pixelVal_in_0_3;
      end else if (8'h9a == _T_14[7:0]) begin
        image_0_154 <= io_pixelVal_in_0_2;
      end else if (8'h9a == _T_11[7:0]) begin
        image_0_154 <= io_pixelVal_in_0_1;
      end else if (8'h9a == _T_7[7:0]) begin
        image_0_154 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_155 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h9b == _T_29[7:0]) begin
        image_0_155 <= io_pixelVal_in_0_7;
      end else if (8'h9b == _T_26[7:0]) begin
        image_0_155 <= io_pixelVal_in_0_6;
      end else if (8'h9b == _T_23[7:0]) begin
        image_0_155 <= io_pixelVal_in_0_5;
      end else if (8'h9b == _T_20[7:0]) begin
        image_0_155 <= io_pixelVal_in_0_4;
      end else if (8'h9b == _T_17[7:0]) begin
        image_0_155 <= io_pixelVal_in_0_3;
      end else if (8'h9b == _T_14[7:0]) begin
        image_0_155 <= io_pixelVal_in_0_2;
      end else if (8'h9b == _T_11[7:0]) begin
        image_0_155 <= io_pixelVal_in_0_1;
      end else if (8'h9b == _T_7[7:0]) begin
        image_0_155 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_156 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h9c == _T_29[7:0]) begin
        image_0_156 <= io_pixelVal_in_0_7;
      end else if (8'h9c == _T_26[7:0]) begin
        image_0_156 <= io_pixelVal_in_0_6;
      end else if (8'h9c == _T_23[7:0]) begin
        image_0_156 <= io_pixelVal_in_0_5;
      end else if (8'h9c == _T_20[7:0]) begin
        image_0_156 <= io_pixelVal_in_0_4;
      end else if (8'h9c == _T_17[7:0]) begin
        image_0_156 <= io_pixelVal_in_0_3;
      end else if (8'h9c == _T_14[7:0]) begin
        image_0_156 <= io_pixelVal_in_0_2;
      end else if (8'h9c == _T_11[7:0]) begin
        image_0_156 <= io_pixelVal_in_0_1;
      end else if (8'h9c == _T_7[7:0]) begin
        image_0_156 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_157 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h9d == _T_29[7:0]) begin
        image_0_157 <= io_pixelVal_in_0_7;
      end else if (8'h9d == _T_26[7:0]) begin
        image_0_157 <= io_pixelVal_in_0_6;
      end else if (8'h9d == _T_23[7:0]) begin
        image_0_157 <= io_pixelVal_in_0_5;
      end else if (8'h9d == _T_20[7:0]) begin
        image_0_157 <= io_pixelVal_in_0_4;
      end else if (8'h9d == _T_17[7:0]) begin
        image_0_157 <= io_pixelVal_in_0_3;
      end else if (8'h9d == _T_14[7:0]) begin
        image_0_157 <= io_pixelVal_in_0_2;
      end else if (8'h9d == _T_11[7:0]) begin
        image_0_157 <= io_pixelVal_in_0_1;
      end else if (8'h9d == _T_7[7:0]) begin
        image_0_157 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_158 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h9e == _T_29[7:0]) begin
        image_0_158 <= io_pixelVal_in_0_7;
      end else if (8'h9e == _T_26[7:0]) begin
        image_0_158 <= io_pixelVal_in_0_6;
      end else if (8'h9e == _T_23[7:0]) begin
        image_0_158 <= io_pixelVal_in_0_5;
      end else if (8'h9e == _T_20[7:0]) begin
        image_0_158 <= io_pixelVal_in_0_4;
      end else if (8'h9e == _T_17[7:0]) begin
        image_0_158 <= io_pixelVal_in_0_3;
      end else if (8'h9e == _T_14[7:0]) begin
        image_0_158 <= io_pixelVal_in_0_2;
      end else if (8'h9e == _T_11[7:0]) begin
        image_0_158 <= io_pixelVal_in_0_1;
      end else if (8'h9e == _T_7[7:0]) begin
        image_0_158 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_159 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h9f == _T_29[7:0]) begin
        image_0_159 <= io_pixelVal_in_0_7;
      end else if (8'h9f == _T_26[7:0]) begin
        image_0_159 <= io_pixelVal_in_0_6;
      end else if (8'h9f == _T_23[7:0]) begin
        image_0_159 <= io_pixelVal_in_0_5;
      end else if (8'h9f == _T_20[7:0]) begin
        image_0_159 <= io_pixelVal_in_0_4;
      end else if (8'h9f == _T_17[7:0]) begin
        image_0_159 <= io_pixelVal_in_0_3;
      end else if (8'h9f == _T_14[7:0]) begin
        image_0_159 <= io_pixelVal_in_0_2;
      end else if (8'h9f == _T_11[7:0]) begin
        image_0_159 <= io_pixelVal_in_0_1;
      end else if (8'h9f == _T_7[7:0]) begin
        image_0_159 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_160 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha0 == _T_29[7:0]) begin
        image_0_160 <= io_pixelVal_in_0_7;
      end else if (8'ha0 == _T_26[7:0]) begin
        image_0_160 <= io_pixelVal_in_0_6;
      end else if (8'ha0 == _T_23[7:0]) begin
        image_0_160 <= io_pixelVal_in_0_5;
      end else if (8'ha0 == _T_20[7:0]) begin
        image_0_160 <= io_pixelVal_in_0_4;
      end else if (8'ha0 == _T_17[7:0]) begin
        image_0_160 <= io_pixelVal_in_0_3;
      end else if (8'ha0 == _T_14[7:0]) begin
        image_0_160 <= io_pixelVal_in_0_2;
      end else if (8'ha0 == _T_11[7:0]) begin
        image_0_160 <= io_pixelVal_in_0_1;
      end else if (8'ha0 == _T_7[7:0]) begin
        image_0_160 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_161 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha1 == _T_29[7:0]) begin
        image_0_161 <= io_pixelVal_in_0_7;
      end else if (8'ha1 == _T_26[7:0]) begin
        image_0_161 <= io_pixelVal_in_0_6;
      end else if (8'ha1 == _T_23[7:0]) begin
        image_0_161 <= io_pixelVal_in_0_5;
      end else if (8'ha1 == _T_20[7:0]) begin
        image_0_161 <= io_pixelVal_in_0_4;
      end else if (8'ha1 == _T_17[7:0]) begin
        image_0_161 <= io_pixelVal_in_0_3;
      end else if (8'ha1 == _T_14[7:0]) begin
        image_0_161 <= io_pixelVal_in_0_2;
      end else if (8'ha1 == _T_11[7:0]) begin
        image_0_161 <= io_pixelVal_in_0_1;
      end else if (8'ha1 == _T_7[7:0]) begin
        image_0_161 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_162 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha2 == _T_29[7:0]) begin
        image_0_162 <= io_pixelVal_in_0_7;
      end else if (8'ha2 == _T_26[7:0]) begin
        image_0_162 <= io_pixelVal_in_0_6;
      end else if (8'ha2 == _T_23[7:0]) begin
        image_0_162 <= io_pixelVal_in_0_5;
      end else if (8'ha2 == _T_20[7:0]) begin
        image_0_162 <= io_pixelVal_in_0_4;
      end else if (8'ha2 == _T_17[7:0]) begin
        image_0_162 <= io_pixelVal_in_0_3;
      end else if (8'ha2 == _T_14[7:0]) begin
        image_0_162 <= io_pixelVal_in_0_2;
      end else if (8'ha2 == _T_11[7:0]) begin
        image_0_162 <= io_pixelVal_in_0_1;
      end else if (8'ha2 == _T_7[7:0]) begin
        image_0_162 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_163 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha3 == _T_29[7:0]) begin
        image_0_163 <= io_pixelVal_in_0_7;
      end else if (8'ha3 == _T_26[7:0]) begin
        image_0_163 <= io_pixelVal_in_0_6;
      end else if (8'ha3 == _T_23[7:0]) begin
        image_0_163 <= io_pixelVal_in_0_5;
      end else if (8'ha3 == _T_20[7:0]) begin
        image_0_163 <= io_pixelVal_in_0_4;
      end else if (8'ha3 == _T_17[7:0]) begin
        image_0_163 <= io_pixelVal_in_0_3;
      end else if (8'ha3 == _T_14[7:0]) begin
        image_0_163 <= io_pixelVal_in_0_2;
      end else if (8'ha3 == _T_11[7:0]) begin
        image_0_163 <= io_pixelVal_in_0_1;
      end else if (8'ha3 == _T_7[7:0]) begin
        image_0_163 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_164 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha4 == _T_29[7:0]) begin
        image_0_164 <= io_pixelVal_in_0_7;
      end else if (8'ha4 == _T_26[7:0]) begin
        image_0_164 <= io_pixelVal_in_0_6;
      end else if (8'ha4 == _T_23[7:0]) begin
        image_0_164 <= io_pixelVal_in_0_5;
      end else if (8'ha4 == _T_20[7:0]) begin
        image_0_164 <= io_pixelVal_in_0_4;
      end else if (8'ha4 == _T_17[7:0]) begin
        image_0_164 <= io_pixelVal_in_0_3;
      end else if (8'ha4 == _T_14[7:0]) begin
        image_0_164 <= io_pixelVal_in_0_2;
      end else if (8'ha4 == _T_11[7:0]) begin
        image_0_164 <= io_pixelVal_in_0_1;
      end else if (8'ha4 == _T_7[7:0]) begin
        image_0_164 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_165 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha5 == _T_29[7:0]) begin
        image_0_165 <= io_pixelVal_in_0_7;
      end else if (8'ha5 == _T_26[7:0]) begin
        image_0_165 <= io_pixelVal_in_0_6;
      end else if (8'ha5 == _T_23[7:0]) begin
        image_0_165 <= io_pixelVal_in_0_5;
      end else if (8'ha5 == _T_20[7:0]) begin
        image_0_165 <= io_pixelVal_in_0_4;
      end else if (8'ha5 == _T_17[7:0]) begin
        image_0_165 <= io_pixelVal_in_0_3;
      end else if (8'ha5 == _T_14[7:0]) begin
        image_0_165 <= io_pixelVal_in_0_2;
      end else if (8'ha5 == _T_11[7:0]) begin
        image_0_165 <= io_pixelVal_in_0_1;
      end else if (8'ha5 == _T_7[7:0]) begin
        image_0_165 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_166 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha6 == _T_29[7:0]) begin
        image_0_166 <= io_pixelVal_in_0_7;
      end else if (8'ha6 == _T_26[7:0]) begin
        image_0_166 <= io_pixelVal_in_0_6;
      end else if (8'ha6 == _T_23[7:0]) begin
        image_0_166 <= io_pixelVal_in_0_5;
      end else if (8'ha6 == _T_20[7:0]) begin
        image_0_166 <= io_pixelVal_in_0_4;
      end else if (8'ha6 == _T_17[7:0]) begin
        image_0_166 <= io_pixelVal_in_0_3;
      end else if (8'ha6 == _T_14[7:0]) begin
        image_0_166 <= io_pixelVal_in_0_2;
      end else if (8'ha6 == _T_11[7:0]) begin
        image_0_166 <= io_pixelVal_in_0_1;
      end else if (8'ha6 == _T_7[7:0]) begin
        image_0_166 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_167 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha7 == _T_29[7:0]) begin
        image_0_167 <= io_pixelVal_in_0_7;
      end else if (8'ha7 == _T_26[7:0]) begin
        image_0_167 <= io_pixelVal_in_0_6;
      end else if (8'ha7 == _T_23[7:0]) begin
        image_0_167 <= io_pixelVal_in_0_5;
      end else if (8'ha7 == _T_20[7:0]) begin
        image_0_167 <= io_pixelVal_in_0_4;
      end else if (8'ha7 == _T_17[7:0]) begin
        image_0_167 <= io_pixelVal_in_0_3;
      end else if (8'ha7 == _T_14[7:0]) begin
        image_0_167 <= io_pixelVal_in_0_2;
      end else if (8'ha7 == _T_11[7:0]) begin
        image_0_167 <= io_pixelVal_in_0_1;
      end else if (8'ha7 == _T_7[7:0]) begin
        image_0_167 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_168 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha8 == _T_29[7:0]) begin
        image_0_168 <= io_pixelVal_in_0_7;
      end else if (8'ha8 == _T_26[7:0]) begin
        image_0_168 <= io_pixelVal_in_0_6;
      end else if (8'ha8 == _T_23[7:0]) begin
        image_0_168 <= io_pixelVal_in_0_5;
      end else if (8'ha8 == _T_20[7:0]) begin
        image_0_168 <= io_pixelVal_in_0_4;
      end else if (8'ha8 == _T_17[7:0]) begin
        image_0_168 <= io_pixelVal_in_0_3;
      end else if (8'ha8 == _T_14[7:0]) begin
        image_0_168 <= io_pixelVal_in_0_2;
      end else if (8'ha8 == _T_11[7:0]) begin
        image_0_168 <= io_pixelVal_in_0_1;
      end else if (8'ha8 == _T_7[7:0]) begin
        image_0_168 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_169 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha9 == _T_29[7:0]) begin
        image_0_169 <= io_pixelVal_in_0_7;
      end else if (8'ha9 == _T_26[7:0]) begin
        image_0_169 <= io_pixelVal_in_0_6;
      end else if (8'ha9 == _T_23[7:0]) begin
        image_0_169 <= io_pixelVal_in_0_5;
      end else if (8'ha9 == _T_20[7:0]) begin
        image_0_169 <= io_pixelVal_in_0_4;
      end else if (8'ha9 == _T_17[7:0]) begin
        image_0_169 <= io_pixelVal_in_0_3;
      end else if (8'ha9 == _T_14[7:0]) begin
        image_0_169 <= io_pixelVal_in_0_2;
      end else if (8'ha9 == _T_11[7:0]) begin
        image_0_169 <= io_pixelVal_in_0_1;
      end else if (8'ha9 == _T_7[7:0]) begin
        image_0_169 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_170 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'haa == _T_29[7:0]) begin
        image_0_170 <= io_pixelVal_in_0_7;
      end else if (8'haa == _T_26[7:0]) begin
        image_0_170 <= io_pixelVal_in_0_6;
      end else if (8'haa == _T_23[7:0]) begin
        image_0_170 <= io_pixelVal_in_0_5;
      end else if (8'haa == _T_20[7:0]) begin
        image_0_170 <= io_pixelVal_in_0_4;
      end else if (8'haa == _T_17[7:0]) begin
        image_0_170 <= io_pixelVal_in_0_3;
      end else if (8'haa == _T_14[7:0]) begin
        image_0_170 <= io_pixelVal_in_0_2;
      end else if (8'haa == _T_11[7:0]) begin
        image_0_170 <= io_pixelVal_in_0_1;
      end else if (8'haa == _T_7[7:0]) begin
        image_0_170 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_171 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hab == _T_29[7:0]) begin
        image_0_171 <= io_pixelVal_in_0_7;
      end else if (8'hab == _T_26[7:0]) begin
        image_0_171 <= io_pixelVal_in_0_6;
      end else if (8'hab == _T_23[7:0]) begin
        image_0_171 <= io_pixelVal_in_0_5;
      end else if (8'hab == _T_20[7:0]) begin
        image_0_171 <= io_pixelVal_in_0_4;
      end else if (8'hab == _T_17[7:0]) begin
        image_0_171 <= io_pixelVal_in_0_3;
      end else if (8'hab == _T_14[7:0]) begin
        image_0_171 <= io_pixelVal_in_0_2;
      end else if (8'hab == _T_11[7:0]) begin
        image_0_171 <= io_pixelVal_in_0_1;
      end else if (8'hab == _T_7[7:0]) begin
        image_0_171 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_172 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hac == _T_29[7:0]) begin
        image_0_172 <= io_pixelVal_in_0_7;
      end else if (8'hac == _T_26[7:0]) begin
        image_0_172 <= io_pixelVal_in_0_6;
      end else if (8'hac == _T_23[7:0]) begin
        image_0_172 <= io_pixelVal_in_0_5;
      end else if (8'hac == _T_20[7:0]) begin
        image_0_172 <= io_pixelVal_in_0_4;
      end else if (8'hac == _T_17[7:0]) begin
        image_0_172 <= io_pixelVal_in_0_3;
      end else if (8'hac == _T_14[7:0]) begin
        image_0_172 <= io_pixelVal_in_0_2;
      end else if (8'hac == _T_11[7:0]) begin
        image_0_172 <= io_pixelVal_in_0_1;
      end else if (8'hac == _T_7[7:0]) begin
        image_0_172 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_173 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'had == _T_29[7:0]) begin
        image_0_173 <= io_pixelVal_in_0_7;
      end else if (8'had == _T_26[7:0]) begin
        image_0_173 <= io_pixelVal_in_0_6;
      end else if (8'had == _T_23[7:0]) begin
        image_0_173 <= io_pixelVal_in_0_5;
      end else if (8'had == _T_20[7:0]) begin
        image_0_173 <= io_pixelVal_in_0_4;
      end else if (8'had == _T_17[7:0]) begin
        image_0_173 <= io_pixelVal_in_0_3;
      end else if (8'had == _T_14[7:0]) begin
        image_0_173 <= io_pixelVal_in_0_2;
      end else if (8'had == _T_11[7:0]) begin
        image_0_173 <= io_pixelVal_in_0_1;
      end else if (8'had == _T_7[7:0]) begin
        image_0_173 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_174 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hae == _T_29[7:0]) begin
        image_0_174 <= io_pixelVal_in_0_7;
      end else if (8'hae == _T_26[7:0]) begin
        image_0_174 <= io_pixelVal_in_0_6;
      end else if (8'hae == _T_23[7:0]) begin
        image_0_174 <= io_pixelVal_in_0_5;
      end else if (8'hae == _T_20[7:0]) begin
        image_0_174 <= io_pixelVal_in_0_4;
      end else if (8'hae == _T_17[7:0]) begin
        image_0_174 <= io_pixelVal_in_0_3;
      end else if (8'hae == _T_14[7:0]) begin
        image_0_174 <= io_pixelVal_in_0_2;
      end else if (8'hae == _T_11[7:0]) begin
        image_0_174 <= io_pixelVal_in_0_1;
      end else if (8'hae == _T_7[7:0]) begin
        image_0_174 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_175 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'haf == _T_29[7:0]) begin
        image_0_175 <= io_pixelVal_in_0_7;
      end else if (8'haf == _T_26[7:0]) begin
        image_0_175 <= io_pixelVal_in_0_6;
      end else if (8'haf == _T_23[7:0]) begin
        image_0_175 <= io_pixelVal_in_0_5;
      end else if (8'haf == _T_20[7:0]) begin
        image_0_175 <= io_pixelVal_in_0_4;
      end else if (8'haf == _T_17[7:0]) begin
        image_0_175 <= io_pixelVal_in_0_3;
      end else if (8'haf == _T_14[7:0]) begin
        image_0_175 <= io_pixelVal_in_0_2;
      end else if (8'haf == _T_11[7:0]) begin
        image_0_175 <= io_pixelVal_in_0_1;
      end else if (8'haf == _T_7[7:0]) begin
        image_0_175 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_176 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb0 == _T_29[7:0]) begin
        image_0_176 <= io_pixelVal_in_0_7;
      end else if (8'hb0 == _T_26[7:0]) begin
        image_0_176 <= io_pixelVal_in_0_6;
      end else if (8'hb0 == _T_23[7:0]) begin
        image_0_176 <= io_pixelVal_in_0_5;
      end else if (8'hb0 == _T_20[7:0]) begin
        image_0_176 <= io_pixelVal_in_0_4;
      end else if (8'hb0 == _T_17[7:0]) begin
        image_0_176 <= io_pixelVal_in_0_3;
      end else if (8'hb0 == _T_14[7:0]) begin
        image_0_176 <= io_pixelVal_in_0_2;
      end else if (8'hb0 == _T_11[7:0]) begin
        image_0_176 <= io_pixelVal_in_0_1;
      end else if (8'hb0 == _T_7[7:0]) begin
        image_0_176 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_177 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb1 == _T_29[7:0]) begin
        image_0_177 <= io_pixelVal_in_0_7;
      end else if (8'hb1 == _T_26[7:0]) begin
        image_0_177 <= io_pixelVal_in_0_6;
      end else if (8'hb1 == _T_23[7:0]) begin
        image_0_177 <= io_pixelVal_in_0_5;
      end else if (8'hb1 == _T_20[7:0]) begin
        image_0_177 <= io_pixelVal_in_0_4;
      end else if (8'hb1 == _T_17[7:0]) begin
        image_0_177 <= io_pixelVal_in_0_3;
      end else if (8'hb1 == _T_14[7:0]) begin
        image_0_177 <= io_pixelVal_in_0_2;
      end else if (8'hb1 == _T_11[7:0]) begin
        image_0_177 <= io_pixelVal_in_0_1;
      end else if (8'hb1 == _T_7[7:0]) begin
        image_0_177 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_178 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb2 == _T_29[7:0]) begin
        image_0_178 <= io_pixelVal_in_0_7;
      end else if (8'hb2 == _T_26[7:0]) begin
        image_0_178 <= io_pixelVal_in_0_6;
      end else if (8'hb2 == _T_23[7:0]) begin
        image_0_178 <= io_pixelVal_in_0_5;
      end else if (8'hb2 == _T_20[7:0]) begin
        image_0_178 <= io_pixelVal_in_0_4;
      end else if (8'hb2 == _T_17[7:0]) begin
        image_0_178 <= io_pixelVal_in_0_3;
      end else if (8'hb2 == _T_14[7:0]) begin
        image_0_178 <= io_pixelVal_in_0_2;
      end else if (8'hb2 == _T_11[7:0]) begin
        image_0_178 <= io_pixelVal_in_0_1;
      end else if (8'hb2 == _T_7[7:0]) begin
        image_0_178 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_179 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb3 == _T_29[7:0]) begin
        image_0_179 <= io_pixelVal_in_0_7;
      end else if (8'hb3 == _T_26[7:0]) begin
        image_0_179 <= io_pixelVal_in_0_6;
      end else if (8'hb3 == _T_23[7:0]) begin
        image_0_179 <= io_pixelVal_in_0_5;
      end else if (8'hb3 == _T_20[7:0]) begin
        image_0_179 <= io_pixelVal_in_0_4;
      end else if (8'hb3 == _T_17[7:0]) begin
        image_0_179 <= io_pixelVal_in_0_3;
      end else if (8'hb3 == _T_14[7:0]) begin
        image_0_179 <= io_pixelVal_in_0_2;
      end else if (8'hb3 == _T_11[7:0]) begin
        image_0_179 <= io_pixelVal_in_0_1;
      end else if (8'hb3 == _T_7[7:0]) begin
        image_0_179 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_180 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb4 == _T_29[7:0]) begin
        image_0_180 <= io_pixelVal_in_0_7;
      end else if (8'hb4 == _T_26[7:0]) begin
        image_0_180 <= io_pixelVal_in_0_6;
      end else if (8'hb4 == _T_23[7:0]) begin
        image_0_180 <= io_pixelVal_in_0_5;
      end else if (8'hb4 == _T_20[7:0]) begin
        image_0_180 <= io_pixelVal_in_0_4;
      end else if (8'hb4 == _T_17[7:0]) begin
        image_0_180 <= io_pixelVal_in_0_3;
      end else if (8'hb4 == _T_14[7:0]) begin
        image_0_180 <= io_pixelVal_in_0_2;
      end else if (8'hb4 == _T_11[7:0]) begin
        image_0_180 <= io_pixelVal_in_0_1;
      end else if (8'hb4 == _T_7[7:0]) begin
        image_0_180 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_181 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb5 == _T_29[7:0]) begin
        image_0_181 <= io_pixelVal_in_0_7;
      end else if (8'hb5 == _T_26[7:0]) begin
        image_0_181 <= io_pixelVal_in_0_6;
      end else if (8'hb5 == _T_23[7:0]) begin
        image_0_181 <= io_pixelVal_in_0_5;
      end else if (8'hb5 == _T_20[7:0]) begin
        image_0_181 <= io_pixelVal_in_0_4;
      end else if (8'hb5 == _T_17[7:0]) begin
        image_0_181 <= io_pixelVal_in_0_3;
      end else if (8'hb5 == _T_14[7:0]) begin
        image_0_181 <= io_pixelVal_in_0_2;
      end else if (8'hb5 == _T_11[7:0]) begin
        image_0_181 <= io_pixelVal_in_0_1;
      end else if (8'hb5 == _T_7[7:0]) begin
        image_0_181 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_182 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb6 == _T_29[7:0]) begin
        image_0_182 <= io_pixelVal_in_0_7;
      end else if (8'hb6 == _T_26[7:0]) begin
        image_0_182 <= io_pixelVal_in_0_6;
      end else if (8'hb6 == _T_23[7:0]) begin
        image_0_182 <= io_pixelVal_in_0_5;
      end else if (8'hb6 == _T_20[7:0]) begin
        image_0_182 <= io_pixelVal_in_0_4;
      end else if (8'hb6 == _T_17[7:0]) begin
        image_0_182 <= io_pixelVal_in_0_3;
      end else if (8'hb6 == _T_14[7:0]) begin
        image_0_182 <= io_pixelVal_in_0_2;
      end else if (8'hb6 == _T_11[7:0]) begin
        image_0_182 <= io_pixelVal_in_0_1;
      end else if (8'hb6 == _T_7[7:0]) begin
        image_0_182 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_183 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb7 == _T_29[7:0]) begin
        image_0_183 <= io_pixelVal_in_0_7;
      end else if (8'hb7 == _T_26[7:0]) begin
        image_0_183 <= io_pixelVal_in_0_6;
      end else if (8'hb7 == _T_23[7:0]) begin
        image_0_183 <= io_pixelVal_in_0_5;
      end else if (8'hb7 == _T_20[7:0]) begin
        image_0_183 <= io_pixelVal_in_0_4;
      end else if (8'hb7 == _T_17[7:0]) begin
        image_0_183 <= io_pixelVal_in_0_3;
      end else if (8'hb7 == _T_14[7:0]) begin
        image_0_183 <= io_pixelVal_in_0_2;
      end else if (8'hb7 == _T_11[7:0]) begin
        image_0_183 <= io_pixelVal_in_0_1;
      end else if (8'hb7 == _T_7[7:0]) begin
        image_0_183 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_184 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb8 == _T_29[7:0]) begin
        image_0_184 <= io_pixelVal_in_0_7;
      end else if (8'hb8 == _T_26[7:0]) begin
        image_0_184 <= io_pixelVal_in_0_6;
      end else if (8'hb8 == _T_23[7:0]) begin
        image_0_184 <= io_pixelVal_in_0_5;
      end else if (8'hb8 == _T_20[7:0]) begin
        image_0_184 <= io_pixelVal_in_0_4;
      end else if (8'hb8 == _T_17[7:0]) begin
        image_0_184 <= io_pixelVal_in_0_3;
      end else if (8'hb8 == _T_14[7:0]) begin
        image_0_184 <= io_pixelVal_in_0_2;
      end else if (8'hb8 == _T_11[7:0]) begin
        image_0_184 <= io_pixelVal_in_0_1;
      end else if (8'hb8 == _T_7[7:0]) begin
        image_0_184 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_185 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb9 == _T_29[7:0]) begin
        image_0_185 <= io_pixelVal_in_0_7;
      end else if (8'hb9 == _T_26[7:0]) begin
        image_0_185 <= io_pixelVal_in_0_6;
      end else if (8'hb9 == _T_23[7:0]) begin
        image_0_185 <= io_pixelVal_in_0_5;
      end else if (8'hb9 == _T_20[7:0]) begin
        image_0_185 <= io_pixelVal_in_0_4;
      end else if (8'hb9 == _T_17[7:0]) begin
        image_0_185 <= io_pixelVal_in_0_3;
      end else if (8'hb9 == _T_14[7:0]) begin
        image_0_185 <= io_pixelVal_in_0_2;
      end else if (8'hb9 == _T_11[7:0]) begin
        image_0_185 <= io_pixelVal_in_0_1;
      end else if (8'hb9 == _T_7[7:0]) begin
        image_0_185 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_186 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hba == _T_29[7:0]) begin
        image_0_186 <= io_pixelVal_in_0_7;
      end else if (8'hba == _T_26[7:0]) begin
        image_0_186 <= io_pixelVal_in_0_6;
      end else if (8'hba == _T_23[7:0]) begin
        image_0_186 <= io_pixelVal_in_0_5;
      end else if (8'hba == _T_20[7:0]) begin
        image_0_186 <= io_pixelVal_in_0_4;
      end else if (8'hba == _T_17[7:0]) begin
        image_0_186 <= io_pixelVal_in_0_3;
      end else if (8'hba == _T_14[7:0]) begin
        image_0_186 <= io_pixelVal_in_0_2;
      end else if (8'hba == _T_11[7:0]) begin
        image_0_186 <= io_pixelVal_in_0_1;
      end else if (8'hba == _T_7[7:0]) begin
        image_0_186 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_187 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hbb == _T_29[7:0]) begin
        image_0_187 <= io_pixelVal_in_0_7;
      end else if (8'hbb == _T_26[7:0]) begin
        image_0_187 <= io_pixelVal_in_0_6;
      end else if (8'hbb == _T_23[7:0]) begin
        image_0_187 <= io_pixelVal_in_0_5;
      end else if (8'hbb == _T_20[7:0]) begin
        image_0_187 <= io_pixelVal_in_0_4;
      end else if (8'hbb == _T_17[7:0]) begin
        image_0_187 <= io_pixelVal_in_0_3;
      end else if (8'hbb == _T_14[7:0]) begin
        image_0_187 <= io_pixelVal_in_0_2;
      end else if (8'hbb == _T_11[7:0]) begin
        image_0_187 <= io_pixelVal_in_0_1;
      end else if (8'hbb == _T_7[7:0]) begin
        image_0_187 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_188 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hbc == _T_29[7:0]) begin
        image_0_188 <= io_pixelVal_in_0_7;
      end else if (8'hbc == _T_26[7:0]) begin
        image_0_188 <= io_pixelVal_in_0_6;
      end else if (8'hbc == _T_23[7:0]) begin
        image_0_188 <= io_pixelVal_in_0_5;
      end else if (8'hbc == _T_20[7:0]) begin
        image_0_188 <= io_pixelVal_in_0_4;
      end else if (8'hbc == _T_17[7:0]) begin
        image_0_188 <= io_pixelVal_in_0_3;
      end else if (8'hbc == _T_14[7:0]) begin
        image_0_188 <= io_pixelVal_in_0_2;
      end else if (8'hbc == _T_11[7:0]) begin
        image_0_188 <= io_pixelVal_in_0_1;
      end else if (8'hbc == _T_7[7:0]) begin
        image_0_188 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_189 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hbd == _T_29[7:0]) begin
        image_0_189 <= io_pixelVal_in_0_7;
      end else if (8'hbd == _T_26[7:0]) begin
        image_0_189 <= io_pixelVal_in_0_6;
      end else if (8'hbd == _T_23[7:0]) begin
        image_0_189 <= io_pixelVal_in_0_5;
      end else if (8'hbd == _T_20[7:0]) begin
        image_0_189 <= io_pixelVal_in_0_4;
      end else if (8'hbd == _T_17[7:0]) begin
        image_0_189 <= io_pixelVal_in_0_3;
      end else if (8'hbd == _T_14[7:0]) begin
        image_0_189 <= io_pixelVal_in_0_2;
      end else if (8'hbd == _T_11[7:0]) begin
        image_0_189 <= io_pixelVal_in_0_1;
      end else if (8'hbd == _T_7[7:0]) begin
        image_0_189 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_190 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hbe == _T_29[7:0]) begin
        image_0_190 <= io_pixelVal_in_0_7;
      end else if (8'hbe == _T_26[7:0]) begin
        image_0_190 <= io_pixelVal_in_0_6;
      end else if (8'hbe == _T_23[7:0]) begin
        image_0_190 <= io_pixelVal_in_0_5;
      end else if (8'hbe == _T_20[7:0]) begin
        image_0_190 <= io_pixelVal_in_0_4;
      end else if (8'hbe == _T_17[7:0]) begin
        image_0_190 <= io_pixelVal_in_0_3;
      end else if (8'hbe == _T_14[7:0]) begin
        image_0_190 <= io_pixelVal_in_0_2;
      end else if (8'hbe == _T_11[7:0]) begin
        image_0_190 <= io_pixelVal_in_0_1;
      end else if (8'hbe == _T_7[7:0]) begin
        image_0_190 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_191 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hbf == _T_29[7:0]) begin
        image_0_191 <= io_pixelVal_in_0_7;
      end else if (8'hbf == _T_26[7:0]) begin
        image_0_191 <= io_pixelVal_in_0_6;
      end else if (8'hbf == _T_23[7:0]) begin
        image_0_191 <= io_pixelVal_in_0_5;
      end else if (8'hbf == _T_20[7:0]) begin
        image_0_191 <= io_pixelVal_in_0_4;
      end else if (8'hbf == _T_17[7:0]) begin
        image_0_191 <= io_pixelVal_in_0_3;
      end else if (8'hbf == _T_14[7:0]) begin
        image_0_191 <= io_pixelVal_in_0_2;
      end else if (8'hbf == _T_11[7:0]) begin
        image_0_191 <= io_pixelVal_in_0_1;
      end else if (8'hbf == _T_7[7:0]) begin
        image_0_191 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_1_0 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h0 == _T_29[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_7;
      end else if (8'h0 == _T_26[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_6;
      end else if (8'h0 == _T_23[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_5;
      end else if (8'h0 == _T_20[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_4;
      end else if (8'h0 == _T_17[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_3;
      end else if (8'h0 == _T_14[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_2;
      end else if (8'h0 == _T_11[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_1;
      end else if (8'h0 == _T_7[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_1 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1 == _T_29[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_7;
      end else if (8'h1 == _T_26[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_6;
      end else if (8'h1 == _T_23[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_5;
      end else if (8'h1 == _T_20[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_4;
      end else if (8'h1 == _T_17[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_3;
      end else if (8'h1 == _T_14[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_2;
      end else if (8'h1 == _T_11[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_1;
      end else if (8'h1 == _T_7[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_2 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2 == _T_29[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_7;
      end else if (8'h2 == _T_26[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_6;
      end else if (8'h2 == _T_23[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_5;
      end else if (8'h2 == _T_20[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_4;
      end else if (8'h2 == _T_17[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_3;
      end else if (8'h2 == _T_14[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_2;
      end else if (8'h2 == _T_11[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_1;
      end else if (8'h2 == _T_7[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_3 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3 == _T_29[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_7;
      end else if (8'h3 == _T_26[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_6;
      end else if (8'h3 == _T_23[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_5;
      end else if (8'h3 == _T_20[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_4;
      end else if (8'h3 == _T_17[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_3;
      end else if (8'h3 == _T_14[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_2;
      end else if (8'h3 == _T_11[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_1;
      end else if (8'h3 == _T_7[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_4 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4 == _T_29[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_7;
      end else if (8'h4 == _T_26[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_6;
      end else if (8'h4 == _T_23[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_5;
      end else if (8'h4 == _T_20[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_4;
      end else if (8'h4 == _T_17[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_3;
      end else if (8'h4 == _T_14[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_2;
      end else if (8'h4 == _T_11[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_1;
      end else if (8'h4 == _T_7[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_5 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5 == _T_29[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_7;
      end else if (8'h5 == _T_26[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_6;
      end else if (8'h5 == _T_23[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_5;
      end else if (8'h5 == _T_20[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_4;
      end else if (8'h5 == _T_17[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_3;
      end else if (8'h5 == _T_14[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_2;
      end else if (8'h5 == _T_11[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_1;
      end else if (8'h5 == _T_7[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_6 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6 == _T_29[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_7;
      end else if (8'h6 == _T_26[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_6;
      end else if (8'h6 == _T_23[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_5;
      end else if (8'h6 == _T_20[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_4;
      end else if (8'h6 == _T_17[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_3;
      end else if (8'h6 == _T_14[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_2;
      end else if (8'h6 == _T_11[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_1;
      end else if (8'h6 == _T_7[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_7 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7 == _T_29[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_7;
      end else if (8'h7 == _T_26[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_6;
      end else if (8'h7 == _T_23[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_5;
      end else if (8'h7 == _T_20[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_4;
      end else if (8'h7 == _T_17[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_3;
      end else if (8'h7 == _T_14[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_2;
      end else if (8'h7 == _T_11[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_1;
      end else if (8'h7 == _T_7[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_8 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8 == _T_29[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_7;
      end else if (8'h8 == _T_26[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_6;
      end else if (8'h8 == _T_23[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_5;
      end else if (8'h8 == _T_20[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_4;
      end else if (8'h8 == _T_17[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_3;
      end else if (8'h8 == _T_14[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_2;
      end else if (8'h8 == _T_11[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_1;
      end else if (8'h8 == _T_7[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_9 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9 == _T_29[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_7;
      end else if (8'h9 == _T_26[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_6;
      end else if (8'h9 == _T_23[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_5;
      end else if (8'h9 == _T_20[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_4;
      end else if (8'h9 == _T_17[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_3;
      end else if (8'h9 == _T_14[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_2;
      end else if (8'h9 == _T_11[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_1;
      end else if (8'h9 == _T_7[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_10 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha == _T_29[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_7;
      end else if (8'ha == _T_26[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_6;
      end else if (8'ha == _T_23[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_5;
      end else if (8'ha == _T_20[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_4;
      end else if (8'ha == _T_17[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_3;
      end else if (8'ha == _T_14[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_2;
      end else if (8'ha == _T_11[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_1;
      end else if (8'ha == _T_7[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_11 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb == _T_29[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_7;
      end else if (8'hb == _T_26[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_6;
      end else if (8'hb == _T_23[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_5;
      end else if (8'hb == _T_20[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_4;
      end else if (8'hb == _T_17[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_3;
      end else if (8'hb == _T_14[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_2;
      end else if (8'hb == _T_11[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_1;
      end else if (8'hb == _T_7[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_12 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc == _T_29[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_7;
      end else if (8'hc == _T_26[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_6;
      end else if (8'hc == _T_23[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_5;
      end else if (8'hc == _T_20[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_4;
      end else if (8'hc == _T_17[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_3;
      end else if (8'hc == _T_14[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_2;
      end else if (8'hc == _T_11[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_1;
      end else if (8'hc == _T_7[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_13 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd == _T_29[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_7;
      end else if (8'hd == _T_26[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_6;
      end else if (8'hd == _T_23[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_5;
      end else if (8'hd == _T_20[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_4;
      end else if (8'hd == _T_17[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_3;
      end else if (8'hd == _T_14[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_2;
      end else if (8'hd == _T_11[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_1;
      end else if (8'hd == _T_7[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_14 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he == _T_29[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_7;
      end else if (8'he == _T_26[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_6;
      end else if (8'he == _T_23[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_5;
      end else if (8'he == _T_20[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_4;
      end else if (8'he == _T_17[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_3;
      end else if (8'he == _T_14[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_2;
      end else if (8'he == _T_11[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_1;
      end else if (8'he == _T_7[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_15 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf == _T_29[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_7;
      end else if (8'hf == _T_26[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_6;
      end else if (8'hf == _T_23[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_5;
      end else if (8'hf == _T_20[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_4;
      end else if (8'hf == _T_17[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_3;
      end else if (8'hf == _T_14[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_2;
      end else if (8'hf == _T_11[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_1;
      end else if (8'hf == _T_7[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_16 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h10 == _T_29[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_7;
      end else if (8'h10 == _T_26[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_6;
      end else if (8'h10 == _T_23[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_5;
      end else if (8'h10 == _T_20[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_4;
      end else if (8'h10 == _T_17[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_3;
      end else if (8'h10 == _T_14[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_2;
      end else if (8'h10 == _T_11[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_1;
      end else if (8'h10 == _T_7[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_17 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h11 == _T_29[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_7;
      end else if (8'h11 == _T_26[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_6;
      end else if (8'h11 == _T_23[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_5;
      end else if (8'h11 == _T_20[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_4;
      end else if (8'h11 == _T_17[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_3;
      end else if (8'h11 == _T_14[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_2;
      end else if (8'h11 == _T_11[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_1;
      end else if (8'h11 == _T_7[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_18 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h12 == _T_29[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_7;
      end else if (8'h12 == _T_26[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_6;
      end else if (8'h12 == _T_23[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_5;
      end else if (8'h12 == _T_20[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_4;
      end else if (8'h12 == _T_17[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_3;
      end else if (8'h12 == _T_14[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_2;
      end else if (8'h12 == _T_11[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_1;
      end else if (8'h12 == _T_7[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_19 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h13 == _T_29[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_7;
      end else if (8'h13 == _T_26[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_6;
      end else if (8'h13 == _T_23[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_5;
      end else if (8'h13 == _T_20[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_4;
      end else if (8'h13 == _T_17[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_3;
      end else if (8'h13 == _T_14[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_2;
      end else if (8'h13 == _T_11[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_1;
      end else if (8'h13 == _T_7[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_20 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h14 == _T_29[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_7;
      end else if (8'h14 == _T_26[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_6;
      end else if (8'h14 == _T_23[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_5;
      end else if (8'h14 == _T_20[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_4;
      end else if (8'h14 == _T_17[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_3;
      end else if (8'h14 == _T_14[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_2;
      end else if (8'h14 == _T_11[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_1;
      end else if (8'h14 == _T_7[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_21 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h15 == _T_29[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_7;
      end else if (8'h15 == _T_26[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_6;
      end else if (8'h15 == _T_23[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_5;
      end else if (8'h15 == _T_20[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_4;
      end else if (8'h15 == _T_17[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_3;
      end else if (8'h15 == _T_14[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_2;
      end else if (8'h15 == _T_11[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_1;
      end else if (8'h15 == _T_7[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_22 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h16 == _T_29[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_7;
      end else if (8'h16 == _T_26[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_6;
      end else if (8'h16 == _T_23[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_5;
      end else if (8'h16 == _T_20[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_4;
      end else if (8'h16 == _T_17[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_3;
      end else if (8'h16 == _T_14[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_2;
      end else if (8'h16 == _T_11[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_1;
      end else if (8'h16 == _T_7[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_23 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h17 == _T_29[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_7;
      end else if (8'h17 == _T_26[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_6;
      end else if (8'h17 == _T_23[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_5;
      end else if (8'h17 == _T_20[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_4;
      end else if (8'h17 == _T_17[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_3;
      end else if (8'h17 == _T_14[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_2;
      end else if (8'h17 == _T_11[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_1;
      end else if (8'h17 == _T_7[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_24 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h18 == _T_29[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_7;
      end else if (8'h18 == _T_26[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_6;
      end else if (8'h18 == _T_23[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_5;
      end else if (8'h18 == _T_20[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_4;
      end else if (8'h18 == _T_17[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_3;
      end else if (8'h18 == _T_14[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_2;
      end else if (8'h18 == _T_11[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_1;
      end else if (8'h18 == _T_7[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_25 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h19 == _T_29[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_7;
      end else if (8'h19 == _T_26[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_6;
      end else if (8'h19 == _T_23[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_5;
      end else if (8'h19 == _T_20[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_4;
      end else if (8'h19 == _T_17[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_3;
      end else if (8'h19 == _T_14[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_2;
      end else if (8'h19 == _T_11[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_1;
      end else if (8'h19 == _T_7[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_26 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1a == _T_29[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_7;
      end else if (8'h1a == _T_26[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_6;
      end else if (8'h1a == _T_23[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_5;
      end else if (8'h1a == _T_20[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_4;
      end else if (8'h1a == _T_17[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_3;
      end else if (8'h1a == _T_14[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_2;
      end else if (8'h1a == _T_11[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_1;
      end else if (8'h1a == _T_7[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_27 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1b == _T_29[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_7;
      end else if (8'h1b == _T_26[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_6;
      end else if (8'h1b == _T_23[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_5;
      end else if (8'h1b == _T_20[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_4;
      end else if (8'h1b == _T_17[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_3;
      end else if (8'h1b == _T_14[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_2;
      end else if (8'h1b == _T_11[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_1;
      end else if (8'h1b == _T_7[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_28 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1c == _T_29[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_7;
      end else if (8'h1c == _T_26[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_6;
      end else if (8'h1c == _T_23[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_5;
      end else if (8'h1c == _T_20[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_4;
      end else if (8'h1c == _T_17[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_3;
      end else if (8'h1c == _T_14[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_2;
      end else if (8'h1c == _T_11[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_1;
      end else if (8'h1c == _T_7[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_29 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1d == _T_29[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_7;
      end else if (8'h1d == _T_26[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_6;
      end else if (8'h1d == _T_23[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_5;
      end else if (8'h1d == _T_20[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_4;
      end else if (8'h1d == _T_17[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_3;
      end else if (8'h1d == _T_14[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_2;
      end else if (8'h1d == _T_11[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_1;
      end else if (8'h1d == _T_7[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_30 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1e == _T_29[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_7;
      end else if (8'h1e == _T_26[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_6;
      end else if (8'h1e == _T_23[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_5;
      end else if (8'h1e == _T_20[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_4;
      end else if (8'h1e == _T_17[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_3;
      end else if (8'h1e == _T_14[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_2;
      end else if (8'h1e == _T_11[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_1;
      end else if (8'h1e == _T_7[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_31 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1f == _T_29[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_7;
      end else if (8'h1f == _T_26[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_6;
      end else if (8'h1f == _T_23[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_5;
      end else if (8'h1f == _T_20[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_4;
      end else if (8'h1f == _T_17[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_3;
      end else if (8'h1f == _T_14[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_2;
      end else if (8'h1f == _T_11[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_1;
      end else if (8'h1f == _T_7[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_32 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h20 == _T_29[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_7;
      end else if (8'h20 == _T_26[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_6;
      end else if (8'h20 == _T_23[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_5;
      end else if (8'h20 == _T_20[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_4;
      end else if (8'h20 == _T_17[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_3;
      end else if (8'h20 == _T_14[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_2;
      end else if (8'h20 == _T_11[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_1;
      end else if (8'h20 == _T_7[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_33 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h21 == _T_29[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_7;
      end else if (8'h21 == _T_26[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_6;
      end else if (8'h21 == _T_23[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_5;
      end else if (8'h21 == _T_20[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_4;
      end else if (8'h21 == _T_17[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_3;
      end else if (8'h21 == _T_14[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_2;
      end else if (8'h21 == _T_11[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_1;
      end else if (8'h21 == _T_7[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_34 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h22 == _T_29[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_7;
      end else if (8'h22 == _T_26[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_6;
      end else if (8'h22 == _T_23[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_5;
      end else if (8'h22 == _T_20[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_4;
      end else if (8'h22 == _T_17[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_3;
      end else if (8'h22 == _T_14[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_2;
      end else if (8'h22 == _T_11[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_1;
      end else if (8'h22 == _T_7[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_35 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h23 == _T_29[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_7;
      end else if (8'h23 == _T_26[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_6;
      end else if (8'h23 == _T_23[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_5;
      end else if (8'h23 == _T_20[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_4;
      end else if (8'h23 == _T_17[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_3;
      end else if (8'h23 == _T_14[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_2;
      end else if (8'h23 == _T_11[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_1;
      end else if (8'h23 == _T_7[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_36 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h24 == _T_29[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_7;
      end else if (8'h24 == _T_26[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_6;
      end else if (8'h24 == _T_23[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_5;
      end else if (8'h24 == _T_20[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_4;
      end else if (8'h24 == _T_17[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_3;
      end else if (8'h24 == _T_14[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_2;
      end else if (8'h24 == _T_11[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_1;
      end else if (8'h24 == _T_7[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_37 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h25 == _T_29[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_7;
      end else if (8'h25 == _T_26[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_6;
      end else if (8'h25 == _T_23[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_5;
      end else if (8'h25 == _T_20[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_4;
      end else if (8'h25 == _T_17[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_3;
      end else if (8'h25 == _T_14[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_2;
      end else if (8'h25 == _T_11[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_1;
      end else if (8'h25 == _T_7[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_38 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h26 == _T_29[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_7;
      end else if (8'h26 == _T_26[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_6;
      end else if (8'h26 == _T_23[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_5;
      end else if (8'h26 == _T_20[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_4;
      end else if (8'h26 == _T_17[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_3;
      end else if (8'h26 == _T_14[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_2;
      end else if (8'h26 == _T_11[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_1;
      end else if (8'h26 == _T_7[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_39 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h27 == _T_29[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_7;
      end else if (8'h27 == _T_26[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_6;
      end else if (8'h27 == _T_23[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_5;
      end else if (8'h27 == _T_20[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_4;
      end else if (8'h27 == _T_17[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_3;
      end else if (8'h27 == _T_14[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_2;
      end else if (8'h27 == _T_11[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_1;
      end else if (8'h27 == _T_7[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_40 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h28 == _T_29[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_7;
      end else if (8'h28 == _T_26[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_6;
      end else if (8'h28 == _T_23[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_5;
      end else if (8'h28 == _T_20[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_4;
      end else if (8'h28 == _T_17[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_3;
      end else if (8'h28 == _T_14[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_2;
      end else if (8'h28 == _T_11[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_1;
      end else if (8'h28 == _T_7[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_41 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h29 == _T_29[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_7;
      end else if (8'h29 == _T_26[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_6;
      end else if (8'h29 == _T_23[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_5;
      end else if (8'h29 == _T_20[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_4;
      end else if (8'h29 == _T_17[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_3;
      end else if (8'h29 == _T_14[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_2;
      end else if (8'h29 == _T_11[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_1;
      end else if (8'h29 == _T_7[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_42 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2a == _T_29[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_7;
      end else if (8'h2a == _T_26[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_6;
      end else if (8'h2a == _T_23[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_5;
      end else if (8'h2a == _T_20[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_4;
      end else if (8'h2a == _T_17[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_3;
      end else if (8'h2a == _T_14[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_2;
      end else if (8'h2a == _T_11[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_1;
      end else if (8'h2a == _T_7[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_43 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2b == _T_29[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_7;
      end else if (8'h2b == _T_26[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_6;
      end else if (8'h2b == _T_23[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_5;
      end else if (8'h2b == _T_20[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_4;
      end else if (8'h2b == _T_17[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_3;
      end else if (8'h2b == _T_14[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_2;
      end else if (8'h2b == _T_11[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_1;
      end else if (8'h2b == _T_7[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_44 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2c == _T_29[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_7;
      end else if (8'h2c == _T_26[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_6;
      end else if (8'h2c == _T_23[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_5;
      end else if (8'h2c == _T_20[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_4;
      end else if (8'h2c == _T_17[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_3;
      end else if (8'h2c == _T_14[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_2;
      end else if (8'h2c == _T_11[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_1;
      end else if (8'h2c == _T_7[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_45 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2d == _T_29[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_7;
      end else if (8'h2d == _T_26[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_6;
      end else if (8'h2d == _T_23[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_5;
      end else if (8'h2d == _T_20[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_4;
      end else if (8'h2d == _T_17[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_3;
      end else if (8'h2d == _T_14[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_2;
      end else if (8'h2d == _T_11[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_1;
      end else if (8'h2d == _T_7[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_46 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2e == _T_29[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_7;
      end else if (8'h2e == _T_26[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_6;
      end else if (8'h2e == _T_23[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_5;
      end else if (8'h2e == _T_20[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_4;
      end else if (8'h2e == _T_17[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_3;
      end else if (8'h2e == _T_14[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_2;
      end else if (8'h2e == _T_11[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_1;
      end else if (8'h2e == _T_7[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_47 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2f == _T_29[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_7;
      end else if (8'h2f == _T_26[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_6;
      end else if (8'h2f == _T_23[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_5;
      end else if (8'h2f == _T_20[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_4;
      end else if (8'h2f == _T_17[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_3;
      end else if (8'h2f == _T_14[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_2;
      end else if (8'h2f == _T_11[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_1;
      end else if (8'h2f == _T_7[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_48 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h30 == _T_29[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_7;
      end else if (8'h30 == _T_26[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_6;
      end else if (8'h30 == _T_23[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_5;
      end else if (8'h30 == _T_20[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_4;
      end else if (8'h30 == _T_17[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_3;
      end else if (8'h30 == _T_14[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_2;
      end else if (8'h30 == _T_11[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_1;
      end else if (8'h30 == _T_7[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_49 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h31 == _T_29[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_7;
      end else if (8'h31 == _T_26[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_6;
      end else if (8'h31 == _T_23[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_5;
      end else if (8'h31 == _T_20[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_4;
      end else if (8'h31 == _T_17[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_3;
      end else if (8'h31 == _T_14[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_2;
      end else if (8'h31 == _T_11[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_1;
      end else if (8'h31 == _T_7[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_50 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h32 == _T_29[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_7;
      end else if (8'h32 == _T_26[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_6;
      end else if (8'h32 == _T_23[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_5;
      end else if (8'h32 == _T_20[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_4;
      end else if (8'h32 == _T_17[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_3;
      end else if (8'h32 == _T_14[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_2;
      end else if (8'h32 == _T_11[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_1;
      end else if (8'h32 == _T_7[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_51 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h33 == _T_29[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_7;
      end else if (8'h33 == _T_26[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_6;
      end else if (8'h33 == _T_23[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_5;
      end else if (8'h33 == _T_20[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_4;
      end else if (8'h33 == _T_17[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_3;
      end else if (8'h33 == _T_14[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_2;
      end else if (8'h33 == _T_11[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_1;
      end else if (8'h33 == _T_7[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_52 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h34 == _T_29[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_7;
      end else if (8'h34 == _T_26[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_6;
      end else if (8'h34 == _T_23[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_5;
      end else if (8'h34 == _T_20[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_4;
      end else if (8'h34 == _T_17[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_3;
      end else if (8'h34 == _T_14[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_2;
      end else if (8'h34 == _T_11[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_1;
      end else if (8'h34 == _T_7[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_53 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h35 == _T_29[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_7;
      end else if (8'h35 == _T_26[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_6;
      end else if (8'h35 == _T_23[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_5;
      end else if (8'h35 == _T_20[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_4;
      end else if (8'h35 == _T_17[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_3;
      end else if (8'h35 == _T_14[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_2;
      end else if (8'h35 == _T_11[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_1;
      end else if (8'h35 == _T_7[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_54 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h36 == _T_29[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_7;
      end else if (8'h36 == _T_26[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_6;
      end else if (8'h36 == _T_23[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_5;
      end else if (8'h36 == _T_20[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_4;
      end else if (8'h36 == _T_17[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_3;
      end else if (8'h36 == _T_14[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_2;
      end else if (8'h36 == _T_11[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_1;
      end else if (8'h36 == _T_7[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_55 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h37 == _T_29[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_7;
      end else if (8'h37 == _T_26[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_6;
      end else if (8'h37 == _T_23[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_5;
      end else if (8'h37 == _T_20[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_4;
      end else if (8'h37 == _T_17[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_3;
      end else if (8'h37 == _T_14[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_2;
      end else if (8'h37 == _T_11[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_1;
      end else if (8'h37 == _T_7[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_56 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h38 == _T_29[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_7;
      end else if (8'h38 == _T_26[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_6;
      end else if (8'h38 == _T_23[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_5;
      end else if (8'h38 == _T_20[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_4;
      end else if (8'h38 == _T_17[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_3;
      end else if (8'h38 == _T_14[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_2;
      end else if (8'h38 == _T_11[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_1;
      end else if (8'h38 == _T_7[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_57 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h39 == _T_29[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_7;
      end else if (8'h39 == _T_26[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_6;
      end else if (8'h39 == _T_23[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_5;
      end else if (8'h39 == _T_20[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_4;
      end else if (8'h39 == _T_17[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_3;
      end else if (8'h39 == _T_14[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_2;
      end else if (8'h39 == _T_11[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_1;
      end else if (8'h39 == _T_7[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_58 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3a == _T_29[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_7;
      end else if (8'h3a == _T_26[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_6;
      end else if (8'h3a == _T_23[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_5;
      end else if (8'h3a == _T_20[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_4;
      end else if (8'h3a == _T_17[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_3;
      end else if (8'h3a == _T_14[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_2;
      end else if (8'h3a == _T_11[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_1;
      end else if (8'h3a == _T_7[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_59 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3b == _T_29[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_7;
      end else if (8'h3b == _T_26[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_6;
      end else if (8'h3b == _T_23[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_5;
      end else if (8'h3b == _T_20[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_4;
      end else if (8'h3b == _T_17[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_3;
      end else if (8'h3b == _T_14[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_2;
      end else if (8'h3b == _T_11[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_1;
      end else if (8'h3b == _T_7[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_60 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3c == _T_29[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_7;
      end else if (8'h3c == _T_26[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_6;
      end else if (8'h3c == _T_23[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_5;
      end else if (8'h3c == _T_20[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_4;
      end else if (8'h3c == _T_17[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_3;
      end else if (8'h3c == _T_14[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_2;
      end else if (8'h3c == _T_11[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_1;
      end else if (8'h3c == _T_7[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_61 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3d == _T_29[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_7;
      end else if (8'h3d == _T_26[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_6;
      end else if (8'h3d == _T_23[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_5;
      end else if (8'h3d == _T_20[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_4;
      end else if (8'h3d == _T_17[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_3;
      end else if (8'h3d == _T_14[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_2;
      end else if (8'h3d == _T_11[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_1;
      end else if (8'h3d == _T_7[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_62 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3e == _T_29[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_7;
      end else if (8'h3e == _T_26[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_6;
      end else if (8'h3e == _T_23[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_5;
      end else if (8'h3e == _T_20[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_4;
      end else if (8'h3e == _T_17[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_3;
      end else if (8'h3e == _T_14[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_2;
      end else if (8'h3e == _T_11[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_1;
      end else if (8'h3e == _T_7[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_63 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3f == _T_29[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_7;
      end else if (8'h3f == _T_26[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_6;
      end else if (8'h3f == _T_23[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_5;
      end else if (8'h3f == _T_20[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_4;
      end else if (8'h3f == _T_17[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_3;
      end else if (8'h3f == _T_14[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_2;
      end else if (8'h3f == _T_11[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_1;
      end else if (8'h3f == _T_7[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_64 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h40 == _T_29[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_7;
      end else if (8'h40 == _T_26[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_6;
      end else if (8'h40 == _T_23[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_5;
      end else if (8'h40 == _T_20[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_4;
      end else if (8'h40 == _T_17[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_3;
      end else if (8'h40 == _T_14[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_2;
      end else if (8'h40 == _T_11[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_1;
      end else if (8'h40 == _T_7[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_65 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h41 == _T_29[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_7;
      end else if (8'h41 == _T_26[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_6;
      end else if (8'h41 == _T_23[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_5;
      end else if (8'h41 == _T_20[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_4;
      end else if (8'h41 == _T_17[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_3;
      end else if (8'h41 == _T_14[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_2;
      end else if (8'h41 == _T_11[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_1;
      end else if (8'h41 == _T_7[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_66 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h42 == _T_29[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_7;
      end else if (8'h42 == _T_26[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_6;
      end else if (8'h42 == _T_23[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_5;
      end else if (8'h42 == _T_20[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_4;
      end else if (8'h42 == _T_17[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_3;
      end else if (8'h42 == _T_14[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_2;
      end else if (8'h42 == _T_11[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_1;
      end else if (8'h42 == _T_7[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_67 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h43 == _T_29[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_7;
      end else if (8'h43 == _T_26[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_6;
      end else if (8'h43 == _T_23[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_5;
      end else if (8'h43 == _T_20[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_4;
      end else if (8'h43 == _T_17[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_3;
      end else if (8'h43 == _T_14[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_2;
      end else if (8'h43 == _T_11[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_1;
      end else if (8'h43 == _T_7[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_68 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h44 == _T_29[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_7;
      end else if (8'h44 == _T_26[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_6;
      end else if (8'h44 == _T_23[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_5;
      end else if (8'h44 == _T_20[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_4;
      end else if (8'h44 == _T_17[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_3;
      end else if (8'h44 == _T_14[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_2;
      end else if (8'h44 == _T_11[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_1;
      end else if (8'h44 == _T_7[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_69 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h45 == _T_29[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_7;
      end else if (8'h45 == _T_26[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_6;
      end else if (8'h45 == _T_23[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_5;
      end else if (8'h45 == _T_20[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_4;
      end else if (8'h45 == _T_17[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_3;
      end else if (8'h45 == _T_14[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_2;
      end else if (8'h45 == _T_11[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_1;
      end else if (8'h45 == _T_7[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_70 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h46 == _T_29[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_7;
      end else if (8'h46 == _T_26[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_6;
      end else if (8'h46 == _T_23[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_5;
      end else if (8'h46 == _T_20[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_4;
      end else if (8'h46 == _T_17[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_3;
      end else if (8'h46 == _T_14[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_2;
      end else if (8'h46 == _T_11[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_1;
      end else if (8'h46 == _T_7[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_71 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h47 == _T_29[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_7;
      end else if (8'h47 == _T_26[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_6;
      end else if (8'h47 == _T_23[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_5;
      end else if (8'h47 == _T_20[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_4;
      end else if (8'h47 == _T_17[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_3;
      end else if (8'h47 == _T_14[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_2;
      end else if (8'h47 == _T_11[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_1;
      end else if (8'h47 == _T_7[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_72 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h48 == _T_29[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_7;
      end else if (8'h48 == _T_26[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_6;
      end else if (8'h48 == _T_23[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_5;
      end else if (8'h48 == _T_20[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_4;
      end else if (8'h48 == _T_17[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_3;
      end else if (8'h48 == _T_14[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_2;
      end else if (8'h48 == _T_11[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_1;
      end else if (8'h48 == _T_7[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_73 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h49 == _T_29[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_7;
      end else if (8'h49 == _T_26[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_6;
      end else if (8'h49 == _T_23[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_5;
      end else if (8'h49 == _T_20[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_4;
      end else if (8'h49 == _T_17[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_3;
      end else if (8'h49 == _T_14[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_2;
      end else if (8'h49 == _T_11[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_1;
      end else if (8'h49 == _T_7[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_74 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4a == _T_29[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_7;
      end else if (8'h4a == _T_26[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_6;
      end else if (8'h4a == _T_23[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_5;
      end else if (8'h4a == _T_20[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_4;
      end else if (8'h4a == _T_17[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_3;
      end else if (8'h4a == _T_14[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_2;
      end else if (8'h4a == _T_11[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_1;
      end else if (8'h4a == _T_7[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_75 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4b == _T_29[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_7;
      end else if (8'h4b == _T_26[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_6;
      end else if (8'h4b == _T_23[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_5;
      end else if (8'h4b == _T_20[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_4;
      end else if (8'h4b == _T_17[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_3;
      end else if (8'h4b == _T_14[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_2;
      end else if (8'h4b == _T_11[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_1;
      end else if (8'h4b == _T_7[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_76 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4c == _T_29[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_7;
      end else if (8'h4c == _T_26[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_6;
      end else if (8'h4c == _T_23[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_5;
      end else if (8'h4c == _T_20[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_4;
      end else if (8'h4c == _T_17[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_3;
      end else if (8'h4c == _T_14[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_2;
      end else if (8'h4c == _T_11[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_1;
      end else if (8'h4c == _T_7[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_77 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4d == _T_29[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_7;
      end else if (8'h4d == _T_26[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_6;
      end else if (8'h4d == _T_23[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_5;
      end else if (8'h4d == _T_20[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_4;
      end else if (8'h4d == _T_17[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_3;
      end else if (8'h4d == _T_14[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_2;
      end else if (8'h4d == _T_11[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_1;
      end else if (8'h4d == _T_7[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_78 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4e == _T_29[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_7;
      end else if (8'h4e == _T_26[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_6;
      end else if (8'h4e == _T_23[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_5;
      end else if (8'h4e == _T_20[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_4;
      end else if (8'h4e == _T_17[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_3;
      end else if (8'h4e == _T_14[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_2;
      end else if (8'h4e == _T_11[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_1;
      end else if (8'h4e == _T_7[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_79 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4f == _T_29[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_7;
      end else if (8'h4f == _T_26[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_6;
      end else if (8'h4f == _T_23[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_5;
      end else if (8'h4f == _T_20[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_4;
      end else if (8'h4f == _T_17[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_3;
      end else if (8'h4f == _T_14[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_2;
      end else if (8'h4f == _T_11[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_1;
      end else if (8'h4f == _T_7[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_80 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h50 == _T_29[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_7;
      end else if (8'h50 == _T_26[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_6;
      end else if (8'h50 == _T_23[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_5;
      end else if (8'h50 == _T_20[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_4;
      end else if (8'h50 == _T_17[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_3;
      end else if (8'h50 == _T_14[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_2;
      end else if (8'h50 == _T_11[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_1;
      end else if (8'h50 == _T_7[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_81 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h51 == _T_29[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_7;
      end else if (8'h51 == _T_26[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_6;
      end else if (8'h51 == _T_23[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_5;
      end else if (8'h51 == _T_20[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_4;
      end else if (8'h51 == _T_17[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_3;
      end else if (8'h51 == _T_14[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_2;
      end else if (8'h51 == _T_11[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_1;
      end else if (8'h51 == _T_7[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_82 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h52 == _T_29[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_7;
      end else if (8'h52 == _T_26[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_6;
      end else if (8'h52 == _T_23[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_5;
      end else if (8'h52 == _T_20[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_4;
      end else if (8'h52 == _T_17[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_3;
      end else if (8'h52 == _T_14[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_2;
      end else if (8'h52 == _T_11[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_1;
      end else if (8'h52 == _T_7[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_83 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h53 == _T_29[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_7;
      end else if (8'h53 == _T_26[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_6;
      end else if (8'h53 == _T_23[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_5;
      end else if (8'h53 == _T_20[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_4;
      end else if (8'h53 == _T_17[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_3;
      end else if (8'h53 == _T_14[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_2;
      end else if (8'h53 == _T_11[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_1;
      end else if (8'h53 == _T_7[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_84 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h54 == _T_29[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_7;
      end else if (8'h54 == _T_26[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_6;
      end else if (8'h54 == _T_23[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_5;
      end else if (8'h54 == _T_20[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_4;
      end else if (8'h54 == _T_17[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_3;
      end else if (8'h54 == _T_14[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_2;
      end else if (8'h54 == _T_11[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_1;
      end else if (8'h54 == _T_7[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_85 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h55 == _T_29[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_7;
      end else if (8'h55 == _T_26[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_6;
      end else if (8'h55 == _T_23[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_5;
      end else if (8'h55 == _T_20[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_4;
      end else if (8'h55 == _T_17[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_3;
      end else if (8'h55 == _T_14[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_2;
      end else if (8'h55 == _T_11[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_1;
      end else if (8'h55 == _T_7[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_86 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h56 == _T_29[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_7;
      end else if (8'h56 == _T_26[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_6;
      end else if (8'h56 == _T_23[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_5;
      end else if (8'h56 == _T_20[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_4;
      end else if (8'h56 == _T_17[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_3;
      end else if (8'h56 == _T_14[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_2;
      end else if (8'h56 == _T_11[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_1;
      end else if (8'h56 == _T_7[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_87 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h57 == _T_29[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_7;
      end else if (8'h57 == _T_26[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_6;
      end else if (8'h57 == _T_23[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_5;
      end else if (8'h57 == _T_20[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_4;
      end else if (8'h57 == _T_17[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_3;
      end else if (8'h57 == _T_14[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_2;
      end else if (8'h57 == _T_11[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_1;
      end else if (8'h57 == _T_7[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_88 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h58 == _T_29[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_7;
      end else if (8'h58 == _T_26[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_6;
      end else if (8'h58 == _T_23[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_5;
      end else if (8'h58 == _T_20[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_4;
      end else if (8'h58 == _T_17[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_3;
      end else if (8'h58 == _T_14[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_2;
      end else if (8'h58 == _T_11[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_1;
      end else if (8'h58 == _T_7[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_89 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h59 == _T_29[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_7;
      end else if (8'h59 == _T_26[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_6;
      end else if (8'h59 == _T_23[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_5;
      end else if (8'h59 == _T_20[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_4;
      end else if (8'h59 == _T_17[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_3;
      end else if (8'h59 == _T_14[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_2;
      end else if (8'h59 == _T_11[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_1;
      end else if (8'h59 == _T_7[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_90 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5a == _T_29[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_7;
      end else if (8'h5a == _T_26[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_6;
      end else if (8'h5a == _T_23[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_5;
      end else if (8'h5a == _T_20[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_4;
      end else if (8'h5a == _T_17[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_3;
      end else if (8'h5a == _T_14[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_2;
      end else if (8'h5a == _T_11[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_1;
      end else if (8'h5a == _T_7[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_91 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5b == _T_29[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_7;
      end else if (8'h5b == _T_26[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_6;
      end else if (8'h5b == _T_23[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_5;
      end else if (8'h5b == _T_20[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_4;
      end else if (8'h5b == _T_17[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_3;
      end else if (8'h5b == _T_14[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_2;
      end else if (8'h5b == _T_11[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_1;
      end else if (8'h5b == _T_7[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_92 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5c == _T_29[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_7;
      end else if (8'h5c == _T_26[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_6;
      end else if (8'h5c == _T_23[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_5;
      end else if (8'h5c == _T_20[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_4;
      end else if (8'h5c == _T_17[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_3;
      end else if (8'h5c == _T_14[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_2;
      end else if (8'h5c == _T_11[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_1;
      end else if (8'h5c == _T_7[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_93 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5d == _T_29[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_7;
      end else if (8'h5d == _T_26[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_6;
      end else if (8'h5d == _T_23[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_5;
      end else if (8'h5d == _T_20[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_4;
      end else if (8'h5d == _T_17[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_3;
      end else if (8'h5d == _T_14[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_2;
      end else if (8'h5d == _T_11[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_1;
      end else if (8'h5d == _T_7[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_94 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5e == _T_29[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_7;
      end else if (8'h5e == _T_26[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_6;
      end else if (8'h5e == _T_23[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_5;
      end else if (8'h5e == _T_20[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_4;
      end else if (8'h5e == _T_17[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_3;
      end else if (8'h5e == _T_14[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_2;
      end else if (8'h5e == _T_11[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_1;
      end else if (8'h5e == _T_7[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_95 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5f == _T_29[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_7;
      end else if (8'h5f == _T_26[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_6;
      end else if (8'h5f == _T_23[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_5;
      end else if (8'h5f == _T_20[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_4;
      end else if (8'h5f == _T_17[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_3;
      end else if (8'h5f == _T_14[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_2;
      end else if (8'h5f == _T_11[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_1;
      end else if (8'h5f == _T_7[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_96 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h60 == _T_29[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_7;
      end else if (8'h60 == _T_26[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_6;
      end else if (8'h60 == _T_23[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_5;
      end else if (8'h60 == _T_20[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_4;
      end else if (8'h60 == _T_17[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_3;
      end else if (8'h60 == _T_14[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_2;
      end else if (8'h60 == _T_11[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_1;
      end else if (8'h60 == _T_7[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_97 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h61 == _T_29[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_7;
      end else if (8'h61 == _T_26[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_6;
      end else if (8'h61 == _T_23[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_5;
      end else if (8'h61 == _T_20[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_4;
      end else if (8'h61 == _T_17[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_3;
      end else if (8'h61 == _T_14[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_2;
      end else if (8'h61 == _T_11[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_1;
      end else if (8'h61 == _T_7[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_98 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h62 == _T_29[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_7;
      end else if (8'h62 == _T_26[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_6;
      end else if (8'h62 == _T_23[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_5;
      end else if (8'h62 == _T_20[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_4;
      end else if (8'h62 == _T_17[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_3;
      end else if (8'h62 == _T_14[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_2;
      end else if (8'h62 == _T_11[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_1;
      end else if (8'h62 == _T_7[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_99 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h63 == _T_29[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_7;
      end else if (8'h63 == _T_26[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_6;
      end else if (8'h63 == _T_23[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_5;
      end else if (8'h63 == _T_20[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_4;
      end else if (8'h63 == _T_17[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_3;
      end else if (8'h63 == _T_14[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_2;
      end else if (8'h63 == _T_11[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_1;
      end else if (8'h63 == _T_7[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_100 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h64 == _T_29[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_7;
      end else if (8'h64 == _T_26[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_6;
      end else if (8'h64 == _T_23[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_5;
      end else if (8'h64 == _T_20[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_4;
      end else if (8'h64 == _T_17[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_3;
      end else if (8'h64 == _T_14[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_2;
      end else if (8'h64 == _T_11[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_1;
      end else if (8'h64 == _T_7[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_101 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h65 == _T_29[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_7;
      end else if (8'h65 == _T_26[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_6;
      end else if (8'h65 == _T_23[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_5;
      end else if (8'h65 == _T_20[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_4;
      end else if (8'h65 == _T_17[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_3;
      end else if (8'h65 == _T_14[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_2;
      end else if (8'h65 == _T_11[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_1;
      end else if (8'h65 == _T_7[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_102 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h66 == _T_29[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_7;
      end else if (8'h66 == _T_26[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_6;
      end else if (8'h66 == _T_23[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_5;
      end else if (8'h66 == _T_20[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_4;
      end else if (8'h66 == _T_17[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_3;
      end else if (8'h66 == _T_14[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_2;
      end else if (8'h66 == _T_11[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_1;
      end else if (8'h66 == _T_7[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_103 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h67 == _T_29[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_7;
      end else if (8'h67 == _T_26[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_6;
      end else if (8'h67 == _T_23[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_5;
      end else if (8'h67 == _T_20[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_4;
      end else if (8'h67 == _T_17[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_3;
      end else if (8'h67 == _T_14[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_2;
      end else if (8'h67 == _T_11[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_1;
      end else if (8'h67 == _T_7[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_104 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h68 == _T_29[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_7;
      end else if (8'h68 == _T_26[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_6;
      end else if (8'h68 == _T_23[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_5;
      end else if (8'h68 == _T_20[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_4;
      end else if (8'h68 == _T_17[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_3;
      end else if (8'h68 == _T_14[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_2;
      end else if (8'h68 == _T_11[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_1;
      end else if (8'h68 == _T_7[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_105 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h69 == _T_29[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_7;
      end else if (8'h69 == _T_26[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_6;
      end else if (8'h69 == _T_23[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_5;
      end else if (8'h69 == _T_20[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_4;
      end else if (8'h69 == _T_17[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_3;
      end else if (8'h69 == _T_14[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_2;
      end else if (8'h69 == _T_11[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_1;
      end else if (8'h69 == _T_7[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_106 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6a == _T_29[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_7;
      end else if (8'h6a == _T_26[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_6;
      end else if (8'h6a == _T_23[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_5;
      end else if (8'h6a == _T_20[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_4;
      end else if (8'h6a == _T_17[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_3;
      end else if (8'h6a == _T_14[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_2;
      end else if (8'h6a == _T_11[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_1;
      end else if (8'h6a == _T_7[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_107 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6b == _T_29[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_7;
      end else if (8'h6b == _T_26[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_6;
      end else if (8'h6b == _T_23[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_5;
      end else if (8'h6b == _T_20[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_4;
      end else if (8'h6b == _T_17[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_3;
      end else if (8'h6b == _T_14[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_2;
      end else if (8'h6b == _T_11[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_1;
      end else if (8'h6b == _T_7[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_108 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6c == _T_29[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_7;
      end else if (8'h6c == _T_26[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_6;
      end else if (8'h6c == _T_23[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_5;
      end else if (8'h6c == _T_20[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_4;
      end else if (8'h6c == _T_17[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_3;
      end else if (8'h6c == _T_14[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_2;
      end else if (8'h6c == _T_11[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_1;
      end else if (8'h6c == _T_7[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_109 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6d == _T_29[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_7;
      end else if (8'h6d == _T_26[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_6;
      end else if (8'h6d == _T_23[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_5;
      end else if (8'h6d == _T_20[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_4;
      end else if (8'h6d == _T_17[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_3;
      end else if (8'h6d == _T_14[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_2;
      end else if (8'h6d == _T_11[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_1;
      end else if (8'h6d == _T_7[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_110 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6e == _T_29[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_7;
      end else if (8'h6e == _T_26[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_6;
      end else if (8'h6e == _T_23[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_5;
      end else if (8'h6e == _T_20[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_4;
      end else if (8'h6e == _T_17[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_3;
      end else if (8'h6e == _T_14[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_2;
      end else if (8'h6e == _T_11[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_1;
      end else if (8'h6e == _T_7[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_111 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6f == _T_29[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_7;
      end else if (8'h6f == _T_26[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_6;
      end else if (8'h6f == _T_23[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_5;
      end else if (8'h6f == _T_20[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_4;
      end else if (8'h6f == _T_17[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_3;
      end else if (8'h6f == _T_14[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_2;
      end else if (8'h6f == _T_11[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_1;
      end else if (8'h6f == _T_7[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_112 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h70 == _T_29[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_7;
      end else if (8'h70 == _T_26[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_6;
      end else if (8'h70 == _T_23[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_5;
      end else if (8'h70 == _T_20[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_4;
      end else if (8'h70 == _T_17[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_3;
      end else if (8'h70 == _T_14[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_2;
      end else if (8'h70 == _T_11[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_1;
      end else if (8'h70 == _T_7[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_113 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h71 == _T_29[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_7;
      end else if (8'h71 == _T_26[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_6;
      end else if (8'h71 == _T_23[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_5;
      end else if (8'h71 == _T_20[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_4;
      end else if (8'h71 == _T_17[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_3;
      end else if (8'h71 == _T_14[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_2;
      end else if (8'h71 == _T_11[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_1;
      end else if (8'h71 == _T_7[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_114 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h72 == _T_29[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_7;
      end else if (8'h72 == _T_26[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_6;
      end else if (8'h72 == _T_23[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_5;
      end else if (8'h72 == _T_20[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_4;
      end else if (8'h72 == _T_17[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_3;
      end else if (8'h72 == _T_14[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_2;
      end else if (8'h72 == _T_11[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_1;
      end else if (8'h72 == _T_7[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_115 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h73 == _T_29[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_7;
      end else if (8'h73 == _T_26[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_6;
      end else if (8'h73 == _T_23[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_5;
      end else if (8'h73 == _T_20[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_4;
      end else if (8'h73 == _T_17[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_3;
      end else if (8'h73 == _T_14[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_2;
      end else if (8'h73 == _T_11[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_1;
      end else if (8'h73 == _T_7[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_116 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h74 == _T_29[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_7;
      end else if (8'h74 == _T_26[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_6;
      end else if (8'h74 == _T_23[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_5;
      end else if (8'h74 == _T_20[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_4;
      end else if (8'h74 == _T_17[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_3;
      end else if (8'h74 == _T_14[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_2;
      end else if (8'h74 == _T_11[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_1;
      end else if (8'h74 == _T_7[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_117 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h75 == _T_29[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_7;
      end else if (8'h75 == _T_26[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_6;
      end else if (8'h75 == _T_23[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_5;
      end else if (8'h75 == _T_20[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_4;
      end else if (8'h75 == _T_17[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_3;
      end else if (8'h75 == _T_14[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_2;
      end else if (8'h75 == _T_11[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_1;
      end else if (8'h75 == _T_7[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_118 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h76 == _T_29[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_7;
      end else if (8'h76 == _T_26[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_6;
      end else if (8'h76 == _T_23[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_5;
      end else if (8'h76 == _T_20[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_4;
      end else if (8'h76 == _T_17[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_3;
      end else if (8'h76 == _T_14[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_2;
      end else if (8'h76 == _T_11[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_1;
      end else if (8'h76 == _T_7[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_119 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h77 == _T_29[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_7;
      end else if (8'h77 == _T_26[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_6;
      end else if (8'h77 == _T_23[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_5;
      end else if (8'h77 == _T_20[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_4;
      end else if (8'h77 == _T_17[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_3;
      end else if (8'h77 == _T_14[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_2;
      end else if (8'h77 == _T_11[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_1;
      end else if (8'h77 == _T_7[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_120 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h78 == _T_29[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_7;
      end else if (8'h78 == _T_26[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_6;
      end else if (8'h78 == _T_23[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_5;
      end else if (8'h78 == _T_20[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_4;
      end else if (8'h78 == _T_17[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_3;
      end else if (8'h78 == _T_14[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_2;
      end else if (8'h78 == _T_11[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_1;
      end else if (8'h78 == _T_7[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_121 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h79 == _T_29[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_7;
      end else if (8'h79 == _T_26[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_6;
      end else if (8'h79 == _T_23[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_5;
      end else if (8'h79 == _T_20[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_4;
      end else if (8'h79 == _T_17[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_3;
      end else if (8'h79 == _T_14[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_2;
      end else if (8'h79 == _T_11[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_1;
      end else if (8'h79 == _T_7[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_122 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7a == _T_29[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_7;
      end else if (8'h7a == _T_26[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_6;
      end else if (8'h7a == _T_23[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_5;
      end else if (8'h7a == _T_20[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_4;
      end else if (8'h7a == _T_17[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_3;
      end else if (8'h7a == _T_14[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_2;
      end else if (8'h7a == _T_11[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_1;
      end else if (8'h7a == _T_7[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_123 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7b == _T_29[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_7;
      end else if (8'h7b == _T_26[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_6;
      end else if (8'h7b == _T_23[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_5;
      end else if (8'h7b == _T_20[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_4;
      end else if (8'h7b == _T_17[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_3;
      end else if (8'h7b == _T_14[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_2;
      end else if (8'h7b == _T_11[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_1;
      end else if (8'h7b == _T_7[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_124 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7c == _T_29[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_7;
      end else if (8'h7c == _T_26[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_6;
      end else if (8'h7c == _T_23[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_5;
      end else if (8'h7c == _T_20[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_4;
      end else if (8'h7c == _T_17[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_3;
      end else if (8'h7c == _T_14[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_2;
      end else if (8'h7c == _T_11[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_1;
      end else if (8'h7c == _T_7[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_125 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7d == _T_29[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_7;
      end else if (8'h7d == _T_26[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_6;
      end else if (8'h7d == _T_23[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_5;
      end else if (8'h7d == _T_20[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_4;
      end else if (8'h7d == _T_17[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_3;
      end else if (8'h7d == _T_14[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_2;
      end else if (8'h7d == _T_11[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_1;
      end else if (8'h7d == _T_7[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_126 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7e == _T_29[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_7;
      end else if (8'h7e == _T_26[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_6;
      end else if (8'h7e == _T_23[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_5;
      end else if (8'h7e == _T_20[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_4;
      end else if (8'h7e == _T_17[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_3;
      end else if (8'h7e == _T_14[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_2;
      end else if (8'h7e == _T_11[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_1;
      end else if (8'h7e == _T_7[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_127 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7f == _T_29[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_7;
      end else if (8'h7f == _T_26[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_6;
      end else if (8'h7f == _T_23[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_5;
      end else if (8'h7f == _T_20[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_4;
      end else if (8'h7f == _T_17[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_3;
      end else if (8'h7f == _T_14[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_2;
      end else if (8'h7f == _T_11[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_1;
      end else if (8'h7f == _T_7[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_128 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h80 == _T_29[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_7;
      end else if (8'h80 == _T_26[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_6;
      end else if (8'h80 == _T_23[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_5;
      end else if (8'h80 == _T_20[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_4;
      end else if (8'h80 == _T_17[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_3;
      end else if (8'h80 == _T_14[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_2;
      end else if (8'h80 == _T_11[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_1;
      end else if (8'h80 == _T_7[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_129 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h81 == _T_29[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_7;
      end else if (8'h81 == _T_26[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_6;
      end else if (8'h81 == _T_23[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_5;
      end else if (8'h81 == _T_20[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_4;
      end else if (8'h81 == _T_17[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_3;
      end else if (8'h81 == _T_14[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_2;
      end else if (8'h81 == _T_11[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_1;
      end else if (8'h81 == _T_7[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_130 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h82 == _T_29[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_7;
      end else if (8'h82 == _T_26[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_6;
      end else if (8'h82 == _T_23[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_5;
      end else if (8'h82 == _T_20[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_4;
      end else if (8'h82 == _T_17[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_3;
      end else if (8'h82 == _T_14[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_2;
      end else if (8'h82 == _T_11[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_1;
      end else if (8'h82 == _T_7[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_131 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h83 == _T_29[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_7;
      end else if (8'h83 == _T_26[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_6;
      end else if (8'h83 == _T_23[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_5;
      end else if (8'h83 == _T_20[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_4;
      end else if (8'h83 == _T_17[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_3;
      end else if (8'h83 == _T_14[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_2;
      end else if (8'h83 == _T_11[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_1;
      end else if (8'h83 == _T_7[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_132 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h84 == _T_29[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_7;
      end else if (8'h84 == _T_26[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_6;
      end else if (8'h84 == _T_23[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_5;
      end else if (8'h84 == _T_20[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_4;
      end else if (8'h84 == _T_17[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_3;
      end else if (8'h84 == _T_14[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_2;
      end else if (8'h84 == _T_11[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_1;
      end else if (8'h84 == _T_7[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_133 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h85 == _T_29[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_7;
      end else if (8'h85 == _T_26[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_6;
      end else if (8'h85 == _T_23[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_5;
      end else if (8'h85 == _T_20[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_4;
      end else if (8'h85 == _T_17[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_3;
      end else if (8'h85 == _T_14[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_2;
      end else if (8'h85 == _T_11[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_1;
      end else if (8'h85 == _T_7[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_134 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h86 == _T_29[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_7;
      end else if (8'h86 == _T_26[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_6;
      end else if (8'h86 == _T_23[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_5;
      end else if (8'h86 == _T_20[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_4;
      end else if (8'h86 == _T_17[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_3;
      end else if (8'h86 == _T_14[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_2;
      end else if (8'h86 == _T_11[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_1;
      end else if (8'h86 == _T_7[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_135 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h87 == _T_29[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_7;
      end else if (8'h87 == _T_26[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_6;
      end else if (8'h87 == _T_23[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_5;
      end else if (8'h87 == _T_20[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_4;
      end else if (8'h87 == _T_17[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_3;
      end else if (8'h87 == _T_14[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_2;
      end else if (8'h87 == _T_11[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_1;
      end else if (8'h87 == _T_7[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_136 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h88 == _T_29[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_7;
      end else if (8'h88 == _T_26[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_6;
      end else if (8'h88 == _T_23[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_5;
      end else if (8'h88 == _T_20[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_4;
      end else if (8'h88 == _T_17[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_3;
      end else if (8'h88 == _T_14[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_2;
      end else if (8'h88 == _T_11[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_1;
      end else if (8'h88 == _T_7[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_137 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h89 == _T_29[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_7;
      end else if (8'h89 == _T_26[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_6;
      end else if (8'h89 == _T_23[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_5;
      end else if (8'h89 == _T_20[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_4;
      end else if (8'h89 == _T_17[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_3;
      end else if (8'h89 == _T_14[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_2;
      end else if (8'h89 == _T_11[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_1;
      end else if (8'h89 == _T_7[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_138 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8a == _T_29[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_7;
      end else if (8'h8a == _T_26[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_6;
      end else if (8'h8a == _T_23[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_5;
      end else if (8'h8a == _T_20[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_4;
      end else if (8'h8a == _T_17[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_3;
      end else if (8'h8a == _T_14[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_2;
      end else if (8'h8a == _T_11[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_1;
      end else if (8'h8a == _T_7[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_139 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8b == _T_29[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_7;
      end else if (8'h8b == _T_26[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_6;
      end else if (8'h8b == _T_23[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_5;
      end else if (8'h8b == _T_20[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_4;
      end else if (8'h8b == _T_17[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_3;
      end else if (8'h8b == _T_14[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_2;
      end else if (8'h8b == _T_11[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_1;
      end else if (8'h8b == _T_7[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_140 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8c == _T_29[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_7;
      end else if (8'h8c == _T_26[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_6;
      end else if (8'h8c == _T_23[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_5;
      end else if (8'h8c == _T_20[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_4;
      end else if (8'h8c == _T_17[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_3;
      end else if (8'h8c == _T_14[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_2;
      end else if (8'h8c == _T_11[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_1;
      end else if (8'h8c == _T_7[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_141 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8d == _T_29[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_7;
      end else if (8'h8d == _T_26[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_6;
      end else if (8'h8d == _T_23[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_5;
      end else if (8'h8d == _T_20[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_4;
      end else if (8'h8d == _T_17[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_3;
      end else if (8'h8d == _T_14[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_2;
      end else if (8'h8d == _T_11[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_1;
      end else if (8'h8d == _T_7[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_142 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8e == _T_29[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_7;
      end else if (8'h8e == _T_26[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_6;
      end else if (8'h8e == _T_23[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_5;
      end else if (8'h8e == _T_20[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_4;
      end else if (8'h8e == _T_17[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_3;
      end else if (8'h8e == _T_14[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_2;
      end else if (8'h8e == _T_11[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_1;
      end else if (8'h8e == _T_7[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_143 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8f == _T_29[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_7;
      end else if (8'h8f == _T_26[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_6;
      end else if (8'h8f == _T_23[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_5;
      end else if (8'h8f == _T_20[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_4;
      end else if (8'h8f == _T_17[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_3;
      end else if (8'h8f == _T_14[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_2;
      end else if (8'h8f == _T_11[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_1;
      end else if (8'h8f == _T_7[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_144 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h90 == _T_29[7:0]) begin
        image_1_144 <= io_pixelVal_in_1_7;
      end else if (8'h90 == _T_26[7:0]) begin
        image_1_144 <= io_pixelVal_in_1_6;
      end else if (8'h90 == _T_23[7:0]) begin
        image_1_144 <= io_pixelVal_in_1_5;
      end else if (8'h90 == _T_20[7:0]) begin
        image_1_144 <= io_pixelVal_in_1_4;
      end else if (8'h90 == _T_17[7:0]) begin
        image_1_144 <= io_pixelVal_in_1_3;
      end else if (8'h90 == _T_14[7:0]) begin
        image_1_144 <= io_pixelVal_in_1_2;
      end else if (8'h90 == _T_11[7:0]) begin
        image_1_144 <= io_pixelVal_in_1_1;
      end else if (8'h90 == _T_7[7:0]) begin
        image_1_144 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_145 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h91 == _T_29[7:0]) begin
        image_1_145 <= io_pixelVal_in_1_7;
      end else if (8'h91 == _T_26[7:0]) begin
        image_1_145 <= io_pixelVal_in_1_6;
      end else if (8'h91 == _T_23[7:0]) begin
        image_1_145 <= io_pixelVal_in_1_5;
      end else if (8'h91 == _T_20[7:0]) begin
        image_1_145 <= io_pixelVal_in_1_4;
      end else if (8'h91 == _T_17[7:0]) begin
        image_1_145 <= io_pixelVal_in_1_3;
      end else if (8'h91 == _T_14[7:0]) begin
        image_1_145 <= io_pixelVal_in_1_2;
      end else if (8'h91 == _T_11[7:0]) begin
        image_1_145 <= io_pixelVal_in_1_1;
      end else if (8'h91 == _T_7[7:0]) begin
        image_1_145 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_146 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h92 == _T_29[7:0]) begin
        image_1_146 <= io_pixelVal_in_1_7;
      end else if (8'h92 == _T_26[7:0]) begin
        image_1_146 <= io_pixelVal_in_1_6;
      end else if (8'h92 == _T_23[7:0]) begin
        image_1_146 <= io_pixelVal_in_1_5;
      end else if (8'h92 == _T_20[7:0]) begin
        image_1_146 <= io_pixelVal_in_1_4;
      end else if (8'h92 == _T_17[7:0]) begin
        image_1_146 <= io_pixelVal_in_1_3;
      end else if (8'h92 == _T_14[7:0]) begin
        image_1_146 <= io_pixelVal_in_1_2;
      end else if (8'h92 == _T_11[7:0]) begin
        image_1_146 <= io_pixelVal_in_1_1;
      end else if (8'h92 == _T_7[7:0]) begin
        image_1_146 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_147 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h93 == _T_29[7:0]) begin
        image_1_147 <= io_pixelVal_in_1_7;
      end else if (8'h93 == _T_26[7:0]) begin
        image_1_147 <= io_pixelVal_in_1_6;
      end else if (8'h93 == _T_23[7:0]) begin
        image_1_147 <= io_pixelVal_in_1_5;
      end else if (8'h93 == _T_20[7:0]) begin
        image_1_147 <= io_pixelVal_in_1_4;
      end else if (8'h93 == _T_17[7:0]) begin
        image_1_147 <= io_pixelVal_in_1_3;
      end else if (8'h93 == _T_14[7:0]) begin
        image_1_147 <= io_pixelVal_in_1_2;
      end else if (8'h93 == _T_11[7:0]) begin
        image_1_147 <= io_pixelVal_in_1_1;
      end else if (8'h93 == _T_7[7:0]) begin
        image_1_147 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_148 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h94 == _T_29[7:0]) begin
        image_1_148 <= io_pixelVal_in_1_7;
      end else if (8'h94 == _T_26[7:0]) begin
        image_1_148 <= io_pixelVal_in_1_6;
      end else if (8'h94 == _T_23[7:0]) begin
        image_1_148 <= io_pixelVal_in_1_5;
      end else if (8'h94 == _T_20[7:0]) begin
        image_1_148 <= io_pixelVal_in_1_4;
      end else if (8'h94 == _T_17[7:0]) begin
        image_1_148 <= io_pixelVal_in_1_3;
      end else if (8'h94 == _T_14[7:0]) begin
        image_1_148 <= io_pixelVal_in_1_2;
      end else if (8'h94 == _T_11[7:0]) begin
        image_1_148 <= io_pixelVal_in_1_1;
      end else if (8'h94 == _T_7[7:0]) begin
        image_1_148 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_149 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h95 == _T_29[7:0]) begin
        image_1_149 <= io_pixelVal_in_1_7;
      end else if (8'h95 == _T_26[7:0]) begin
        image_1_149 <= io_pixelVal_in_1_6;
      end else if (8'h95 == _T_23[7:0]) begin
        image_1_149 <= io_pixelVal_in_1_5;
      end else if (8'h95 == _T_20[7:0]) begin
        image_1_149 <= io_pixelVal_in_1_4;
      end else if (8'h95 == _T_17[7:0]) begin
        image_1_149 <= io_pixelVal_in_1_3;
      end else if (8'h95 == _T_14[7:0]) begin
        image_1_149 <= io_pixelVal_in_1_2;
      end else if (8'h95 == _T_11[7:0]) begin
        image_1_149 <= io_pixelVal_in_1_1;
      end else if (8'h95 == _T_7[7:0]) begin
        image_1_149 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_150 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h96 == _T_29[7:0]) begin
        image_1_150 <= io_pixelVal_in_1_7;
      end else if (8'h96 == _T_26[7:0]) begin
        image_1_150 <= io_pixelVal_in_1_6;
      end else if (8'h96 == _T_23[7:0]) begin
        image_1_150 <= io_pixelVal_in_1_5;
      end else if (8'h96 == _T_20[7:0]) begin
        image_1_150 <= io_pixelVal_in_1_4;
      end else if (8'h96 == _T_17[7:0]) begin
        image_1_150 <= io_pixelVal_in_1_3;
      end else if (8'h96 == _T_14[7:0]) begin
        image_1_150 <= io_pixelVal_in_1_2;
      end else if (8'h96 == _T_11[7:0]) begin
        image_1_150 <= io_pixelVal_in_1_1;
      end else if (8'h96 == _T_7[7:0]) begin
        image_1_150 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_151 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h97 == _T_29[7:0]) begin
        image_1_151 <= io_pixelVal_in_1_7;
      end else if (8'h97 == _T_26[7:0]) begin
        image_1_151 <= io_pixelVal_in_1_6;
      end else if (8'h97 == _T_23[7:0]) begin
        image_1_151 <= io_pixelVal_in_1_5;
      end else if (8'h97 == _T_20[7:0]) begin
        image_1_151 <= io_pixelVal_in_1_4;
      end else if (8'h97 == _T_17[7:0]) begin
        image_1_151 <= io_pixelVal_in_1_3;
      end else if (8'h97 == _T_14[7:0]) begin
        image_1_151 <= io_pixelVal_in_1_2;
      end else if (8'h97 == _T_11[7:0]) begin
        image_1_151 <= io_pixelVal_in_1_1;
      end else if (8'h97 == _T_7[7:0]) begin
        image_1_151 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_152 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h98 == _T_29[7:0]) begin
        image_1_152 <= io_pixelVal_in_1_7;
      end else if (8'h98 == _T_26[7:0]) begin
        image_1_152 <= io_pixelVal_in_1_6;
      end else if (8'h98 == _T_23[7:0]) begin
        image_1_152 <= io_pixelVal_in_1_5;
      end else if (8'h98 == _T_20[7:0]) begin
        image_1_152 <= io_pixelVal_in_1_4;
      end else if (8'h98 == _T_17[7:0]) begin
        image_1_152 <= io_pixelVal_in_1_3;
      end else if (8'h98 == _T_14[7:0]) begin
        image_1_152 <= io_pixelVal_in_1_2;
      end else if (8'h98 == _T_11[7:0]) begin
        image_1_152 <= io_pixelVal_in_1_1;
      end else if (8'h98 == _T_7[7:0]) begin
        image_1_152 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_153 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h99 == _T_29[7:0]) begin
        image_1_153 <= io_pixelVal_in_1_7;
      end else if (8'h99 == _T_26[7:0]) begin
        image_1_153 <= io_pixelVal_in_1_6;
      end else if (8'h99 == _T_23[7:0]) begin
        image_1_153 <= io_pixelVal_in_1_5;
      end else if (8'h99 == _T_20[7:0]) begin
        image_1_153 <= io_pixelVal_in_1_4;
      end else if (8'h99 == _T_17[7:0]) begin
        image_1_153 <= io_pixelVal_in_1_3;
      end else if (8'h99 == _T_14[7:0]) begin
        image_1_153 <= io_pixelVal_in_1_2;
      end else if (8'h99 == _T_11[7:0]) begin
        image_1_153 <= io_pixelVal_in_1_1;
      end else if (8'h99 == _T_7[7:0]) begin
        image_1_153 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_154 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9a == _T_29[7:0]) begin
        image_1_154 <= io_pixelVal_in_1_7;
      end else if (8'h9a == _T_26[7:0]) begin
        image_1_154 <= io_pixelVal_in_1_6;
      end else if (8'h9a == _T_23[7:0]) begin
        image_1_154 <= io_pixelVal_in_1_5;
      end else if (8'h9a == _T_20[7:0]) begin
        image_1_154 <= io_pixelVal_in_1_4;
      end else if (8'h9a == _T_17[7:0]) begin
        image_1_154 <= io_pixelVal_in_1_3;
      end else if (8'h9a == _T_14[7:0]) begin
        image_1_154 <= io_pixelVal_in_1_2;
      end else if (8'h9a == _T_11[7:0]) begin
        image_1_154 <= io_pixelVal_in_1_1;
      end else if (8'h9a == _T_7[7:0]) begin
        image_1_154 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_155 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9b == _T_29[7:0]) begin
        image_1_155 <= io_pixelVal_in_1_7;
      end else if (8'h9b == _T_26[7:0]) begin
        image_1_155 <= io_pixelVal_in_1_6;
      end else if (8'h9b == _T_23[7:0]) begin
        image_1_155 <= io_pixelVal_in_1_5;
      end else if (8'h9b == _T_20[7:0]) begin
        image_1_155 <= io_pixelVal_in_1_4;
      end else if (8'h9b == _T_17[7:0]) begin
        image_1_155 <= io_pixelVal_in_1_3;
      end else if (8'h9b == _T_14[7:0]) begin
        image_1_155 <= io_pixelVal_in_1_2;
      end else if (8'h9b == _T_11[7:0]) begin
        image_1_155 <= io_pixelVal_in_1_1;
      end else if (8'h9b == _T_7[7:0]) begin
        image_1_155 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_156 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9c == _T_29[7:0]) begin
        image_1_156 <= io_pixelVal_in_1_7;
      end else if (8'h9c == _T_26[7:0]) begin
        image_1_156 <= io_pixelVal_in_1_6;
      end else if (8'h9c == _T_23[7:0]) begin
        image_1_156 <= io_pixelVal_in_1_5;
      end else if (8'h9c == _T_20[7:0]) begin
        image_1_156 <= io_pixelVal_in_1_4;
      end else if (8'h9c == _T_17[7:0]) begin
        image_1_156 <= io_pixelVal_in_1_3;
      end else if (8'h9c == _T_14[7:0]) begin
        image_1_156 <= io_pixelVal_in_1_2;
      end else if (8'h9c == _T_11[7:0]) begin
        image_1_156 <= io_pixelVal_in_1_1;
      end else if (8'h9c == _T_7[7:0]) begin
        image_1_156 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_157 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9d == _T_29[7:0]) begin
        image_1_157 <= io_pixelVal_in_1_7;
      end else if (8'h9d == _T_26[7:0]) begin
        image_1_157 <= io_pixelVal_in_1_6;
      end else if (8'h9d == _T_23[7:0]) begin
        image_1_157 <= io_pixelVal_in_1_5;
      end else if (8'h9d == _T_20[7:0]) begin
        image_1_157 <= io_pixelVal_in_1_4;
      end else if (8'h9d == _T_17[7:0]) begin
        image_1_157 <= io_pixelVal_in_1_3;
      end else if (8'h9d == _T_14[7:0]) begin
        image_1_157 <= io_pixelVal_in_1_2;
      end else if (8'h9d == _T_11[7:0]) begin
        image_1_157 <= io_pixelVal_in_1_1;
      end else if (8'h9d == _T_7[7:0]) begin
        image_1_157 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_158 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9e == _T_29[7:0]) begin
        image_1_158 <= io_pixelVal_in_1_7;
      end else if (8'h9e == _T_26[7:0]) begin
        image_1_158 <= io_pixelVal_in_1_6;
      end else if (8'h9e == _T_23[7:0]) begin
        image_1_158 <= io_pixelVal_in_1_5;
      end else if (8'h9e == _T_20[7:0]) begin
        image_1_158 <= io_pixelVal_in_1_4;
      end else if (8'h9e == _T_17[7:0]) begin
        image_1_158 <= io_pixelVal_in_1_3;
      end else if (8'h9e == _T_14[7:0]) begin
        image_1_158 <= io_pixelVal_in_1_2;
      end else if (8'h9e == _T_11[7:0]) begin
        image_1_158 <= io_pixelVal_in_1_1;
      end else if (8'h9e == _T_7[7:0]) begin
        image_1_158 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_159 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9f == _T_29[7:0]) begin
        image_1_159 <= io_pixelVal_in_1_7;
      end else if (8'h9f == _T_26[7:0]) begin
        image_1_159 <= io_pixelVal_in_1_6;
      end else if (8'h9f == _T_23[7:0]) begin
        image_1_159 <= io_pixelVal_in_1_5;
      end else if (8'h9f == _T_20[7:0]) begin
        image_1_159 <= io_pixelVal_in_1_4;
      end else if (8'h9f == _T_17[7:0]) begin
        image_1_159 <= io_pixelVal_in_1_3;
      end else if (8'h9f == _T_14[7:0]) begin
        image_1_159 <= io_pixelVal_in_1_2;
      end else if (8'h9f == _T_11[7:0]) begin
        image_1_159 <= io_pixelVal_in_1_1;
      end else if (8'h9f == _T_7[7:0]) begin
        image_1_159 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_160 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha0 == _T_29[7:0]) begin
        image_1_160 <= io_pixelVal_in_1_7;
      end else if (8'ha0 == _T_26[7:0]) begin
        image_1_160 <= io_pixelVal_in_1_6;
      end else if (8'ha0 == _T_23[7:0]) begin
        image_1_160 <= io_pixelVal_in_1_5;
      end else if (8'ha0 == _T_20[7:0]) begin
        image_1_160 <= io_pixelVal_in_1_4;
      end else if (8'ha0 == _T_17[7:0]) begin
        image_1_160 <= io_pixelVal_in_1_3;
      end else if (8'ha0 == _T_14[7:0]) begin
        image_1_160 <= io_pixelVal_in_1_2;
      end else if (8'ha0 == _T_11[7:0]) begin
        image_1_160 <= io_pixelVal_in_1_1;
      end else if (8'ha0 == _T_7[7:0]) begin
        image_1_160 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_161 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha1 == _T_29[7:0]) begin
        image_1_161 <= io_pixelVal_in_1_7;
      end else if (8'ha1 == _T_26[7:0]) begin
        image_1_161 <= io_pixelVal_in_1_6;
      end else if (8'ha1 == _T_23[7:0]) begin
        image_1_161 <= io_pixelVal_in_1_5;
      end else if (8'ha1 == _T_20[7:0]) begin
        image_1_161 <= io_pixelVal_in_1_4;
      end else if (8'ha1 == _T_17[7:0]) begin
        image_1_161 <= io_pixelVal_in_1_3;
      end else if (8'ha1 == _T_14[7:0]) begin
        image_1_161 <= io_pixelVal_in_1_2;
      end else if (8'ha1 == _T_11[7:0]) begin
        image_1_161 <= io_pixelVal_in_1_1;
      end else if (8'ha1 == _T_7[7:0]) begin
        image_1_161 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_162 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha2 == _T_29[7:0]) begin
        image_1_162 <= io_pixelVal_in_1_7;
      end else if (8'ha2 == _T_26[7:0]) begin
        image_1_162 <= io_pixelVal_in_1_6;
      end else if (8'ha2 == _T_23[7:0]) begin
        image_1_162 <= io_pixelVal_in_1_5;
      end else if (8'ha2 == _T_20[7:0]) begin
        image_1_162 <= io_pixelVal_in_1_4;
      end else if (8'ha2 == _T_17[7:0]) begin
        image_1_162 <= io_pixelVal_in_1_3;
      end else if (8'ha2 == _T_14[7:0]) begin
        image_1_162 <= io_pixelVal_in_1_2;
      end else if (8'ha2 == _T_11[7:0]) begin
        image_1_162 <= io_pixelVal_in_1_1;
      end else if (8'ha2 == _T_7[7:0]) begin
        image_1_162 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_163 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha3 == _T_29[7:0]) begin
        image_1_163 <= io_pixelVal_in_1_7;
      end else if (8'ha3 == _T_26[7:0]) begin
        image_1_163 <= io_pixelVal_in_1_6;
      end else if (8'ha3 == _T_23[7:0]) begin
        image_1_163 <= io_pixelVal_in_1_5;
      end else if (8'ha3 == _T_20[7:0]) begin
        image_1_163 <= io_pixelVal_in_1_4;
      end else if (8'ha3 == _T_17[7:0]) begin
        image_1_163 <= io_pixelVal_in_1_3;
      end else if (8'ha3 == _T_14[7:0]) begin
        image_1_163 <= io_pixelVal_in_1_2;
      end else if (8'ha3 == _T_11[7:0]) begin
        image_1_163 <= io_pixelVal_in_1_1;
      end else if (8'ha3 == _T_7[7:0]) begin
        image_1_163 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_164 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha4 == _T_29[7:0]) begin
        image_1_164 <= io_pixelVal_in_1_7;
      end else if (8'ha4 == _T_26[7:0]) begin
        image_1_164 <= io_pixelVal_in_1_6;
      end else if (8'ha4 == _T_23[7:0]) begin
        image_1_164 <= io_pixelVal_in_1_5;
      end else if (8'ha4 == _T_20[7:0]) begin
        image_1_164 <= io_pixelVal_in_1_4;
      end else if (8'ha4 == _T_17[7:0]) begin
        image_1_164 <= io_pixelVal_in_1_3;
      end else if (8'ha4 == _T_14[7:0]) begin
        image_1_164 <= io_pixelVal_in_1_2;
      end else if (8'ha4 == _T_11[7:0]) begin
        image_1_164 <= io_pixelVal_in_1_1;
      end else if (8'ha4 == _T_7[7:0]) begin
        image_1_164 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_165 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha5 == _T_29[7:0]) begin
        image_1_165 <= io_pixelVal_in_1_7;
      end else if (8'ha5 == _T_26[7:0]) begin
        image_1_165 <= io_pixelVal_in_1_6;
      end else if (8'ha5 == _T_23[7:0]) begin
        image_1_165 <= io_pixelVal_in_1_5;
      end else if (8'ha5 == _T_20[7:0]) begin
        image_1_165 <= io_pixelVal_in_1_4;
      end else if (8'ha5 == _T_17[7:0]) begin
        image_1_165 <= io_pixelVal_in_1_3;
      end else if (8'ha5 == _T_14[7:0]) begin
        image_1_165 <= io_pixelVal_in_1_2;
      end else if (8'ha5 == _T_11[7:0]) begin
        image_1_165 <= io_pixelVal_in_1_1;
      end else if (8'ha5 == _T_7[7:0]) begin
        image_1_165 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_166 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha6 == _T_29[7:0]) begin
        image_1_166 <= io_pixelVal_in_1_7;
      end else if (8'ha6 == _T_26[7:0]) begin
        image_1_166 <= io_pixelVal_in_1_6;
      end else if (8'ha6 == _T_23[7:0]) begin
        image_1_166 <= io_pixelVal_in_1_5;
      end else if (8'ha6 == _T_20[7:0]) begin
        image_1_166 <= io_pixelVal_in_1_4;
      end else if (8'ha6 == _T_17[7:0]) begin
        image_1_166 <= io_pixelVal_in_1_3;
      end else if (8'ha6 == _T_14[7:0]) begin
        image_1_166 <= io_pixelVal_in_1_2;
      end else if (8'ha6 == _T_11[7:0]) begin
        image_1_166 <= io_pixelVal_in_1_1;
      end else if (8'ha6 == _T_7[7:0]) begin
        image_1_166 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_167 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha7 == _T_29[7:0]) begin
        image_1_167 <= io_pixelVal_in_1_7;
      end else if (8'ha7 == _T_26[7:0]) begin
        image_1_167 <= io_pixelVal_in_1_6;
      end else if (8'ha7 == _T_23[7:0]) begin
        image_1_167 <= io_pixelVal_in_1_5;
      end else if (8'ha7 == _T_20[7:0]) begin
        image_1_167 <= io_pixelVal_in_1_4;
      end else if (8'ha7 == _T_17[7:0]) begin
        image_1_167 <= io_pixelVal_in_1_3;
      end else if (8'ha7 == _T_14[7:0]) begin
        image_1_167 <= io_pixelVal_in_1_2;
      end else if (8'ha7 == _T_11[7:0]) begin
        image_1_167 <= io_pixelVal_in_1_1;
      end else if (8'ha7 == _T_7[7:0]) begin
        image_1_167 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_168 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha8 == _T_29[7:0]) begin
        image_1_168 <= io_pixelVal_in_1_7;
      end else if (8'ha8 == _T_26[7:0]) begin
        image_1_168 <= io_pixelVal_in_1_6;
      end else if (8'ha8 == _T_23[7:0]) begin
        image_1_168 <= io_pixelVal_in_1_5;
      end else if (8'ha8 == _T_20[7:0]) begin
        image_1_168 <= io_pixelVal_in_1_4;
      end else if (8'ha8 == _T_17[7:0]) begin
        image_1_168 <= io_pixelVal_in_1_3;
      end else if (8'ha8 == _T_14[7:0]) begin
        image_1_168 <= io_pixelVal_in_1_2;
      end else if (8'ha8 == _T_11[7:0]) begin
        image_1_168 <= io_pixelVal_in_1_1;
      end else if (8'ha8 == _T_7[7:0]) begin
        image_1_168 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_169 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha9 == _T_29[7:0]) begin
        image_1_169 <= io_pixelVal_in_1_7;
      end else if (8'ha9 == _T_26[7:0]) begin
        image_1_169 <= io_pixelVal_in_1_6;
      end else if (8'ha9 == _T_23[7:0]) begin
        image_1_169 <= io_pixelVal_in_1_5;
      end else if (8'ha9 == _T_20[7:0]) begin
        image_1_169 <= io_pixelVal_in_1_4;
      end else if (8'ha9 == _T_17[7:0]) begin
        image_1_169 <= io_pixelVal_in_1_3;
      end else if (8'ha9 == _T_14[7:0]) begin
        image_1_169 <= io_pixelVal_in_1_2;
      end else if (8'ha9 == _T_11[7:0]) begin
        image_1_169 <= io_pixelVal_in_1_1;
      end else if (8'ha9 == _T_7[7:0]) begin
        image_1_169 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_170 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'haa == _T_29[7:0]) begin
        image_1_170 <= io_pixelVal_in_1_7;
      end else if (8'haa == _T_26[7:0]) begin
        image_1_170 <= io_pixelVal_in_1_6;
      end else if (8'haa == _T_23[7:0]) begin
        image_1_170 <= io_pixelVal_in_1_5;
      end else if (8'haa == _T_20[7:0]) begin
        image_1_170 <= io_pixelVal_in_1_4;
      end else if (8'haa == _T_17[7:0]) begin
        image_1_170 <= io_pixelVal_in_1_3;
      end else if (8'haa == _T_14[7:0]) begin
        image_1_170 <= io_pixelVal_in_1_2;
      end else if (8'haa == _T_11[7:0]) begin
        image_1_170 <= io_pixelVal_in_1_1;
      end else if (8'haa == _T_7[7:0]) begin
        image_1_170 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_171 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hab == _T_29[7:0]) begin
        image_1_171 <= io_pixelVal_in_1_7;
      end else if (8'hab == _T_26[7:0]) begin
        image_1_171 <= io_pixelVal_in_1_6;
      end else if (8'hab == _T_23[7:0]) begin
        image_1_171 <= io_pixelVal_in_1_5;
      end else if (8'hab == _T_20[7:0]) begin
        image_1_171 <= io_pixelVal_in_1_4;
      end else if (8'hab == _T_17[7:0]) begin
        image_1_171 <= io_pixelVal_in_1_3;
      end else if (8'hab == _T_14[7:0]) begin
        image_1_171 <= io_pixelVal_in_1_2;
      end else if (8'hab == _T_11[7:0]) begin
        image_1_171 <= io_pixelVal_in_1_1;
      end else if (8'hab == _T_7[7:0]) begin
        image_1_171 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_172 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hac == _T_29[7:0]) begin
        image_1_172 <= io_pixelVal_in_1_7;
      end else if (8'hac == _T_26[7:0]) begin
        image_1_172 <= io_pixelVal_in_1_6;
      end else if (8'hac == _T_23[7:0]) begin
        image_1_172 <= io_pixelVal_in_1_5;
      end else if (8'hac == _T_20[7:0]) begin
        image_1_172 <= io_pixelVal_in_1_4;
      end else if (8'hac == _T_17[7:0]) begin
        image_1_172 <= io_pixelVal_in_1_3;
      end else if (8'hac == _T_14[7:0]) begin
        image_1_172 <= io_pixelVal_in_1_2;
      end else if (8'hac == _T_11[7:0]) begin
        image_1_172 <= io_pixelVal_in_1_1;
      end else if (8'hac == _T_7[7:0]) begin
        image_1_172 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_173 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'had == _T_29[7:0]) begin
        image_1_173 <= io_pixelVal_in_1_7;
      end else if (8'had == _T_26[7:0]) begin
        image_1_173 <= io_pixelVal_in_1_6;
      end else if (8'had == _T_23[7:0]) begin
        image_1_173 <= io_pixelVal_in_1_5;
      end else if (8'had == _T_20[7:0]) begin
        image_1_173 <= io_pixelVal_in_1_4;
      end else if (8'had == _T_17[7:0]) begin
        image_1_173 <= io_pixelVal_in_1_3;
      end else if (8'had == _T_14[7:0]) begin
        image_1_173 <= io_pixelVal_in_1_2;
      end else if (8'had == _T_11[7:0]) begin
        image_1_173 <= io_pixelVal_in_1_1;
      end else if (8'had == _T_7[7:0]) begin
        image_1_173 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_174 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hae == _T_29[7:0]) begin
        image_1_174 <= io_pixelVal_in_1_7;
      end else if (8'hae == _T_26[7:0]) begin
        image_1_174 <= io_pixelVal_in_1_6;
      end else if (8'hae == _T_23[7:0]) begin
        image_1_174 <= io_pixelVal_in_1_5;
      end else if (8'hae == _T_20[7:0]) begin
        image_1_174 <= io_pixelVal_in_1_4;
      end else if (8'hae == _T_17[7:0]) begin
        image_1_174 <= io_pixelVal_in_1_3;
      end else if (8'hae == _T_14[7:0]) begin
        image_1_174 <= io_pixelVal_in_1_2;
      end else if (8'hae == _T_11[7:0]) begin
        image_1_174 <= io_pixelVal_in_1_1;
      end else if (8'hae == _T_7[7:0]) begin
        image_1_174 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_175 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'haf == _T_29[7:0]) begin
        image_1_175 <= io_pixelVal_in_1_7;
      end else if (8'haf == _T_26[7:0]) begin
        image_1_175 <= io_pixelVal_in_1_6;
      end else if (8'haf == _T_23[7:0]) begin
        image_1_175 <= io_pixelVal_in_1_5;
      end else if (8'haf == _T_20[7:0]) begin
        image_1_175 <= io_pixelVal_in_1_4;
      end else if (8'haf == _T_17[7:0]) begin
        image_1_175 <= io_pixelVal_in_1_3;
      end else if (8'haf == _T_14[7:0]) begin
        image_1_175 <= io_pixelVal_in_1_2;
      end else if (8'haf == _T_11[7:0]) begin
        image_1_175 <= io_pixelVal_in_1_1;
      end else if (8'haf == _T_7[7:0]) begin
        image_1_175 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_176 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb0 == _T_29[7:0]) begin
        image_1_176 <= io_pixelVal_in_1_7;
      end else if (8'hb0 == _T_26[7:0]) begin
        image_1_176 <= io_pixelVal_in_1_6;
      end else if (8'hb0 == _T_23[7:0]) begin
        image_1_176 <= io_pixelVal_in_1_5;
      end else if (8'hb0 == _T_20[7:0]) begin
        image_1_176 <= io_pixelVal_in_1_4;
      end else if (8'hb0 == _T_17[7:0]) begin
        image_1_176 <= io_pixelVal_in_1_3;
      end else if (8'hb0 == _T_14[7:0]) begin
        image_1_176 <= io_pixelVal_in_1_2;
      end else if (8'hb0 == _T_11[7:0]) begin
        image_1_176 <= io_pixelVal_in_1_1;
      end else if (8'hb0 == _T_7[7:0]) begin
        image_1_176 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_177 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb1 == _T_29[7:0]) begin
        image_1_177 <= io_pixelVal_in_1_7;
      end else if (8'hb1 == _T_26[7:0]) begin
        image_1_177 <= io_pixelVal_in_1_6;
      end else if (8'hb1 == _T_23[7:0]) begin
        image_1_177 <= io_pixelVal_in_1_5;
      end else if (8'hb1 == _T_20[7:0]) begin
        image_1_177 <= io_pixelVal_in_1_4;
      end else if (8'hb1 == _T_17[7:0]) begin
        image_1_177 <= io_pixelVal_in_1_3;
      end else if (8'hb1 == _T_14[7:0]) begin
        image_1_177 <= io_pixelVal_in_1_2;
      end else if (8'hb1 == _T_11[7:0]) begin
        image_1_177 <= io_pixelVal_in_1_1;
      end else if (8'hb1 == _T_7[7:0]) begin
        image_1_177 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_178 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb2 == _T_29[7:0]) begin
        image_1_178 <= io_pixelVal_in_1_7;
      end else if (8'hb2 == _T_26[7:0]) begin
        image_1_178 <= io_pixelVal_in_1_6;
      end else if (8'hb2 == _T_23[7:0]) begin
        image_1_178 <= io_pixelVal_in_1_5;
      end else if (8'hb2 == _T_20[7:0]) begin
        image_1_178 <= io_pixelVal_in_1_4;
      end else if (8'hb2 == _T_17[7:0]) begin
        image_1_178 <= io_pixelVal_in_1_3;
      end else if (8'hb2 == _T_14[7:0]) begin
        image_1_178 <= io_pixelVal_in_1_2;
      end else if (8'hb2 == _T_11[7:0]) begin
        image_1_178 <= io_pixelVal_in_1_1;
      end else if (8'hb2 == _T_7[7:0]) begin
        image_1_178 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_179 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb3 == _T_29[7:0]) begin
        image_1_179 <= io_pixelVal_in_1_7;
      end else if (8'hb3 == _T_26[7:0]) begin
        image_1_179 <= io_pixelVal_in_1_6;
      end else if (8'hb3 == _T_23[7:0]) begin
        image_1_179 <= io_pixelVal_in_1_5;
      end else if (8'hb3 == _T_20[7:0]) begin
        image_1_179 <= io_pixelVal_in_1_4;
      end else if (8'hb3 == _T_17[7:0]) begin
        image_1_179 <= io_pixelVal_in_1_3;
      end else if (8'hb3 == _T_14[7:0]) begin
        image_1_179 <= io_pixelVal_in_1_2;
      end else if (8'hb3 == _T_11[7:0]) begin
        image_1_179 <= io_pixelVal_in_1_1;
      end else if (8'hb3 == _T_7[7:0]) begin
        image_1_179 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_180 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb4 == _T_29[7:0]) begin
        image_1_180 <= io_pixelVal_in_1_7;
      end else if (8'hb4 == _T_26[7:0]) begin
        image_1_180 <= io_pixelVal_in_1_6;
      end else if (8'hb4 == _T_23[7:0]) begin
        image_1_180 <= io_pixelVal_in_1_5;
      end else if (8'hb4 == _T_20[7:0]) begin
        image_1_180 <= io_pixelVal_in_1_4;
      end else if (8'hb4 == _T_17[7:0]) begin
        image_1_180 <= io_pixelVal_in_1_3;
      end else if (8'hb4 == _T_14[7:0]) begin
        image_1_180 <= io_pixelVal_in_1_2;
      end else if (8'hb4 == _T_11[7:0]) begin
        image_1_180 <= io_pixelVal_in_1_1;
      end else if (8'hb4 == _T_7[7:0]) begin
        image_1_180 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_181 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb5 == _T_29[7:0]) begin
        image_1_181 <= io_pixelVal_in_1_7;
      end else if (8'hb5 == _T_26[7:0]) begin
        image_1_181 <= io_pixelVal_in_1_6;
      end else if (8'hb5 == _T_23[7:0]) begin
        image_1_181 <= io_pixelVal_in_1_5;
      end else if (8'hb5 == _T_20[7:0]) begin
        image_1_181 <= io_pixelVal_in_1_4;
      end else if (8'hb5 == _T_17[7:0]) begin
        image_1_181 <= io_pixelVal_in_1_3;
      end else if (8'hb5 == _T_14[7:0]) begin
        image_1_181 <= io_pixelVal_in_1_2;
      end else if (8'hb5 == _T_11[7:0]) begin
        image_1_181 <= io_pixelVal_in_1_1;
      end else if (8'hb5 == _T_7[7:0]) begin
        image_1_181 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_182 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb6 == _T_29[7:0]) begin
        image_1_182 <= io_pixelVal_in_1_7;
      end else if (8'hb6 == _T_26[7:0]) begin
        image_1_182 <= io_pixelVal_in_1_6;
      end else if (8'hb6 == _T_23[7:0]) begin
        image_1_182 <= io_pixelVal_in_1_5;
      end else if (8'hb6 == _T_20[7:0]) begin
        image_1_182 <= io_pixelVal_in_1_4;
      end else if (8'hb6 == _T_17[7:0]) begin
        image_1_182 <= io_pixelVal_in_1_3;
      end else if (8'hb6 == _T_14[7:0]) begin
        image_1_182 <= io_pixelVal_in_1_2;
      end else if (8'hb6 == _T_11[7:0]) begin
        image_1_182 <= io_pixelVal_in_1_1;
      end else if (8'hb6 == _T_7[7:0]) begin
        image_1_182 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_183 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb7 == _T_29[7:0]) begin
        image_1_183 <= io_pixelVal_in_1_7;
      end else if (8'hb7 == _T_26[7:0]) begin
        image_1_183 <= io_pixelVal_in_1_6;
      end else if (8'hb7 == _T_23[7:0]) begin
        image_1_183 <= io_pixelVal_in_1_5;
      end else if (8'hb7 == _T_20[7:0]) begin
        image_1_183 <= io_pixelVal_in_1_4;
      end else if (8'hb7 == _T_17[7:0]) begin
        image_1_183 <= io_pixelVal_in_1_3;
      end else if (8'hb7 == _T_14[7:0]) begin
        image_1_183 <= io_pixelVal_in_1_2;
      end else if (8'hb7 == _T_11[7:0]) begin
        image_1_183 <= io_pixelVal_in_1_1;
      end else if (8'hb7 == _T_7[7:0]) begin
        image_1_183 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_184 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb8 == _T_29[7:0]) begin
        image_1_184 <= io_pixelVal_in_1_7;
      end else if (8'hb8 == _T_26[7:0]) begin
        image_1_184 <= io_pixelVal_in_1_6;
      end else if (8'hb8 == _T_23[7:0]) begin
        image_1_184 <= io_pixelVal_in_1_5;
      end else if (8'hb8 == _T_20[7:0]) begin
        image_1_184 <= io_pixelVal_in_1_4;
      end else if (8'hb8 == _T_17[7:0]) begin
        image_1_184 <= io_pixelVal_in_1_3;
      end else if (8'hb8 == _T_14[7:0]) begin
        image_1_184 <= io_pixelVal_in_1_2;
      end else if (8'hb8 == _T_11[7:0]) begin
        image_1_184 <= io_pixelVal_in_1_1;
      end else if (8'hb8 == _T_7[7:0]) begin
        image_1_184 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_185 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb9 == _T_29[7:0]) begin
        image_1_185 <= io_pixelVal_in_1_7;
      end else if (8'hb9 == _T_26[7:0]) begin
        image_1_185 <= io_pixelVal_in_1_6;
      end else if (8'hb9 == _T_23[7:0]) begin
        image_1_185 <= io_pixelVal_in_1_5;
      end else if (8'hb9 == _T_20[7:0]) begin
        image_1_185 <= io_pixelVal_in_1_4;
      end else if (8'hb9 == _T_17[7:0]) begin
        image_1_185 <= io_pixelVal_in_1_3;
      end else if (8'hb9 == _T_14[7:0]) begin
        image_1_185 <= io_pixelVal_in_1_2;
      end else if (8'hb9 == _T_11[7:0]) begin
        image_1_185 <= io_pixelVal_in_1_1;
      end else if (8'hb9 == _T_7[7:0]) begin
        image_1_185 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_186 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hba == _T_29[7:0]) begin
        image_1_186 <= io_pixelVal_in_1_7;
      end else if (8'hba == _T_26[7:0]) begin
        image_1_186 <= io_pixelVal_in_1_6;
      end else if (8'hba == _T_23[7:0]) begin
        image_1_186 <= io_pixelVal_in_1_5;
      end else if (8'hba == _T_20[7:0]) begin
        image_1_186 <= io_pixelVal_in_1_4;
      end else if (8'hba == _T_17[7:0]) begin
        image_1_186 <= io_pixelVal_in_1_3;
      end else if (8'hba == _T_14[7:0]) begin
        image_1_186 <= io_pixelVal_in_1_2;
      end else if (8'hba == _T_11[7:0]) begin
        image_1_186 <= io_pixelVal_in_1_1;
      end else if (8'hba == _T_7[7:0]) begin
        image_1_186 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_187 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbb == _T_29[7:0]) begin
        image_1_187 <= io_pixelVal_in_1_7;
      end else if (8'hbb == _T_26[7:0]) begin
        image_1_187 <= io_pixelVal_in_1_6;
      end else if (8'hbb == _T_23[7:0]) begin
        image_1_187 <= io_pixelVal_in_1_5;
      end else if (8'hbb == _T_20[7:0]) begin
        image_1_187 <= io_pixelVal_in_1_4;
      end else if (8'hbb == _T_17[7:0]) begin
        image_1_187 <= io_pixelVal_in_1_3;
      end else if (8'hbb == _T_14[7:0]) begin
        image_1_187 <= io_pixelVal_in_1_2;
      end else if (8'hbb == _T_11[7:0]) begin
        image_1_187 <= io_pixelVal_in_1_1;
      end else if (8'hbb == _T_7[7:0]) begin
        image_1_187 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_188 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbc == _T_29[7:0]) begin
        image_1_188 <= io_pixelVal_in_1_7;
      end else if (8'hbc == _T_26[7:0]) begin
        image_1_188 <= io_pixelVal_in_1_6;
      end else if (8'hbc == _T_23[7:0]) begin
        image_1_188 <= io_pixelVal_in_1_5;
      end else if (8'hbc == _T_20[7:0]) begin
        image_1_188 <= io_pixelVal_in_1_4;
      end else if (8'hbc == _T_17[7:0]) begin
        image_1_188 <= io_pixelVal_in_1_3;
      end else if (8'hbc == _T_14[7:0]) begin
        image_1_188 <= io_pixelVal_in_1_2;
      end else if (8'hbc == _T_11[7:0]) begin
        image_1_188 <= io_pixelVal_in_1_1;
      end else if (8'hbc == _T_7[7:0]) begin
        image_1_188 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_189 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbd == _T_29[7:0]) begin
        image_1_189 <= io_pixelVal_in_1_7;
      end else if (8'hbd == _T_26[7:0]) begin
        image_1_189 <= io_pixelVal_in_1_6;
      end else if (8'hbd == _T_23[7:0]) begin
        image_1_189 <= io_pixelVal_in_1_5;
      end else if (8'hbd == _T_20[7:0]) begin
        image_1_189 <= io_pixelVal_in_1_4;
      end else if (8'hbd == _T_17[7:0]) begin
        image_1_189 <= io_pixelVal_in_1_3;
      end else if (8'hbd == _T_14[7:0]) begin
        image_1_189 <= io_pixelVal_in_1_2;
      end else if (8'hbd == _T_11[7:0]) begin
        image_1_189 <= io_pixelVal_in_1_1;
      end else if (8'hbd == _T_7[7:0]) begin
        image_1_189 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_190 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbe == _T_29[7:0]) begin
        image_1_190 <= io_pixelVal_in_1_7;
      end else if (8'hbe == _T_26[7:0]) begin
        image_1_190 <= io_pixelVal_in_1_6;
      end else if (8'hbe == _T_23[7:0]) begin
        image_1_190 <= io_pixelVal_in_1_5;
      end else if (8'hbe == _T_20[7:0]) begin
        image_1_190 <= io_pixelVal_in_1_4;
      end else if (8'hbe == _T_17[7:0]) begin
        image_1_190 <= io_pixelVal_in_1_3;
      end else if (8'hbe == _T_14[7:0]) begin
        image_1_190 <= io_pixelVal_in_1_2;
      end else if (8'hbe == _T_11[7:0]) begin
        image_1_190 <= io_pixelVal_in_1_1;
      end else if (8'hbe == _T_7[7:0]) begin
        image_1_190 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_191 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbf == _T_29[7:0]) begin
        image_1_191 <= io_pixelVal_in_1_7;
      end else if (8'hbf == _T_26[7:0]) begin
        image_1_191 <= io_pixelVal_in_1_6;
      end else if (8'hbf == _T_23[7:0]) begin
        image_1_191 <= io_pixelVal_in_1_5;
      end else if (8'hbf == _T_20[7:0]) begin
        image_1_191 <= io_pixelVal_in_1_4;
      end else if (8'hbf == _T_17[7:0]) begin
        image_1_191 <= io_pixelVal_in_1_3;
      end else if (8'hbf == _T_14[7:0]) begin
        image_1_191 <= io_pixelVal_in_1_2;
      end else if (8'hbf == _T_11[7:0]) begin
        image_1_191 <= io_pixelVal_in_1_1;
      end else if (8'hbf == _T_7[7:0]) begin
        image_1_191 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_2_0 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h0 == _T_29[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_7;
      end else if (8'h0 == _T_26[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_6;
      end else if (8'h0 == _T_23[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_5;
      end else if (8'h0 == _T_20[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_4;
      end else if (8'h0 == _T_17[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_3;
      end else if (8'h0 == _T_14[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_2;
      end else if (8'h0 == _T_11[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_1;
      end else if (8'h0 == _T_7[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_1 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1 == _T_29[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_7;
      end else if (8'h1 == _T_26[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_6;
      end else if (8'h1 == _T_23[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_5;
      end else if (8'h1 == _T_20[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_4;
      end else if (8'h1 == _T_17[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_3;
      end else if (8'h1 == _T_14[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_2;
      end else if (8'h1 == _T_11[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_1;
      end else if (8'h1 == _T_7[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_2 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2 == _T_29[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_7;
      end else if (8'h2 == _T_26[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_6;
      end else if (8'h2 == _T_23[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_5;
      end else if (8'h2 == _T_20[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_4;
      end else if (8'h2 == _T_17[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_3;
      end else if (8'h2 == _T_14[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_2;
      end else if (8'h2 == _T_11[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_1;
      end else if (8'h2 == _T_7[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_3 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3 == _T_29[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_7;
      end else if (8'h3 == _T_26[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_6;
      end else if (8'h3 == _T_23[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_5;
      end else if (8'h3 == _T_20[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_4;
      end else if (8'h3 == _T_17[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_3;
      end else if (8'h3 == _T_14[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_2;
      end else if (8'h3 == _T_11[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_1;
      end else if (8'h3 == _T_7[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_4 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4 == _T_29[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_7;
      end else if (8'h4 == _T_26[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_6;
      end else if (8'h4 == _T_23[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_5;
      end else if (8'h4 == _T_20[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_4;
      end else if (8'h4 == _T_17[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_3;
      end else if (8'h4 == _T_14[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_2;
      end else if (8'h4 == _T_11[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_1;
      end else if (8'h4 == _T_7[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_5 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5 == _T_29[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_7;
      end else if (8'h5 == _T_26[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_6;
      end else if (8'h5 == _T_23[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_5;
      end else if (8'h5 == _T_20[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_4;
      end else if (8'h5 == _T_17[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_3;
      end else if (8'h5 == _T_14[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_2;
      end else if (8'h5 == _T_11[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_1;
      end else if (8'h5 == _T_7[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_6 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6 == _T_29[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_7;
      end else if (8'h6 == _T_26[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_6;
      end else if (8'h6 == _T_23[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_5;
      end else if (8'h6 == _T_20[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_4;
      end else if (8'h6 == _T_17[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_3;
      end else if (8'h6 == _T_14[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_2;
      end else if (8'h6 == _T_11[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_1;
      end else if (8'h6 == _T_7[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_7 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7 == _T_29[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_7;
      end else if (8'h7 == _T_26[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_6;
      end else if (8'h7 == _T_23[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_5;
      end else if (8'h7 == _T_20[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_4;
      end else if (8'h7 == _T_17[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_3;
      end else if (8'h7 == _T_14[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_2;
      end else if (8'h7 == _T_11[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_1;
      end else if (8'h7 == _T_7[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_8 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8 == _T_29[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_7;
      end else if (8'h8 == _T_26[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_6;
      end else if (8'h8 == _T_23[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_5;
      end else if (8'h8 == _T_20[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_4;
      end else if (8'h8 == _T_17[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_3;
      end else if (8'h8 == _T_14[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_2;
      end else if (8'h8 == _T_11[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_1;
      end else if (8'h8 == _T_7[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_9 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9 == _T_29[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_7;
      end else if (8'h9 == _T_26[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_6;
      end else if (8'h9 == _T_23[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_5;
      end else if (8'h9 == _T_20[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_4;
      end else if (8'h9 == _T_17[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_3;
      end else if (8'h9 == _T_14[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_2;
      end else if (8'h9 == _T_11[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_1;
      end else if (8'h9 == _T_7[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_10 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha == _T_29[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_7;
      end else if (8'ha == _T_26[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_6;
      end else if (8'ha == _T_23[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_5;
      end else if (8'ha == _T_20[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_4;
      end else if (8'ha == _T_17[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_3;
      end else if (8'ha == _T_14[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_2;
      end else if (8'ha == _T_11[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_1;
      end else if (8'ha == _T_7[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_11 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb == _T_29[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_7;
      end else if (8'hb == _T_26[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_6;
      end else if (8'hb == _T_23[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_5;
      end else if (8'hb == _T_20[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_4;
      end else if (8'hb == _T_17[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_3;
      end else if (8'hb == _T_14[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_2;
      end else if (8'hb == _T_11[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_1;
      end else if (8'hb == _T_7[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_12 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc == _T_29[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_7;
      end else if (8'hc == _T_26[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_6;
      end else if (8'hc == _T_23[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_5;
      end else if (8'hc == _T_20[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_4;
      end else if (8'hc == _T_17[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_3;
      end else if (8'hc == _T_14[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_2;
      end else if (8'hc == _T_11[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_1;
      end else if (8'hc == _T_7[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_13 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd == _T_29[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_7;
      end else if (8'hd == _T_26[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_6;
      end else if (8'hd == _T_23[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_5;
      end else if (8'hd == _T_20[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_4;
      end else if (8'hd == _T_17[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_3;
      end else if (8'hd == _T_14[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_2;
      end else if (8'hd == _T_11[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_1;
      end else if (8'hd == _T_7[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_14 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he == _T_29[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_7;
      end else if (8'he == _T_26[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_6;
      end else if (8'he == _T_23[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_5;
      end else if (8'he == _T_20[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_4;
      end else if (8'he == _T_17[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_3;
      end else if (8'he == _T_14[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_2;
      end else if (8'he == _T_11[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_1;
      end else if (8'he == _T_7[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_15 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf == _T_29[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_7;
      end else if (8'hf == _T_26[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_6;
      end else if (8'hf == _T_23[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_5;
      end else if (8'hf == _T_20[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_4;
      end else if (8'hf == _T_17[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_3;
      end else if (8'hf == _T_14[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_2;
      end else if (8'hf == _T_11[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_1;
      end else if (8'hf == _T_7[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_16 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h10 == _T_29[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_7;
      end else if (8'h10 == _T_26[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_6;
      end else if (8'h10 == _T_23[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_5;
      end else if (8'h10 == _T_20[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_4;
      end else if (8'h10 == _T_17[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_3;
      end else if (8'h10 == _T_14[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_2;
      end else if (8'h10 == _T_11[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_1;
      end else if (8'h10 == _T_7[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_17 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h11 == _T_29[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_7;
      end else if (8'h11 == _T_26[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_6;
      end else if (8'h11 == _T_23[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_5;
      end else if (8'h11 == _T_20[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_4;
      end else if (8'h11 == _T_17[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_3;
      end else if (8'h11 == _T_14[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_2;
      end else if (8'h11 == _T_11[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_1;
      end else if (8'h11 == _T_7[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_18 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h12 == _T_29[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_7;
      end else if (8'h12 == _T_26[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_6;
      end else if (8'h12 == _T_23[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_5;
      end else if (8'h12 == _T_20[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_4;
      end else if (8'h12 == _T_17[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_3;
      end else if (8'h12 == _T_14[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_2;
      end else if (8'h12 == _T_11[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_1;
      end else if (8'h12 == _T_7[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_19 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h13 == _T_29[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_7;
      end else if (8'h13 == _T_26[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_6;
      end else if (8'h13 == _T_23[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_5;
      end else if (8'h13 == _T_20[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_4;
      end else if (8'h13 == _T_17[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_3;
      end else if (8'h13 == _T_14[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_2;
      end else if (8'h13 == _T_11[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_1;
      end else if (8'h13 == _T_7[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_20 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h14 == _T_29[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_7;
      end else if (8'h14 == _T_26[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_6;
      end else if (8'h14 == _T_23[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_5;
      end else if (8'h14 == _T_20[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_4;
      end else if (8'h14 == _T_17[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_3;
      end else if (8'h14 == _T_14[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_2;
      end else if (8'h14 == _T_11[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_1;
      end else if (8'h14 == _T_7[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_21 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h15 == _T_29[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_7;
      end else if (8'h15 == _T_26[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_6;
      end else if (8'h15 == _T_23[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_5;
      end else if (8'h15 == _T_20[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_4;
      end else if (8'h15 == _T_17[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_3;
      end else if (8'h15 == _T_14[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_2;
      end else if (8'h15 == _T_11[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_1;
      end else if (8'h15 == _T_7[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_22 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h16 == _T_29[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_7;
      end else if (8'h16 == _T_26[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_6;
      end else if (8'h16 == _T_23[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_5;
      end else if (8'h16 == _T_20[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_4;
      end else if (8'h16 == _T_17[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_3;
      end else if (8'h16 == _T_14[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_2;
      end else if (8'h16 == _T_11[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_1;
      end else if (8'h16 == _T_7[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_23 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h17 == _T_29[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_7;
      end else if (8'h17 == _T_26[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_6;
      end else if (8'h17 == _T_23[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_5;
      end else if (8'h17 == _T_20[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_4;
      end else if (8'h17 == _T_17[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_3;
      end else if (8'h17 == _T_14[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_2;
      end else if (8'h17 == _T_11[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_1;
      end else if (8'h17 == _T_7[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_24 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h18 == _T_29[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_7;
      end else if (8'h18 == _T_26[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_6;
      end else if (8'h18 == _T_23[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_5;
      end else if (8'h18 == _T_20[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_4;
      end else if (8'h18 == _T_17[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_3;
      end else if (8'h18 == _T_14[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_2;
      end else if (8'h18 == _T_11[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_1;
      end else if (8'h18 == _T_7[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_25 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h19 == _T_29[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_7;
      end else if (8'h19 == _T_26[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_6;
      end else if (8'h19 == _T_23[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_5;
      end else if (8'h19 == _T_20[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_4;
      end else if (8'h19 == _T_17[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_3;
      end else if (8'h19 == _T_14[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_2;
      end else if (8'h19 == _T_11[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_1;
      end else if (8'h19 == _T_7[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_26 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1a == _T_29[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_7;
      end else if (8'h1a == _T_26[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_6;
      end else if (8'h1a == _T_23[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_5;
      end else if (8'h1a == _T_20[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_4;
      end else if (8'h1a == _T_17[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_3;
      end else if (8'h1a == _T_14[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_2;
      end else if (8'h1a == _T_11[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_1;
      end else if (8'h1a == _T_7[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_27 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1b == _T_29[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_7;
      end else if (8'h1b == _T_26[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_6;
      end else if (8'h1b == _T_23[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_5;
      end else if (8'h1b == _T_20[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_4;
      end else if (8'h1b == _T_17[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_3;
      end else if (8'h1b == _T_14[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_2;
      end else if (8'h1b == _T_11[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_1;
      end else if (8'h1b == _T_7[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_28 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1c == _T_29[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_7;
      end else if (8'h1c == _T_26[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_6;
      end else if (8'h1c == _T_23[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_5;
      end else if (8'h1c == _T_20[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_4;
      end else if (8'h1c == _T_17[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_3;
      end else if (8'h1c == _T_14[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_2;
      end else if (8'h1c == _T_11[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_1;
      end else if (8'h1c == _T_7[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_29 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1d == _T_29[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_7;
      end else if (8'h1d == _T_26[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_6;
      end else if (8'h1d == _T_23[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_5;
      end else if (8'h1d == _T_20[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_4;
      end else if (8'h1d == _T_17[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_3;
      end else if (8'h1d == _T_14[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_2;
      end else if (8'h1d == _T_11[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_1;
      end else if (8'h1d == _T_7[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_30 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1e == _T_29[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_7;
      end else if (8'h1e == _T_26[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_6;
      end else if (8'h1e == _T_23[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_5;
      end else if (8'h1e == _T_20[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_4;
      end else if (8'h1e == _T_17[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_3;
      end else if (8'h1e == _T_14[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_2;
      end else if (8'h1e == _T_11[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_1;
      end else if (8'h1e == _T_7[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_31 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1f == _T_29[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_7;
      end else if (8'h1f == _T_26[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_6;
      end else if (8'h1f == _T_23[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_5;
      end else if (8'h1f == _T_20[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_4;
      end else if (8'h1f == _T_17[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_3;
      end else if (8'h1f == _T_14[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_2;
      end else if (8'h1f == _T_11[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_1;
      end else if (8'h1f == _T_7[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_32 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h20 == _T_29[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_7;
      end else if (8'h20 == _T_26[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_6;
      end else if (8'h20 == _T_23[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_5;
      end else if (8'h20 == _T_20[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_4;
      end else if (8'h20 == _T_17[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_3;
      end else if (8'h20 == _T_14[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_2;
      end else if (8'h20 == _T_11[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_1;
      end else if (8'h20 == _T_7[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_33 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h21 == _T_29[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_7;
      end else if (8'h21 == _T_26[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_6;
      end else if (8'h21 == _T_23[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_5;
      end else if (8'h21 == _T_20[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_4;
      end else if (8'h21 == _T_17[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_3;
      end else if (8'h21 == _T_14[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_2;
      end else if (8'h21 == _T_11[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_1;
      end else if (8'h21 == _T_7[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_34 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h22 == _T_29[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_7;
      end else if (8'h22 == _T_26[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_6;
      end else if (8'h22 == _T_23[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_5;
      end else if (8'h22 == _T_20[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_4;
      end else if (8'h22 == _T_17[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_3;
      end else if (8'h22 == _T_14[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_2;
      end else if (8'h22 == _T_11[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_1;
      end else if (8'h22 == _T_7[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_35 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h23 == _T_29[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_7;
      end else if (8'h23 == _T_26[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_6;
      end else if (8'h23 == _T_23[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_5;
      end else if (8'h23 == _T_20[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_4;
      end else if (8'h23 == _T_17[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_3;
      end else if (8'h23 == _T_14[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_2;
      end else if (8'h23 == _T_11[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_1;
      end else if (8'h23 == _T_7[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_36 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h24 == _T_29[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_7;
      end else if (8'h24 == _T_26[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_6;
      end else if (8'h24 == _T_23[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_5;
      end else if (8'h24 == _T_20[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_4;
      end else if (8'h24 == _T_17[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_3;
      end else if (8'h24 == _T_14[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_2;
      end else if (8'h24 == _T_11[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_1;
      end else if (8'h24 == _T_7[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_37 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h25 == _T_29[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_7;
      end else if (8'h25 == _T_26[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_6;
      end else if (8'h25 == _T_23[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_5;
      end else if (8'h25 == _T_20[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_4;
      end else if (8'h25 == _T_17[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_3;
      end else if (8'h25 == _T_14[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_2;
      end else if (8'h25 == _T_11[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_1;
      end else if (8'h25 == _T_7[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_38 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h26 == _T_29[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_7;
      end else if (8'h26 == _T_26[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_6;
      end else if (8'h26 == _T_23[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_5;
      end else if (8'h26 == _T_20[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_4;
      end else if (8'h26 == _T_17[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_3;
      end else if (8'h26 == _T_14[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_2;
      end else if (8'h26 == _T_11[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_1;
      end else if (8'h26 == _T_7[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_39 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h27 == _T_29[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_7;
      end else if (8'h27 == _T_26[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_6;
      end else if (8'h27 == _T_23[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_5;
      end else if (8'h27 == _T_20[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_4;
      end else if (8'h27 == _T_17[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_3;
      end else if (8'h27 == _T_14[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_2;
      end else if (8'h27 == _T_11[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_1;
      end else if (8'h27 == _T_7[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_40 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h28 == _T_29[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_7;
      end else if (8'h28 == _T_26[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_6;
      end else if (8'h28 == _T_23[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_5;
      end else if (8'h28 == _T_20[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_4;
      end else if (8'h28 == _T_17[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_3;
      end else if (8'h28 == _T_14[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_2;
      end else if (8'h28 == _T_11[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_1;
      end else if (8'h28 == _T_7[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_41 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h29 == _T_29[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_7;
      end else if (8'h29 == _T_26[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_6;
      end else if (8'h29 == _T_23[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_5;
      end else if (8'h29 == _T_20[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_4;
      end else if (8'h29 == _T_17[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_3;
      end else if (8'h29 == _T_14[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_2;
      end else if (8'h29 == _T_11[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_1;
      end else if (8'h29 == _T_7[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_42 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2a == _T_29[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_7;
      end else if (8'h2a == _T_26[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_6;
      end else if (8'h2a == _T_23[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_5;
      end else if (8'h2a == _T_20[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_4;
      end else if (8'h2a == _T_17[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_3;
      end else if (8'h2a == _T_14[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_2;
      end else if (8'h2a == _T_11[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_1;
      end else if (8'h2a == _T_7[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_43 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2b == _T_29[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_7;
      end else if (8'h2b == _T_26[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_6;
      end else if (8'h2b == _T_23[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_5;
      end else if (8'h2b == _T_20[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_4;
      end else if (8'h2b == _T_17[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_3;
      end else if (8'h2b == _T_14[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_2;
      end else if (8'h2b == _T_11[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_1;
      end else if (8'h2b == _T_7[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_44 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2c == _T_29[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_7;
      end else if (8'h2c == _T_26[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_6;
      end else if (8'h2c == _T_23[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_5;
      end else if (8'h2c == _T_20[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_4;
      end else if (8'h2c == _T_17[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_3;
      end else if (8'h2c == _T_14[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_2;
      end else if (8'h2c == _T_11[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_1;
      end else if (8'h2c == _T_7[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_45 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2d == _T_29[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_7;
      end else if (8'h2d == _T_26[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_6;
      end else if (8'h2d == _T_23[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_5;
      end else if (8'h2d == _T_20[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_4;
      end else if (8'h2d == _T_17[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_3;
      end else if (8'h2d == _T_14[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_2;
      end else if (8'h2d == _T_11[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_1;
      end else if (8'h2d == _T_7[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_46 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2e == _T_29[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_7;
      end else if (8'h2e == _T_26[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_6;
      end else if (8'h2e == _T_23[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_5;
      end else if (8'h2e == _T_20[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_4;
      end else if (8'h2e == _T_17[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_3;
      end else if (8'h2e == _T_14[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_2;
      end else if (8'h2e == _T_11[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_1;
      end else if (8'h2e == _T_7[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_47 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2f == _T_29[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_7;
      end else if (8'h2f == _T_26[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_6;
      end else if (8'h2f == _T_23[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_5;
      end else if (8'h2f == _T_20[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_4;
      end else if (8'h2f == _T_17[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_3;
      end else if (8'h2f == _T_14[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_2;
      end else if (8'h2f == _T_11[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_1;
      end else if (8'h2f == _T_7[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_48 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h30 == _T_29[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_7;
      end else if (8'h30 == _T_26[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_6;
      end else if (8'h30 == _T_23[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_5;
      end else if (8'h30 == _T_20[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_4;
      end else if (8'h30 == _T_17[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_3;
      end else if (8'h30 == _T_14[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_2;
      end else if (8'h30 == _T_11[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_1;
      end else if (8'h30 == _T_7[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_49 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h31 == _T_29[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_7;
      end else if (8'h31 == _T_26[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_6;
      end else if (8'h31 == _T_23[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_5;
      end else if (8'h31 == _T_20[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_4;
      end else if (8'h31 == _T_17[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_3;
      end else if (8'h31 == _T_14[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_2;
      end else if (8'h31 == _T_11[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_1;
      end else if (8'h31 == _T_7[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_50 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h32 == _T_29[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_7;
      end else if (8'h32 == _T_26[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_6;
      end else if (8'h32 == _T_23[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_5;
      end else if (8'h32 == _T_20[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_4;
      end else if (8'h32 == _T_17[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_3;
      end else if (8'h32 == _T_14[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_2;
      end else if (8'h32 == _T_11[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_1;
      end else if (8'h32 == _T_7[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_51 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h33 == _T_29[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_7;
      end else if (8'h33 == _T_26[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_6;
      end else if (8'h33 == _T_23[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_5;
      end else if (8'h33 == _T_20[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_4;
      end else if (8'h33 == _T_17[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_3;
      end else if (8'h33 == _T_14[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_2;
      end else if (8'h33 == _T_11[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_1;
      end else if (8'h33 == _T_7[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_52 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h34 == _T_29[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_7;
      end else if (8'h34 == _T_26[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_6;
      end else if (8'h34 == _T_23[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_5;
      end else if (8'h34 == _T_20[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_4;
      end else if (8'h34 == _T_17[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_3;
      end else if (8'h34 == _T_14[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_2;
      end else if (8'h34 == _T_11[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_1;
      end else if (8'h34 == _T_7[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_53 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h35 == _T_29[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_7;
      end else if (8'h35 == _T_26[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_6;
      end else if (8'h35 == _T_23[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_5;
      end else if (8'h35 == _T_20[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_4;
      end else if (8'h35 == _T_17[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_3;
      end else if (8'h35 == _T_14[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_2;
      end else if (8'h35 == _T_11[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_1;
      end else if (8'h35 == _T_7[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_54 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h36 == _T_29[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_7;
      end else if (8'h36 == _T_26[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_6;
      end else if (8'h36 == _T_23[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_5;
      end else if (8'h36 == _T_20[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_4;
      end else if (8'h36 == _T_17[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_3;
      end else if (8'h36 == _T_14[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_2;
      end else if (8'h36 == _T_11[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_1;
      end else if (8'h36 == _T_7[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_55 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h37 == _T_29[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_7;
      end else if (8'h37 == _T_26[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_6;
      end else if (8'h37 == _T_23[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_5;
      end else if (8'h37 == _T_20[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_4;
      end else if (8'h37 == _T_17[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_3;
      end else if (8'h37 == _T_14[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_2;
      end else if (8'h37 == _T_11[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_1;
      end else if (8'h37 == _T_7[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_56 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h38 == _T_29[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_7;
      end else if (8'h38 == _T_26[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_6;
      end else if (8'h38 == _T_23[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_5;
      end else if (8'h38 == _T_20[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_4;
      end else if (8'h38 == _T_17[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_3;
      end else if (8'h38 == _T_14[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_2;
      end else if (8'h38 == _T_11[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_1;
      end else if (8'h38 == _T_7[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_57 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h39 == _T_29[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_7;
      end else if (8'h39 == _T_26[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_6;
      end else if (8'h39 == _T_23[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_5;
      end else if (8'h39 == _T_20[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_4;
      end else if (8'h39 == _T_17[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_3;
      end else if (8'h39 == _T_14[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_2;
      end else if (8'h39 == _T_11[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_1;
      end else if (8'h39 == _T_7[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_58 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3a == _T_29[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_7;
      end else if (8'h3a == _T_26[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_6;
      end else if (8'h3a == _T_23[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_5;
      end else if (8'h3a == _T_20[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_4;
      end else if (8'h3a == _T_17[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_3;
      end else if (8'h3a == _T_14[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_2;
      end else if (8'h3a == _T_11[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_1;
      end else if (8'h3a == _T_7[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_59 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3b == _T_29[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_7;
      end else if (8'h3b == _T_26[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_6;
      end else if (8'h3b == _T_23[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_5;
      end else if (8'h3b == _T_20[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_4;
      end else if (8'h3b == _T_17[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_3;
      end else if (8'h3b == _T_14[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_2;
      end else if (8'h3b == _T_11[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_1;
      end else if (8'h3b == _T_7[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_60 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3c == _T_29[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_7;
      end else if (8'h3c == _T_26[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_6;
      end else if (8'h3c == _T_23[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_5;
      end else if (8'h3c == _T_20[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_4;
      end else if (8'h3c == _T_17[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_3;
      end else if (8'h3c == _T_14[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_2;
      end else if (8'h3c == _T_11[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_1;
      end else if (8'h3c == _T_7[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_61 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3d == _T_29[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_7;
      end else if (8'h3d == _T_26[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_6;
      end else if (8'h3d == _T_23[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_5;
      end else if (8'h3d == _T_20[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_4;
      end else if (8'h3d == _T_17[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_3;
      end else if (8'h3d == _T_14[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_2;
      end else if (8'h3d == _T_11[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_1;
      end else if (8'h3d == _T_7[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_62 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3e == _T_29[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_7;
      end else if (8'h3e == _T_26[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_6;
      end else if (8'h3e == _T_23[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_5;
      end else if (8'h3e == _T_20[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_4;
      end else if (8'h3e == _T_17[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_3;
      end else if (8'h3e == _T_14[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_2;
      end else if (8'h3e == _T_11[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_1;
      end else if (8'h3e == _T_7[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_63 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3f == _T_29[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_7;
      end else if (8'h3f == _T_26[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_6;
      end else if (8'h3f == _T_23[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_5;
      end else if (8'h3f == _T_20[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_4;
      end else if (8'h3f == _T_17[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_3;
      end else if (8'h3f == _T_14[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_2;
      end else if (8'h3f == _T_11[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_1;
      end else if (8'h3f == _T_7[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_64 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h40 == _T_29[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_7;
      end else if (8'h40 == _T_26[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_6;
      end else if (8'h40 == _T_23[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_5;
      end else if (8'h40 == _T_20[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_4;
      end else if (8'h40 == _T_17[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_3;
      end else if (8'h40 == _T_14[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_2;
      end else if (8'h40 == _T_11[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_1;
      end else if (8'h40 == _T_7[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_65 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h41 == _T_29[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_7;
      end else if (8'h41 == _T_26[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_6;
      end else if (8'h41 == _T_23[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_5;
      end else if (8'h41 == _T_20[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_4;
      end else if (8'h41 == _T_17[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_3;
      end else if (8'h41 == _T_14[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_2;
      end else if (8'h41 == _T_11[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_1;
      end else if (8'h41 == _T_7[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_66 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h42 == _T_29[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_7;
      end else if (8'h42 == _T_26[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_6;
      end else if (8'h42 == _T_23[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_5;
      end else if (8'h42 == _T_20[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_4;
      end else if (8'h42 == _T_17[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_3;
      end else if (8'h42 == _T_14[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_2;
      end else if (8'h42 == _T_11[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_1;
      end else if (8'h42 == _T_7[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_67 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h43 == _T_29[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_7;
      end else if (8'h43 == _T_26[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_6;
      end else if (8'h43 == _T_23[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_5;
      end else if (8'h43 == _T_20[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_4;
      end else if (8'h43 == _T_17[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_3;
      end else if (8'h43 == _T_14[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_2;
      end else if (8'h43 == _T_11[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_1;
      end else if (8'h43 == _T_7[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_68 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h44 == _T_29[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_7;
      end else if (8'h44 == _T_26[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_6;
      end else if (8'h44 == _T_23[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_5;
      end else if (8'h44 == _T_20[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_4;
      end else if (8'h44 == _T_17[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_3;
      end else if (8'h44 == _T_14[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_2;
      end else if (8'h44 == _T_11[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_1;
      end else if (8'h44 == _T_7[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_69 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h45 == _T_29[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_7;
      end else if (8'h45 == _T_26[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_6;
      end else if (8'h45 == _T_23[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_5;
      end else if (8'h45 == _T_20[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_4;
      end else if (8'h45 == _T_17[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_3;
      end else if (8'h45 == _T_14[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_2;
      end else if (8'h45 == _T_11[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_1;
      end else if (8'h45 == _T_7[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_70 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h46 == _T_29[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_7;
      end else if (8'h46 == _T_26[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_6;
      end else if (8'h46 == _T_23[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_5;
      end else if (8'h46 == _T_20[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_4;
      end else if (8'h46 == _T_17[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_3;
      end else if (8'h46 == _T_14[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_2;
      end else if (8'h46 == _T_11[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_1;
      end else if (8'h46 == _T_7[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_71 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h47 == _T_29[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_7;
      end else if (8'h47 == _T_26[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_6;
      end else if (8'h47 == _T_23[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_5;
      end else if (8'h47 == _T_20[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_4;
      end else if (8'h47 == _T_17[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_3;
      end else if (8'h47 == _T_14[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_2;
      end else if (8'h47 == _T_11[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_1;
      end else if (8'h47 == _T_7[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_72 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h48 == _T_29[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_7;
      end else if (8'h48 == _T_26[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_6;
      end else if (8'h48 == _T_23[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_5;
      end else if (8'h48 == _T_20[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_4;
      end else if (8'h48 == _T_17[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_3;
      end else if (8'h48 == _T_14[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_2;
      end else if (8'h48 == _T_11[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_1;
      end else if (8'h48 == _T_7[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_73 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h49 == _T_29[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_7;
      end else if (8'h49 == _T_26[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_6;
      end else if (8'h49 == _T_23[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_5;
      end else if (8'h49 == _T_20[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_4;
      end else if (8'h49 == _T_17[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_3;
      end else if (8'h49 == _T_14[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_2;
      end else if (8'h49 == _T_11[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_1;
      end else if (8'h49 == _T_7[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_74 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4a == _T_29[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_7;
      end else if (8'h4a == _T_26[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_6;
      end else if (8'h4a == _T_23[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_5;
      end else if (8'h4a == _T_20[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_4;
      end else if (8'h4a == _T_17[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_3;
      end else if (8'h4a == _T_14[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_2;
      end else if (8'h4a == _T_11[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_1;
      end else if (8'h4a == _T_7[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_75 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4b == _T_29[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_7;
      end else if (8'h4b == _T_26[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_6;
      end else if (8'h4b == _T_23[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_5;
      end else if (8'h4b == _T_20[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_4;
      end else if (8'h4b == _T_17[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_3;
      end else if (8'h4b == _T_14[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_2;
      end else if (8'h4b == _T_11[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_1;
      end else if (8'h4b == _T_7[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_76 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4c == _T_29[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_7;
      end else if (8'h4c == _T_26[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_6;
      end else if (8'h4c == _T_23[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_5;
      end else if (8'h4c == _T_20[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_4;
      end else if (8'h4c == _T_17[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_3;
      end else if (8'h4c == _T_14[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_2;
      end else if (8'h4c == _T_11[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_1;
      end else if (8'h4c == _T_7[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_77 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4d == _T_29[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_7;
      end else if (8'h4d == _T_26[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_6;
      end else if (8'h4d == _T_23[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_5;
      end else if (8'h4d == _T_20[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_4;
      end else if (8'h4d == _T_17[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_3;
      end else if (8'h4d == _T_14[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_2;
      end else if (8'h4d == _T_11[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_1;
      end else if (8'h4d == _T_7[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_78 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4e == _T_29[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_7;
      end else if (8'h4e == _T_26[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_6;
      end else if (8'h4e == _T_23[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_5;
      end else if (8'h4e == _T_20[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_4;
      end else if (8'h4e == _T_17[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_3;
      end else if (8'h4e == _T_14[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_2;
      end else if (8'h4e == _T_11[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_1;
      end else if (8'h4e == _T_7[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_79 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4f == _T_29[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_7;
      end else if (8'h4f == _T_26[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_6;
      end else if (8'h4f == _T_23[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_5;
      end else if (8'h4f == _T_20[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_4;
      end else if (8'h4f == _T_17[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_3;
      end else if (8'h4f == _T_14[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_2;
      end else if (8'h4f == _T_11[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_1;
      end else if (8'h4f == _T_7[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_80 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h50 == _T_29[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_7;
      end else if (8'h50 == _T_26[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_6;
      end else if (8'h50 == _T_23[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_5;
      end else if (8'h50 == _T_20[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_4;
      end else if (8'h50 == _T_17[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_3;
      end else if (8'h50 == _T_14[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_2;
      end else if (8'h50 == _T_11[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_1;
      end else if (8'h50 == _T_7[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_81 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h51 == _T_29[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_7;
      end else if (8'h51 == _T_26[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_6;
      end else if (8'h51 == _T_23[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_5;
      end else if (8'h51 == _T_20[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_4;
      end else if (8'h51 == _T_17[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_3;
      end else if (8'h51 == _T_14[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_2;
      end else if (8'h51 == _T_11[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_1;
      end else if (8'h51 == _T_7[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_82 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h52 == _T_29[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_7;
      end else if (8'h52 == _T_26[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_6;
      end else if (8'h52 == _T_23[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_5;
      end else if (8'h52 == _T_20[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_4;
      end else if (8'h52 == _T_17[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_3;
      end else if (8'h52 == _T_14[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_2;
      end else if (8'h52 == _T_11[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_1;
      end else if (8'h52 == _T_7[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_83 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h53 == _T_29[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_7;
      end else if (8'h53 == _T_26[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_6;
      end else if (8'h53 == _T_23[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_5;
      end else if (8'h53 == _T_20[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_4;
      end else if (8'h53 == _T_17[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_3;
      end else if (8'h53 == _T_14[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_2;
      end else if (8'h53 == _T_11[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_1;
      end else if (8'h53 == _T_7[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_84 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h54 == _T_29[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_7;
      end else if (8'h54 == _T_26[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_6;
      end else if (8'h54 == _T_23[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_5;
      end else if (8'h54 == _T_20[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_4;
      end else if (8'h54 == _T_17[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_3;
      end else if (8'h54 == _T_14[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_2;
      end else if (8'h54 == _T_11[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_1;
      end else if (8'h54 == _T_7[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_85 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h55 == _T_29[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_7;
      end else if (8'h55 == _T_26[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_6;
      end else if (8'h55 == _T_23[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_5;
      end else if (8'h55 == _T_20[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_4;
      end else if (8'h55 == _T_17[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_3;
      end else if (8'h55 == _T_14[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_2;
      end else if (8'h55 == _T_11[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_1;
      end else if (8'h55 == _T_7[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_86 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h56 == _T_29[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_7;
      end else if (8'h56 == _T_26[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_6;
      end else if (8'h56 == _T_23[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_5;
      end else if (8'h56 == _T_20[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_4;
      end else if (8'h56 == _T_17[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_3;
      end else if (8'h56 == _T_14[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_2;
      end else if (8'h56 == _T_11[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_1;
      end else if (8'h56 == _T_7[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_87 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h57 == _T_29[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_7;
      end else if (8'h57 == _T_26[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_6;
      end else if (8'h57 == _T_23[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_5;
      end else if (8'h57 == _T_20[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_4;
      end else if (8'h57 == _T_17[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_3;
      end else if (8'h57 == _T_14[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_2;
      end else if (8'h57 == _T_11[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_1;
      end else if (8'h57 == _T_7[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_88 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h58 == _T_29[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_7;
      end else if (8'h58 == _T_26[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_6;
      end else if (8'h58 == _T_23[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_5;
      end else if (8'h58 == _T_20[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_4;
      end else if (8'h58 == _T_17[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_3;
      end else if (8'h58 == _T_14[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_2;
      end else if (8'h58 == _T_11[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_1;
      end else if (8'h58 == _T_7[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_89 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h59 == _T_29[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_7;
      end else if (8'h59 == _T_26[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_6;
      end else if (8'h59 == _T_23[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_5;
      end else if (8'h59 == _T_20[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_4;
      end else if (8'h59 == _T_17[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_3;
      end else if (8'h59 == _T_14[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_2;
      end else if (8'h59 == _T_11[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_1;
      end else if (8'h59 == _T_7[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_90 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5a == _T_29[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_7;
      end else if (8'h5a == _T_26[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_6;
      end else if (8'h5a == _T_23[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_5;
      end else if (8'h5a == _T_20[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_4;
      end else if (8'h5a == _T_17[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_3;
      end else if (8'h5a == _T_14[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_2;
      end else if (8'h5a == _T_11[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_1;
      end else if (8'h5a == _T_7[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_91 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5b == _T_29[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_7;
      end else if (8'h5b == _T_26[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_6;
      end else if (8'h5b == _T_23[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_5;
      end else if (8'h5b == _T_20[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_4;
      end else if (8'h5b == _T_17[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_3;
      end else if (8'h5b == _T_14[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_2;
      end else if (8'h5b == _T_11[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_1;
      end else if (8'h5b == _T_7[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_92 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5c == _T_29[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_7;
      end else if (8'h5c == _T_26[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_6;
      end else if (8'h5c == _T_23[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_5;
      end else if (8'h5c == _T_20[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_4;
      end else if (8'h5c == _T_17[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_3;
      end else if (8'h5c == _T_14[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_2;
      end else if (8'h5c == _T_11[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_1;
      end else if (8'h5c == _T_7[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_93 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5d == _T_29[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_7;
      end else if (8'h5d == _T_26[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_6;
      end else if (8'h5d == _T_23[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_5;
      end else if (8'h5d == _T_20[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_4;
      end else if (8'h5d == _T_17[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_3;
      end else if (8'h5d == _T_14[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_2;
      end else if (8'h5d == _T_11[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_1;
      end else if (8'h5d == _T_7[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_94 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5e == _T_29[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_7;
      end else if (8'h5e == _T_26[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_6;
      end else if (8'h5e == _T_23[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_5;
      end else if (8'h5e == _T_20[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_4;
      end else if (8'h5e == _T_17[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_3;
      end else if (8'h5e == _T_14[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_2;
      end else if (8'h5e == _T_11[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_1;
      end else if (8'h5e == _T_7[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_95 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5f == _T_29[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_7;
      end else if (8'h5f == _T_26[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_6;
      end else if (8'h5f == _T_23[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_5;
      end else if (8'h5f == _T_20[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_4;
      end else if (8'h5f == _T_17[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_3;
      end else if (8'h5f == _T_14[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_2;
      end else if (8'h5f == _T_11[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_1;
      end else if (8'h5f == _T_7[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_96 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h60 == _T_29[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_7;
      end else if (8'h60 == _T_26[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_6;
      end else if (8'h60 == _T_23[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_5;
      end else if (8'h60 == _T_20[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_4;
      end else if (8'h60 == _T_17[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_3;
      end else if (8'h60 == _T_14[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_2;
      end else if (8'h60 == _T_11[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_1;
      end else if (8'h60 == _T_7[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_97 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h61 == _T_29[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_7;
      end else if (8'h61 == _T_26[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_6;
      end else if (8'h61 == _T_23[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_5;
      end else if (8'h61 == _T_20[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_4;
      end else if (8'h61 == _T_17[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_3;
      end else if (8'h61 == _T_14[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_2;
      end else if (8'h61 == _T_11[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_1;
      end else if (8'h61 == _T_7[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_98 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h62 == _T_29[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_7;
      end else if (8'h62 == _T_26[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_6;
      end else if (8'h62 == _T_23[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_5;
      end else if (8'h62 == _T_20[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_4;
      end else if (8'h62 == _T_17[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_3;
      end else if (8'h62 == _T_14[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_2;
      end else if (8'h62 == _T_11[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_1;
      end else if (8'h62 == _T_7[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_99 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h63 == _T_29[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_7;
      end else if (8'h63 == _T_26[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_6;
      end else if (8'h63 == _T_23[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_5;
      end else if (8'h63 == _T_20[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_4;
      end else if (8'h63 == _T_17[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_3;
      end else if (8'h63 == _T_14[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_2;
      end else if (8'h63 == _T_11[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_1;
      end else if (8'h63 == _T_7[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_100 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h64 == _T_29[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_7;
      end else if (8'h64 == _T_26[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_6;
      end else if (8'h64 == _T_23[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_5;
      end else if (8'h64 == _T_20[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_4;
      end else if (8'h64 == _T_17[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_3;
      end else if (8'h64 == _T_14[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_2;
      end else if (8'h64 == _T_11[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_1;
      end else if (8'h64 == _T_7[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_101 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h65 == _T_29[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_7;
      end else if (8'h65 == _T_26[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_6;
      end else if (8'h65 == _T_23[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_5;
      end else if (8'h65 == _T_20[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_4;
      end else if (8'h65 == _T_17[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_3;
      end else if (8'h65 == _T_14[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_2;
      end else if (8'h65 == _T_11[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_1;
      end else if (8'h65 == _T_7[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_102 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h66 == _T_29[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_7;
      end else if (8'h66 == _T_26[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_6;
      end else if (8'h66 == _T_23[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_5;
      end else if (8'h66 == _T_20[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_4;
      end else if (8'h66 == _T_17[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_3;
      end else if (8'h66 == _T_14[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_2;
      end else if (8'h66 == _T_11[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_1;
      end else if (8'h66 == _T_7[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_103 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h67 == _T_29[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_7;
      end else if (8'h67 == _T_26[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_6;
      end else if (8'h67 == _T_23[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_5;
      end else if (8'h67 == _T_20[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_4;
      end else if (8'h67 == _T_17[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_3;
      end else if (8'h67 == _T_14[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_2;
      end else if (8'h67 == _T_11[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_1;
      end else if (8'h67 == _T_7[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_104 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h68 == _T_29[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_7;
      end else if (8'h68 == _T_26[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_6;
      end else if (8'h68 == _T_23[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_5;
      end else if (8'h68 == _T_20[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_4;
      end else if (8'h68 == _T_17[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_3;
      end else if (8'h68 == _T_14[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_2;
      end else if (8'h68 == _T_11[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_1;
      end else if (8'h68 == _T_7[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_105 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h69 == _T_29[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_7;
      end else if (8'h69 == _T_26[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_6;
      end else if (8'h69 == _T_23[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_5;
      end else if (8'h69 == _T_20[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_4;
      end else if (8'h69 == _T_17[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_3;
      end else if (8'h69 == _T_14[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_2;
      end else if (8'h69 == _T_11[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_1;
      end else if (8'h69 == _T_7[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_106 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6a == _T_29[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_7;
      end else if (8'h6a == _T_26[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_6;
      end else if (8'h6a == _T_23[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_5;
      end else if (8'h6a == _T_20[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_4;
      end else if (8'h6a == _T_17[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_3;
      end else if (8'h6a == _T_14[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_2;
      end else if (8'h6a == _T_11[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_1;
      end else if (8'h6a == _T_7[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_107 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6b == _T_29[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_7;
      end else if (8'h6b == _T_26[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_6;
      end else if (8'h6b == _T_23[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_5;
      end else if (8'h6b == _T_20[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_4;
      end else if (8'h6b == _T_17[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_3;
      end else if (8'h6b == _T_14[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_2;
      end else if (8'h6b == _T_11[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_1;
      end else if (8'h6b == _T_7[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_108 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6c == _T_29[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_7;
      end else if (8'h6c == _T_26[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_6;
      end else if (8'h6c == _T_23[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_5;
      end else if (8'h6c == _T_20[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_4;
      end else if (8'h6c == _T_17[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_3;
      end else if (8'h6c == _T_14[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_2;
      end else if (8'h6c == _T_11[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_1;
      end else if (8'h6c == _T_7[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_109 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6d == _T_29[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_7;
      end else if (8'h6d == _T_26[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_6;
      end else if (8'h6d == _T_23[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_5;
      end else if (8'h6d == _T_20[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_4;
      end else if (8'h6d == _T_17[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_3;
      end else if (8'h6d == _T_14[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_2;
      end else if (8'h6d == _T_11[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_1;
      end else if (8'h6d == _T_7[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_110 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6e == _T_29[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_7;
      end else if (8'h6e == _T_26[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_6;
      end else if (8'h6e == _T_23[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_5;
      end else if (8'h6e == _T_20[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_4;
      end else if (8'h6e == _T_17[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_3;
      end else if (8'h6e == _T_14[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_2;
      end else if (8'h6e == _T_11[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_1;
      end else if (8'h6e == _T_7[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_111 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6f == _T_29[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_7;
      end else if (8'h6f == _T_26[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_6;
      end else if (8'h6f == _T_23[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_5;
      end else if (8'h6f == _T_20[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_4;
      end else if (8'h6f == _T_17[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_3;
      end else if (8'h6f == _T_14[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_2;
      end else if (8'h6f == _T_11[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_1;
      end else if (8'h6f == _T_7[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_112 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h70 == _T_29[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_7;
      end else if (8'h70 == _T_26[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_6;
      end else if (8'h70 == _T_23[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_5;
      end else if (8'h70 == _T_20[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_4;
      end else if (8'h70 == _T_17[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_3;
      end else if (8'h70 == _T_14[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_2;
      end else if (8'h70 == _T_11[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_1;
      end else if (8'h70 == _T_7[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_113 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h71 == _T_29[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_7;
      end else if (8'h71 == _T_26[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_6;
      end else if (8'h71 == _T_23[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_5;
      end else if (8'h71 == _T_20[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_4;
      end else if (8'h71 == _T_17[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_3;
      end else if (8'h71 == _T_14[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_2;
      end else if (8'h71 == _T_11[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_1;
      end else if (8'h71 == _T_7[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_114 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h72 == _T_29[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_7;
      end else if (8'h72 == _T_26[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_6;
      end else if (8'h72 == _T_23[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_5;
      end else if (8'h72 == _T_20[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_4;
      end else if (8'h72 == _T_17[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_3;
      end else if (8'h72 == _T_14[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_2;
      end else if (8'h72 == _T_11[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_1;
      end else if (8'h72 == _T_7[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_115 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h73 == _T_29[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_7;
      end else if (8'h73 == _T_26[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_6;
      end else if (8'h73 == _T_23[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_5;
      end else if (8'h73 == _T_20[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_4;
      end else if (8'h73 == _T_17[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_3;
      end else if (8'h73 == _T_14[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_2;
      end else if (8'h73 == _T_11[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_1;
      end else if (8'h73 == _T_7[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_116 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h74 == _T_29[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_7;
      end else if (8'h74 == _T_26[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_6;
      end else if (8'h74 == _T_23[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_5;
      end else if (8'h74 == _T_20[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_4;
      end else if (8'h74 == _T_17[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_3;
      end else if (8'h74 == _T_14[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_2;
      end else if (8'h74 == _T_11[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_1;
      end else if (8'h74 == _T_7[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_117 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h75 == _T_29[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_7;
      end else if (8'h75 == _T_26[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_6;
      end else if (8'h75 == _T_23[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_5;
      end else if (8'h75 == _T_20[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_4;
      end else if (8'h75 == _T_17[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_3;
      end else if (8'h75 == _T_14[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_2;
      end else if (8'h75 == _T_11[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_1;
      end else if (8'h75 == _T_7[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_118 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h76 == _T_29[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_7;
      end else if (8'h76 == _T_26[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_6;
      end else if (8'h76 == _T_23[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_5;
      end else if (8'h76 == _T_20[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_4;
      end else if (8'h76 == _T_17[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_3;
      end else if (8'h76 == _T_14[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_2;
      end else if (8'h76 == _T_11[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_1;
      end else if (8'h76 == _T_7[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_119 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h77 == _T_29[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_7;
      end else if (8'h77 == _T_26[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_6;
      end else if (8'h77 == _T_23[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_5;
      end else if (8'h77 == _T_20[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_4;
      end else if (8'h77 == _T_17[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_3;
      end else if (8'h77 == _T_14[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_2;
      end else if (8'h77 == _T_11[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_1;
      end else if (8'h77 == _T_7[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_120 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h78 == _T_29[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_7;
      end else if (8'h78 == _T_26[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_6;
      end else if (8'h78 == _T_23[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_5;
      end else if (8'h78 == _T_20[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_4;
      end else if (8'h78 == _T_17[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_3;
      end else if (8'h78 == _T_14[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_2;
      end else if (8'h78 == _T_11[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_1;
      end else if (8'h78 == _T_7[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_121 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h79 == _T_29[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_7;
      end else if (8'h79 == _T_26[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_6;
      end else if (8'h79 == _T_23[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_5;
      end else if (8'h79 == _T_20[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_4;
      end else if (8'h79 == _T_17[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_3;
      end else if (8'h79 == _T_14[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_2;
      end else if (8'h79 == _T_11[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_1;
      end else if (8'h79 == _T_7[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_122 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7a == _T_29[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_7;
      end else if (8'h7a == _T_26[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_6;
      end else if (8'h7a == _T_23[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_5;
      end else if (8'h7a == _T_20[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_4;
      end else if (8'h7a == _T_17[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_3;
      end else if (8'h7a == _T_14[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_2;
      end else if (8'h7a == _T_11[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_1;
      end else if (8'h7a == _T_7[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_123 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7b == _T_29[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_7;
      end else if (8'h7b == _T_26[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_6;
      end else if (8'h7b == _T_23[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_5;
      end else if (8'h7b == _T_20[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_4;
      end else if (8'h7b == _T_17[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_3;
      end else if (8'h7b == _T_14[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_2;
      end else if (8'h7b == _T_11[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_1;
      end else if (8'h7b == _T_7[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_124 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7c == _T_29[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_7;
      end else if (8'h7c == _T_26[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_6;
      end else if (8'h7c == _T_23[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_5;
      end else if (8'h7c == _T_20[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_4;
      end else if (8'h7c == _T_17[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_3;
      end else if (8'h7c == _T_14[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_2;
      end else if (8'h7c == _T_11[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_1;
      end else if (8'h7c == _T_7[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_125 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7d == _T_29[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_7;
      end else if (8'h7d == _T_26[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_6;
      end else if (8'h7d == _T_23[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_5;
      end else if (8'h7d == _T_20[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_4;
      end else if (8'h7d == _T_17[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_3;
      end else if (8'h7d == _T_14[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_2;
      end else if (8'h7d == _T_11[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_1;
      end else if (8'h7d == _T_7[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_126 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7e == _T_29[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_7;
      end else if (8'h7e == _T_26[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_6;
      end else if (8'h7e == _T_23[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_5;
      end else if (8'h7e == _T_20[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_4;
      end else if (8'h7e == _T_17[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_3;
      end else if (8'h7e == _T_14[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_2;
      end else if (8'h7e == _T_11[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_1;
      end else if (8'h7e == _T_7[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_127 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7f == _T_29[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_7;
      end else if (8'h7f == _T_26[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_6;
      end else if (8'h7f == _T_23[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_5;
      end else if (8'h7f == _T_20[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_4;
      end else if (8'h7f == _T_17[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_3;
      end else if (8'h7f == _T_14[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_2;
      end else if (8'h7f == _T_11[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_1;
      end else if (8'h7f == _T_7[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_128 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h80 == _T_29[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_7;
      end else if (8'h80 == _T_26[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_6;
      end else if (8'h80 == _T_23[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_5;
      end else if (8'h80 == _T_20[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_4;
      end else if (8'h80 == _T_17[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_3;
      end else if (8'h80 == _T_14[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_2;
      end else if (8'h80 == _T_11[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_1;
      end else if (8'h80 == _T_7[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_129 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h81 == _T_29[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_7;
      end else if (8'h81 == _T_26[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_6;
      end else if (8'h81 == _T_23[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_5;
      end else if (8'h81 == _T_20[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_4;
      end else if (8'h81 == _T_17[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_3;
      end else if (8'h81 == _T_14[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_2;
      end else if (8'h81 == _T_11[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_1;
      end else if (8'h81 == _T_7[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_130 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h82 == _T_29[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_7;
      end else if (8'h82 == _T_26[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_6;
      end else if (8'h82 == _T_23[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_5;
      end else if (8'h82 == _T_20[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_4;
      end else if (8'h82 == _T_17[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_3;
      end else if (8'h82 == _T_14[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_2;
      end else if (8'h82 == _T_11[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_1;
      end else if (8'h82 == _T_7[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_131 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h83 == _T_29[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_7;
      end else if (8'h83 == _T_26[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_6;
      end else if (8'h83 == _T_23[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_5;
      end else if (8'h83 == _T_20[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_4;
      end else if (8'h83 == _T_17[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_3;
      end else if (8'h83 == _T_14[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_2;
      end else if (8'h83 == _T_11[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_1;
      end else if (8'h83 == _T_7[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_132 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h84 == _T_29[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_7;
      end else if (8'h84 == _T_26[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_6;
      end else if (8'h84 == _T_23[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_5;
      end else if (8'h84 == _T_20[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_4;
      end else if (8'h84 == _T_17[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_3;
      end else if (8'h84 == _T_14[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_2;
      end else if (8'h84 == _T_11[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_1;
      end else if (8'h84 == _T_7[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_133 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h85 == _T_29[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_7;
      end else if (8'h85 == _T_26[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_6;
      end else if (8'h85 == _T_23[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_5;
      end else if (8'h85 == _T_20[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_4;
      end else if (8'h85 == _T_17[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_3;
      end else if (8'h85 == _T_14[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_2;
      end else if (8'h85 == _T_11[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_1;
      end else if (8'h85 == _T_7[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_134 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h86 == _T_29[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_7;
      end else if (8'h86 == _T_26[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_6;
      end else if (8'h86 == _T_23[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_5;
      end else if (8'h86 == _T_20[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_4;
      end else if (8'h86 == _T_17[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_3;
      end else if (8'h86 == _T_14[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_2;
      end else if (8'h86 == _T_11[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_1;
      end else if (8'h86 == _T_7[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_135 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h87 == _T_29[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_7;
      end else if (8'h87 == _T_26[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_6;
      end else if (8'h87 == _T_23[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_5;
      end else if (8'h87 == _T_20[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_4;
      end else if (8'h87 == _T_17[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_3;
      end else if (8'h87 == _T_14[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_2;
      end else if (8'h87 == _T_11[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_1;
      end else if (8'h87 == _T_7[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_136 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h88 == _T_29[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_7;
      end else if (8'h88 == _T_26[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_6;
      end else if (8'h88 == _T_23[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_5;
      end else if (8'h88 == _T_20[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_4;
      end else if (8'h88 == _T_17[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_3;
      end else if (8'h88 == _T_14[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_2;
      end else if (8'h88 == _T_11[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_1;
      end else if (8'h88 == _T_7[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_137 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h89 == _T_29[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_7;
      end else if (8'h89 == _T_26[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_6;
      end else if (8'h89 == _T_23[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_5;
      end else if (8'h89 == _T_20[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_4;
      end else if (8'h89 == _T_17[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_3;
      end else if (8'h89 == _T_14[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_2;
      end else if (8'h89 == _T_11[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_1;
      end else if (8'h89 == _T_7[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_138 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8a == _T_29[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_7;
      end else if (8'h8a == _T_26[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_6;
      end else if (8'h8a == _T_23[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_5;
      end else if (8'h8a == _T_20[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_4;
      end else if (8'h8a == _T_17[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_3;
      end else if (8'h8a == _T_14[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_2;
      end else if (8'h8a == _T_11[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_1;
      end else if (8'h8a == _T_7[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_139 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8b == _T_29[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_7;
      end else if (8'h8b == _T_26[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_6;
      end else if (8'h8b == _T_23[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_5;
      end else if (8'h8b == _T_20[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_4;
      end else if (8'h8b == _T_17[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_3;
      end else if (8'h8b == _T_14[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_2;
      end else if (8'h8b == _T_11[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_1;
      end else if (8'h8b == _T_7[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_140 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8c == _T_29[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_7;
      end else if (8'h8c == _T_26[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_6;
      end else if (8'h8c == _T_23[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_5;
      end else if (8'h8c == _T_20[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_4;
      end else if (8'h8c == _T_17[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_3;
      end else if (8'h8c == _T_14[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_2;
      end else if (8'h8c == _T_11[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_1;
      end else if (8'h8c == _T_7[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_141 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8d == _T_29[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_7;
      end else if (8'h8d == _T_26[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_6;
      end else if (8'h8d == _T_23[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_5;
      end else if (8'h8d == _T_20[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_4;
      end else if (8'h8d == _T_17[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_3;
      end else if (8'h8d == _T_14[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_2;
      end else if (8'h8d == _T_11[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_1;
      end else if (8'h8d == _T_7[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_142 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8e == _T_29[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_7;
      end else if (8'h8e == _T_26[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_6;
      end else if (8'h8e == _T_23[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_5;
      end else if (8'h8e == _T_20[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_4;
      end else if (8'h8e == _T_17[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_3;
      end else if (8'h8e == _T_14[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_2;
      end else if (8'h8e == _T_11[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_1;
      end else if (8'h8e == _T_7[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_143 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8f == _T_29[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_7;
      end else if (8'h8f == _T_26[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_6;
      end else if (8'h8f == _T_23[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_5;
      end else if (8'h8f == _T_20[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_4;
      end else if (8'h8f == _T_17[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_3;
      end else if (8'h8f == _T_14[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_2;
      end else if (8'h8f == _T_11[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_1;
      end else if (8'h8f == _T_7[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_144 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h90 == _T_29[7:0]) begin
        image_2_144 <= io_pixelVal_in_2_7;
      end else if (8'h90 == _T_26[7:0]) begin
        image_2_144 <= io_pixelVal_in_2_6;
      end else if (8'h90 == _T_23[7:0]) begin
        image_2_144 <= io_pixelVal_in_2_5;
      end else if (8'h90 == _T_20[7:0]) begin
        image_2_144 <= io_pixelVal_in_2_4;
      end else if (8'h90 == _T_17[7:0]) begin
        image_2_144 <= io_pixelVal_in_2_3;
      end else if (8'h90 == _T_14[7:0]) begin
        image_2_144 <= io_pixelVal_in_2_2;
      end else if (8'h90 == _T_11[7:0]) begin
        image_2_144 <= io_pixelVal_in_2_1;
      end else if (8'h90 == _T_7[7:0]) begin
        image_2_144 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_145 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h91 == _T_29[7:0]) begin
        image_2_145 <= io_pixelVal_in_2_7;
      end else if (8'h91 == _T_26[7:0]) begin
        image_2_145 <= io_pixelVal_in_2_6;
      end else if (8'h91 == _T_23[7:0]) begin
        image_2_145 <= io_pixelVal_in_2_5;
      end else if (8'h91 == _T_20[7:0]) begin
        image_2_145 <= io_pixelVal_in_2_4;
      end else if (8'h91 == _T_17[7:0]) begin
        image_2_145 <= io_pixelVal_in_2_3;
      end else if (8'h91 == _T_14[7:0]) begin
        image_2_145 <= io_pixelVal_in_2_2;
      end else if (8'h91 == _T_11[7:0]) begin
        image_2_145 <= io_pixelVal_in_2_1;
      end else if (8'h91 == _T_7[7:0]) begin
        image_2_145 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_146 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h92 == _T_29[7:0]) begin
        image_2_146 <= io_pixelVal_in_2_7;
      end else if (8'h92 == _T_26[7:0]) begin
        image_2_146 <= io_pixelVal_in_2_6;
      end else if (8'h92 == _T_23[7:0]) begin
        image_2_146 <= io_pixelVal_in_2_5;
      end else if (8'h92 == _T_20[7:0]) begin
        image_2_146 <= io_pixelVal_in_2_4;
      end else if (8'h92 == _T_17[7:0]) begin
        image_2_146 <= io_pixelVal_in_2_3;
      end else if (8'h92 == _T_14[7:0]) begin
        image_2_146 <= io_pixelVal_in_2_2;
      end else if (8'h92 == _T_11[7:0]) begin
        image_2_146 <= io_pixelVal_in_2_1;
      end else if (8'h92 == _T_7[7:0]) begin
        image_2_146 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_147 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h93 == _T_29[7:0]) begin
        image_2_147 <= io_pixelVal_in_2_7;
      end else if (8'h93 == _T_26[7:0]) begin
        image_2_147 <= io_pixelVal_in_2_6;
      end else if (8'h93 == _T_23[7:0]) begin
        image_2_147 <= io_pixelVal_in_2_5;
      end else if (8'h93 == _T_20[7:0]) begin
        image_2_147 <= io_pixelVal_in_2_4;
      end else if (8'h93 == _T_17[7:0]) begin
        image_2_147 <= io_pixelVal_in_2_3;
      end else if (8'h93 == _T_14[7:0]) begin
        image_2_147 <= io_pixelVal_in_2_2;
      end else if (8'h93 == _T_11[7:0]) begin
        image_2_147 <= io_pixelVal_in_2_1;
      end else if (8'h93 == _T_7[7:0]) begin
        image_2_147 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_148 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h94 == _T_29[7:0]) begin
        image_2_148 <= io_pixelVal_in_2_7;
      end else if (8'h94 == _T_26[7:0]) begin
        image_2_148 <= io_pixelVal_in_2_6;
      end else if (8'h94 == _T_23[7:0]) begin
        image_2_148 <= io_pixelVal_in_2_5;
      end else if (8'h94 == _T_20[7:0]) begin
        image_2_148 <= io_pixelVal_in_2_4;
      end else if (8'h94 == _T_17[7:0]) begin
        image_2_148 <= io_pixelVal_in_2_3;
      end else if (8'h94 == _T_14[7:0]) begin
        image_2_148 <= io_pixelVal_in_2_2;
      end else if (8'h94 == _T_11[7:0]) begin
        image_2_148 <= io_pixelVal_in_2_1;
      end else if (8'h94 == _T_7[7:0]) begin
        image_2_148 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_149 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h95 == _T_29[7:0]) begin
        image_2_149 <= io_pixelVal_in_2_7;
      end else if (8'h95 == _T_26[7:0]) begin
        image_2_149 <= io_pixelVal_in_2_6;
      end else if (8'h95 == _T_23[7:0]) begin
        image_2_149 <= io_pixelVal_in_2_5;
      end else if (8'h95 == _T_20[7:0]) begin
        image_2_149 <= io_pixelVal_in_2_4;
      end else if (8'h95 == _T_17[7:0]) begin
        image_2_149 <= io_pixelVal_in_2_3;
      end else if (8'h95 == _T_14[7:0]) begin
        image_2_149 <= io_pixelVal_in_2_2;
      end else if (8'h95 == _T_11[7:0]) begin
        image_2_149 <= io_pixelVal_in_2_1;
      end else if (8'h95 == _T_7[7:0]) begin
        image_2_149 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_150 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h96 == _T_29[7:0]) begin
        image_2_150 <= io_pixelVal_in_2_7;
      end else if (8'h96 == _T_26[7:0]) begin
        image_2_150 <= io_pixelVal_in_2_6;
      end else if (8'h96 == _T_23[7:0]) begin
        image_2_150 <= io_pixelVal_in_2_5;
      end else if (8'h96 == _T_20[7:0]) begin
        image_2_150 <= io_pixelVal_in_2_4;
      end else if (8'h96 == _T_17[7:0]) begin
        image_2_150 <= io_pixelVal_in_2_3;
      end else if (8'h96 == _T_14[7:0]) begin
        image_2_150 <= io_pixelVal_in_2_2;
      end else if (8'h96 == _T_11[7:0]) begin
        image_2_150 <= io_pixelVal_in_2_1;
      end else if (8'h96 == _T_7[7:0]) begin
        image_2_150 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_151 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h97 == _T_29[7:0]) begin
        image_2_151 <= io_pixelVal_in_2_7;
      end else if (8'h97 == _T_26[7:0]) begin
        image_2_151 <= io_pixelVal_in_2_6;
      end else if (8'h97 == _T_23[7:0]) begin
        image_2_151 <= io_pixelVal_in_2_5;
      end else if (8'h97 == _T_20[7:0]) begin
        image_2_151 <= io_pixelVal_in_2_4;
      end else if (8'h97 == _T_17[7:0]) begin
        image_2_151 <= io_pixelVal_in_2_3;
      end else if (8'h97 == _T_14[7:0]) begin
        image_2_151 <= io_pixelVal_in_2_2;
      end else if (8'h97 == _T_11[7:0]) begin
        image_2_151 <= io_pixelVal_in_2_1;
      end else if (8'h97 == _T_7[7:0]) begin
        image_2_151 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_152 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h98 == _T_29[7:0]) begin
        image_2_152 <= io_pixelVal_in_2_7;
      end else if (8'h98 == _T_26[7:0]) begin
        image_2_152 <= io_pixelVal_in_2_6;
      end else if (8'h98 == _T_23[7:0]) begin
        image_2_152 <= io_pixelVal_in_2_5;
      end else if (8'h98 == _T_20[7:0]) begin
        image_2_152 <= io_pixelVal_in_2_4;
      end else if (8'h98 == _T_17[7:0]) begin
        image_2_152 <= io_pixelVal_in_2_3;
      end else if (8'h98 == _T_14[7:0]) begin
        image_2_152 <= io_pixelVal_in_2_2;
      end else if (8'h98 == _T_11[7:0]) begin
        image_2_152 <= io_pixelVal_in_2_1;
      end else if (8'h98 == _T_7[7:0]) begin
        image_2_152 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_153 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h99 == _T_29[7:0]) begin
        image_2_153 <= io_pixelVal_in_2_7;
      end else if (8'h99 == _T_26[7:0]) begin
        image_2_153 <= io_pixelVal_in_2_6;
      end else if (8'h99 == _T_23[7:0]) begin
        image_2_153 <= io_pixelVal_in_2_5;
      end else if (8'h99 == _T_20[7:0]) begin
        image_2_153 <= io_pixelVal_in_2_4;
      end else if (8'h99 == _T_17[7:0]) begin
        image_2_153 <= io_pixelVal_in_2_3;
      end else if (8'h99 == _T_14[7:0]) begin
        image_2_153 <= io_pixelVal_in_2_2;
      end else if (8'h99 == _T_11[7:0]) begin
        image_2_153 <= io_pixelVal_in_2_1;
      end else if (8'h99 == _T_7[7:0]) begin
        image_2_153 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_154 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9a == _T_29[7:0]) begin
        image_2_154 <= io_pixelVal_in_2_7;
      end else if (8'h9a == _T_26[7:0]) begin
        image_2_154 <= io_pixelVal_in_2_6;
      end else if (8'h9a == _T_23[7:0]) begin
        image_2_154 <= io_pixelVal_in_2_5;
      end else if (8'h9a == _T_20[7:0]) begin
        image_2_154 <= io_pixelVal_in_2_4;
      end else if (8'h9a == _T_17[7:0]) begin
        image_2_154 <= io_pixelVal_in_2_3;
      end else if (8'h9a == _T_14[7:0]) begin
        image_2_154 <= io_pixelVal_in_2_2;
      end else if (8'h9a == _T_11[7:0]) begin
        image_2_154 <= io_pixelVal_in_2_1;
      end else if (8'h9a == _T_7[7:0]) begin
        image_2_154 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_155 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9b == _T_29[7:0]) begin
        image_2_155 <= io_pixelVal_in_2_7;
      end else if (8'h9b == _T_26[7:0]) begin
        image_2_155 <= io_pixelVal_in_2_6;
      end else if (8'h9b == _T_23[7:0]) begin
        image_2_155 <= io_pixelVal_in_2_5;
      end else if (8'h9b == _T_20[7:0]) begin
        image_2_155 <= io_pixelVal_in_2_4;
      end else if (8'h9b == _T_17[7:0]) begin
        image_2_155 <= io_pixelVal_in_2_3;
      end else if (8'h9b == _T_14[7:0]) begin
        image_2_155 <= io_pixelVal_in_2_2;
      end else if (8'h9b == _T_11[7:0]) begin
        image_2_155 <= io_pixelVal_in_2_1;
      end else if (8'h9b == _T_7[7:0]) begin
        image_2_155 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_156 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9c == _T_29[7:0]) begin
        image_2_156 <= io_pixelVal_in_2_7;
      end else if (8'h9c == _T_26[7:0]) begin
        image_2_156 <= io_pixelVal_in_2_6;
      end else if (8'h9c == _T_23[7:0]) begin
        image_2_156 <= io_pixelVal_in_2_5;
      end else if (8'h9c == _T_20[7:0]) begin
        image_2_156 <= io_pixelVal_in_2_4;
      end else if (8'h9c == _T_17[7:0]) begin
        image_2_156 <= io_pixelVal_in_2_3;
      end else if (8'h9c == _T_14[7:0]) begin
        image_2_156 <= io_pixelVal_in_2_2;
      end else if (8'h9c == _T_11[7:0]) begin
        image_2_156 <= io_pixelVal_in_2_1;
      end else if (8'h9c == _T_7[7:0]) begin
        image_2_156 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_157 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9d == _T_29[7:0]) begin
        image_2_157 <= io_pixelVal_in_2_7;
      end else if (8'h9d == _T_26[7:0]) begin
        image_2_157 <= io_pixelVal_in_2_6;
      end else if (8'h9d == _T_23[7:0]) begin
        image_2_157 <= io_pixelVal_in_2_5;
      end else if (8'h9d == _T_20[7:0]) begin
        image_2_157 <= io_pixelVal_in_2_4;
      end else if (8'h9d == _T_17[7:0]) begin
        image_2_157 <= io_pixelVal_in_2_3;
      end else if (8'h9d == _T_14[7:0]) begin
        image_2_157 <= io_pixelVal_in_2_2;
      end else if (8'h9d == _T_11[7:0]) begin
        image_2_157 <= io_pixelVal_in_2_1;
      end else if (8'h9d == _T_7[7:0]) begin
        image_2_157 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_158 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9e == _T_29[7:0]) begin
        image_2_158 <= io_pixelVal_in_2_7;
      end else if (8'h9e == _T_26[7:0]) begin
        image_2_158 <= io_pixelVal_in_2_6;
      end else if (8'h9e == _T_23[7:0]) begin
        image_2_158 <= io_pixelVal_in_2_5;
      end else if (8'h9e == _T_20[7:0]) begin
        image_2_158 <= io_pixelVal_in_2_4;
      end else if (8'h9e == _T_17[7:0]) begin
        image_2_158 <= io_pixelVal_in_2_3;
      end else if (8'h9e == _T_14[7:0]) begin
        image_2_158 <= io_pixelVal_in_2_2;
      end else if (8'h9e == _T_11[7:0]) begin
        image_2_158 <= io_pixelVal_in_2_1;
      end else if (8'h9e == _T_7[7:0]) begin
        image_2_158 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_159 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9f == _T_29[7:0]) begin
        image_2_159 <= io_pixelVal_in_2_7;
      end else if (8'h9f == _T_26[7:0]) begin
        image_2_159 <= io_pixelVal_in_2_6;
      end else if (8'h9f == _T_23[7:0]) begin
        image_2_159 <= io_pixelVal_in_2_5;
      end else if (8'h9f == _T_20[7:0]) begin
        image_2_159 <= io_pixelVal_in_2_4;
      end else if (8'h9f == _T_17[7:0]) begin
        image_2_159 <= io_pixelVal_in_2_3;
      end else if (8'h9f == _T_14[7:0]) begin
        image_2_159 <= io_pixelVal_in_2_2;
      end else if (8'h9f == _T_11[7:0]) begin
        image_2_159 <= io_pixelVal_in_2_1;
      end else if (8'h9f == _T_7[7:0]) begin
        image_2_159 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_160 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha0 == _T_29[7:0]) begin
        image_2_160 <= io_pixelVal_in_2_7;
      end else if (8'ha0 == _T_26[7:0]) begin
        image_2_160 <= io_pixelVal_in_2_6;
      end else if (8'ha0 == _T_23[7:0]) begin
        image_2_160 <= io_pixelVal_in_2_5;
      end else if (8'ha0 == _T_20[7:0]) begin
        image_2_160 <= io_pixelVal_in_2_4;
      end else if (8'ha0 == _T_17[7:0]) begin
        image_2_160 <= io_pixelVal_in_2_3;
      end else if (8'ha0 == _T_14[7:0]) begin
        image_2_160 <= io_pixelVal_in_2_2;
      end else if (8'ha0 == _T_11[7:0]) begin
        image_2_160 <= io_pixelVal_in_2_1;
      end else if (8'ha0 == _T_7[7:0]) begin
        image_2_160 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_161 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha1 == _T_29[7:0]) begin
        image_2_161 <= io_pixelVal_in_2_7;
      end else if (8'ha1 == _T_26[7:0]) begin
        image_2_161 <= io_pixelVal_in_2_6;
      end else if (8'ha1 == _T_23[7:0]) begin
        image_2_161 <= io_pixelVal_in_2_5;
      end else if (8'ha1 == _T_20[7:0]) begin
        image_2_161 <= io_pixelVal_in_2_4;
      end else if (8'ha1 == _T_17[7:0]) begin
        image_2_161 <= io_pixelVal_in_2_3;
      end else if (8'ha1 == _T_14[7:0]) begin
        image_2_161 <= io_pixelVal_in_2_2;
      end else if (8'ha1 == _T_11[7:0]) begin
        image_2_161 <= io_pixelVal_in_2_1;
      end else if (8'ha1 == _T_7[7:0]) begin
        image_2_161 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_162 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha2 == _T_29[7:0]) begin
        image_2_162 <= io_pixelVal_in_2_7;
      end else if (8'ha2 == _T_26[7:0]) begin
        image_2_162 <= io_pixelVal_in_2_6;
      end else if (8'ha2 == _T_23[7:0]) begin
        image_2_162 <= io_pixelVal_in_2_5;
      end else if (8'ha2 == _T_20[7:0]) begin
        image_2_162 <= io_pixelVal_in_2_4;
      end else if (8'ha2 == _T_17[7:0]) begin
        image_2_162 <= io_pixelVal_in_2_3;
      end else if (8'ha2 == _T_14[7:0]) begin
        image_2_162 <= io_pixelVal_in_2_2;
      end else if (8'ha2 == _T_11[7:0]) begin
        image_2_162 <= io_pixelVal_in_2_1;
      end else if (8'ha2 == _T_7[7:0]) begin
        image_2_162 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_163 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha3 == _T_29[7:0]) begin
        image_2_163 <= io_pixelVal_in_2_7;
      end else if (8'ha3 == _T_26[7:0]) begin
        image_2_163 <= io_pixelVal_in_2_6;
      end else if (8'ha3 == _T_23[7:0]) begin
        image_2_163 <= io_pixelVal_in_2_5;
      end else if (8'ha3 == _T_20[7:0]) begin
        image_2_163 <= io_pixelVal_in_2_4;
      end else if (8'ha3 == _T_17[7:0]) begin
        image_2_163 <= io_pixelVal_in_2_3;
      end else if (8'ha3 == _T_14[7:0]) begin
        image_2_163 <= io_pixelVal_in_2_2;
      end else if (8'ha3 == _T_11[7:0]) begin
        image_2_163 <= io_pixelVal_in_2_1;
      end else if (8'ha3 == _T_7[7:0]) begin
        image_2_163 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_164 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha4 == _T_29[7:0]) begin
        image_2_164 <= io_pixelVal_in_2_7;
      end else if (8'ha4 == _T_26[7:0]) begin
        image_2_164 <= io_pixelVal_in_2_6;
      end else if (8'ha4 == _T_23[7:0]) begin
        image_2_164 <= io_pixelVal_in_2_5;
      end else if (8'ha4 == _T_20[7:0]) begin
        image_2_164 <= io_pixelVal_in_2_4;
      end else if (8'ha4 == _T_17[7:0]) begin
        image_2_164 <= io_pixelVal_in_2_3;
      end else if (8'ha4 == _T_14[7:0]) begin
        image_2_164 <= io_pixelVal_in_2_2;
      end else if (8'ha4 == _T_11[7:0]) begin
        image_2_164 <= io_pixelVal_in_2_1;
      end else if (8'ha4 == _T_7[7:0]) begin
        image_2_164 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_165 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha5 == _T_29[7:0]) begin
        image_2_165 <= io_pixelVal_in_2_7;
      end else if (8'ha5 == _T_26[7:0]) begin
        image_2_165 <= io_pixelVal_in_2_6;
      end else if (8'ha5 == _T_23[7:0]) begin
        image_2_165 <= io_pixelVal_in_2_5;
      end else if (8'ha5 == _T_20[7:0]) begin
        image_2_165 <= io_pixelVal_in_2_4;
      end else if (8'ha5 == _T_17[7:0]) begin
        image_2_165 <= io_pixelVal_in_2_3;
      end else if (8'ha5 == _T_14[7:0]) begin
        image_2_165 <= io_pixelVal_in_2_2;
      end else if (8'ha5 == _T_11[7:0]) begin
        image_2_165 <= io_pixelVal_in_2_1;
      end else if (8'ha5 == _T_7[7:0]) begin
        image_2_165 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_166 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha6 == _T_29[7:0]) begin
        image_2_166 <= io_pixelVal_in_2_7;
      end else if (8'ha6 == _T_26[7:0]) begin
        image_2_166 <= io_pixelVal_in_2_6;
      end else if (8'ha6 == _T_23[7:0]) begin
        image_2_166 <= io_pixelVal_in_2_5;
      end else if (8'ha6 == _T_20[7:0]) begin
        image_2_166 <= io_pixelVal_in_2_4;
      end else if (8'ha6 == _T_17[7:0]) begin
        image_2_166 <= io_pixelVal_in_2_3;
      end else if (8'ha6 == _T_14[7:0]) begin
        image_2_166 <= io_pixelVal_in_2_2;
      end else if (8'ha6 == _T_11[7:0]) begin
        image_2_166 <= io_pixelVal_in_2_1;
      end else if (8'ha6 == _T_7[7:0]) begin
        image_2_166 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_167 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha7 == _T_29[7:0]) begin
        image_2_167 <= io_pixelVal_in_2_7;
      end else if (8'ha7 == _T_26[7:0]) begin
        image_2_167 <= io_pixelVal_in_2_6;
      end else if (8'ha7 == _T_23[7:0]) begin
        image_2_167 <= io_pixelVal_in_2_5;
      end else if (8'ha7 == _T_20[7:0]) begin
        image_2_167 <= io_pixelVal_in_2_4;
      end else if (8'ha7 == _T_17[7:0]) begin
        image_2_167 <= io_pixelVal_in_2_3;
      end else if (8'ha7 == _T_14[7:0]) begin
        image_2_167 <= io_pixelVal_in_2_2;
      end else if (8'ha7 == _T_11[7:0]) begin
        image_2_167 <= io_pixelVal_in_2_1;
      end else if (8'ha7 == _T_7[7:0]) begin
        image_2_167 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_168 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha8 == _T_29[7:0]) begin
        image_2_168 <= io_pixelVal_in_2_7;
      end else if (8'ha8 == _T_26[7:0]) begin
        image_2_168 <= io_pixelVal_in_2_6;
      end else if (8'ha8 == _T_23[7:0]) begin
        image_2_168 <= io_pixelVal_in_2_5;
      end else if (8'ha8 == _T_20[7:0]) begin
        image_2_168 <= io_pixelVal_in_2_4;
      end else if (8'ha8 == _T_17[7:0]) begin
        image_2_168 <= io_pixelVal_in_2_3;
      end else if (8'ha8 == _T_14[7:0]) begin
        image_2_168 <= io_pixelVal_in_2_2;
      end else if (8'ha8 == _T_11[7:0]) begin
        image_2_168 <= io_pixelVal_in_2_1;
      end else if (8'ha8 == _T_7[7:0]) begin
        image_2_168 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_169 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha9 == _T_29[7:0]) begin
        image_2_169 <= io_pixelVal_in_2_7;
      end else if (8'ha9 == _T_26[7:0]) begin
        image_2_169 <= io_pixelVal_in_2_6;
      end else if (8'ha9 == _T_23[7:0]) begin
        image_2_169 <= io_pixelVal_in_2_5;
      end else if (8'ha9 == _T_20[7:0]) begin
        image_2_169 <= io_pixelVal_in_2_4;
      end else if (8'ha9 == _T_17[7:0]) begin
        image_2_169 <= io_pixelVal_in_2_3;
      end else if (8'ha9 == _T_14[7:0]) begin
        image_2_169 <= io_pixelVal_in_2_2;
      end else if (8'ha9 == _T_11[7:0]) begin
        image_2_169 <= io_pixelVal_in_2_1;
      end else if (8'ha9 == _T_7[7:0]) begin
        image_2_169 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_170 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'haa == _T_29[7:0]) begin
        image_2_170 <= io_pixelVal_in_2_7;
      end else if (8'haa == _T_26[7:0]) begin
        image_2_170 <= io_pixelVal_in_2_6;
      end else if (8'haa == _T_23[7:0]) begin
        image_2_170 <= io_pixelVal_in_2_5;
      end else if (8'haa == _T_20[7:0]) begin
        image_2_170 <= io_pixelVal_in_2_4;
      end else if (8'haa == _T_17[7:0]) begin
        image_2_170 <= io_pixelVal_in_2_3;
      end else if (8'haa == _T_14[7:0]) begin
        image_2_170 <= io_pixelVal_in_2_2;
      end else if (8'haa == _T_11[7:0]) begin
        image_2_170 <= io_pixelVal_in_2_1;
      end else if (8'haa == _T_7[7:0]) begin
        image_2_170 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_171 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hab == _T_29[7:0]) begin
        image_2_171 <= io_pixelVal_in_2_7;
      end else if (8'hab == _T_26[7:0]) begin
        image_2_171 <= io_pixelVal_in_2_6;
      end else if (8'hab == _T_23[7:0]) begin
        image_2_171 <= io_pixelVal_in_2_5;
      end else if (8'hab == _T_20[7:0]) begin
        image_2_171 <= io_pixelVal_in_2_4;
      end else if (8'hab == _T_17[7:0]) begin
        image_2_171 <= io_pixelVal_in_2_3;
      end else if (8'hab == _T_14[7:0]) begin
        image_2_171 <= io_pixelVal_in_2_2;
      end else if (8'hab == _T_11[7:0]) begin
        image_2_171 <= io_pixelVal_in_2_1;
      end else if (8'hab == _T_7[7:0]) begin
        image_2_171 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_172 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hac == _T_29[7:0]) begin
        image_2_172 <= io_pixelVal_in_2_7;
      end else if (8'hac == _T_26[7:0]) begin
        image_2_172 <= io_pixelVal_in_2_6;
      end else if (8'hac == _T_23[7:0]) begin
        image_2_172 <= io_pixelVal_in_2_5;
      end else if (8'hac == _T_20[7:0]) begin
        image_2_172 <= io_pixelVal_in_2_4;
      end else if (8'hac == _T_17[7:0]) begin
        image_2_172 <= io_pixelVal_in_2_3;
      end else if (8'hac == _T_14[7:0]) begin
        image_2_172 <= io_pixelVal_in_2_2;
      end else if (8'hac == _T_11[7:0]) begin
        image_2_172 <= io_pixelVal_in_2_1;
      end else if (8'hac == _T_7[7:0]) begin
        image_2_172 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_173 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'had == _T_29[7:0]) begin
        image_2_173 <= io_pixelVal_in_2_7;
      end else if (8'had == _T_26[7:0]) begin
        image_2_173 <= io_pixelVal_in_2_6;
      end else if (8'had == _T_23[7:0]) begin
        image_2_173 <= io_pixelVal_in_2_5;
      end else if (8'had == _T_20[7:0]) begin
        image_2_173 <= io_pixelVal_in_2_4;
      end else if (8'had == _T_17[7:0]) begin
        image_2_173 <= io_pixelVal_in_2_3;
      end else if (8'had == _T_14[7:0]) begin
        image_2_173 <= io_pixelVal_in_2_2;
      end else if (8'had == _T_11[7:0]) begin
        image_2_173 <= io_pixelVal_in_2_1;
      end else if (8'had == _T_7[7:0]) begin
        image_2_173 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_174 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hae == _T_29[7:0]) begin
        image_2_174 <= io_pixelVal_in_2_7;
      end else if (8'hae == _T_26[7:0]) begin
        image_2_174 <= io_pixelVal_in_2_6;
      end else if (8'hae == _T_23[7:0]) begin
        image_2_174 <= io_pixelVal_in_2_5;
      end else if (8'hae == _T_20[7:0]) begin
        image_2_174 <= io_pixelVal_in_2_4;
      end else if (8'hae == _T_17[7:0]) begin
        image_2_174 <= io_pixelVal_in_2_3;
      end else if (8'hae == _T_14[7:0]) begin
        image_2_174 <= io_pixelVal_in_2_2;
      end else if (8'hae == _T_11[7:0]) begin
        image_2_174 <= io_pixelVal_in_2_1;
      end else if (8'hae == _T_7[7:0]) begin
        image_2_174 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_175 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'haf == _T_29[7:0]) begin
        image_2_175 <= io_pixelVal_in_2_7;
      end else if (8'haf == _T_26[7:0]) begin
        image_2_175 <= io_pixelVal_in_2_6;
      end else if (8'haf == _T_23[7:0]) begin
        image_2_175 <= io_pixelVal_in_2_5;
      end else if (8'haf == _T_20[7:0]) begin
        image_2_175 <= io_pixelVal_in_2_4;
      end else if (8'haf == _T_17[7:0]) begin
        image_2_175 <= io_pixelVal_in_2_3;
      end else if (8'haf == _T_14[7:0]) begin
        image_2_175 <= io_pixelVal_in_2_2;
      end else if (8'haf == _T_11[7:0]) begin
        image_2_175 <= io_pixelVal_in_2_1;
      end else if (8'haf == _T_7[7:0]) begin
        image_2_175 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_176 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb0 == _T_29[7:0]) begin
        image_2_176 <= io_pixelVal_in_2_7;
      end else if (8'hb0 == _T_26[7:0]) begin
        image_2_176 <= io_pixelVal_in_2_6;
      end else if (8'hb0 == _T_23[7:0]) begin
        image_2_176 <= io_pixelVal_in_2_5;
      end else if (8'hb0 == _T_20[7:0]) begin
        image_2_176 <= io_pixelVal_in_2_4;
      end else if (8'hb0 == _T_17[7:0]) begin
        image_2_176 <= io_pixelVal_in_2_3;
      end else if (8'hb0 == _T_14[7:0]) begin
        image_2_176 <= io_pixelVal_in_2_2;
      end else if (8'hb0 == _T_11[7:0]) begin
        image_2_176 <= io_pixelVal_in_2_1;
      end else if (8'hb0 == _T_7[7:0]) begin
        image_2_176 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_177 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb1 == _T_29[7:0]) begin
        image_2_177 <= io_pixelVal_in_2_7;
      end else if (8'hb1 == _T_26[7:0]) begin
        image_2_177 <= io_pixelVal_in_2_6;
      end else if (8'hb1 == _T_23[7:0]) begin
        image_2_177 <= io_pixelVal_in_2_5;
      end else if (8'hb1 == _T_20[7:0]) begin
        image_2_177 <= io_pixelVal_in_2_4;
      end else if (8'hb1 == _T_17[7:0]) begin
        image_2_177 <= io_pixelVal_in_2_3;
      end else if (8'hb1 == _T_14[7:0]) begin
        image_2_177 <= io_pixelVal_in_2_2;
      end else if (8'hb1 == _T_11[7:0]) begin
        image_2_177 <= io_pixelVal_in_2_1;
      end else if (8'hb1 == _T_7[7:0]) begin
        image_2_177 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_178 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb2 == _T_29[7:0]) begin
        image_2_178 <= io_pixelVal_in_2_7;
      end else if (8'hb2 == _T_26[7:0]) begin
        image_2_178 <= io_pixelVal_in_2_6;
      end else if (8'hb2 == _T_23[7:0]) begin
        image_2_178 <= io_pixelVal_in_2_5;
      end else if (8'hb2 == _T_20[7:0]) begin
        image_2_178 <= io_pixelVal_in_2_4;
      end else if (8'hb2 == _T_17[7:0]) begin
        image_2_178 <= io_pixelVal_in_2_3;
      end else if (8'hb2 == _T_14[7:0]) begin
        image_2_178 <= io_pixelVal_in_2_2;
      end else if (8'hb2 == _T_11[7:0]) begin
        image_2_178 <= io_pixelVal_in_2_1;
      end else if (8'hb2 == _T_7[7:0]) begin
        image_2_178 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_179 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb3 == _T_29[7:0]) begin
        image_2_179 <= io_pixelVal_in_2_7;
      end else if (8'hb3 == _T_26[7:0]) begin
        image_2_179 <= io_pixelVal_in_2_6;
      end else if (8'hb3 == _T_23[7:0]) begin
        image_2_179 <= io_pixelVal_in_2_5;
      end else if (8'hb3 == _T_20[7:0]) begin
        image_2_179 <= io_pixelVal_in_2_4;
      end else if (8'hb3 == _T_17[7:0]) begin
        image_2_179 <= io_pixelVal_in_2_3;
      end else if (8'hb3 == _T_14[7:0]) begin
        image_2_179 <= io_pixelVal_in_2_2;
      end else if (8'hb3 == _T_11[7:0]) begin
        image_2_179 <= io_pixelVal_in_2_1;
      end else if (8'hb3 == _T_7[7:0]) begin
        image_2_179 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_180 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb4 == _T_29[7:0]) begin
        image_2_180 <= io_pixelVal_in_2_7;
      end else if (8'hb4 == _T_26[7:0]) begin
        image_2_180 <= io_pixelVal_in_2_6;
      end else if (8'hb4 == _T_23[7:0]) begin
        image_2_180 <= io_pixelVal_in_2_5;
      end else if (8'hb4 == _T_20[7:0]) begin
        image_2_180 <= io_pixelVal_in_2_4;
      end else if (8'hb4 == _T_17[7:0]) begin
        image_2_180 <= io_pixelVal_in_2_3;
      end else if (8'hb4 == _T_14[7:0]) begin
        image_2_180 <= io_pixelVal_in_2_2;
      end else if (8'hb4 == _T_11[7:0]) begin
        image_2_180 <= io_pixelVal_in_2_1;
      end else if (8'hb4 == _T_7[7:0]) begin
        image_2_180 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_181 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb5 == _T_29[7:0]) begin
        image_2_181 <= io_pixelVal_in_2_7;
      end else if (8'hb5 == _T_26[7:0]) begin
        image_2_181 <= io_pixelVal_in_2_6;
      end else if (8'hb5 == _T_23[7:0]) begin
        image_2_181 <= io_pixelVal_in_2_5;
      end else if (8'hb5 == _T_20[7:0]) begin
        image_2_181 <= io_pixelVal_in_2_4;
      end else if (8'hb5 == _T_17[7:0]) begin
        image_2_181 <= io_pixelVal_in_2_3;
      end else if (8'hb5 == _T_14[7:0]) begin
        image_2_181 <= io_pixelVal_in_2_2;
      end else if (8'hb5 == _T_11[7:0]) begin
        image_2_181 <= io_pixelVal_in_2_1;
      end else if (8'hb5 == _T_7[7:0]) begin
        image_2_181 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_182 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb6 == _T_29[7:0]) begin
        image_2_182 <= io_pixelVal_in_2_7;
      end else if (8'hb6 == _T_26[7:0]) begin
        image_2_182 <= io_pixelVal_in_2_6;
      end else if (8'hb6 == _T_23[7:0]) begin
        image_2_182 <= io_pixelVal_in_2_5;
      end else if (8'hb6 == _T_20[7:0]) begin
        image_2_182 <= io_pixelVal_in_2_4;
      end else if (8'hb6 == _T_17[7:0]) begin
        image_2_182 <= io_pixelVal_in_2_3;
      end else if (8'hb6 == _T_14[7:0]) begin
        image_2_182 <= io_pixelVal_in_2_2;
      end else if (8'hb6 == _T_11[7:0]) begin
        image_2_182 <= io_pixelVal_in_2_1;
      end else if (8'hb6 == _T_7[7:0]) begin
        image_2_182 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_183 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb7 == _T_29[7:0]) begin
        image_2_183 <= io_pixelVal_in_2_7;
      end else if (8'hb7 == _T_26[7:0]) begin
        image_2_183 <= io_pixelVal_in_2_6;
      end else if (8'hb7 == _T_23[7:0]) begin
        image_2_183 <= io_pixelVal_in_2_5;
      end else if (8'hb7 == _T_20[7:0]) begin
        image_2_183 <= io_pixelVal_in_2_4;
      end else if (8'hb7 == _T_17[7:0]) begin
        image_2_183 <= io_pixelVal_in_2_3;
      end else if (8'hb7 == _T_14[7:0]) begin
        image_2_183 <= io_pixelVal_in_2_2;
      end else if (8'hb7 == _T_11[7:0]) begin
        image_2_183 <= io_pixelVal_in_2_1;
      end else if (8'hb7 == _T_7[7:0]) begin
        image_2_183 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_184 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb8 == _T_29[7:0]) begin
        image_2_184 <= io_pixelVal_in_2_7;
      end else if (8'hb8 == _T_26[7:0]) begin
        image_2_184 <= io_pixelVal_in_2_6;
      end else if (8'hb8 == _T_23[7:0]) begin
        image_2_184 <= io_pixelVal_in_2_5;
      end else if (8'hb8 == _T_20[7:0]) begin
        image_2_184 <= io_pixelVal_in_2_4;
      end else if (8'hb8 == _T_17[7:0]) begin
        image_2_184 <= io_pixelVal_in_2_3;
      end else if (8'hb8 == _T_14[7:0]) begin
        image_2_184 <= io_pixelVal_in_2_2;
      end else if (8'hb8 == _T_11[7:0]) begin
        image_2_184 <= io_pixelVal_in_2_1;
      end else if (8'hb8 == _T_7[7:0]) begin
        image_2_184 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_185 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb9 == _T_29[7:0]) begin
        image_2_185 <= io_pixelVal_in_2_7;
      end else if (8'hb9 == _T_26[7:0]) begin
        image_2_185 <= io_pixelVal_in_2_6;
      end else if (8'hb9 == _T_23[7:0]) begin
        image_2_185 <= io_pixelVal_in_2_5;
      end else if (8'hb9 == _T_20[7:0]) begin
        image_2_185 <= io_pixelVal_in_2_4;
      end else if (8'hb9 == _T_17[7:0]) begin
        image_2_185 <= io_pixelVal_in_2_3;
      end else if (8'hb9 == _T_14[7:0]) begin
        image_2_185 <= io_pixelVal_in_2_2;
      end else if (8'hb9 == _T_11[7:0]) begin
        image_2_185 <= io_pixelVal_in_2_1;
      end else if (8'hb9 == _T_7[7:0]) begin
        image_2_185 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_186 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hba == _T_29[7:0]) begin
        image_2_186 <= io_pixelVal_in_2_7;
      end else if (8'hba == _T_26[7:0]) begin
        image_2_186 <= io_pixelVal_in_2_6;
      end else if (8'hba == _T_23[7:0]) begin
        image_2_186 <= io_pixelVal_in_2_5;
      end else if (8'hba == _T_20[7:0]) begin
        image_2_186 <= io_pixelVal_in_2_4;
      end else if (8'hba == _T_17[7:0]) begin
        image_2_186 <= io_pixelVal_in_2_3;
      end else if (8'hba == _T_14[7:0]) begin
        image_2_186 <= io_pixelVal_in_2_2;
      end else if (8'hba == _T_11[7:0]) begin
        image_2_186 <= io_pixelVal_in_2_1;
      end else if (8'hba == _T_7[7:0]) begin
        image_2_186 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_187 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbb == _T_29[7:0]) begin
        image_2_187 <= io_pixelVal_in_2_7;
      end else if (8'hbb == _T_26[7:0]) begin
        image_2_187 <= io_pixelVal_in_2_6;
      end else if (8'hbb == _T_23[7:0]) begin
        image_2_187 <= io_pixelVal_in_2_5;
      end else if (8'hbb == _T_20[7:0]) begin
        image_2_187 <= io_pixelVal_in_2_4;
      end else if (8'hbb == _T_17[7:0]) begin
        image_2_187 <= io_pixelVal_in_2_3;
      end else if (8'hbb == _T_14[7:0]) begin
        image_2_187 <= io_pixelVal_in_2_2;
      end else if (8'hbb == _T_11[7:0]) begin
        image_2_187 <= io_pixelVal_in_2_1;
      end else if (8'hbb == _T_7[7:0]) begin
        image_2_187 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_188 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbc == _T_29[7:0]) begin
        image_2_188 <= io_pixelVal_in_2_7;
      end else if (8'hbc == _T_26[7:0]) begin
        image_2_188 <= io_pixelVal_in_2_6;
      end else if (8'hbc == _T_23[7:0]) begin
        image_2_188 <= io_pixelVal_in_2_5;
      end else if (8'hbc == _T_20[7:0]) begin
        image_2_188 <= io_pixelVal_in_2_4;
      end else if (8'hbc == _T_17[7:0]) begin
        image_2_188 <= io_pixelVal_in_2_3;
      end else if (8'hbc == _T_14[7:0]) begin
        image_2_188 <= io_pixelVal_in_2_2;
      end else if (8'hbc == _T_11[7:0]) begin
        image_2_188 <= io_pixelVal_in_2_1;
      end else if (8'hbc == _T_7[7:0]) begin
        image_2_188 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_189 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbd == _T_29[7:0]) begin
        image_2_189 <= io_pixelVal_in_2_7;
      end else if (8'hbd == _T_26[7:0]) begin
        image_2_189 <= io_pixelVal_in_2_6;
      end else if (8'hbd == _T_23[7:0]) begin
        image_2_189 <= io_pixelVal_in_2_5;
      end else if (8'hbd == _T_20[7:0]) begin
        image_2_189 <= io_pixelVal_in_2_4;
      end else if (8'hbd == _T_17[7:0]) begin
        image_2_189 <= io_pixelVal_in_2_3;
      end else if (8'hbd == _T_14[7:0]) begin
        image_2_189 <= io_pixelVal_in_2_2;
      end else if (8'hbd == _T_11[7:0]) begin
        image_2_189 <= io_pixelVal_in_2_1;
      end else if (8'hbd == _T_7[7:0]) begin
        image_2_189 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_190 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbe == _T_29[7:0]) begin
        image_2_190 <= io_pixelVal_in_2_7;
      end else if (8'hbe == _T_26[7:0]) begin
        image_2_190 <= io_pixelVal_in_2_6;
      end else if (8'hbe == _T_23[7:0]) begin
        image_2_190 <= io_pixelVal_in_2_5;
      end else if (8'hbe == _T_20[7:0]) begin
        image_2_190 <= io_pixelVal_in_2_4;
      end else if (8'hbe == _T_17[7:0]) begin
        image_2_190 <= io_pixelVal_in_2_3;
      end else if (8'hbe == _T_14[7:0]) begin
        image_2_190 <= io_pixelVal_in_2_2;
      end else if (8'hbe == _T_11[7:0]) begin
        image_2_190 <= io_pixelVal_in_2_1;
      end else if (8'hbe == _T_7[7:0]) begin
        image_2_190 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_191 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbf == _T_29[7:0]) begin
        image_2_191 <= io_pixelVal_in_2_7;
      end else if (8'hbf == _T_26[7:0]) begin
        image_2_191 <= io_pixelVal_in_2_6;
      end else if (8'hbf == _T_23[7:0]) begin
        image_2_191 <= io_pixelVal_in_2_5;
      end else if (8'hbf == _T_20[7:0]) begin
        image_2_191 <= io_pixelVal_in_2_4;
      end else if (8'hbf == _T_17[7:0]) begin
        image_2_191 <= io_pixelVal_in_2_3;
      end else if (8'hbf == _T_14[7:0]) begin
        image_2_191 <= io_pixelVal_in_2_2;
      end else if (8'hbf == _T_11[7:0]) begin
        image_2_191 <= io_pixelVal_in_2_1;
      end else if (8'hbf == _T_7[7:0]) begin
        image_2_191 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      pixelIndex <= 32'h0;
    end else if (_T_90) begin
      pixelIndex <= 32'h0;
    end else begin
      pixelIndex <= _T_88;
    end
  end
endmodule
module ImageProcessing(
  input         clock,
  input         reset,
  input  [5:0]  io_SPI_filterIndex,
  input         io_SPI_invert,
  input         io_SPI_distort,
  input  [10:0] io_rowIndex,
  input  [10:0] io_colIndex,
  output [3:0]  io_pixelVal_out_0,
  output [3:0]  io_pixelVal_out_1,
  output [3:0]  io_pixelVal_out_2
);
  wire  filter_clock; // @[ImageProcessing.scala 22:22]
  wire  filter_reset; // @[ImageProcessing.scala 22:22]
  wire [5:0] filter_io_SPI_filterIndex; // @[ImageProcessing.scala 22:22]
  wire  filter_io_SPI_distort; // @[ImageProcessing.scala 22:22]
  wire [3:0] filter_io_pixelVal_out_0_0; // @[ImageProcessing.scala 22:22]
  wire [3:0] filter_io_pixelVal_out_0_1; // @[ImageProcessing.scala 22:22]
  wire [3:0] filter_io_pixelVal_out_0_2; // @[ImageProcessing.scala 22:22]
  wire [3:0] filter_io_pixelVal_out_0_3; // @[ImageProcessing.scala 22:22]
  wire [3:0] filter_io_pixelVal_out_0_4; // @[ImageProcessing.scala 22:22]
  wire [3:0] filter_io_pixelVal_out_0_5; // @[ImageProcessing.scala 22:22]
  wire [3:0] filter_io_pixelVal_out_0_6; // @[ImageProcessing.scala 22:22]
  wire [3:0] filter_io_pixelVal_out_0_7; // @[ImageProcessing.scala 22:22]
  wire [3:0] filter_io_pixelVal_out_1_0; // @[ImageProcessing.scala 22:22]
  wire [3:0] filter_io_pixelVal_out_1_1; // @[ImageProcessing.scala 22:22]
  wire [3:0] filter_io_pixelVal_out_1_2; // @[ImageProcessing.scala 22:22]
  wire [3:0] filter_io_pixelVal_out_1_3; // @[ImageProcessing.scala 22:22]
  wire [3:0] filter_io_pixelVal_out_1_4; // @[ImageProcessing.scala 22:22]
  wire [3:0] filter_io_pixelVal_out_1_5; // @[ImageProcessing.scala 22:22]
  wire [3:0] filter_io_pixelVal_out_1_6; // @[ImageProcessing.scala 22:22]
  wire [3:0] filter_io_pixelVal_out_1_7; // @[ImageProcessing.scala 22:22]
  wire [3:0] filter_io_pixelVal_out_2_0; // @[ImageProcessing.scala 22:22]
  wire [3:0] filter_io_pixelVal_out_2_1; // @[ImageProcessing.scala 22:22]
  wire [3:0] filter_io_pixelVal_out_2_2; // @[ImageProcessing.scala 22:22]
  wire [3:0] filter_io_pixelVal_out_2_3; // @[ImageProcessing.scala 22:22]
  wire [3:0] filter_io_pixelVal_out_2_4; // @[ImageProcessing.scala 22:22]
  wire [3:0] filter_io_pixelVal_out_2_5; // @[ImageProcessing.scala 22:22]
  wire [3:0] filter_io_pixelVal_out_2_6; // @[ImageProcessing.scala 22:22]
  wire [3:0] filter_io_pixelVal_out_2_7; // @[ImageProcessing.scala 22:22]
  wire  filter_io_valid_out; // @[ImageProcessing.scala 22:22]
  wire  videoBuffer_clock; // @[ImageProcessing.scala 23:27]
  wire  videoBuffer_reset; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_0; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_1; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_2; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_3; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_4; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_5; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_6; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_7; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_0; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_1; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_2; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_3; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_4; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_5; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_6; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_7; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_0; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_1; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_2; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_3; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_4; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_5; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_6; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_7; // @[ImageProcessing.scala 23:27]
  wire  videoBuffer_io_valid_in; // @[ImageProcessing.scala 23:27]
  wire [10:0] videoBuffer_io_rowIndex; // @[ImageProcessing.scala 23:27]
  wire [10:0] videoBuffer_io_colIndex; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_out_0; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_out_1; // @[ImageProcessing.scala 23:27]
  wire [3:0] videoBuffer_io_pixelVal_out_2; // @[ImageProcessing.scala 23:27]
  Filter filter ( // @[ImageProcessing.scala 22:22]
    .clock(filter_clock),
    .reset(filter_reset),
    .io_SPI_filterIndex(filter_io_SPI_filterIndex),
    .io_SPI_distort(filter_io_SPI_distort),
    .io_pixelVal_out_0_0(filter_io_pixelVal_out_0_0),
    .io_pixelVal_out_0_1(filter_io_pixelVal_out_0_1),
    .io_pixelVal_out_0_2(filter_io_pixelVal_out_0_2),
    .io_pixelVal_out_0_3(filter_io_pixelVal_out_0_3),
    .io_pixelVal_out_0_4(filter_io_pixelVal_out_0_4),
    .io_pixelVal_out_0_5(filter_io_pixelVal_out_0_5),
    .io_pixelVal_out_0_6(filter_io_pixelVal_out_0_6),
    .io_pixelVal_out_0_7(filter_io_pixelVal_out_0_7),
    .io_pixelVal_out_1_0(filter_io_pixelVal_out_1_0),
    .io_pixelVal_out_1_1(filter_io_pixelVal_out_1_1),
    .io_pixelVal_out_1_2(filter_io_pixelVal_out_1_2),
    .io_pixelVal_out_1_3(filter_io_pixelVal_out_1_3),
    .io_pixelVal_out_1_4(filter_io_pixelVal_out_1_4),
    .io_pixelVal_out_1_5(filter_io_pixelVal_out_1_5),
    .io_pixelVal_out_1_6(filter_io_pixelVal_out_1_6),
    .io_pixelVal_out_1_7(filter_io_pixelVal_out_1_7),
    .io_pixelVal_out_2_0(filter_io_pixelVal_out_2_0),
    .io_pixelVal_out_2_1(filter_io_pixelVal_out_2_1),
    .io_pixelVal_out_2_2(filter_io_pixelVal_out_2_2),
    .io_pixelVal_out_2_3(filter_io_pixelVal_out_2_3),
    .io_pixelVal_out_2_4(filter_io_pixelVal_out_2_4),
    .io_pixelVal_out_2_5(filter_io_pixelVal_out_2_5),
    .io_pixelVal_out_2_6(filter_io_pixelVal_out_2_6),
    .io_pixelVal_out_2_7(filter_io_pixelVal_out_2_7),
    .io_valid_out(filter_io_valid_out)
  );
  VideoBuffer videoBuffer ( // @[ImageProcessing.scala 23:27]
    .clock(videoBuffer_clock),
    .reset(videoBuffer_reset),
    .io_pixelVal_in_0_0(videoBuffer_io_pixelVal_in_0_0),
    .io_pixelVal_in_0_1(videoBuffer_io_pixelVal_in_0_1),
    .io_pixelVal_in_0_2(videoBuffer_io_pixelVal_in_0_2),
    .io_pixelVal_in_0_3(videoBuffer_io_pixelVal_in_0_3),
    .io_pixelVal_in_0_4(videoBuffer_io_pixelVal_in_0_4),
    .io_pixelVal_in_0_5(videoBuffer_io_pixelVal_in_0_5),
    .io_pixelVal_in_0_6(videoBuffer_io_pixelVal_in_0_6),
    .io_pixelVal_in_0_7(videoBuffer_io_pixelVal_in_0_7),
    .io_pixelVal_in_1_0(videoBuffer_io_pixelVal_in_1_0),
    .io_pixelVal_in_1_1(videoBuffer_io_pixelVal_in_1_1),
    .io_pixelVal_in_1_2(videoBuffer_io_pixelVal_in_1_2),
    .io_pixelVal_in_1_3(videoBuffer_io_pixelVal_in_1_3),
    .io_pixelVal_in_1_4(videoBuffer_io_pixelVal_in_1_4),
    .io_pixelVal_in_1_5(videoBuffer_io_pixelVal_in_1_5),
    .io_pixelVal_in_1_6(videoBuffer_io_pixelVal_in_1_6),
    .io_pixelVal_in_1_7(videoBuffer_io_pixelVal_in_1_7),
    .io_pixelVal_in_2_0(videoBuffer_io_pixelVal_in_2_0),
    .io_pixelVal_in_2_1(videoBuffer_io_pixelVal_in_2_1),
    .io_pixelVal_in_2_2(videoBuffer_io_pixelVal_in_2_2),
    .io_pixelVal_in_2_3(videoBuffer_io_pixelVal_in_2_3),
    .io_pixelVal_in_2_4(videoBuffer_io_pixelVal_in_2_4),
    .io_pixelVal_in_2_5(videoBuffer_io_pixelVal_in_2_5),
    .io_pixelVal_in_2_6(videoBuffer_io_pixelVal_in_2_6),
    .io_pixelVal_in_2_7(videoBuffer_io_pixelVal_in_2_7),
    .io_valid_in(videoBuffer_io_valid_in),
    .io_rowIndex(videoBuffer_io_rowIndex),
    .io_colIndex(videoBuffer_io_colIndex),
    .io_pixelVal_out_0(videoBuffer_io_pixelVal_out_0),
    .io_pixelVal_out_1(videoBuffer_io_pixelVal_out_1),
    .io_pixelVal_out_2(videoBuffer_io_pixelVal_out_2)
  );
  assign io_pixelVal_out_0 = videoBuffer_io_pixelVal_out_0; // @[ImageProcessing.scala 35:25 ImageProcessing.scala 35:25 ImageProcessing.scala 35:25 ImageProcessing.scala 35:25 ImageProcessing.scala 35:25 ImageProcessing.scala 35:25 ImageProcessing.scala 35:25 ImageProcessing.scala 35:25]
  assign io_pixelVal_out_1 = videoBuffer_io_pixelVal_out_1; // @[ImageProcessing.scala 35:25 ImageProcessing.scala 35:25 ImageProcessing.scala 35:25 ImageProcessing.scala 35:25 ImageProcessing.scala 35:25 ImageProcessing.scala 35:25 ImageProcessing.scala 35:25 ImageProcessing.scala 35:25]
  assign io_pixelVal_out_2 = videoBuffer_io_pixelVal_out_2; // @[ImageProcessing.scala 35:25 ImageProcessing.scala 35:25 ImageProcessing.scala 35:25 ImageProcessing.scala 35:25 ImageProcessing.scala 35:25 ImageProcessing.scala 35:25 ImageProcessing.scala 35:25 ImageProcessing.scala 35:25]
  assign filter_clock = clock;
  assign filter_reset = reset;
  assign filter_io_SPI_filterIndex = io_SPI_filterIndex; // @[ImageProcessing.scala 28:29]
  assign filter_io_SPI_distort = io_SPI_distort; // @[ImageProcessing.scala 30:29]
  assign videoBuffer_clock = clock;
  assign videoBuffer_reset = reset;
  assign videoBuffer_io_pixelVal_in_0_0 = filter_io_pixelVal_out_0_0; // @[ImageProcessing.scala 34:39]
  assign videoBuffer_io_pixelVal_in_0_1 = filter_io_pixelVal_out_0_1; // @[ImageProcessing.scala 34:39]
  assign videoBuffer_io_pixelVal_in_0_2 = filter_io_pixelVal_out_0_2; // @[ImageProcessing.scala 34:39]
  assign videoBuffer_io_pixelVal_in_0_3 = filter_io_pixelVal_out_0_3; // @[ImageProcessing.scala 34:39]
  assign videoBuffer_io_pixelVal_in_0_4 = filter_io_pixelVal_out_0_4; // @[ImageProcessing.scala 34:39]
  assign videoBuffer_io_pixelVal_in_0_5 = filter_io_pixelVal_out_0_5; // @[ImageProcessing.scala 34:39]
  assign videoBuffer_io_pixelVal_in_0_6 = filter_io_pixelVal_out_0_6; // @[ImageProcessing.scala 34:39]
  assign videoBuffer_io_pixelVal_in_0_7 = filter_io_pixelVal_out_0_7; // @[ImageProcessing.scala 34:39]
  assign videoBuffer_io_pixelVal_in_1_0 = filter_io_pixelVal_out_1_0; // @[ImageProcessing.scala 34:39]
  assign videoBuffer_io_pixelVal_in_1_1 = filter_io_pixelVal_out_1_1; // @[ImageProcessing.scala 34:39]
  assign videoBuffer_io_pixelVal_in_1_2 = filter_io_pixelVal_out_1_2; // @[ImageProcessing.scala 34:39]
  assign videoBuffer_io_pixelVal_in_1_3 = filter_io_pixelVal_out_1_3; // @[ImageProcessing.scala 34:39]
  assign videoBuffer_io_pixelVal_in_1_4 = filter_io_pixelVal_out_1_4; // @[ImageProcessing.scala 34:39]
  assign videoBuffer_io_pixelVal_in_1_5 = filter_io_pixelVal_out_1_5; // @[ImageProcessing.scala 34:39]
  assign videoBuffer_io_pixelVal_in_1_6 = filter_io_pixelVal_out_1_6; // @[ImageProcessing.scala 34:39]
  assign videoBuffer_io_pixelVal_in_1_7 = filter_io_pixelVal_out_1_7; // @[ImageProcessing.scala 34:39]
  assign videoBuffer_io_pixelVal_in_2_0 = filter_io_pixelVal_out_2_0; // @[ImageProcessing.scala 34:39]
  assign videoBuffer_io_pixelVal_in_2_1 = filter_io_pixelVal_out_2_1; // @[ImageProcessing.scala 34:39]
  assign videoBuffer_io_pixelVal_in_2_2 = filter_io_pixelVal_out_2_2; // @[ImageProcessing.scala 34:39]
  assign videoBuffer_io_pixelVal_in_2_3 = filter_io_pixelVal_out_2_3; // @[ImageProcessing.scala 34:39]
  assign videoBuffer_io_pixelVal_in_2_4 = filter_io_pixelVal_out_2_4; // @[ImageProcessing.scala 34:39]
  assign videoBuffer_io_pixelVal_in_2_5 = filter_io_pixelVal_out_2_5; // @[ImageProcessing.scala 34:39]
  assign videoBuffer_io_pixelVal_in_2_6 = filter_io_pixelVal_out_2_6; // @[ImageProcessing.scala 34:39]
  assign videoBuffer_io_pixelVal_in_2_7 = filter_io_pixelVal_out_2_7; // @[ImageProcessing.scala 34:39]
  assign videoBuffer_io_valid_in = filter_io_valid_out; // @[ImageProcessing.scala 38:27]
  assign videoBuffer_io_rowIndex = io_rowIndex; // @[ImageProcessing.scala 25:27]
  assign videoBuffer_io_colIndex = io_colIndex; // @[ImageProcessing.scala 26:27]
endmodule
