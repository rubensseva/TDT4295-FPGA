module VideoBuffer(
  input         clock,
  input         reset,
  input  [3:0]  io_pixelVal_in_0,
  input  [3:0]  io_pixelVal_in_1,
  input  [3:0]  io_pixelVal_in_2,
  input  [3:0]  io_pixelVal_in_3,
  input  [3:0]  io_pixelVal_in_4,
  input  [3:0]  io_pixelVal_in_5,
  input  [3:0]  io_pixelVal_in_6,
  input  [3:0]  io_pixelVal_in_7,
  input         io_valid_in,
  input  [10:0] io_rowIndex,
  input  [10:0] io_colIndex,
  output [3:0]  io_pixelVal_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] image_0; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_1; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_2; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_3; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_4; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_5; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_6; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_7; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_8; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_9; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_10; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_11; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_12; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_13; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_14; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_15; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_16; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_17; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_18; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_19; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_20; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_21; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_22; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_23; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_24; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_25; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_26; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_27; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_28; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_29; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_30; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_31; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_32; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_33; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_34; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_35; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_36; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_37; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_38; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_39; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_40; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_41; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_42; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_43; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_44; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_45; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_46; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_47; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_48; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_49; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_50; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_51; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_52; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_53; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_54; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_55; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_56; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_57; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_58; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_59; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_60; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_61; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_62; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_63; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_64; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_65; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_66; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_67; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_68; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_69; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_70; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_71; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_72; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_73; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_74; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_75; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_76; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_77; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_78; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_79; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_80; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_81; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_82; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_83; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_84; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_85; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_86; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_87; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_88; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_89; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_90; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_91; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_92; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_93; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_94; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_95; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_96; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_97; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_98; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_99; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_100; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_101; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_102; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_103; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_104; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_105; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_106; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_107; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_108; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_109; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_110; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_111; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_112; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_113; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_114; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_115; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_116; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_117; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_118; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_119; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_120; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_121; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_122; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_123; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_124; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_125; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_126; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_127; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_128; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_129; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_130; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_131; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_132; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_133; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_134; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_135; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_136; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_137; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_138; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_139; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_140; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_141; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_142; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_143; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_144; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_145; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_146; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_147; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_148; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_149; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_150; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_151; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_152; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_153; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_154; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_155; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_156; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_157; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_158; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_159; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_160; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_161; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_162; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_163; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_164; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_165; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_166; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_167; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_168; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_169; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_170; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_171; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_172; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_173; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_174; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_175; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_176; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_177; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_178; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_179; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_180; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_181; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_182; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_183; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_184; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_185; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_186; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_187; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_188; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_189; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_190; // @[VideoBuffer.scala 20:24]
  reg [3:0] image_191; // @[VideoBuffer.scala 20:24]
  wire [15:0] _T_1 = io_rowIndex * 11'h10; // @[VideoBuffer.scala 35:46]
  wire [15:0] _GEN_1922 = {{5'd0}, io_colIndex}; // @[VideoBuffer.scala 35:61]
  wire [15:0] _T_3 = _T_1 + _GEN_1922; // @[VideoBuffer.scala 35:61]
  wire [3:0] _GEN_1 = 8'h1 == _T_3[7:0] ? image_1 : image_0; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_2 = 8'h2 == _T_3[7:0] ? image_2 : _GEN_1; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_3 = 8'h3 == _T_3[7:0] ? image_3 : _GEN_2; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_4 = 8'h4 == _T_3[7:0] ? image_4 : _GEN_3; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_5 = 8'h5 == _T_3[7:0] ? image_5 : _GEN_4; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_6 = 8'h6 == _T_3[7:0] ? image_6 : _GEN_5; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_7 = 8'h7 == _T_3[7:0] ? image_7 : _GEN_6; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_8 = 8'h8 == _T_3[7:0] ? image_8 : _GEN_7; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_9 = 8'h9 == _T_3[7:0] ? image_9 : _GEN_8; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_10 = 8'ha == _T_3[7:0] ? image_10 : _GEN_9; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_11 = 8'hb == _T_3[7:0] ? image_11 : _GEN_10; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_12 = 8'hc == _T_3[7:0] ? image_12 : _GEN_11; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_13 = 8'hd == _T_3[7:0] ? image_13 : _GEN_12; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_14 = 8'he == _T_3[7:0] ? image_14 : _GEN_13; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_15 = 8'hf == _T_3[7:0] ? image_15 : _GEN_14; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_16 = 8'h10 == _T_3[7:0] ? image_16 : _GEN_15; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_17 = 8'h11 == _T_3[7:0] ? image_17 : _GEN_16; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_18 = 8'h12 == _T_3[7:0] ? image_18 : _GEN_17; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_19 = 8'h13 == _T_3[7:0] ? image_19 : _GEN_18; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_20 = 8'h14 == _T_3[7:0] ? image_20 : _GEN_19; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_21 = 8'h15 == _T_3[7:0] ? image_21 : _GEN_20; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_22 = 8'h16 == _T_3[7:0] ? image_22 : _GEN_21; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_23 = 8'h17 == _T_3[7:0] ? image_23 : _GEN_22; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_24 = 8'h18 == _T_3[7:0] ? image_24 : _GEN_23; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_25 = 8'h19 == _T_3[7:0] ? image_25 : _GEN_24; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_26 = 8'h1a == _T_3[7:0] ? image_26 : _GEN_25; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_27 = 8'h1b == _T_3[7:0] ? image_27 : _GEN_26; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_28 = 8'h1c == _T_3[7:0] ? image_28 : _GEN_27; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_29 = 8'h1d == _T_3[7:0] ? image_29 : _GEN_28; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_30 = 8'h1e == _T_3[7:0] ? image_30 : _GEN_29; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_31 = 8'h1f == _T_3[7:0] ? image_31 : _GEN_30; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_32 = 8'h20 == _T_3[7:0] ? image_32 : _GEN_31; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_33 = 8'h21 == _T_3[7:0] ? image_33 : _GEN_32; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_34 = 8'h22 == _T_3[7:0] ? image_34 : _GEN_33; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_35 = 8'h23 == _T_3[7:0] ? image_35 : _GEN_34; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_36 = 8'h24 == _T_3[7:0] ? image_36 : _GEN_35; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_37 = 8'h25 == _T_3[7:0] ? image_37 : _GEN_36; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_38 = 8'h26 == _T_3[7:0] ? image_38 : _GEN_37; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_39 = 8'h27 == _T_3[7:0] ? image_39 : _GEN_38; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_40 = 8'h28 == _T_3[7:0] ? image_40 : _GEN_39; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_41 = 8'h29 == _T_3[7:0] ? image_41 : _GEN_40; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_42 = 8'h2a == _T_3[7:0] ? image_42 : _GEN_41; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_43 = 8'h2b == _T_3[7:0] ? image_43 : _GEN_42; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_44 = 8'h2c == _T_3[7:0] ? image_44 : _GEN_43; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_45 = 8'h2d == _T_3[7:0] ? image_45 : _GEN_44; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_46 = 8'h2e == _T_3[7:0] ? image_46 : _GEN_45; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_47 = 8'h2f == _T_3[7:0] ? image_47 : _GEN_46; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_48 = 8'h30 == _T_3[7:0] ? image_48 : _GEN_47; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_49 = 8'h31 == _T_3[7:0] ? image_49 : _GEN_48; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_50 = 8'h32 == _T_3[7:0] ? image_50 : _GEN_49; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_51 = 8'h33 == _T_3[7:0] ? image_51 : _GEN_50; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_52 = 8'h34 == _T_3[7:0] ? image_52 : _GEN_51; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_53 = 8'h35 == _T_3[7:0] ? image_53 : _GEN_52; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_54 = 8'h36 == _T_3[7:0] ? image_54 : _GEN_53; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_55 = 8'h37 == _T_3[7:0] ? image_55 : _GEN_54; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_56 = 8'h38 == _T_3[7:0] ? image_56 : _GEN_55; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_57 = 8'h39 == _T_3[7:0] ? image_57 : _GEN_56; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_58 = 8'h3a == _T_3[7:0] ? image_58 : _GEN_57; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_59 = 8'h3b == _T_3[7:0] ? image_59 : _GEN_58; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_60 = 8'h3c == _T_3[7:0] ? image_60 : _GEN_59; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_61 = 8'h3d == _T_3[7:0] ? image_61 : _GEN_60; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_62 = 8'h3e == _T_3[7:0] ? image_62 : _GEN_61; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_63 = 8'h3f == _T_3[7:0] ? image_63 : _GEN_62; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_64 = 8'h40 == _T_3[7:0] ? image_64 : _GEN_63; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_65 = 8'h41 == _T_3[7:0] ? image_65 : _GEN_64; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_66 = 8'h42 == _T_3[7:0] ? image_66 : _GEN_65; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_67 = 8'h43 == _T_3[7:0] ? image_67 : _GEN_66; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_68 = 8'h44 == _T_3[7:0] ? image_68 : _GEN_67; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_69 = 8'h45 == _T_3[7:0] ? image_69 : _GEN_68; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_70 = 8'h46 == _T_3[7:0] ? image_70 : _GEN_69; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_71 = 8'h47 == _T_3[7:0] ? image_71 : _GEN_70; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_72 = 8'h48 == _T_3[7:0] ? image_72 : _GEN_71; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_73 = 8'h49 == _T_3[7:0] ? image_73 : _GEN_72; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_74 = 8'h4a == _T_3[7:0] ? image_74 : _GEN_73; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_75 = 8'h4b == _T_3[7:0] ? image_75 : _GEN_74; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_76 = 8'h4c == _T_3[7:0] ? image_76 : _GEN_75; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_77 = 8'h4d == _T_3[7:0] ? image_77 : _GEN_76; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_78 = 8'h4e == _T_3[7:0] ? image_78 : _GEN_77; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_79 = 8'h4f == _T_3[7:0] ? image_79 : _GEN_78; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_80 = 8'h50 == _T_3[7:0] ? image_80 : _GEN_79; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_81 = 8'h51 == _T_3[7:0] ? image_81 : _GEN_80; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_82 = 8'h52 == _T_3[7:0] ? image_82 : _GEN_81; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_83 = 8'h53 == _T_3[7:0] ? image_83 : _GEN_82; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_84 = 8'h54 == _T_3[7:0] ? image_84 : _GEN_83; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_85 = 8'h55 == _T_3[7:0] ? image_85 : _GEN_84; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_86 = 8'h56 == _T_3[7:0] ? image_86 : _GEN_85; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_87 = 8'h57 == _T_3[7:0] ? image_87 : _GEN_86; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_88 = 8'h58 == _T_3[7:0] ? image_88 : _GEN_87; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_89 = 8'h59 == _T_3[7:0] ? image_89 : _GEN_88; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_90 = 8'h5a == _T_3[7:0] ? image_90 : _GEN_89; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_91 = 8'h5b == _T_3[7:0] ? image_91 : _GEN_90; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_92 = 8'h5c == _T_3[7:0] ? image_92 : _GEN_91; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_93 = 8'h5d == _T_3[7:0] ? image_93 : _GEN_92; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_94 = 8'h5e == _T_3[7:0] ? image_94 : _GEN_93; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_95 = 8'h5f == _T_3[7:0] ? image_95 : _GEN_94; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_96 = 8'h60 == _T_3[7:0] ? image_96 : _GEN_95; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_97 = 8'h61 == _T_3[7:0] ? image_97 : _GEN_96; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_98 = 8'h62 == _T_3[7:0] ? image_98 : _GEN_97; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_99 = 8'h63 == _T_3[7:0] ? image_99 : _GEN_98; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_100 = 8'h64 == _T_3[7:0] ? image_100 : _GEN_99; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_101 = 8'h65 == _T_3[7:0] ? image_101 : _GEN_100; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_102 = 8'h66 == _T_3[7:0] ? image_102 : _GEN_101; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_103 = 8'h67 == _T_3[7:0] ? image_103 : _GEN_102; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_104 = 8'h68 == _T_3[7:0] ? image_104 : _GEN_103; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_105 = 8'h69 == _T_3[7:0] ? image_105 : _GEN_104; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_106 = 8'h6a == _T_3[7:0] ? image_106 : _GEN_105; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_107 = 8'h6b == _T_3[7:0] ? image_107 : _GEN_106; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_108 = 8'h6c == _T_3[7:0] ? image_108 : _GEN_107; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_109 = 8'h6d == _T_3[7:0] ? image_109 : _GEN_108; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_110 = 8'h6e == _T_3[7:0] ? image_110 : _GEN_109; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_111 = 8'h6f == _T_3[7:0] ? image_111 : _GEN_110; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_112 = 8'h70 == _T_3[7:0] ? image_112 : _GEN_111; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_113 = 8'h71 == _T_3[7:0] ? image_113 : _GEN_112; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_114 = 8'h72 == _T_3[7:0] ? image_114 : _GEN_113; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_115 = 8'h73 == _T_3[7:0] ? image_115 : _GEN_114; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_116 = 8'h74 == _T_3[7:0] ? image_116 : _GEN_115; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_117 = 8'h75 == _T_3[7:0] ? image_117 : _GEN_116; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_118 = 8'h76 == _T_3[7:0] ? image_118 : _GEN_117; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_119 = 8'h77 == _T_3[7:0] ? image_119 : _GEN_118; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_120 = 8'h78 == _T_3[7:0] ? image_120 : _GEN_119; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_121 = 8'h79 == _T_3[7:0] ? image_121 : _GEN_120; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_122 = 8'h7a == _T_3[7:0] ? image_122 : _GEN_121; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_123 = 8'h7b == _T_3[7:0] ? image_123 : _GEN_122; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_124 = 8'h7c == _T_3[7:0] ? image_124 : _GEN_123; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_125 = 8'h7d == _T_3[7:0] ? image_125 : _GEN_124; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_126 = 8'h7e == _T_3[7:0] ? image_126 : _GEN_125; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_127 = 8'h7f == _T_3[7:0] ? image_127 : _GEN_126; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_128 = 8'h80 == _T_3[7:0] ? image_128 : _GEN_127; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_129 = 8'h81 == _T_3[7:0] ? image_129 : _GEN_128; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_130 = 8'h82 == _T_3[7:0] ? image_130 : _GEN_129; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_131 = 8'h83 == _T_3[7:0] ? image_131 : _GEN_130; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_132 = 8'h84 == _T_3[7:0] ? image_132 : _GEN_131; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_133 = 8'h85 == _T_3[7:0] ? image_133 : _GEN_132; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_134 = 8'h86 == _T_3[7:0] ? image_134 : _GEN_133; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_135 = 8'h87 == _T_3[7:0] ? image_135 : _GEN_134; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_136 = 8'h88 == _T_3[7:0] ? image_136 : _GEN_135; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_137 = 8'h89 == _T_3[7:0] ? image_137 : _GEN_136; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_138 = 8'h8a == _T_3[7:0] ? image_138 : _GEN_137; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_139 = 8'h8b == _T_3[7:0] ? image_139 : _GEN_138; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_140 = 8'h8c == _T_3[7:0] ? image_140 : _GEN_139; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_141 = 8'h8d == _T_3[7:0] ? image_141 : _GEN_140; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_142 = 8'h8e == _T_3[7:0] ? image_142 : _GEN_141; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_143 = 8'h8f == _T_3[7:0] ? image_143 : _GEN_142; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_144 = 8'h90 == _T_3[7:0] ? image_144 : _GEN_143; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_145 = 8'h91 == _T_3[7:0] ? image_145 : _GEN_144; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_146 = 8'h92 == _T_3[7:0] ? image_146 : _GEN_145; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_147 = 8'h93 == _T_3[7:0] ? image_147 : _GEN_146; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_148 = 8'h94 == _T_3[7:0] ? image_148 : _GEN_147; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_149 = 8'h95 == _T_3[7:0] ? image_149 : _GEN_148; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_150 = 8'h96 == _T_3[7:0] ? image_150 : _GEN_149; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_151 = 8'h97 == _T_3[7:0] ? image_151 : _GEN_150; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_152 = 8'h98 == _T_3[7:0] ? image_152 : _GEN_151; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_153 = 8'h99 == _T_3[7:0] ? image_153 : _GEN_152; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_154 = 8'h9a == _T_3[7:0] ? image_154 : _GEN_153; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_155 = 8'h9b == _T_3[7:0] ? image_155 : _GEN_154; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_156 = 8'h9c == _T_3[7:0] ? image_156 : _GEN_155; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_157 = 8'h9d == _T_3[7:0] ? image_157 : _GEN_156; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_158 = 8'h9e == _T_3[7:0] ? image_158 : _GEN_157; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_159 = 8'h9f == _T_3[7:0] ? image_159 : _GEN_158; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_160 = 8'ha0 == _T_3[7:0] ? image_160 : _GEN_159; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_161 = 8'ha1 == _T_3[7:0] ? image_161 : _GEN_160; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_162 = 8'ha2 == _T_3[7:0] ? image_162 : _GEN_161; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_163 = 8'ha3 == _T_3[7:0] ? image_163 : _GEN_162; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_164 = 8'ha4 == _T_3[7:0] ? image_164 : _GEN_163; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_165 = 8'ha5 == _T_3[7:0] ? image_165 : _GEN_164; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_166 = 8'ha6 == _T_3[7:0] ? image_166 : _GEN_165; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_167 = 8'ha7 == _T_3[7:0] ? image_167 : _GEN_166; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_168 = 8'ha8 == _T_3[7:0] ? image_168 : _GEN_167; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_169 = 8'ha9 == _T_3[7:0] ? image_169 : _GEN_168; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_170 = 8'haa == _T_3[7:0] ? image_170 : _GEN_169; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_171 = 8'hab == _T_3[7:0] ? image_171 : _GEN_170; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_172 = 8'hac == _T_3[7:0] ? image_172 : _GEN_171; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_173 = 8'had == _T_3[7:0] ? image_173 : _GEN_172; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_174 = 8'hae == _T_3[7:0] ? image_174 : _GEN_173; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_175 = 8'haf == _T_3[7:0] ? image_175 : _GEN_174; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_176 = 8'hb0 == _T_3[7:0] ? image_176 : _GEN_175; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_177 = 8'hb1 == _T_3[7:0] ? image_177 : _GEN_176; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_178 = 8'hb2 == _T_3[7:0] ? image_178 : _GEN_177; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_179 = 8'hb3 == _T_3[7:0] ? image_179 : _GEN_178; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_180 = 8'hb4 == _T_3[7:0] ? image_180 : _GEN_179; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_181 = 8'hb5 == _T_3[7:0] ? image_181 : _GEN_180; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_182 = 8'hb6 == _T_3[7:0] ? image_182 : _GEN_181; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_183 = 8'hb7 == _T_3[7:0] ? image_183 : _GEN_182; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_184 = 8'hb8 == _T_3[7:0] ? image_184 : _GEN_183; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_185 = 8'hb9 == _T_3[7:0] ? image_185 : _GEN_184; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_186 = 8'hba == _T_3[7:0] ? image_186 : _GEN_185; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_187 = 8'hbb == _T_3[7:0] ? image_187 : _GEN_186; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_188 = 8'hbc == _T_3[7:0] ? image_188 : _GEN_187; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_189 = 8'hbd == _T_3[7:0] ? image_189 : _GEN_188; // @[VideoBuffer.scala 35:25]
  wire [3:0] _GEN_190 = 8'hbe == _T_3[7:0] ? image_190 : _GEN_189; // @[VideoBuffer.scala 35:25]
  reg [31:0] pixelIndex; // @[VideoBuffer.scala 37:33]
  wire [32:0] _T_5 = {{1'd0}, pixelIndex}; // @[VideoBuffer.scala 41:42]
  wire [31:0] _T_9 = pixelIndex + 32'h1; // @[VideoBuffer.scala 41:42]
  wire [31:0] _T_12 = pixelIndex + 32'h2; // @[VideoBuffer.scala 41:42]
  wire [31:0] _T_15 = pixelIndex + 32'h3; // @[VideoBuffer.scala 41:42]
  wire [31:0] _T_18 = pixelIndex + 32'h4; // @[VideoBuffer.scala 41:42]
  wire [31:0] _T_21 = pixelIndex + 32'h5; // @[VideoBuffer.scala 41:42]
  wire [31:0] _T_24 = pixelIndex + 32'h6; // @[VideoBuffer.scala 41:42]
  wire [31:0] _T_27 = pixelIndex + 32'h7; // @[VideoBuffer.scala 41:42]
  wire [31:0] _T_30 = pixelIndex + 32'h8; // @[VideoBuffer.scala 43:42]
  wire [8:0] _T_31 = 5'h10 * 5'hc; // @[VideoBuffer.scala 44:42]
  wire [31:0] _GEN_1923 = {{23'd0}, _T_31}; // @[VideoBuffer.scala 44:25]
  wire  _T_32 = pixelIndex == _GEN_1923; // @[VideoBuffer.scala 44:25]
  assign io_pixelVal_out = 8'hbf == _T_3[7:0] ? image_191 : _GEN_190; // @[VideoBuffer.scala 35:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  image_0 = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  image_1 = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  image_2 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  image_3 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  image_4 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  image_5 = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  image_6 = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  image_7 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  image_8 = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  image_9 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  image_10 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  image_11 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  image_12 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  image_13 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  image_14 = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  image_15 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  image_16 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  image_17 = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  image_18 = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  image_19 = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  image_20 = _RAND_20[3:0];
  _RAND_21 = {1{`RANDOM}};
  image_21 = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  image_22 = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  image_23 = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  image_24 = _RAND_24[3:0];
  _RAND_25 = {1{`RANDOM}};
  image_25 = _RAND_25[3:0];
  _RAND_26 = {1{`RANDOM}};
  image_26 = _RAND_26[3:0];
  _RAND_27 = {1{`RANDOM}};
  image_27 = _RAND_27[3:0];
  _RAND_28 = {1{`RANDOM}};
  image_28 = _RAND_28[3:0];
  _RAND_29 = {1{`RANDOM}};
  image_29 = _RAND_29[3:0];
  _RAND_30 = {1{`RANDOM}};
  image_30 = _RAND_30[3:0];
  _RAND_31 = {1{`RANDOM}};
  image_31 = _RAND_31[3:0];
  _RAND_32 = {1{`RANDOM}};
  image_32 = _RAND_32[3:0];
  _RAND_33 = {1{`RANDOM}};
  image_33 = _RAND_33[3:0];
  _RAND_34 = {1{`RANDOM}};
  image_34 = _RAND_34[3:0];
  _RAND_35 = {1{`RANDOM}};
  image_35 = _RAND_35[3:0];
  _RAND_36 = {1{`RANDOM}};
  image_36 = _RAND_36[3:0];
  _RAND_37 = {1{`RANDOM}};
  image_37 = _RAND_37[3:0];
  _RAND_38 = {1{`RANDOM}};
  image_38 = _RAND_38[3:0];
  _RAND_39 = {1{`RANDOM}};
  image_39 = _RAND_39[3:0];
  _RAND_40 = {1{`RANDOM}};
  image_40 = _RAND_40[3:0];
  _RAND_41 = {1{`RANDOM}};
  image_41 = _RAND_41[3:0];
  _RAND_42 = {1{`RANDOM}};
  image_42 = _RAND_42[3:0];
  _RAND_43 = {1{`RANDOM}};
  image_43 = _RAND_43[3:0];
  _RAND_44 = {1{`RANDOM}};
  image_44 = _RAND_44[3:0];
  _RAND_45 = {1{`RANDOM}};
  image_45 = _RAND_45[3:0];
  _RAND_46 = {1{`RANDOM}};
  image_46 = _RAND_46[3:0];
  _RAND_47 = {1{`RANDOM}};
  image_47 = _RAND_47[3:0];
  _RAND_48 = {1{`RANDOM}};
  image_48 = _RAND_48[3:0];
  _RAND_49 = {1{`RANDOM}};
  image_49 = _RAND_49[3:0];
  _RAND_50 = {1{`RANDOM}};
  image_50 = _RAND_50[3:0];
  _RAND_51 = {1{`RANDOM}};
  image_51 = _RAND_51[3:0];
  _RAND_52 = {1{`RANDOM}};
  image_52 = _RAND_52[3:0];
  _RAND_53 = {1{`RANDOM}};
  image_53 = _RAND_53[3:0];
  _RAND_54 = {1{`RANDOM}};
  image_54 = _RAND_54[3:0];
  _RAND_55 = {1{`RANDOM}};
  image_55 = _RAND_55[3:0];
  _RAND_56 = {1{`RANDOM}};
  image_56 = _RAND_56[3:0];
  _RAND_57 = {1{`RANDOM}};
  image_57 = _RAND_57[3:0];
  _RAND_58 = {1{`RANDOM}};
  image_58 = _RAND_58[3:0];
  _RAND_59 = {1{`RANDOM}};
  image_59 = _RAND_59[3:0];
  _RAND_60 = {1{`RANDOM}};
  image_60 = _RAND_60[3:0];
  _RAND_61 = {1{`RANDOM}};
  image_61 = _RAND_61[3:0];
  _RAND_62 = {1{`RANDOM}};
  image_62 = _RAND_62[3:0];
  _RAND_63 = {1{`RANDOM}};
  image_63 = _RAND_63[3:0];
  _RAND_64 = {1{`RANDOM}};
  image_64 = _RAND_64[3:0];
  _RAND_65 = {1{`RANDOM}};
  image_65 = _RAND_65[3:0];
  _RAND_66 = {1{`RANDOM}};
  image_66 = _RAND_66[3:0];
  _RAND_67 = {1{`RANDOM}};
  image_67 = _RAND_67[3:0];
  _RAND_68 = {1{`RANDOM}};
  image_68 = _RAND_68[3:0];
  _RAND_69 = {1{`RANDOM}};
  image_69 = _RAND_69[3:0];
  _RAND_70 = {1{`RANDOM}};
  image_70 = _RAND_70[3:0];
  _RAND_71 = {1{`RANDOM}};
  image_71 = _RAND_71[3:0];
  _RAND_72 = {1{`RANDOM}};
  image_72 = _RAND_72[3:0];
  _RAND_73 = {1{`RANDOM}};
  image_73 = _RAND_73[3:0];
  _RAND_74 = {1{`RANDOM}};
  image_74 = _RAND_74[3:0];
  _RAND_75 = {1{`RANDOM}};
  image_75 = _RAND_75[3:0];
  _RAND_76 = {1{`RANDOM}};
  image_76 = _RAND_76[3:0];
  _RAND_77 = {1{`RANDOM}};
  image_77 = _RAND_77[3:0];
  _RAND_78 = {1{`RANDOM}};
  image_78 = _RAND_78[3:0];
  _RAND_79 = {1{`RANDOM}};
  image_79 = _RAND_79[3:0];
  _RAND_80 = {1{`RANDOM}};
  image_80 = _RAND_80[3:0];
  _RAND_81 = {1{`RANDOM}};
  image_81 = _RAND_81[3:0];
  _RAND_82 = {1{`RANDOM}};
  image_82 = _RAND_82[3:0];
  _RAND_83 = {1{`RANDOM}};
  image_83 = _RAND_83[3:0];
  _RAND_84 = {1{`RANDOM}};
  image_84 = _RAND_84[3:0];
  _RAND_85 = {1{`RANDOM}};
  image_85 = _RAND_85[3:0];
  _RAND_86 = {1{`RANDOM}};
  image_86 = _RAND_86[3:0];
  _RAND_87 = {1{`RANDOM}};
  image_87 = _RAND_87[3:0];
  _RAND_88 = {1{`RANDOM}};
  image_88 = _RAND_88[3:0];
  _RAND_89 = {1{`RANDOM}};
  image_89 = _RAND_89[3:0];
  _RAND_90 = {1{`RANDOM}};
  image_90 = _RAND_90[3:0];
  _RAND_91 = {1{`RANDOM}};
  image_91 = _RAND_91[3:0];
  _RAND_92 = {1{`RANDOM}};
  image_92 = _RAND_92[3:0];
  _RAND_93 = {1{`RANDOM}};
  image_93 = _RAND_93[3:0];
  _RAND_94 = {1{`RANDOM}};
  image_94 = _RAND_94[3:0];
  _RAND_95 = {1{`RANDOM}};
  image_95 = _RAND_95[3:0];
  _RAND_96 = {1{`RANDOM}};
  image_96 = _RAND_96[3:0];
  _RAND_97 = {1{`RANDOM}};
  image_97 = _RAND_97[3:0];
  _RAND_98 = {1{`RANDOM}};
  image_98 = _RAND_98[3:0];
  _RAND_99 = {1{`RANDOM}};
  image_99 = _RAND_99[3:0];
  _RAND_100 = {1{`RANDOM}};
  image_100 = _RAND_100[3:0];
  _RAND_101 = {1{`RANDOM}};
  image_101 = _RAND_101[3:0];
  _RAND_102 = {1{`RANDOM}};
  image_102 = _RAND_102[3:0];
  _RAND_103 = {1{`RANDOM}};
  image_103 = _RAND_103[3:0];
  _RAND_104 = {1{`RANDOM}};
  image_104 = _RAND_104[3:0];
  _RAND_105 = {1{`RANDOM}};
  image_105 = _RAND_105[3:0];
  _RAND_106 = {1{`RANDOM}};
  image_106 = _RAND_106[3:0];
  _RAND_107 = {1{`RANDOM}};
  image_107 = _RAND_107[3:0];
  _RAND_108 = {1{`RANDOM}};
  image_108 = _RAND_108[3:0];
  _RAND_109 = {1{`RANDOM}};
  image_109 = _RAND_109[3:0];
  _RAND_110 = {1{`RANDOM}};
  image_110 = _RAND_110[3:0];
  _RAND_111 = {1{`RANDOM}};
  image_111 = _RAND_111[3:0];
  _RAND_112 = {1{`RANDOM}};
  image_112 = _RAND_112[3:0];
  _RAND_113 = {1{`RANDOM}};
  image_113 = _RAND_113[3:0];
  _RAND_114 = {1{`RANDOM}};
  image_114 = _RAND_114[3:0];
  _RAND_115 = {1{`RANDOM}};
  image_115 = _RAND_115[3:0];
  _RAND_116 = {1{`RANDOM}};
  image_116 = _RAND_116[3:0];
  _RAND_117 = {1{`RANDOM}};
  image_117 = _RAND_117[3:0];
  _RAND_118 = {1{`RANDOM}};
  image_118 = _RAND_118[3:0];
  _RAND_119 = {1{`RANDOM}};
  image_119 = _RAND_119[3:0];
  _RAND_120 = {1{`RANDOM}};
  image_120 = _RAND_120[3:0];
  _RAND_121 = {1{`RANDOM}};
  image_121 = _RAND_121[3:0];
  _RAND_122 = {1{`RANDOM}};
  image_122 = _RAND_122[3:0];
  _RAND_123 = {1{`RANDOM}};
  image_123 = _RAND_123[3:0];
  _RAND_124 = {1{`RANDOM}};
  image_124 = _RAND_124[3:0];
  _RAND_125 = {1{`RANDOM}};
  image_125 = _RAND_125[3:0];
  _RAND_126 = {1{`RANDOM}};
  image_126 = _RAND_126[3:0];
  _RAND_127 = {1{`RANDOM}};
  image_127 = _RAND_127[3:0];
  _RAND_128 = {1{`RANDOM}};
  image_128 = _RAND_128[3:0];
  _RAND_129 = {1{`RANDOM}};
  image_129 = _RAND_129[3:0];
  _RAND_130 = {1{`RANDOM}};
  image_130 = _RAND_130[3:0];
  _RAND_131 = {1{`RANDOM}};
  image_131 = _RAND_131[3:0];
  _RAND_132 = {1{`RANDOM}};
  image_132 = _RAND_132[3:0];
  _RAND_133 = {1{`RANDOM}};
  image_133 = _RAND_133[3:0];
  _RAND_134 = {1{`RANDOM}};
  image_134 = _RAND_134[3:0];
  _RAND_135 = {1{`RANDOM}};
  image_135 = _RAND_135[3:0];
  _RAND_136 = {1{`RANDOM}};
  image_136 = _RAND_136[3:0];
  _RAND_137 = {1{`RANDOM}};
  image_137 = _RAND_137[3:0];
  _RAND_138 = {1{`RANDOM}};
  image_138 = _RAND_138[3:0];
  _RAND_139 = {1{`RANDOM}};
  image_139 = _RAND_139[3:0];
  _RAND_140 = {1{`RANDOM}};
  image_140 = _RAND_140[3:0];
  _RAND_141 = {1{`RANDOM}};
  image_141 = _RAND_141[3:0];
  _RAND_142 = {1{`RANDOM}};
  image_142 = _RAND_142[3:0];
  _RAND_143 = {1{`RANDOM}};
  image_143 = _RAND_143[3:0];
  _RAND_144 = {1{`RANDOM}};
  image_144 = _RAND_144[3:0];
  _RAND_145 = {1{`RANDOM}};
  image_145 = _RAND_145[3:0];
  _RAND_146 = {1{`RANDOM}};
  image_146 = _RAND_146[3:0];
  _RAND_147 = {1{`RANDOM}};
  image_147 = _RAND_147[3:0];
  _RAND_148 = {1{`RANDOM}};
  image_148 = _RAND_148[3:0];
  _RAND_149 = {1{`RANDOM}};
  image_149 = _RAND_149[3:0];
  _RAND_150 = {1{`RANDOM}};
  image_150 = _RAND_150[3:0];
  _RAND_151 = {1{`RANDOM}};
  image_151 = _RAND_151[3:0];
  _RAND_152 = {1{`RANDOM}};
  image_152 = _RAND_152[3:0];
  _RAND_153 = {1{`RANDOM}};
  image_153 = _RAND_153[3:0];
  _RAND_154 = {1{`RANDOM}};
  image_154 = _RAND_154[3:0];
  _RAND_155 = {1{`RANDOM}};
  image_155 = _RAND_155[3:0];
  _RAND_156 = {1{`RANDOM}};
  image_156 = _RAND_156[3:0];
  _RAND_157 = {1{`RANDOM}};
  image_157 = _RAND_157[3:0];
  _RAND_158 = {1{`RANDOM}};
  image_158 = _RAND_158[3:0];
  _RAND_159 = {1{`RANDOM}};
  image_159 = _RAND_159[3:0];
  _RAND_160 = {1{`RANDOM}};
  image_160 = _RAND_160[3:0];
  _RAND_161 = {1{`RANDOM}};
  image_161 = _RAND_161[3:0];
  _RAND_162 = {1{`RANDOM}};
  image_162 = _RAND_162[3:0];
  _RAND_163 = {1{`RANDOM}};
  image_163 = _RAND_163[3:0];
  _RAND_164 = {1{`RANDOM}};
  image_164 = _RAND_164[3:0];
  _RAND_165 = {1{`RANDOM}};
  image_165 = _RAND_165[3:0];
  _RAND_166 = {1{`RANDOM}};
  image_166 = _RAND_166[3:0];
  _RAND_167 = {1{`RANDOM}};
  image_167 = _RAND_167[3:0];
  _RAND_168 = {1{`RANDOM}};
  image_168 = _RAND_168[3:0];
  _RAND_169 = {1{`RANDOM}};
  image_169 = _RAND_169[3:0];
  _RAND_170 = {1{`RANDOM}};
  image_170 = _RAND_170[3:0];
  _RAND_171 = {1{`RANDOM}};
  image_171 = _RAND_171[3:0];
  _RAND_172 = {1{`RANDOM}};
  image_172 = _RAND_172[3:0];
  _RAND_173 = {1{`RANDOM}};
  image_173 = _RAND_173[3:0];
  _RAND_174 = {1{`RANDOM}};
  image_174 = _RAND_174[3:0];
  _RAND_175 = {1{`RANDOM}};
  image_175 = _RAND_175[3:0];
  _RAND_176 = {1{`RANDOM}};
  image_176 = _RAND_176[3:0];
  _RAND_177 = {1{`RANDOM}};
  image_177 = _RAND_177[3:0];
  _RAND_178 = {1{`RANDOM}};
  image_178 = _RAND_178[3:0];
  _RAND_179 = {1{`RANDOM}};
  image_179 = _RAND_179[3:0];
  _RAND_180 = {1{`RANDOM}};
  image_180 = _RAND_180[3:0];
  _RAND_181 = {1{`RANDOM}};
  image_181 = _RAND_181[3:0];
  _RAND_182 = {1{`RANDOM}};
  image_182 = _RAND_182[3:0];
  _RAND_183 = {1{`RANDOM}};
  image_183 = _RAND_183[3:0];
  _RAND_184 = {1{`RANDOM}};
  image_184 = _RAND_184[3:0];
  _RAND_185 = {1{`RANDOM}};
  image_185 = _RAND_185[3:0];
  _RAND_186 = {1{`RANDOM}};
  image_186 = _RAND_186[3:0];
  _RAND_187 = {1{`RANDOM}};
  image_187 = _RAND_187[3:0];
  _RAND_188 = {1{`RANDOM}};
  image_188 = _RAND_188[3:0];
  _RAND_189 = {1{`RANDOM}};
  image_189 = _RAND_189[3:0];
  _RAND_190 = {1{`RANDOM}};
  image_190 = _RAND_190[3:0];
  _RAND_191 = {1{`RANDOM}};
  image_191 = _RAND_191[3:0];
  _RAND_192 = {1{`RANDOM}};
  pixelIndex = _RAND_192[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      image_0 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h0 == _T_27[7:0]) begin
        image_0 <= io_pixelVal_in_7;
      end else if (8'h0 == _T_24[7:0]) begin
        image_0 <= io_pixelVal_in_6;
      end else if (8'h0 == _T_21[7:0]) begin
        image_0 <= io_pixelVal_in_5;
      end else if (8'h0 == _T_18[7:0]) begin
        image_0 <= io_pixelVal_in_4;
      end else if (8'h0 == _T_15[7:0]) begin
        image_0 <= io_pixelVal_in_3;
      end else if (8'h0 == _T_12[7:0]) begin
        image_0 <= io_pixelVal_in_2;
      end else if (8'h0 == _T_9[7:0]) begin
        image_0 <= io_pixelVal_in_1;
      end else if (8'h0 == _T_5[7:0]) begin
        image_0 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_1 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1 == _T_27[7:0]) begin
        image_1 <= io_pixelVal_in_7;
      end else if (8'h1 == _T_24[7:0]) begin
        image_1 <= io_pixelVal_in_6;
      end else if (8'h1 == _T_21[7:0]) begin
        image_1 <= io_pixelVal_in_5;
      end else if (8'h1 == _T_18[7:0]) begin
        image_1 <= io_pixelVal_in_4;
      end else if (8'h1 == _T_15[7:0]) begin
        image_1 <= io_pixelVal_in_3;
      end else if (8'h1 == _T_12[7:0]) begin
        image_1 <= io_pixelVal_in_2;
      end else if (8'h1 == _T_9[7:0]) begin
        image_1 <= io_pixelVal_in_1;
      end else if (8'h1 == _T_5[7:0]) begin
        image_1 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_2 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h2 == _T_27[7:0]) begin
        image_2 <= io_pixelVal_in_7;
      end else if (8'h2 == _T_24[7:0]) begin
        image_2 <= io_pixelVal_in_6;
      end else if (8'h2 == _T_21[7:0]) begin
        image_2 <= io_pixelVal_in_5;
      end else if (8'h2 == _T_18[7:0]) begin
        image_2 <= io_pixelVal_in_4;
      end else if (8'h2 == _T_15[7:0]) begin
        image_2 <= io_pixelVal_in_3;
      end else if (8'h2 == _T_12[7:0]) begin
        image_2 <= io_pixelVal_in_2;
      end else if (8'h2 == _T_9[7:0]) begin
        image_2 <= io_pixelVal_in_1;
      end else if (8'h2 == _T_5[7:0]) begin
        image_2 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_3 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h3 == _T_27[7:0]) begin
        image_3 <= io_pixelVal_in_7;
      end else if (8'h3 == _T_24[7:0]) begin
        image_3 <= io_pixelVal_in_6;
      end else if (8'h3 == _T_21[7:0]) begin
        image_3 <= io_pixelVal_in_5;
      end else if (8'h3 == _T_18[7:0]) begin
        image_3 <= io_pixelVal_in_4;
      end else if (8'h3 == _T_15[7:0]) begin
        image_3 <= io_pixelVal_in_3;
      end else if (8'h3 == _T_12[7:0]) begin
        image_3 <= io_pixelVal_in_2;
      end else if (8'h3 == _T_9[7:0]) begin
        image_3 <= io_pixelVal_in_1;
      end else if (8'h3 == _T_5[7:0]) begin
        image_3 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_4 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h4 == _T_27[7:0]) begin
        image_4 <= io_pixelVal_in_7;
      end else if (8'h4 == _T_24[7:0]) begin
        image_4 <= io_pixelVal_in_6;
      end else if (8'h4 == _T_21[7:0]) begin
        image_4 <= io_pixelVal_in_5;
      end else if (8'h4 == _T_18[7:0]) begin
        image_4 <= io_pixelVal_in_4;
      end else if (8'h4 == _T_15[7:0]) begin
        image_4 <= io_pixelVal_in_3;
      end else if (8'h4 == _T_12[7:0]) begin
        image_4 <= io_pixelVal_in_2;
      end else if (8'h4 == _T_9[7:0]) begin
        image_4 <= io_pixelVal_in_1;
      end else if (8'h4 == _T_5[7:0]) begin
        image_4 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_5 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h5 == _T_27[7:0]) begin
        image_5 <= io_pixelVal_in_7;
      end else if (8'h5 == _T_24[7:0]) begin
        image_5 <= io_pixelVal_in_6;
      end else if (8'h5 == _T_21[7:0]) begin
        image_5 <= io_pixelVal_in_5;
      end else if (8'h5 == _T_18[7:0]) begin
        image_5 <= io_pixelVal_in_4;
      end else if (8'h5 == _T_15[7:0]) begin
        image_5 <= io_pixelVal_in_3;
      end else if (8'h5 == _T_12[7:0]) begin
        image_5 <= io_pixelVal_in_2;
      end else if (8'h5 == _T_9[7:0]) begin
        image_5 <= io_pixelVal_in_1;
      end else if (8'h5 == _T_5[7:0]) begin
        image_5 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_6 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h6 == _T_27[7:0]) begin
        image_6 <= io_pixelVal_in_7;
      end else if (8'h6 == _T_24[7:0]) begin
        image_6 <= io_pixelVal_in_6;
      end else if (8'h6 == _T_21[7:0]) begin
        image_6 <= io_pixelVal_in_5;
      end else if (8'h6 == _T_18[7:0]) begin
        image_6 <= io_pixelVal_in_4;
      end else if (8'h6 == _T_15[7:0]) begin
        image_6 <= io_pixelVal_in_3;
      end else if (8'h6 == _T_12[7:0]) begin
        image_6 <= io_pixelVal_in_2;
      end else if (8'h6 == _T_9[7:0]) begin
        image_6 <= io_pixelVal_in_1;
      end else if (8'h6 == _T_5[7:0]) begin
        image_6 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_7 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h7 == _T_27[7:0]) begin
        image_7 <= io_pixelVal_in_7;
      end else if (8'h7 == _T_24[7:0]) begin
        image_7 <= io_pixelVal_in_6;
      end else if (8'h7 == _T_21[7:0]) begin
        image_7 <= io_pixelVal_in_5;
      end else if (8'h7 == _T_18[7:0]) begin
        image_7 <= io_pixelVal_in_4;
      end else if (8'h7 == _T_15[7:0]) begin
        image_7 <= io_pixelVal_in_3;
      end else if (8'h7 == _T_12[7:0]) begin
        image_7 <= io_pixelVal_in_2;
      end else if (8'h7 == _T_9[7:0]) begin
        image_7 <= io_pixelVal_in_1;
      end else if (8'h7 == _T_5[7:0]) begin
        image_7 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_8 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h8 == _T_27[7:0]) begin
        image_8 <= io_pixelVal_in_7;
      end else if (8'h8 == _T_24[7:0]) begin
        image_8 <= io_pixelVal_in_6;
      end else if (8'h8 == _T_21[7:0]) begin
        image_8 <= io_pixelVal_in_5;
      end else if (8'h8 == _T_18[7:0]) begin
        image_8 <= io_pixelVal_in_4;
      end else if (8'h8 == _T_15[7:0]) begin
        image_8 <= io_pixelVal_in_3;
      end else if (8'h8 == _T_12[7:0]) begin
        image_8 <= io_pixelVal_in_2;
      end else if (8'h8 == _T_9[7:0]) begin
        image_8 <= io_pixelVal_in_1;
      end else if (8'h8 == _T_5[7:0]) begin
        image_8 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_9 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h9 == _T_27[7:0]) begin
        image_9 <= io_pixelVal_in_7;
      end else if (8'h9 == _T_24[7:0]) begin
        image_9 <= io_pixelVal_in_6;
      end else if (8'h9 == _T_21[7:0]) begin
        image_9 <= io_pixelVal_in_5;
      end else if (8'h9 == _T_18[7:0]) begin
        image_9 <= io_pixelVal_in_4;
      end else if (8'h9 == _T_15[7:0]) begin
        image_9 <= io_pixelVal_in_3;
      end else if (8'h9 == _T_12[7:0]) begin
        image_9 <= io_pixelVal_in_2;
      end else if (8'h9 == _T_9[7:0]) begin
        image_9 <= io_pixelVal_in_1;
      end else if (8'h9 == _T_5[7:0]) begin
        image_9 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_10 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'ha == _T_27[7:0]) begin
        image_10 <= io_pixelVal_in_7;
      end else if (8'ha == _T_24[7:0]) begin
        image_10 <= io_pixelVal_in_6;
      end else if (8'ha == _T_21[7:0]) begin
        image_10 <= io_pixelVal_in_5;
      end else if (8'ha == _T_18[7:0]) begin
        image_10 <= io_pixelVal_in_4;
      end else if (8'ha == _T_15[7:0]) begin
        image_10 <= io_pixelVal_in_3;
      end else if (8'ha == _T_12[7:0]) begin
        image_10 <= io_pixelVal_in_2;
      end else if (8'ha == _T_9[7:0]) begin
        image_10 <= io_pixelVal_in_1;
      end else if (8'ha == _T_5[7:0]) begin
        image_10 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_11 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'hb == _T_27[7:0]) begin
        image_11 <= io_pixelVal_in_7;
      end else if (8'hb == _T_24[7:0]) begin
        image_11 <= io_pixelVal_in_6;
      end else if (8'hb == _T_21[7:0]) begin
        image_11 <= io_pixelVal_in_5;
      end else if (8'hb == _T_18[7:0]) begin
        image_11 <= io_pixelVal_in_4;
      end else if (8'hb == _T_15[7:0]) begin
        image_11 <= io_pixelVal_in_3;
      end else if (8'hb == _T_12[7:0]) begin
        image_11 <= io_pixelVal_in_2;
      end else if (8'hb == _T_9[7:0]) begin
        image_11 <= io_pixelVal_in_1;
      end else if (8'hb == _T_5[7:0]) begin
        image_11 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_12 <= 4'h4;
    end else if (io_valid_in) begin
      if (8'hc == _T_27[7:0]) begin
        image_12 <= io_pixelVal_in_7;
      end else if (8'hc == _T_24[7:0]) begin
        image_12 <= io_pixelVal_in_6;
      end else if (8'hc == _T_21[7:0]) begin
        image_12 <= io_pixelVal_in_5;
      end else if (8'hc == _T_18[7:0]) begin
        image_12 <= io_pixelVal_in_4;
      end else if (8'hc == _T_15[7:0]) begin
        image_12 <= io_pixelVal_in_3;
      end else if (8'hc == _T_12[7:0]) begin
        image_12 <= io_pixelVal_in_2;
      end else if (8'hc == _T_9[7:0]) begin
        image_12 <= io_pixelVal_in_1;
      end else if (8'hc == _T_5[7:0]) begin
        image_12 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_13 <= 4'h1;
    end else if (io_valid_in) begin
      if (8'hd == _T_27[7:0]) begin
        image_13 <= io_pixelVal_in_7;
      end else if (8'hd == _T_24[7:0]) begin
        image_13 <= io_pixelVal_in_6;
      end else if (8'hd == _T_21[7:0]) begin
        image_13 <= io_pixelVal_in_5;
      end else if (8'hd == _T_18[7:0]) begin
        image_13 <= io_pixelVal_in_4;
      end else if (8'hd == _T_15[7:0]) begin
        image_13 <= io_pixelVal_in_3;
      end else if (8'hd == _T_12[7:0]) begin
        image_13 <= io_pixelVal_in_2;
      end else if (8'hd == _T_9[7:0]) begin
        image_13 <= io_pixelVal_in_1;
      end else if (8'hd == _T_5[7:0]) begin
        image_13 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_14 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he == _T_27[7:0]) begin
        image_14 <= io_pixelVal_in_7;
      end else if (8'he == _T_24[7:0]) begin
        image_14 <= io_pixelVal_in_6;
      end else if (8'he == _T_21[7:0]) begin
        image_14 <= io_pixelVal_in_5;
      end else if (8'he == _T_18[7:0]) begin
        image_14 <= io_pixelVal_in_4;
      end else if (8'he == _T_15[7:0]) begin
        image_14 <= io_pixelVal_in_3;
      end else if (8'he == _T_12[7:0]) begin
        image_14 <= io_pixelVal_in_2;
      end else if (8'he == _T_9[7:0]) begin
        image_14 <= io_pixelVal_in_1;
      end else if (8'he == _T_5[7:0]) begin
        image_14 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_15 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf == _T_27[7:0]) begin
        image_15 <= io_pixelVal_in_7;
      end else if (8'hf == _T_24[7:0]) begin
        image_15 <= io_pixelVal_in_6;
      end else if (8'hf == _T_21[7:0]) begin
        image_15 <= io_pixelVal_in_5;
      end else if (8'hf == _T_18[7:0]) begin
        image_15 <= io_pixelVal_in_4;
      end else if (8'hf == _T_15[7:0]) begin
        image_15 <= io_pixelVal_in_3;
      end else if (8'hf == _T_12[7:0]) begin
        image_15 <= io_pixelVal_in_2;
      end else if (8'hf == _T_9[7:0]) begin
        image_15 <= io_pixelVal_in_1;
      end else if (8'hf == _T_5[7:0]) begin
        image_15 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_16 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h10 == _T_27[7:0]) begin
        image_16 <= io_pixelVal_in_7;
      end else if (8'h10 == _T_24[7:0]) begin
        image_16 <= io_pixelVal_in_6;
      end else if (8'h10 == _T_21[7:0]) begin
        image_16 <= io_pixelVal_in_5;
      end else if (8'h10 == _T_18[7:0]) begin
        image_16 <= io_pixelVal_in_4;
      end else if (8'h10 == _T_15[7:0]) begin
        image_16 <= io_pixelVal_in_3;
      end else if (8'h10 == _T_12[7:0]) begin
        image_16 <= io_pixelVal_in_2;
      end else if (8'h10 == _T_9[7:0]) begin
        image_16 <= io_pixelVal_in_1;
      end else if (8'h10 == _T_5[7:0]) begin
        image_16 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_17 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h11 == _T_27[7:0]) begin
        image_17 <= io_pixelVal_in_7;
      end else if (8'h11 == _T_24[7:0]) begin
        image_17 <= io_pixelVal_in_6;
      end else if (8'h11 == _T_21[7:0]) begin
        image_17 <= io_pixelVal_in_5;
      end else if (8'h11 == _T_18[7:0]) begin
        image_17 <= io_pixelVal_in_4;
      end else if (8'h11 == _T_15[7:0]) begin
        image_17 <= io_pixelVal_in_3;
      end else if (8'h11 == _T_12[7:0]) begin
        image_17 <= io_pixelVal_in_2;
      end else if (8'h11 == _T_9[7:0]) begin
        image_17 <= io_pixelVal_in_1;
      end else if (8'h11 == _T_5[7:0]) begin
        image_17 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_18 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h12 == _T_27[7:0]) begin
        image_18 <= io_pixelVal_in_7;
      end else if (8'h12 == _T_24[7:0]) begin
        image_18 <= io_pixelVal_in_6;
      end else if (8'h12 == _T_21[7:0]) begin
        image_18 <= io_pixelVal_in_5;
      end else if (8'h12 == _T_18[7:0]) begin
        image_18 <= io_pixelVal_in_4;
      end else if (8'h12 == _T_15[7:0]) begin
        image_18 <= io_pixelVal_in_3;
      end else if (8'h12 == _T_12[7:0]) begin
        image_18 <= io_pixelVal_in_2;
      end else if (8'h12 == _T_9[7:0]) begin
        image_18 <= io_pixelVal_in_1;
      end else if (8'h12 == _T_5[7:0]) begin
        image_18 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_19 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h13 == _T_27[7:0]) begin
        image_19 <= io_pixelVal_in_7;
      end else if (8'h13 == _T_24[7:0]) begin
        image_19 <= io_pixelVal_in_6;
      end else if (8'h13 == _T_21[7:0]) begin
        image_19 <= io_pixelVal_in_5;
      end else if (8'h13 == _T_18[7:0]) begin
        image_19 <= io_pixelVal_in_4;
      end else if (8'h13 == _T_15[7:0]) begin
        image_19 <= io_pixelVal_in_3;
      end else if (8'h13 == _T_12[7:0]) begin
        image_19 <= io_pixelVal_in_2;
      end else if (8'h13 == _T_9[7:0]) begin
        image_19 <= io_pixelVal_in_1;
      end else if (8'h13 == _T_5[7:0]) begin
        image_19 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_20 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h14 == _T_27[7:0]) begin
        image_20 <= io_pixelVal_in_7;
      end else if (8'h14 == _T_24[7:0]) begin
        image_20 <= io_pixelVal_in_6;
      end else if (8'h14 == _T_21[7:0]) begin
        image_20 <= io_pixelVal_in_5;
      end else if (8'h14 == _T_18[7:0]) begin
        image_20 <= io_pixelVal_in_4;
      end else if (8'h14 == _T_15[7:0]) begin
        image_20 <= io_pixelVal_in_3;
      end else if (8'h14 == _T_12[7:0]) begin
        image_20 <= io_pixelVal_in_2;
      end else if (8'h14 == _T_9[7:0]) begin
        image_20 <= io_pixelVal_in_1;
      end else if (8'h14 == _T_5[7:0]) begin
        image_20 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_21 <= 4'h7;
    end else if (io_valid_in) begin
      if (8'h15 == _T_27[7:0]) begin
        image_21 <= io_pixelVal_in_7;
      end else if (8'h15 == _T_24[7:0]) begin
        image_21 <= io_pixelVal_in_6;
      end else if (8'h15 == _T_21[7:0]) begin
        image_21 <= io_pixelVal_in_5;
      end else if (8'h15 == _T_18[7:0]) begin
        image_21 <= io_pixelVal_in_4;
      end else if (8'h15 == _T_15[7:0]) begin
        image_21 <= io_pixelVal_in_3;
      end else if (8'h15 == _T_12[7:0]) begin
        image_21 <= io_pixelVal_in_2;
      end else if (8'h15 == _T_9[7:0]) begin
        image_21 <= io_pixelVal_in_1;
      end else if (8'h15 == _T_5[7:0]) begin
        image_21 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_22 <= 4'ha;
    end else if (io_valid_in) begin
      if (8'h16 == _T_27[7:0]) begin
        image_22 <= io_pixelVal_in_7;
      end else if (8'h16 == _T_24[7:0]) begin
        image_22 <= io_pixelVal_in_6;
      end else if (8'h16 == _T_21[7:0]) begin
        image_22 <= io_pixelVal_in_5;
      end else if (8'h16 == _T_18[7:0]) begin
        image_22 <= io_pixelVal_in_4;
      end else if (8'h16 == _T_15[7:0]) begin
        image_22 <= io_pixelVal_in_3;
      end else if (8'h16 == _T_12[7:0]) begin
        image_22 <= io_pixelVal_in_2;
      end else if (8'h16 == _T_9[7:0]) begin
        image_22 <= io_pixelVal_in_1;
      end else if (8'h16 == _T_5[7:0]) begin
        image_22 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_23 <= 4'hb;
    end else if (io_valid_in) begin
      if (8'h17 == _T_27[7:0]) begin
        image_23 <= io_pixelVal_in_7;
      end else if (8'h17 == _T_24[7:0]) begin
        image_23 <= io_pixelVal_in_6;
      end else if (8'h17 == _T_21[7:0]) begin
        image_23 <= io_pixelVal_in_5;
      end else if (8'h17 == _T_18[7:0]) begin
        image_23 <= io_pixelVal_in_4;
      end else if (8'h17 == _T_15[7:0]) begin
        image_23 <= io_pixelVal_in_3;
      end else if (8'h17 == _T_12[7:0]) begin
        image_23 <= io_pixelVal_in_2;
      end else if (8'h17 == _T_9[7:0]) begin
        image_23 <= io_pixelVal_in_1;
      end else if (8'h17 == _T_5[7:0]) begin
        image_23 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_24 <= 4'h9;
    end else if (io_valid_in) begin
      if (8'h18 == _T_27[7:0]) begin
        image_24 <= io_pixelVal_in_7;
      end else if (8'h18 == _T_24[7:0]) begin
        image_24 <= io_pixelVal_in_6;
      end else if (8'h18 == _T_21[7:0]) begin
        image_24 <= io_pixelVal_in_5;
      end else if (8'h18 == _T_18[7:0]) begin
        image_24 <= io_pixelVal_in_4;
      end else if (8'h18 == _T_15[7:0]) begin
        image_24 <= io_pixelVal_in_3;
      end else if (8'h18 == _T_12[7:0]) begin
        image_24 <= io_pixelVal_in_2;
      end else if (8'h18 == _T_9[7:0]) begin
        image_24 <= io_pixelVal_in_1;
      end else if (8'h18 == _T_5[7:0]) begin
        image_24 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_25 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h19 == _T_27[7:0]) begin
        image_25 <= io_pixelVal_in_7;
      end else if (8'h19 == _T_24[7:0]) begin
        image_25 <= io_pixelVal_in_6;
      end else if (8'h19 == _T_21[7:0]) begin
        image_25 <= io_pixelVal_in_5;
      end else if (8'h19 == _T_18[7:0]) begin
        image_25 <= io_pixelVal_in_4;
      end else if (8'h19 == _T_15[7:0]) begin
        image_25 <= io_pixelVal_in_3;
      end else if (8'h19 == _T_12[7:0]) begin
        image_25 <= io_pixelVal_in_2;
      end else if (8'h19 == _T_9[7:0]) begin
        image_25 <= io_pixelVal_in_1;
      end else if (8'h19 == _T_5[7:0]) begin
        image_25 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_26 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h1a == _T_27[7:0]) begin
        image_26 <= io_pixelVal_in_7;
      end else if (8'h1a == _T_24[7:0]) begin
        image_26 <= io_pixelVal_in_6;
      end else if (8'h1a == _T_21[7:0]) begin
        image_26 <= io_pixelVal_in_5;
      end else if (8'h1a == _T_18[7:0]) begin
        image_26 <= io_pixelVal_in_4;
      end else if (8'h1a == _T_15[7:0]) begin
        image_26 <= io_pixelVal_in_3;
      end else if (8'h1a == _T_12[7:0]) begin
        image_26 <= io_pixelVal_in_2;
      end else if (8'h1a == _T_9[7:0]) begin
        image_26 <= io_pixelVal_in_1;
      end else if (8'h1a == _T_5[7:0]) begin
        image_26 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_27 <= 4'ha;
    end else if (io_valid_in) begin
      if (8'h1b == _T_27[7:0]) begin
        image_27 <= io_pixelVal_in_7;
      end else if (8'h1b == _T_24[7:0]) begin
        image_27 <= io_pixelVal_in_6;
      end else if (8'h1b == _T_21[7:0]) begin
        image_27 <= io_pixelVal_in_5;
      end else if (8'h1b == _T_18[7:0]) begin
        image_27 <= io_pixelVal_in_4;
      end else if (8'h1b == _T_15[7:0]) begin
        image_27 <= io_pixelVal_in_3;
      end else if (8'h1b == _T_12[7:0]) begin
        image_27 <= io_pixelVal_in_2;
      end else if (8'h1b == _T_9[7:0]) begin
        image_27 <= io_pixelVal_in_1;
      end else if (8'h1b == _T_5[7:0]) begin
        image_27 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_28 <= 4'hd;
    end else if (io_valid_in) begin
      if (8'h1c == _T_27[7:0]) begin
        image_28 <= io_pixelVal_in_7;
      end else if (8'h1c == _T_24[7:0]) begin
        image_28 <= io_pixelVal_in_6;
      end else if (8'h1c == _T_21[7:0]) begin
        image_28 <= io_pixelVal_in_5;
      end else if (8'h1c == _T_18[7:0]) begin
        image_28 <= io_pixelVal_in_4;
      end else if (8'h1c == _T_15[7:0]) begin
        image_28 <= io_pixelVal_in_3;
      end else if (8'h1c == _T_12[7:0]) begin
        image_28 <= io_pixelVal_in_2;
      end else if (8'h1c == _T_9[7:0]) begin
        image_28 <= io_pixelVal_in_1;
      end else if (8'h1c == _T_5[7:0]) begin
        image_28 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_29 <= 4'hc;
    end else if (io_valid_in) begin
      if (8'h1d == _T_27[7:0]) begin
        image_29 <= io_pixelVal_in_7;
      end else if (8'h1d == _T_24[7:0]) begin
        image_29 <= io_pixelVal_in_6;
      end else if (8'h1d == _T_21[7:0]) begin
        image_29 <= io_pixelVal_in_5;
      end else if (8'h1d == _T_18[7:0]) begin
        image_29 <= io_pixelVal_in_4;
      end else if (8'h1d == _T_15[7:0]) begin
        image_29 <= io_pixelVal_in_3;
      end else if (8'h1d == _T_12[7:0]) begin
        image_29 <= io_pixelVal_in_2;
      end else if (8'h1d == _T_9[7:0]) begin
        image_29 <= io_pixelVal_in_1;
      end else if (8'h1d == _T_5[7:0]) begin
        image_29 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_30 <= 4'ha;
    end else if (io_valid_in) begin
      if (8'h1e == _T_27[7:0]) begin
        image_30 <= io_pixelVal_in_7;
      end else if (8'h1e == _T_24[7:0]) begin
        image_30 <= io_pixelVal_in_6;
      end else if (8'h1e == _T_21[7:0]) begin
        image_30 <= io_pixelVal_in_5;
      end else if (8'h1e == _T_18[7:0]) begin
        image_30 <= io_pixelVal_in_4;
      end else if (8'h1e == _T_15[7:0]) begin
        image_30 <= io_pixelVal_in_3;
      end else if (8'h1e == _T_12[7:0]) begin
        image_30 <= io_pixelVal_in_2;
      end else if (8'h1e == _T_9[7:0]) begin
        image_30 <= io_pixelVal_in_1;
      end else if (8'h1e == _T_5[7:0]) begin
        image_30 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_31 <= 4'h1;
    end else if (io_valid_in) begin
      if (8'h1f == _T_27[7:0]) begin
        image_31 <= io_pixelVal_in_7;
      end else if (8'h1f == _T_24[7:0]) begin
        image_31 <= io_pixelVal_in_6;
      end else if (8'h1f == _T_21[7:0]) begin
        image_31 <= io_pixelVal_in_5;
      end else if (8'h1f == _T_18[7:0]) begin
        image_31 <= io_pixelVal_in_4;
      end else if (8'h1f == _T_15[7:0]) begin
        image_31 <= io_pixelVal_in_3;
      end else if (8'h1f == _T_12[7:0]) begin
        image_31 <= io_pixelVal_in_2;
      end else if (8'h1f == _T_9[7:0]) begin
        image_31 <= io_pixelVal_in_1;
      end else if (8'h1f == _T_5[7:0]) begin
        image_31 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_32 <= 4'h4;
    end else if (io_valid_in) begin
      if (8'h20 == _T_27[7:0]) begin
        image_32 <= io_pixelVal_in_7;
      end else if (8'h20 == _T_24[7:0]) begin
        image_32 <= io_pixelVal_in_6;
      end else if (8'h20 == _T_21[7:0]) begin
        image_32 <= io_pixelVal_in_5;
      end else if (8'h20 == _T_18[7:0]) begin
        image_32 <= io_pixelVal_in_4;
      end else if (8'h20 == _T_15[7:0]) begin
        image_32 <= io_pixelVal_in_3;
      end else if (8'h20 == _T_12[7:0]) begin
        image_32 <= io_pixelVal_in_2;
      end else if (8'h20 == _T_9[7:0]) begin
        image_32 <= io_pixelVal_in_1;
      end else if (8'h20 == _T_5[7:0]) begin
        image_32 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_33 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h21 == _T_27[7:0]) begin
        image_33 <= io_pixelVal_in_7;
      end else if (8'h21 == _T_24[7:0]) begin
        image_33 <= io_pixelVal_in_6;
      end else if (8'h21 == _T_21[7:0]) begin
        image_33 <= io_pixelVal_in_5;
      end else if (8'h21 == _T_18[7:0]) begin
        image_33 <= io_pixelVal_in_4;
      end else if (8'h21 == _T_15[7:0]) begin
        image_33 <= io_pixelVal_in_3;
      end else if (8'h21 == _T_12[7:0]) begin
        image_33 <= io_pixelVal_in_2;
      end else if (8'h21 == _T_9[7:0]) begin
        image_33 <= io_pixelVal_in_1;
      end else if (8'h21 == _T_5[7:0]) begin
        image_33 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_34 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h22 == _T_27[7:0]) begin
        image_34 <= io_pixelVal_in_7;
      end else if (8'h22 == _T_24[7:0]) begin
        image_34 <= io_pixelVal_in_6;
      end else if (8'h22 == _T_21[7:0]) begin
        image_34 <= io_pixelVal_in_5;
      end else if (8'h22 == _T_18[7:0]) begin
        image_34 <= io_pixelVal_in_4;
      end else if (8'h22 == _T_15[7:0]) begin
        image_34 <= io_pixelVal_in_3;
      end else if (8'h22 == _T_12[7:0]) begin
        image_34 <= io_pixelVal_in_2;
      end else if (8'h22 == _T_9[7:0]) begin
        image_34 <= io_pixelVal_in_1;
      end else if (8'h22 == _T_5[7:0]) begin
        image_34 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_35 <= 4'h7;
    end else if (io_valid_in) begin
      if (8'h23 == _T_27[7:0]) begin
        image_35 <= io_pixelVal_in_7;
      end else if (8'h23 == _T_24[7:0]) begin
        image_35 <= io_pixelVal_in_6;
      end else if (8'h23 == _T_21[7:0]) begin
        image_35 <= io_pixelVal_in_5;
      end else if (8'h23 == _T_18[7:0]) begin
        image_35 <= io_pixelVal_in_4;
      end else if (8'h23 == _T_15[7:0]) begin
        image_35 <= io_pixelVal_in_3;
      end else if (8'h23 == _T_12[7:0]) begin
        image_35 <= io_pixelVal_in_2;
      end else if (8'h23 == _T_9[7:0]) begin
        image_35 <= io_pixelVal_in_1;
      end else if (8'h23 == _T_5[7:0]) begin
        image_35 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_36 <= 4'hb;
    end else if (io_valid_in) begin
      if (8'h24 == _T_27[7:0]) begin
        image_36 <= io_pixelVal_in_7;
      end else if (8'h24 == _T_24[7:0]) begin
        image_36 <= io_pixelVal_in_6;
      end else if (8'h24 == _T_21[7:0]) begin
        image_36 <= io_pixelVal_in_5;
      end else if (8'h24 == _T_18[7:0]) begin
        image_36 <= io_pixelVal_in_4;
      end else if (8'h24 == _T_15[7:0]) begin
        image_36 <= io_pixelVal_in_3;
      end else if (8'h24 == _T_12[7:0]) begin
        image_36 <= io_pixelVal_in_2;
      end else if (8'h24 == _T_9[7:0]) begin
        image_36 <= io_pixelVal_in_1;
      end else if (8'h24 == _T_5[7:0]) begin
        image_36 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_37 <= 4'he;
    end else if (io_valid_in) begin
      if (8'h25 == _T_27[7:0]) begin
        image_37 <= io_pixelVal_in_7;
      end else if (8'h25 == _T_24[7:0]) begin
        image_37 <= io_pixelVal_in_6;
      end else if (8'h25 == _T_21[7:0]) begin
        image_37 <= io_pixelVal_in_5;
      end else if (8'h25 == _T_18[7:0]) begin
        image_37 <= io_pixelVal_in_4;
      end else if (8'h25 == _T_15[7:0]) begin
        image_37 <= io_pixelVal_in_3;
      end else if (8'h25 == _T_12[7:0]) begin
        image_37 <= io_pixelVal_in_2;
      end else if (8'h25 == _T_9[7:0]) begin
        image_37 <= io_pixelVal_in_1;
      end else if (8'h25 == _T_5[7:0]) begin
        image_37 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_38 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h26 == _T_27[7:0]) begin
        image_38 <= io_pixelVal_in_7;
      end else if (8'h26 == _T_24[7:0]) begin
        image_38 <= io_pixelVal_in_6;
      end else if (8'h26 == _T_21[7:0]) begin
        image_38 <= io_pixelVal_in_5;
      end else if (8'h26 == _T_18[7:0]) begin
        image_38 <= io_pixelVal_in_4;
      end else if (8'h26 == _T_15[7:0]) begin
        image_38 <= io_pixelVal_in_3;
      end else if (8'h26 == _T_12[7:0]) begin
        image_38 <= io_pixelVal_in_2;
      end else if (8'h26 == _T_9[7:0]) begin
        image_38 <= io_pixelVal_in_1;
      end else if (8'h26 == _T_5[7:0]) begin
        image_38 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_39 <= 4'hc;
    end else if (io_valid_in) begin
      if (8'h27 == _T_27[7:0]) begin
        image_39 <= io_pixelVal_in_7;
      end else if (8'h27 == _T_24[7:0]) begin
        image_39 <= io_pixelVal_in_6;
      end else if (8'h27 == _T_21[7:0]) begin
        image_39 <= io_pixelVal_in_5;
      end else if (8'h27 == _T_18[7:0]) begin
        image_39 <= io_pixelVal_in_4;
      end else if (8'h27 == _T_15[7:0]) begin
        image_39 <= io_pixelVal_in_3;
      end else if (8'h27 == _T_12[7:0]) begin
        image_39 <= io_pixelVal_in_2;
      end else if (8'h27 == _T_9[7:0]) begin
        image_39 <= io_pixelVal_in_1;
      end else if (8'h27 == _T_5[7:0]) begin
        image_39 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_40 <= 4'h7;
    end else if (io_valid_in) begin
      if (8'h28 == _T_27[7:0]) begin
        image_40 <= io_pixelVal_in_7;
      end else if (8'h28 == _T_24[7:0]) begin
        image_40 <= io_pixelVal_in_6;
      end else if (8'h28 == _T_21[7:0]) begin
        image_40 <= io_pixelVal_in_5;
      end else if (8'h28 == _T_18[7:0]) begin
        image_40 <= io_pixelVal_in_4;
      end else if (8'h28 == _T_15[7:0]) begin
        image_40 <= io_pixelVal_in_3;
      end else if (8'h28 == _T_12[7:0]) begin
        image_40 <= io_pixelVal_in_2;
      end else if (8'h28 == _T_9[7:0]) begin
        image_40 <= io_pixelVal_in_1;
      end else if (8'h28 == _T_5[7:0]) begin
        image_40 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_41 <= 4'h8;
    end else if (io_valid_in) begin
      if (8'h29 == _T_27[7:0]) begin
        image_41 <= io_pixelVal_in_7;
      end else if (8'h29 == _T_24[7:0]) begin
        image_41 <= io_pixelVal_in_6;
      end else if (8'h29 == _T_21[7:0]) begin
        image_41 <= io_pixelVal_in_5;
      end else if (8'h29 == _T_18[7:0]) begin
        image_41 <= io_pixelVal_in_4;
      end else if (8'h29 == _T_15[7:0]) begin
        image_41 <= io_pixelVal_in_3;
      end else if (8'h29 == _T_12[7:0]) begin
        image_41 <= io_pixelVal_in_2;
      end else if (8'h29 == _T_9[7:0]) begin
        image_41 <= io_pixelVal_in_1;
      end else if (8'h29 == _T_5[7:0]) begin
        image_41 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_42 <= 4'hc;
    end else if (io_valid_in) begin
      if (8'h2a == _T_27[7:0]) begin
        image_42 <= io_pixelVal_in_7;
      end else if (8'h2a == _T_24[7:0]) begin
        image_42 <= io_pixelVal_in_6;
      end else if (8'h2a == _T_21[7:0]) begin
        image_42 <= io_pixelVal_in_5;
      end else if (8'h2a == _T_18[7:0]) begin
        image_42 <= io_pixelVal_in_4;
      end else if (8'h2a == _T_15[7:0]) begin
        image_42 <= io_pixelVal_in_3;
      end else if (8'h2a == _T_12[7:0]) begin
        image_42 <= io_pixelVal_in_2;
      end else if (8'h2a == _T_9[7:0]) begin
        image_42 <= io_pixelVal_in_1;
      end else if (8'h2a == _T_5[7:0]) begin
        image_42 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_43 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2b == _T_27[7:0]) begin
        image_43 <= io_pixelVal_in_7;
      end else if (8'h2b == _T_24[7:0]) begin
        image_43 <= io_pixelVal_in_6;
      end else if (8'h2b == _T_21[7:0]) begin
        image_43 <= io_pixelVal_in_5;
      end else if (8'h2b == _T_18[7:0]) begin
        image_43 <= io_pixelVal_in_4;
      end else if (8'h2b == _T_15[7:0]) begin
        image_43 <= io_pixelVal_in_3;
      end else if (8'h2b == _T_12[7:0]) begin
        image_43 <= io_pixelVal_in_2;
      end else if (8'h2b == _T_9[7:0]) begin
        image_43 <= io_pixelVal_in_1;
      end else if (8'h2b == _T_5[7:0]) begin
        image_43 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_44 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2c == _T_27[7:0]) begin
        image_44 <= io_pixelVal_in_7;
      end else if (8'h2c == _T_24[7:0]) begin
        image_44 <= io_pixelVal_in_6;
      end else if (8'h2c == _T_21[7:0]) begin
        image_44 <= io_pixelVal_in_5;
      end else if (8'h2c == _T_18[7:0]) begin
        image_44 <= io_pixelVal_in_4;
      end else if (8'h2c == _T_15[7:0]) begin
        image_44 <= io_pixelVal_in_3;
      end else if (8'h2c == _T_12[7:0]) begin
        image_44 <= io_pixelVal_in_2;
      end else if (8'h2c == _T_9[7:0]) begin
        image_44 <= io_pixelVal_in_1;
      end else if (8'h2c == _T_5[7:0]) begin
        image_44 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_45 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h2d == _T_27[7:0]) begin
        image_45 <= io_pixelVal_in_7;
      end else if (8'h2d == _T_24[7:0]) begin
        image_45 <= io_pixelVal_in_6;
      end else if (8'h2d == _T_21[7:0]) begin
        image_45 <= io_pixelVal_in_5;
      end else if (8'h2d == _T_18[7:0]) begin
        image_45 <= io_pixelVal_in_4;
      end else if (8'h2d == _T_15[7:0]) begin
        image_45 <= io_pixelVal_in_3;
      end else if (8'h2d == _T_12[7:0]) begin
        image_45 <= io_pixelVal_in_2;
      end else if (8'h2d == _T_9[7:0]) begin
        image_45 <= io_pixelVal_in_1;
      end else if (8'h2d == _T_5[7:0]) begin
        image_45 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_46 <= 4'h8;
    end else if (io_valid_in) begin
      if (8'h2e == _T_27[7:0]) begin
        image_46 <= io_pixelVal_in_7;
      end else if (8'h2e == _T_24[7:0]) begin
        image_46 <= io_pixelVal_in_6;
      end else if (8'h2e == _T_21[7:0]) begin
        image_46 <= io_pixelVal_in_5;
      end else if (8'h2e == _T_18[7:0]) begin
        image_46 <= io_pixelVal_in_4;
      end else if (8'h2e == _T_15[7:0]) begin
        image_46 <= io_pixelVal_in_3;
      end else if (8'h2e == _T_12[7:0]) begin
        image_46 <= io_pixelVal_in_2;
      end else if (8'h2e == _T_9[7:0]) begin
        image_46 <= io_pixelVal_in_1;
      end else if (8'h2e == _T_5[7:0]) begin
        image_46 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_47 <= 4'hb;
    end else if (io_valid_in) begin
      if (8'h2f == _T_27[7:0]) begin
        image_47 <= io_pixelVal_in_7;
      end else if (8'h2f == _T_24[7:0]) begin
        image_47 <= io_pixelVal_in_6;
      end else if (8'h2f == _T_21[7:0]) begin
        image_47 <= io_pixelVal_in_5;
      end else if (8'h2f == _T_18[7:0]) begin
        image_47 <= io_pixelVal_in_4;
      end else if (8'h2f == _T_15[7:0]) begin
        image_47 <= io_pixelVal_in_3;
      end else if (8'h2f == _T_12[7:0]) begin
        image_47 <= io_pixelVal_in_2;
      end else if (8'h2f == _T_9[7:0]) begin
        image_47 <= io_pixelVal_in_1;
      end else if (8'h2f == _T_5[7:0]) begin
        image_47 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_48 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h30 == _T_27[7:0]) begin
        image_48 <= io_pixelVal_in_7;
      end else if (8'h30 == _T_24[7:0]) begin
        image_48 <= io_pixelVal_in_6;
      end else if (8'h30 == _T_21[7:0]) begin
        image_48 <= io_pixelVal_in_5;
      end else if (8'h30 == _T_18[7:0]) begin
        image_48 <= io_pixelVal_in_4;
      end else if (8'h30 == _T_15[7:0]) begin
        image_48 <= io_pixelVal_in_3;
      end else if (8'h30 == _T_12[7:0]) begin
        image_48 <= io_pixelVal_in_2;
      end else if (8'h30 == _T_9[7:0]) begin
        image_48 <= io_pixelVal_in_1;
      end else if (8'h30 == _T_5[7:0]) begin
        image_48 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_49 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h31 == _T_27[7:0]) begin
        image_49 <= io_pixelVal_in_7;
      end else if (8'h31 == _T_24[7:0]) begin
        image_49 <= io_pixelVal_in_6;
      end else if (8'h31 == _T_21[7:0]) begin
        image_49 <= io_pixelVal_in_5;
      end else if (8'h31 == _T_18[7:0]) begin
        image_49 <= io_pixelVal_in_4;
      end else if (8'h31 == _T_15[7:0]) begin
        image_49 <= io_pixelVal_in_3;
      end else if (8'h31 == _T_12[7:0]) begin
        image_49 <= io_pixelVal_in_2;
      end else if (8'h31 == _T_9[7:0]) begin
        image_49 <= io_pixelVal_in_1;
      end else if (8'h31 == _T_5[7:0]) begin
        image_49 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_50 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h32 == _T_27[7:0]) begin
        image_50 <= io_pixelVal_in_7;
      end else if (8'h32 == _T_24[7:0]) begin
        image_50 <= io_pixelVal_in_6;
      end else if (8'h32 == _T_21[7:0]) begin
        image_50 <= io_pixelVal_in_5;
      end else if (8'h32 == _T_18[7:0]) begin
        image_50 <= io_pixelVal_in_4;
      end else if (8'h32 == _T_15[7:0]) begin
        image_50 <= io_pixelVal_in_3;
      end else if (8'h32 == _T_12[7:0]) begin
        image_50 <= io_pixelVal_in_2;
      end else if (8'h32 == _T_9[7:0]) begin
        image_50 <= io_pixelVal_in_1;
      end else if (8'h32 == _T_5[7:0]) begin
        image_50 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_51 <= 4'h8;
    end else if (io_valid_in) begin
      if (8'h33 == _T_27[7:0]) begin
        image_51 <= io_pixelVal_in_7;
      end else if (8'h33 == _T_24[7:0]) begin
        image_51 <= io_pixelVal_in_6;
      end else if (8'h33 == _T_21[7:0]) begin
        image_51 <= io_pixelVal_in_5;
      end else if (8'h33 == _T_18[7:0]) begin
        image_51 <= io_pixelVal_in_4;
      end else if (8'h33 == _T_15[7:0]) begin
        image_51 <= io_pixelVal_in_3;
      end else if (8'h33 == _T_12[7:0]) begin
        image_51 <= io_pixelVal_in_2;
      end else if (8'h33 == _T_9[7:0]) begin
        image_51 <= io_pixelVal_in_1;
      end else if (8'h33 == _T_5[7:0]) begin
        image_51 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_52 <= 4'hc;
    end else if (io_valid_in) begin
      if (8'h34 == _T_27[7:0]) begin
        image_52 <= io_pixelVal_in_7;
      end else if (8'h34 == _T_24[7:0]) begin
        image_52 <= io_pixelVal_in_6;
      end else if (8'h34 == _T_21[7:0]) begin
        image_52 <= io_pixelVal_in_5;
      end else if (8'h34 == _T_18[7:0]) begin
        image_52 <= io_pixelVal_in_4;
      end else if (8'h34 == _T_15[7:0]) begin
        image_52 <= io_pixelVal_in_3;
      end else if (8'h34 == _T_12[7:0]) begin
        image_52 <= io_pixelVal_in_2;
      end else if (8'h34 == _T_9[7:0]) begin
        image_52 <= io_pixelVal_in_1;
      end else if (8'h34 == _T_5[7:0]) begin
        image_52 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_53 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h35 == _T_27[7:0]) begin
        image_53 <= io_pixelVal_in_7;
      end else if (8'h35 == _T_24[7:0]) begin
        image_53 <= io_pixelVal_in_6;
      end else if (8'h35 == _T_21[7:0]) begin
        image_53 <= io_pixelVal_in_5;
      end else if (8'h35 == _T_18[7:0]) begin
        image_53 <= io_pixelVal_in_4;
      end else if (8'h35 == _T_15[7:0]) begin
        image_53 <= io_pixelVal_in_3;
      end else if (8'h35 == _T_12[7:0]) begin
        image_53 <= io_pixelVal_in_2;
      end else if (8'h35 == _T_9[7:0]) begin
        image_53 <= io_pixelVal_in_1;
      end else if (8'h35 == _T_5[7:0]) begin
        image_53 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_54 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h36 == _T_27[7:0]) begin
        image_54 <= io_pixelVal_in_7;
      end else if (8'h36 == _T_24[7:0]) begin
        image_54 <= io_pixelVal_in_6;
      end else if (8'h36 == _T_21[7:0]) begin
        image_54 <= io_pixelVal_in_5;
      end else if (8'h36 == _T_18[7:0]) begin
        image_54 <= io_pixelVal_in_4;
      end else if (8'h36 == _T_15[7:0]) begin
        image_54 <= io_pixelVal_in_3;
      end else if (8'h36 == _T_12[7:0]) begin
        image_54 <= io_pixelVal_in_2;
      end else if (8'h36 == _T_9[7:0]) begin
        image_54 <= io_pixelVal_in_1;
      end else if (8'h36 == _T_5[7:0]) begin
        image_54 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_55 <= 4'hc;
    end else if (io_valid_in) begin
      if (8'h37 == _T_27[7:0]) begin
        image_55 <= io_pixelVal_in_7;
      end else if (8'h37 == _T_24[7:0]) begin
        image_55 <= io_pixelVal_in_6;
      end else if (8'h37 == _T_21[7:0]) begin
        image_55 <= io_pixelVal_in_5;
      end else if (8'h37 == _T_18[7:0]) begin
        image_55 <= io_pixelVal_in_4;
      end else if (8'h37 == _T_15[7:0]) begin
        image_55 <= io_pixelVal_in_3;
      end else if (8'h37 == _T_12[7:0]) begin
        image_55 <= io_pixelVal_in_2;
      end else if (8'h37 == _T_9[7:0]) begin
        image_55 <= io_pixelVal_in_1;
      end else if (8'h37 == _T_5[7:0]) begin
        image_55 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_56 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h38 == _T_27[7:0]) begin
        image_56 <= io_pixelVal_in_7;
      end else if (8'h38 == _T_24[7:0]) begin
        image_56 <= io_pixelVal_in_6;
      end else if (8'h38 == _T_21[7:0]) begin
        image_56 <= io_pixelVal_in_5;
      end else if (8'h38 == _T_18[7:0]) begin
        image_56 <= io_pixelVal_in_4;
      end else if (8'h38 == _T_15[7:0]) begin
        image_56 <= io_pixelVal_in_3;
      end else if (8'h38 == _T_12[7:0]) begin
        image_56 <= io_pixelVal_in_2;
      end else if (8'h38 == _T_9[7:0]) begin
        image_56 <= io_pixelVal_in_1;
      end else if (8'h38 == _T_5[7:0]) begin
        image_56 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_57 <= 4'h8;
    end else if (io_valid_in) begin
      if (8'h39 == _T_27[7:0]) begin
        image_57 <= io_pixelVal_in_7;
      end else if (8'h39 == _T_24[7:0]) begin
        image_57 <= io_pixelVal_in_6;
      end else if (8'h39 == _T_21[7:0]) begin
        image_57 <= io_pixelVal_in_5;
      end else if (8'h39 == _T_18[7:0]) begin
        image_57 <= io_pixelVal_in_4;
      end else if (8'h39 == _T_15[7:0]) begin
        image_57 <= io_pixelVal_in_3;
      end else if (8'h39 == _T_12[7:0]) begin
        image_57 <= io_pixelVal_in_2;
      end else if (8'h39 == _T_9[7:0]) begin
        image_57 <= io_pixelVal_in_1;
      end else if (8'h39 == _T_5[7:0]) begin
        image_57 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_58 <= 4'hb;
    end else if (io_valid_in) begin
      if (8'h3a == _T_27[7:0]) begin
        image_58 <= io_pixelVal_in_7;
      end else if (8'h3a == _T_24[7:0]) begin
        image_58 <= io_pixelVal_in_6;
      end else if (8'h3a == _T_21[7:0]) begin
        image_58 <= io_pixelVal_in_5;
      end else if (8'h3a == _T_18[7:0]) begin
        image_58 <= io_pixelVal_in_4;
      end else if (8'h3a == _T_15[7:0]) begin
        image_58 <= io_pixelVal_in_3;
      end else if (8'h3a == _T_12[7:0]) begin
        image_58 <= io_pixelVal_in_2;
      end else if (8'h3a == _T_9[7:0]) begin
        image_58 <= io_pixelVal_in_1;
      end else if (8'h3a == _T_5[7:0]) begin
        image_58 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_59 <= 4'hd;
    end else if (io_valid_in) begin
      if (8'h3b == _T_27[7:0]) begin
        image_59 <= io_pixelVal_in_7;
      end else if (8'h3b == _T_24[7:0]) begin
        image_59 <= io_pixelVal_in_6;
      end else if (8'h3b == _T_21[7:0]) begin
        image_59 <= io_pixelVal_in_5;
      end else if (8'h3b == _T_18[7:0]) begin
        image_59 <= io_pixelVal_in_4;
      end else if (8'h3b == _T_15[7:0]) begin
        image_59 <= io_pixelVal_in_3;
      end else if (8'h3b == _T_12[7:0]) begin
        image_59 <= io_pixelVal_in_2;
      end else if (8'h3b == _T_9[7:0]) begin
        image_59 <= io_pixelVal_in_1;
      end else if (8'h3b == _T_5[7:0]) begin
        image_59 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_60 <= 4'he;
    end else if (io_valid_in) begin
      if (8'h3c == _T_27[7:0]) begin
        image_60 <= io_pixelVal_in_7;
      end else if (8'h3c == _T_24[7:0]) begin
        image_60 <= io_pixelVal_in_6;
      end else if (8'h3c == _T_21[7:0]) begin
        image_60 <= io_pixelVal_in_5;
      end else if (8'h3c == _T_18[7:0]) begin
        image_60 <= io_pixelVal_in_4;
      end else if (8'h3c == _T_15[7:0]) begin
        image_60 <= io_pixelVal_in_3;
      end else if (8'h3c == _T_12[7:0]) begin
        image_60 <= io_pixelVal_in_2;
      end else if (8'h3c == _T_9[7:0]) begin
        image_60 <= io_pixelVal_in_1;
      end else if (8'h3c == _T_5[7:0]) begin
        image_60 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_61 <= 4'hb;
    end else if (io_valid_in) begin
      if (8'h3d == _T_27[7:0]) begin
        image_61 <= io_pixelVal_in_7;
      end else if (8'h3d == _T_24[7:0]) begin
        image_61 <= io_pixelVal_in_6;
      end else if (8'h3d == _T_21[7:0]) begin
        image_61 <= io_pixelVal_in_5;
      end else if (8'h3d == _T_18[7:0]) begin
        image_61 <= io_pixelVal_in_4;
      end else if (8'h3d == _T_15[7:0]) begin
        image_61 <= io_pixelVal_in_3;
      end else if (8'h3d == _T_12[7:0]) begin
        image_61 <= io_pixelVal_in_2;
      end else if (8'h3d == _T_9[7:0]) begin
        image_61 <= io_pixelVal_in_1;
      end else if (8'h3d == _T_5[7:0]) begin
        image_61 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_62 <= 4'h9;
    end else if (io_valid_in) begin
      if (8'h3e == _T_27[7:0]) begin
        image_62 <= io_pixelVal_in_7;
      end else if (8'h3e == _T_24[7:0]) begin
        image_62 <= io_pixelVal_in_6;
      end else if (8'h3e == _T_21[7:0]) begin
        image_62 <= io_pixelVal_in_5;
      end else if (8'h3e == _T_18[7:0]) begin
        image_62 <= io_pixelVal_in_4;
      end else if (8'h3e == _T_15[7:0]) begin
        image_62 <= io_pixelVal_in_3;
      end else if (8'h3e == _T_12[7:0]) begin
        image_62 <= io_pixelVal_in_2;
      end else if (8'h3e == _T_9[7:0]) begin
        image_62 <= io_pixelVal_in_1;
      end else if (8'h3e == _T_5[7:0]) begin
        image_62 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_63 <= 4'hc;
    end else if (io_valid_in) begin
      if (8'h3f == _T_27[7:0]) begin
        image_63 <= io_pixelVal_in_7;
      end else if (8'h3f == _T_24[7:0]) begin
        image_63 <= io_pixelVal_in_6;
      end else if (8'h3f == _T_21[7:0]) begin
        image_63 <= io_pixelVal_in_5;
      end else if (8'h3f == _T_18[7:0]) begin
        image_63 <= io_pixelVal_in_4;
      end else if (8'h3f == _T_15[7:0]) begin
        image_63 <= io_pixelVal_in_3;
      end else if (8'h3f == _T_12[7:0]) begin
        image_63 <= io_pixelVal_in_2;
      end else if (8'h3f == _T_9[7:0]) begin
        image_63 <= io_pixelVal_in_1;
      end else if (8'h3f == _T_5[7:0]) begin
        image_63 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_64 <= 4'h4;
    end else if (io_valid_in) begin
      if (8'h40 == _T_27[7:0]) begin
        image_64 <= io_pixelVal_in_7;
      end else if (8'h40 == _T_24[7:0]) begin
        image_64 <= io_pixelVal_in_6;
      end else if (8'h40 == _T_21[7:0]) begin
        image_64 <= io_pixelVal_in_5;
      end else if (8'h40 == _T_18[7:0]) begin
        image_64 <= io_pixelVal_in_4;
      end else if (8'h40 == _T_15[7:0]) begin
        image_64 <= io_pixelVal_in_3;
      end else if (8'h40 == _T_12[7:0]) begin
        image_64 <= io_pixelVal_in_2;
      end else if (8'h40 == _T_9[7:0]) begin
        image_64 <= io_pixelVal_in_1;
      end else if (8'h40 == _T_5[7:0]) begin
        image_64 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_65 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h41 == _T_27[7:0]) begin
        image_65 <= io_pixelVal_in_7;
      end else if (8'h41 == _T_24[7:0]) begin
        image_65 <= io_pixelVal_in_6;
      end else if (8'h41 == _T_21[7:0]) begin
        image_65 <= io_pixelVal_in_5;
      end else if (8'h41 == _T_18[7:0]) begin
        image_65 <= io_pixelVal_in_4;
      end else if (8'h41 == _T_15[7:0]) begin
        image_65 <= io_pixelVal_in_3;
      end else if (8'h41 == _T_12[7:0]) begin
        image_65 <= io_pixelVal_in_2;
      end else if (8'h41 == _T_9[7:0]) begin
        image_65 <= io_pixelVal_in_1;
      end else if (8'h41 == _T_5[7:0]) begin
        image_65 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_66 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h42 == _T_27[7:0]) begin
        image_66 <= io_pixelVal_in_7;
      end else if (8'h42 == _T_24[7:0]) begin
        image_66 <= io_pixelVal_in_6;
      end else if (8'h42 == _T_21[7:0]) begin
        image_66 <= io_pixelVal_in_5;
      end else if (8'h42 == _T_18[7:0]) begin
        image_66 <= io_pixelVal_in_4;
      end else if (8'h42 == _T_15[7:0]) begin
        image_66 <= io_pixelVal_in_3;
      end else if (8'h42 == _T_12[7:0]) begin
        image_66 <= io_pixelVal_in_2;
      end else if (8'h42 == _T_9[7:0]) begin
        image_66 <= io_pixelVal_in_1;
      end else if (8'h42 == _T_5[7:0]) begin
        image_66 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_67 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h43 == _T_27[7:0]) begin
        image_67 <= io_pixelVal_in_7;
      end else if (8'h43 == _T_24[7:0]) begin
        image_67 <= io_pixelVal_in_6;
      end else if (8'h43 == _T_21[7:0]) begin
        image_67 <= io_pixelVal_in_5;
      end else if (8'h43 == _T_18[7:0]) begin
        image_67 <= io_pixelVal_in_4;
      end else if (8'h43 == _T_15[7:0]) begin
        image_67 <= io_pixelVal_in_3;
      end else if (8'h43 == _T_12[7:0]) begin
        image_67 <= io_pixelVal_in_2;
      end else if (8'h43 == _T_9[7:0]) begin
        image_67 <= io_pixelVal_in_1;
      end else if (8'h43 == _T_5[7:0]) begin
        image_67 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_68 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h44 == _T_27[7:0]) begin
        image_68 <= io_pixelVal_in_7;
      end else if (8'h44 == _T_24[7:0]) begin
        image_68 <= io_pixelVal_in_6;
      end else if (8'h44 == _T_21[7:0]) begin
        image_68 <= io_pixelVal_in_5;
      end else if (8'h44 == _T_18[7:0]) begin
        image_68 <= io_pixelVal_in_4;
      end else if (8'h44 == _T_15[7:0]) begin
        image_68 <= io_pixelVal_in_3;
      end else if (8'h44 == _T_12[7:0]) begin
        image_68 <= io_pixelVal_in_2;
      end else if (8'h44 == _T_9[7:0]) begin
        image_68 <= io_pixelVal_in_1;
      end else if (8'h44 == _T_5[7:0]) begin
        image_68 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_69 <= 4'h8;
    end else if (io_valid_in) begin
      if (8'h45 == _T_27[7:0]) begin
        image_69 <= io_pixelVal_in_7;
      end else if (8'h45 == _T_24[7:0]) begin
        image_69 <= io_pixelVal_in_6;
      end else if (8'h45 == _T_21[7:0]) begin
        image_69 <= io_pixelVal_in_5;
      end else if (8'h45 == _T_18[7:0]) begin
        image_69 <= io_pixelVal_in_4;
      end else if (8'h45 == _T_15[7:0]) begin
        image_69 <= io_pixelVal_in_3;
      end else if (8'h45 == _T_12[7:0]) begin
        image_69 <= io_pixelVal_in_2;
      end else if (8'h45 == _T_9[7:0]) begin
        image_69 <= io_pixelVal_in_1;
      end else if (8'h45 == _T_5[7:0]) begin
        image_69 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_70 <= 4'hb;
    end else if (io_valid_in) begin
      if (8'h46 == _T_27[7:0]) begin
        image_70 <= io_pixelVal_in_7;
      end else if (8'h46 == _T_24[7:0]) begin
        image_70 <= io_pixelVal_in_6;
      end else if (8'h46 == _T_21[7:0]) begin
        image_70 <= io_pixelVal_in_5;
      end else if (8'h46 == _T_18[7:0]) begin
        image_70 <= io_pixelVal_in_4;
      end else if (8'h46 == _T_15[7:0]) begin
        image_70 <= io_pixelVal_in_3;
      end else if (8'h46 == _T_12[7:0]) begin
        image_70 <= io_pixelVal_in_2;
      end else if (8'h46 == _T_9[7:0]) begin
        image_70 <= io_pixelVal_in_1;
      end else if (8'h46 == _T_5[7:0]) begin
        image_70 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_71 <= 4'hd;
    end else if (io_valid_in) begin
      if (8'h47 == _T_27[7:0]) begin
        image_71 <= io_pixelVal_in_7;
      end else if (8'h47 == _T_24[7:0]) begin
        image_71 <= io_pixelVal_in_6;
      end else if (8'h47 == _T_21[7:0]) begin
        image_71 <= io_pixelVal_in_5;
      end else if (8'h47 == _T_18[7:0]) begin
        image_71 <= io_pixelVal_in_4;
      end else if (8'h47 == _T_15[7:0]) begin
        image_71 <= io_pixelVal_in_3;
      end else if (8'h47 == _T_12[7:0]) begin
        image_71 <= io_pixelVal_in_2;
      end else if (8'h47 == _T_9[7:0]) begin
        image_71 <= io_pixelVal_in_1;
      end else if (8'h47 == _T_5[7:0]) begin
        image_71 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_72 <= 4'hb;
    end else if (io_valid_in) begin
      if (8'h48 == _T_27[7:0]) begin
        image_72 <= io_pixelVal_in_7;
      end else if (8'h48 == _T_24[7:0]) begin
        image_72 <= io_pixelVal_in_6;
      end else if (8'h48 == _T_21[7:0]) begin
        image_72 <= io_pixelVal_in_5;
      end else if (8'h48 == _T_18[7:0]) begin
        image_72 <= io_pixelVal_in_4;
      end else if (8'h48 == _T_15[7:0]) begin
        image_72 <= io_pixelVal_in_3;
      end else if (8'h48 == _T_12[7:0]) begin
        image_72 <= io_pixelVal_in_2;
      end else if (8'h48 == _T_9[7:0]) begin
        image_72 <= io_pixelVal_in_1;
      end else if (8'h48 == _T_5[7:0]) begin
        image_72 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_73 <= 4'ha;
    end else if (io_valid_in) begin
      if (8'h49 == _T_27[7:0]) begin
        image_73 <= io_pixelVal_in_7;
      end else if (8'h49 == _T_24[7:0]) begin
        image_73 <= io_pixelVal_in_6;
      end else if (8'h49 == _T_21[7:0]) begin
        image_73 <= io_pixelVal_in_5;
      end else if (8'h49 == _T_18[7:0]) begin
        image_73 <= io_pixelVal_in_4;
      end else if (8'h49 == _T_15[7:0]) begin
        image_73 <= io_pixelVal_in_3;
      end else if (8'h49 == _T_12[7:0]) begin
        image_73 <= io_pixelVal_in_2;
      end else if (8'h49 == _T_9[7:0]) begin
        image_73 <= io_pixelVal_in_1;
      end else if (8'h49 == _T_5[7:0]) begin
        image_73 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_74 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h4a == _T_27[7:0]) begin
        image_74 <= io_pixelVal_in_7;
      end else if (8'h4a == _T_24[7:0]) begin
        image_74 <= io_pixelVal_in_6;
      end else if (8'h4a == _T_21[7:0]) begin
        image_74 <= io_pixelVal_in_5;
      end else if (8'h4a == _T_18[7:0]) begin
        image_74 <= io_pixelVal_in_4;
      end else if (8'h4a == _T_15[7:0]) begin
        image_74 <= io_pixelVal_in_3;
      end else if (8'h4a == _T_12[7:0]) begin
        image_74 <= io_pixelVal_in_2;
      end else if (8'h4a == _T_9[7:0]) begin
        image_74 <= io_pixelVal_in_1;
      end else if (8'h4a == _T_5[7:0]) begin
        image_74 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_75 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h4b == _T_27[7:0]) begin
        image_75 <= io_pixelVal_in_7;
      end else if (8'h4b == _T_24[7:0]) begin
        image_75 <= io_pixelVal_in_6;
      end else if (8'h4b == _T_21[7:0]) begin
        image_75 <= io_pixelVal_in_5;
      end else if (8'h4b == _T_18[7:0]) begin
        image_75 <= io_pixelVal_in_4;
      end else if (8'h4b == _T_15[7:0]) begin
        image_75 <= io_pixelVal_in_3;
      end else if (8'h4b == _T_12[7:0]) begin
        image_75 <= io_pixelVal_in_2;
      end else if (8'h4b == _T_9[7:0]) begin
        image_75 <= io_pixelVal_in_1;
      end else if (8'h4b == _T_5[7:0]) begin
        image_75 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_76 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h4c == _T_27[7:0]) begin
        image_76 <= io_pixelVal_in_7;
      end else if (8'h4c == _T_24[7:0]) begin
        image_76 <= io_pixelVal_in_6;
      end else if (8'h4c == _T_21[7:0]) begin
        image_76 <= io_pixelVal_in_5;
      end else if (8'h4c == _T_18[7:0]) begin
        image_76 <= io_pixelVal_in_4;
      end else if (8'h4c == _T_15[7:0]) begin
        image_76 <= io_pixelVal_in_3;
      end else if (8'h4c == _T_12[7:0]) begin
        image_76 <= io_pixelVal_in_2;
      end else if (8'h4c == _T_9[7:0]) begin
        image_76 <= io_pixelVal_in_1;
      end else if (8'h4c == _T_5[7:0]) begin
        image_76 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_77 <= 4'h7;
    end else if (io_valid_in) begin
      if (8'h4d == _T_27[7:0]) begin
        image_77 <= io_pixelVal_in_7;
      end else if (8'h4d == _T_24[7:0]) begin
        image_77 <= io_pixelVal_in_6;
      end else if (8'h4d == _T_21[7:0]) begin
        image_77 <= io_pixelVal_in_5;
      end else if (8'h4d == _T_18[7:0]) begin
        image_77 <= io_pixelVal_in_4;
      end else if (8'h4d == _T_15[7:0]) begin
        image_77 <= io_pixelVal_in_3;
      end else if (8'h4d == _T_12[7:0]) begin
        image_77 <= io_pixelVal_in_2;
      end else if (8'h4d == _T_9[7:0]) begin
        image_77 <= io_pixelVal_in_1;
      end else if (8'h4d == _T_5[7:0]) begin
        image_77 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_78 <= 4'h4;
    end else if (io_valid_in) begin
      if (8'h4e == _T_27[7:0]) begin
        image_78 <= io_pixelVal_in_7;
      end else if (8'h4e == _T_24[7:0]) begin
        image_78 <= io_pixelVal_in_6;
      end else if (8'h4e == _T_21[7:0]) begin
        image_78 <= io_pixelVal_in_5;
      end else if (8'h4e == _T_18[7:0]) begin
        image_78 <= io_pixelVal_in_4;
      end else if (8'h4e == _T_15[7:0]) begin
        image_78 <= io_pixelVal_in_3;
      end else if (8'h4e == _T_12[7:0]) begin
        image_78 <= io_pixelVal_in_2;
      end else if (8'h4e == _T_9[7:0]) begin
        image_78 <= io_pixelVal_in_1;
      end else if (8'h4e == _T_5[7:0]) begin
        image_78 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_79 <= 4'h4;
    end else if (io_valid_in) begin
      if (8'h4f == _T_27[7:0]) begin
        image_79 <= io_pixelVal_in_7;
      end else if (8'h4f == _T_24[7:0]) begin
        image_79 <= io_pixelVal_in_6;
      end else if (8'h4f == _T_21[7:0]) begin
        image_79 <= io_pixelVal_in_5;
      end else if (8'h4f == _T_18[7:0]) begin
        image_79 <= io_pixelVal_in_4;
      end else if (8'h4f == _T_15[7:0]) begin
        image_79 <= io_pixelVal_in_3;
      end else if (8'h4f == _T_12[7:0]) begin
        image_79 <= io_pixelVal_in_2;
      end else if (8'h4f == _T_9[7:0]) begin
        image_79 <= io_pixelVal_in_1;
      end else if (8'h4f == _T_5[7:0]) begin
        image_79 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_80 <= 4'h4;
    end else if (io_valid_in) begin
      if (8'h50 == _T_27[7:0]) begin
        image_80 <= io_pixelVal_in_7;
      end else if (8'h50 == _T_24[7:0]) begin
        image_80 <= io_pixelVal_in_6;
      end else if (8'h50 == _T_21[7:0]) begin
        image_80 <= io_pixelVal_in_5;
      end else if (8'h50 == _T_18[7:0]) begin
        image_80 <= io_pixelVal_in_4;
      end else if (8'h50 == _T_15[7:0]) begin
        image_80 <= io_pixelVal_in_3;
      end else if (8'h50 == _T_12[7:0]) begin
        image_80 <= io_pixelVal_in_2;
      end else if (8'h50 == _T_9[7:0]) begin
        image_80 <= io_pixelVal_in_1;
      end else if (8'h50 == _T_5[7:0]) begin
        image_80 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_81 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h51 == _T_27[7:0]) begin
        image_81 <= io_pixelVal_in_7;
      end else if (8'h51 == _T_24[7:0]) begin
        image_81 <= io_pixelVal_in_6;
      end else if (8'h51 == _T_21[7:0]) begin
        image_81 <= io_pixelVal_in_5;
      end else if (8'h51 == _T_18[7:0]) begin
        image_81 <= io_pixelVal_in_4;
      end else if (8'h51 == _T_15[7:0]) begin
        image_81 <= io_pixelVal_in_3;
      end else if (8'h51 == _T_12[7:0]) begin
        image_81 <= io_pixelVal_in_2;
      end else if (8'h51 == _T_9[7:0]) begin
        image_81 <= io_pixelVal_in_1;
      end else if (8'h51 == _T_5[7:0]) begin
        image_81 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_82 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h52 == _T_27[7:0]) begin
        image_82 <= io_pixelVal_in_7;
      end else if (8'h52 == _T_24[7:0]) begin
        image_82 <= io_pixelVal_in_6;
      end else if (8'h52 == _T_21[7:0]) begin
        image_82 <= io_pixelVal_in_5;
      end else if (8'h52 == _T_18[7:0]) begin
        image_82 <= io_pixelVal_in_4;
      end else if (8'h52 == _T_15[7:0]) begin
        image_82 <= io_pixelVal_in_3;
      end else if (8'h52 == _T_12[7:0]) begin
        image_82 <= io_pixelVal_in_2;
      end else if (8'h52 == _T_9[7:0]) begin
        image_82 <= io_pixelVal_in_1;
      end else if (8'h52 == _T_5[7:0]) begin
        image_82 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_83 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h53 == _T_27[7:0]) begin
        image_83 <= io_pixelVal_in_7;
      end else if (8'h53 == _T_24[7:0]) begin
        image_83 <= io_pixelVal_in_6;
      end else if (8'h53 == _T_21[7:0]) begin
        image_83 <= io_pixelVal_in_5;
      end else if (8'h53 == _T_18[7:0]) begin
        image_83 <= io_pixelVal_in_4;
      end else if (8'h53 == _T_15[7:0]) begin
        image_83 <= io_pixelVal_in_3;
      end else if (8'h53 == _T_12[7:0]) begin
        image_83 <= io_pixelVal_in_2;
      end else if (8'h53 == _T_9[7:0]) begin
        image_83 <= io_pixelVal_in_1;
      end else if (8'h53 == _T_5[7:0]) begin
        image_83 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_84 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h54 == _T_27[7:0]) begin
        image_84 <= io_pixelVal_in_7;
      end else if (8'h54 == _T_24[7:0]) begin
        image_84 <= io_pixelVal_in_6;
      end else if (8'h54 == _T_21[7:0]) begin
        image_84 <= io_pixelVal_in_5;
      end else if (8'h54 == _T_18[7:0]) begin
        image_84 <= io_pixelVal_in_4;
      end else if (8'h54 == _T_15[7:0]) begin
        image_84 <= io_pixelVal_in_3;
      end else if (8'h54 == _T_12[7:0]) begin
        image_84 <= io_pixelVal_in_2;
      end else if (8'h54 == _T_9[7:0]) begin
        image_84 <= io_pixelVal_in_1;
      end else if (8'h54 == _T_5[7:0]) begin
        image_84 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_85 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h55 == _T_27[7:0]) begin
        image_85 <= io_pixelVal_in_7;
      end else if (8'h55 == _T_24[7:0]) begin
        image_85 <= io_pixelVal_in_6;
      end else if (8'h55 == _T_21[7:0]) begin
        image_85 <= io_pixelVal_in_5;
      end else if (8'h55 == _T_18[7:0]) begin
        image_85 <= io_pixelVal_in_4;
      end else if (8'h55 == _T_15[7:0]) begin
        image_85 <= io_pixelVal_in_3;
      end else if (8'h55 == _T_12[7:0]) begin
        image_85 <= io_pixelVal_in_2;
      end else if (8'h55 == _T_9[7:0]) begin
        image_85 <= io_pixelVal_in_1;
      end else if (8'h55 == _T_5[7:0]) begin
        image_85 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_86 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h56 == _T_27[7:0]) begin
        image_86 <= io_pixelVal_in_7;
      end else if (8'h56 == _T_24[7:0]) begin
        image_86 <= io_pixelVal_in_6;
      end else if (8'h56 == _T_21[7:0]) begin
        image_86 <= io_pixelVal_in_5;
      end else if (8'h56 == _T_18[7:0]) begin
        image_86 <= io_pixelVal_in_4;
      end else if (8'h56 == _T_15[7:0]) begin
        image_86 <= io_pixelVal_in_3;
      end else if (8'h56 == _T_12[7:0]) begin
        image_86 <= io_pixelVal_in_2;
      end else if (8'h56 == _T_9[7:0]) begin
        image_86 <= io_pixelVal_in_1;
      end else if (8'h56 == _T_5[7:0]) begin
        image_86 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_87 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h57 == _T_27[7:0]) begin
        image_87 <= io_pixelVal_in_7;
      end else if (8'h57 == _T_24[7:0]) begin
        image_87 <= io_pixelVal_in_6;
      end else if (8'h57 == _T_21[7:0]) begin
        image_87 <= io_pixelVal_in_5;
      end else if (8'h57 == _T_18[7:0]) begin
        image_87 <= io_pixelVal_in_4;
      end else if (8'h57 == _T_15[7:0]) begin
        image_87 <= io_pixelVal_in_3;
      end else if (8'h57 == _T_12[7:0]) begin
        image_87 <= io_pixelVal_in_2;
      end else if (8'h57 == _T_9[7:0]) begin
        image_87 <= io_pixelVal_in_1;
      end else if (8'h57 == _T_5[7:0]) begin
        image_87 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_88 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h58 == _T_27[7:0]) begin
        image_88 <= io_pixelVal_in_7;
      end else if (8'h58 == _T_24[7:0]) begin
        image_88 <= io_pixelVal_in_6;
      end else if (8'h58 == _T_21[7:0]) begin
        image_88 <= io_pixelVal_in_5;
      end else if (8'h58 == _T_18[7:0]) begin
        image_88 <= io_pixelVal_in_4;
      end else if (8'h58 == _T_15[7:0]) begin
        image_88 <= io_pixelVal_in_3;
      end else if (8'h58 == _T_12[7:0]) begin
        image_88 <= io_pixelVal_in_2;
      end else if (8'h58 == _T_9[7:0]) begin
        image_88 <= io_pixelVal_in_1;
      end else if (8'h58 == _T_5[7:0]) begin
        image_88 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_89 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h59 == _T_27[7:0]) begin
        image_89 <= io_pixelVal_in_7;
      end else if (8'h59 == _T_24[7:0]) begin
        image_89 <= io_pixelVal_in_6;
      end else if (8'h59 == _T_21[7:0]) begin
        image_89 <= io_pixelVal_in_5;
      end else if (8'h59 == _T_18[7:0]) begin
        image_89 <= io_pixelVal_in_4;
      end else if (8'h59 == _T_15[7:0]) begin
        image_89 <= io_pixelVal_in_3;
      end else if (8'h59 == _T_12[7:0]) begin
        image_89 <= io_pixelVal_in_2;
      end else if (8'h59 == _T_9[7:0]) begin
        image_89 <= io_pixelVal_in_1;
      end else if (8'h59 == _T_5[7:0]) begin
        image_89 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_90 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h5a == _T_27[7:0]) begin
        image_90 <= io_pixelVal_in_7;
      end else if (8'h5a == _T_24[7:0]) begin
        image_90 <= io_pixelVal_in_6;
      end else if (8'h5a == _T_21[7:0]) begin
        image_90 <= io_pixelVal_in_5;
      end else if (8'h5a == _T_18[7:0]) begin
        image_90 <= io_pixelVal_in_4;
      end else if (8'h5a == _T_15[7:0]) begin
        image_90 <= io_pixelVal_in_3;
      end else if (8'h5a == _T_12[7:0]) begin
        image_90 <= io_pixelVal_in_2;
      end else if (8'h5a == _T_9[7:0]) begin
        image_90 <= io_pixelVal_in_1;
      end else if (8'h5a == _T_5[7:0]) begin
        image_90 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_91 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h5b == _T_27[7:0]) begin
        image_91 <= io_pixelVal_in_7;
      end else if (8'h5b == _T_24[7:0]) begin
        image_91 <= io_pixelVal_in_6;
      end else if (8'h5b == _T_21[7:0]) begin
        image_91 <= io_pixelVal_in_5;
      end else if (8'h5b == _T_18[7:0]) begin
        image_91 <= io_pixelVal_in_4;
      end else if (8'h5b == _T_15[7:0]) begin
        image_91 <= io_pixelVal_in_3;
      end else if (8'h5b == _T_12[7:0]) begin
        image_91 <= io_pixelVal_in_2;
      end else if (8'h5b == _T_9[7:0]) begin
        image_91 <= io_pixelVal_in_1;
      end else if (8'h5b == _T_5[7:0]) begin
        image_91 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_92 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h5c == _T_27[7:0]) begin
        image_92 <= io_pixelVal_in_7;
      end else if (8'h5c == _T_24[7:0]) begin
        image_92 <= io_pixelVal_in_6;
      end else if (8'h5c == _T_21[7:0]) begin
        image_92 <= io_pixelVal_in_5;
      end else if (8'h5c == _T_18[7:0]) begin
        image_92 <= io_pixelVal_in_4;
      end else if (8'h5c == _T_15[7:0]) begin
        image_92 <= io_pixelVal_in_3;
      end else if (8'h5c == _T_12[7:0]) begin
        image_92 <= io_pixelVal_in_2;
      end else if (8'h5c == _T_9[7:0]) begin
        image_92 <= io_pixelVal_in_1;
      end else if (8'h5c == _T_5[7:0]) begin
        image_92 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_93 <= 4'h7;
    end else if (io_valid_in) begin
      if (8'h5d == _T_27[7:0]) begin
        image_93 <= io_pixelVal_in_7;
      end else if (8'h5d == _T_24[7:0]) begin
        image_93 <= io_pixelVal_in_6;
      end else if (8'h5d == _T_21[7:0]) begin
        image_93 <= io_pixelVal_in_5;
      end else if (8'h5d == _T_18[7:0]) begin
        image_93 <= io_pixelVal_in_4;
      end else if (8'h5d == _T_15[7:0]) begin
        image_93 <= io_pixelVal_in_3;
      end else if (8'h5d == _T_12[7:0]) begin
        image_93 <= io_pixelVal_in_2;
      end else if (8'h5d == _T_9[7:0]) begin
        image_93 <= io_pixelVal_in_1;
      end else if (8'h5d == _T_5[7:0]) begin
        image_93 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_94 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h5e == _T_27[7:0]) begin
        image_94 <= io_pixelVal_in_7;
      end else if (8'h5e == _T_24[7:0]) begin
        image_94 <= io_pixelVal_in_6;
      end else if (8'h5e == _T_21[7:0]) begin
        image_94 <= io_pixelVal_in_5;
      end else if (8'h5e == _T_18[7:0]) begin
        image_94 <= io_pixelVal_in_4;
      end else if (8'h5e == _T_15[7:0]) begin
        image_94 <= io_pixelVal_in_3;
      end else if (8'h5e == _T_12[7:0]) begin
        image_94 <= io_pixelVal_in_2;
      end else if (8'h5e == _T_9[7:0]) begin
        image_94 <= io_pixelVal_in_1;
      end else if (8'h5e == _T_5[7:0]) begin
        image_94 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_95 <= 4'h4;
    end else if (io_valid_in) begin
      if (8'h5f == _T_27[7:0]) begin
        image_95 <= io_pixelVal_in_7;
      end else if (8'h5f == _T_24[7:0]) begin
        image_95 <= io_pixelVal_in_6;
      end else if (8'h5f == _T_21[7:0]) begin
        image_95 <= io_pixelVal_in_5;
      end else if (8'h5f == _T_18[7:0]) begin
        image_95 <= io_pixelVal_in_4;
      end else if (8'h5f == _T_15[7:0]) begin
        image_95 <= io_pixelVal_in_3;
      end else if (8'h5f == _T_12[7:0]) begin
        image_95 <= io_pixelVal_in_2;
      end else if (8'h5f == _T_9[7:0]) begin
        image_95 <= io_pixelVal_in_1;
      end else if (8'h5f == _T_5[7:0]) begin
        image_95 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_96 <= 4'h4;
    end else if (io_valid_in) begin
      if (8'h60 == _T_27[7:0]) begin
        image_96 <= io_pixelVal_in_7;
      end else if (8'h60 == _T_24[7:0]) begin
        image_96 <= io_pixelVal_in_6;
      end else if (8'h60 == _T_21[7:0]) begin
        image_96 <= io_pixelVal_in_5;
      end else if (8'h60 == _T_18[7:0]) begin
        image_96 <= io_pixelVal_in_4;
      end else if (8'h60 == _T_15[7:0]) begin
        image_96 <= io_pixelVal_in_3;
      end else if (8'h60 == _T_12[7:0]) begin
        image_96 <= io_pixelVal_in_2;
      end else if (8'h60 == _T_9[7:0]) begin
        image_96 <= io_pixelVal_in_1;
      end else if (8'h60 == _T_5[7:0]) begin
        image_96 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_97 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h61 == _T_27[7:0]) begin
        image_97 <= io_pixelVal_in_7;
      end else if (8'h61 == _T_24[7:0]) begin
        image_97 <= io_pixelVal_in_6;
      end else if (8'h61 == _T_21[7:0]) begin
        image_97 <= io_pixelVal_in_5;
      end else if (8'h61 == _T_18[7:0]) begin
        image_97 <= io_pixelVal_in_4;
      end else if (8'h61 == _T_15[7:0]) begin
        image_97 <= io_pixelVal_in_3;
      end else if (8'h61 == _T_12[7:0]) begin
        image_97 <= io_pixelVal_in_2;
      end else if (8'h61 == _T_9[7:0]) begin
        image_97 <= io_pixelVal_in_1;
      end else if (8'h61 == _T_5[7:0]) begin
        image_97 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_98 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h62 == _T_27[7:0]) begin
        image_98 <= io_pixelVal_in_7;
      end else if (8'h62 == _T_24[7:0]) begin
        image_98 <= io_pixelVal_in_6;
      end else if (8'h62 == _T_21[7:0]) begin
        image_98 <= io_pixelVal_in_5;
      end else if (8'h62 == _T_18[7:0]) begin
        image_98 <= io_pixelVal_in_4;
      end else if (8'h62 == _T_15[7:0]) begin
        image_98 <= io_pixelVal_in_3;
      end else if (8'h62 == _T_12[7:0]) begin
        image_98 <= io_pixelVal_in_2;
      end else if (8'h62 == _T_9[7:0]) begin
        image_98 <= io_pixelVal_in_1;
      end else if (8'h62 == _T_5[7:0]) begin
        image_98 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_99 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h63 == _T_27[7:0]) begin
        image_99 <= io_pixelVal_in_7;
      end else if (8'h63 == _T_24[7:0]) begin
        image_99 <= io_pixelVal_in_6;
      end else if (8'h63 == _T_21[7:0]) begin
        image_99 <= io_pixelVal_in_5;
      end else if (8'h63 == _T_18[7:0]) begin
        image_99 <= io_pixelVal_in_4;
      end else if (8'h63 == _T_15[7:0]) begin
        image_99 <= io_pixelVal_in_3;
      end else if (8'h63 == _T_12[7:0]) begin
        image_99 <= io_pixelVal_in_2;
      end else if (8'h63 == _T_9[7:0]) begin
        image_99 <= io_pixelVal_in_1;
      end else if (8'h63 == _T_5[7:0]) begin
        image_99 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_100 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h64 == _T_27[7:0]) begin
        image_100 <= io_pixelVal_in_7;
      end else if (8'h64 == _T_24[7:0]) begin
        image_100 <= io_pixelVal_in_6;
      end else if (8'h64 == _T_21[7:0]) begin
        image_100 <= io_pixelVal_in_5;
      end else if (8'h64 == _T_18[7:0]) begin
        image_100 <= io_pixelVal_in_4;
      end else if (8'h64 == _T_15[7:0]) begin
        image_100 <= io_pixelVal_in_3;
      end else if (8'h64 == _T_12[7:0]) begin
        image_100 <= io_pixelVal_in_2;
      end else if (8'h64 == _T_9[7:0]) begin
        image_100 <= io_pixelVal_in_1;
      end else if (8'h64 == _T_5[7:0]) begin
        image_100 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_101 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h65 == _T_27[7:0]) begin
        image_101 <= io_pixelVal_in_7;
      end else if (8'h65 == _T_24[7:0]) begin
        image_101 <= io_pixelVal_in_6;
      end else if (8'h65 == _T_21[7:0]) begin
        image_101 <= io_pixelVal_in_5;
      end else if (8'h65 == _T_18[7:0]) begin
        image_101 <= io_pixelVal_in_4;
      end else if (8'h65 == _T_15[7:0]) begin
        image_101 <= io_pixelVal_in_3;
      end else if (8'h65 == _T_12[7:0]) begin
        image_101 <= io_pixelVal_in_2;
      end else if (8'h65 == _T_9[7:0]) begin
        image_101 <= io_pixelVal_in_1;
      end else if (8'h65 == _T_5[7:0]) begin
        image_101 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_102 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h66 == _T_27[7:0]) begin
        image_102 <= io_pixelVal_in_7;
      end else if (8'h66 == _T_24[7:0]) begin
        image_102 <= io_pixelVal_in_6;
      end else if (8'h66 == _T_21[7:0]) begin
        image_102 <= io_pixelVal_in_5;
      end else if (8'h66 == _T_18[7:0]) begin
        image_102 <= io_pixelVal_in_4;
      end else if (8'h66 == _T_15[7:0]) begin
        image_102 <= io_pixelVal_in_3;
      end else if (8'h66 == _T_12[7:0]) begin
        image_102 <= io_pixelVal_in_2;
      end else if (8'h66 == _T_9[7:0]) begin
        image_102 <= io_pixelVal_in_1;
      end else if (8'h66 == _T_5[7:0]) begin
        image_102 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_103 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h67 == _T_27[7:0]) begin
        image_103 <= io_pixelVal_in_7;
      end else if (8'h67 == _T_24[7:0]) begin
        image_103 <= io_pixelVal_in_6;
      end else if (8'h67 == _T_21[7:0]) begin
        image_103 <= io_pixelVal_in_5;
      end else if (8'h67 == _T_18[7:0]) begin
        image_103 <= io_pixelVal_in_4;
      end else if (8'h67 == _T_15[7:0]) begin
        image_103 <= io_pixelVal_in_3;
      end else if (8'h67 == _T_12[7:0]) begin
        image_103 <= io_pixelVal_in_2;
      end else if (8'h67 == _T_9[7:0]) begin
        image_103 <= io_pixelVal_in_1;
      end else if (8'h67 == _T_5[7:0]) begin
        image_103 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_104 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h68 == _T_27[7:0]) begin
        image_104 <= io_pixelVal_in_7;
      end else if (8'h68 == _T_24[7:0]) begin
        image_104 <= io_pixelVal_in_6;
      end else if (8'h68 == _T_21[7:0]) begin
        image_104 <= io_pixelVal_in_5;
      end else if (8'h68 == _T_18[7:0]) begin
        image_104 <= io_pixelVal_in_4;
      end else if (8'h68 == _T_15[7:0]) begin
        image_104 <= io_pixelVal_in_3;
      end else if (8'h68 == _T_12[7:0]) begin
        image_104 <= io_pixelVal_in_2;
      end else if (8'h68 == _T_9[7:0]) begin
        image_104 <= io_pixelVal_in_1;
      end else if (8'h68 == _T_5[7:0]) begin
        image_104 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_105 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h69 == _T_27[7:0]) begin
        image_105 <= io_pixelVal_in_7;
      end else if (8'h69 == _T_24[7:0]) begin
        image_105 <= io_pixelVal_in_6;
      end else if (8'h69 == _T_21[7:0]) begin
        image_105 <= io_pixelVal_in_5;
      end else if (8'h69 == _T_18[7:0]) begin
        image_105 <= io_pixelVal_in_4;
      end else if (8'h69 == _T_15[7:0]) begin
        image_105 <= io_pixelVal_in_3;
      end else if (8'h69 == _T_12[7:0]) begin
        image_105 <= io_pixelVal_in_2;
      end else if (8'h69 == _T_9[7:0]) begin
        image_105 <= io_pixelVal_in_1;
      end else if (8'h69 == _T_5[7:0]) begin
        image_105 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_106 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h6a == _T_27[7:0]) begin
        image_106 <= io_pixelVal_in_7;
      end else if (8'h6a == _T_24[7:0]) begin
        image_106 <= io_pixelVal_in_6;
      end else if (8'h6a == _T_21[7:0]) begin
        image_106 <= io_pixelVal_in_5;
      end else if (8'h6a == _T_18[7:0]) begin
        image_106 <= io_pixelVal_in_4;
      end else if (8'h6a == _T_15[7:0]) begin
        image_106 <= io_pixelVal_in_3;
      end else if (8'h6a == _T_12[7:0]) begin
        image_106 <= io_pixelVal_in_2;
      end else if (8'h6a == _T_9[7:0]) begin
        image_106 <= io_pixelVal_in_1;
      end else if (8'h6a == _T_5[7:0]) begin
        image_106 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_107 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h6b == _T_27[7:0]) begin
        image_107 <= io_pixelVal_in_7;
      end else if (8'h6b == _T_24[7:0]) begin
        image_107 <= io_pixelVal_in_6;
      end else if (8'h6b == _T_21[7:0]) begin
        image_107 <= io_pixelVal_in_5;
      end else if (8'h6b == _T_18[7:0]) begin
        image_107 <= io_pixelVal_in_4;
      end else if (8'h6b == _T_15[7:0]) begin
        image_107 <= io_pixelVal_in_3;
      end else if (8'h6b == _T_12[7:0]) begin
        image_107 <= io_pixelVal_in_2;
      end else if (8'h6b == _T_9[7:0]) begin
        image_107 <= io_pixelVal_in_1;
      end else if (8'h6b == _T_5[7:0]) begin
        image_107 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_108 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h6c == _T_27[7:0]) begin
        image_108 <= io_pixelVal_in_7;
      end else if (8'h6c == _T_24[7:0]) begin
        image_108 <= io_pixelVal_in_6;
      end else if (8'h6c == _T_21[7:0]) begin
        image_108 <= io_pixelVal_in_5;
      end else if (8'h6c == _T_18[7:0]) begin
        image_108 <= io_pixelVal_in_4;
      end else if (8'h6c == _T_15[7:0]) begin
        image_108 <= io_pixelVal_in_3;
      end else if (8'h6c == _T_12[7:0]) begin
        image_108 <= io_pixelVal_in_2;
      end else if (8'h6c == _T_9[7:0]) begin
        image_108 <= io_pixelVal_in_1;
      end else if (8'h6c == _T_5[7:0]) begin
        image_108 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_109 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h6d == _T_27[7:0]) begin
        image_109 <= io_pixelVal_in_7;
      end else if (8'h6d == _T_24[7:0]) begin
        image_109 <= io_pixelVal_in_6;
      end else if (8'h6d == _T_21[7:0]) begin
        image_109 <= io_pixelVal_in_5;
      end else if (8'h6d == _T_18[7:0]) begin
        image_109 <= io_pixelVal_in_4;
      end else if (8'h6d == _T_15[7:0]) begin
        image_109 <= io_pixelVal_in_3;
      end else if (8'h6d == _T_12[7:0]) begin
        image_109 <= io_pixelVal_in_2;
      end else if (8'h6d == _T_9[7:0]) begin
        image_109 <= io_pixelVal_in_1;
      end else if (8'h6d == _T_5[7:0]) begin
        image_109 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_110 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h6e == _T_27[7:0]) begin
        image_110 <= io_pixelVal_in_7;
      end else if (8'h6e == _T_24[7:0]) begin
        image_110 <= io_pixelVal_in_6;
      end else if (8'h6e == _T_21[7:0]) begin
        image_110 <= io_pixelVal_in_5;
      end else if (8'h6e == _T_18[7:0]) begin
        image_110 <= io_pixelVal_in_4;
      end else if (8'h6e == _T_15[7:0]) begin
        image_110 <= io_pixelVal_in_3;
      end else if (8'h6e == _T_12[7:0]) begin
        image_110 <= io_pixelVal_in_2;
      end else if (8'h6e == _T_9[7:0]) begin
        image_110 <= io_pixelVal_in_1;
      end else if (8'h6e == _T_5[7:0]) begin
        image_110 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_111 <= 4'h3;
    end else if (io_valid_in) begin
      if (8'h6f == _T_27[7:0]) begin
        image_111 <= io_pixelVal_in_7;
      end else if (8'h6f == _T_24[7:0]) begin
        image_111 <= io_pixelVal_in_6;
      end else if (8'h6f == _T_21[7:0]) begin
        image_111 <= io_pixelVal_in_5;
      end else if (8'h6f == _T_18[7:0]) begin
        image_111 <= io_pixelVal_in_4;
      end else if (8'h6f == _T_15[7:0]) begin
        image_111 <= io_pixelVal_in_3;
      end else if (8'h6f == _T_12[7:0]) begin
        image_111 <= io_pixelVal_in_2;
      end else if (8'h6f == _T_9[7:0]) begin
        image_111 <= io_pixelVal_in_1;
      end else if (8'h6f == _T_5[7:0]) begin
        image_111 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_112 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h70 == _T_27[7:0]) begin
        image_112 <= io_pixelVal_in_7;
      end else if (8'h70 == _T_24[7:0]) begin
        image_112 <= io_pixelVal_in_6;
      end else if (8'h70 == _T_21[7:0]) begin
        image_112 <= io_pixelVal_in_5;
      end else if (8'h70 == _T_18[7:0]) begin
        image_112 <= io_pixelVal_in_4;
      end else if (8'h70 == _T_15[7:0]) begin
        image_112 <= io_pixelVal_in_3;
      end else if (8'h70 == _T_12[7:0]) begin
        image_112 <= io_pixelVal_in_2;
      end else if (8'h70 == _T_9[7:0]) begin
        image_112 <= io_pixelVal_in_1;
      end else if (8'h70 == _T_5[7:0]) begin
        image_112 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_113 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h71 == _T_27[7:0]) begin
        image_113 <= io_pixelVal_in_7;
      end else if (8'h71 == _T_24[7:0]) begin
        image_113 <= io_pixelVal_in_6;
      end else if (8'h71 == _T_21[7:0]) begin
        image_113 <= io_pixelVal_in_5;
      end else if (8'h71 == _T_18[7:0]) begin
        image_113 <= io_pixelVal_in_4;
      end else if (8'h71 == _T_15[7:0]) begin
        image_113 <= io_pixelVal_in_3;
      end else if (8'h71 == _T_12[7:0]) begin
        image_113 <= io_pixelVal_in_2;
      end else if (8'h71 == _T_9[7:0]) begin
        image_113 <= io_pixelVal_in_1;
      end else if (8'h71 == _T_5[7:0]) begin
        image_113 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_114 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h72 == _T_27[7:0]) begin
        image_114 <= io_pixelVal_in_7;
      end else if (8'h72 == _T_24[7:0]) begin
        image_114 <= io_pixelVal_in_6;
      end else if (8'h72 == _T_21[7:0]) begin
        image_114 <= io_pixelVal_in_5;
      end else if (8'h72 == _T_18[7:0]) begin
        image_114 <= io_pixelVal_in_4;
      end else if (8'h72 == _T_15[7:0]) begin
        image_114 <= io_pixelVal_in_3;
      end else if (8'h72 == _T_12[7:0]) begin
        image_114 <= io_pixelVal_in_2;
      end else if (8'h72 == _T_9[7:0]) begin
        image_114 <= io_pixelVal_in_1;
      end else if (8'h72 == _T_5[7:0]) begin
        image_114 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_115 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h73 == _T_27[7:0]) begin
        image_115 <= io_pixelVal_in_7;
      end else if (8'h73 == _T_24[7:0]) begin
        image_115 <= io_pixelVal_in_6;
      end else if (8'h73 == _T_21[7:0]) begin
        image_115 <= io_pixelVal_in_5;
      end else if (8'h73 == _T_18[7:0]) begin
        image_115 <= io_pixelVal_in_4;
      end else if (8'h73 == _T_15[7:0]) begin
        image_115 <= io_pixelVal_in_3;
      end else if (8'h73 == _T_12[7:0]) begin
        image_115 <= io_pixelVal_in_2;
      end else if (8'h73 == _T_9[7:0]) begin
        image_115 <= io_pixelVal_in_1;
      end else if (8'h73 == _T_5[7:0]) begin
        image_115 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_116 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h74 == _T_27[7:0]) begin
        image_116 <= io_pixelVal_in_7;
      end else if (8'h74 == _T_24[7:0]) begin
        image_116 <= io_pixelVal_in_6;
      end else if (8'h74 == _T_21[7:0]) begin
        image_116 <= io_pixelVal_in_5;
      end else if (8'h74 == _T_18[7:0]) begin
        image_116 <= io_pixelVal_in_4;
      end else if (8'h74 == _T_15[7:0]) begin
        image_116 <= io_pixelVal_in_3;
      end else if (8'h74 == _T_12[7:0]) begin
        image_116 <= io_pixelVal_in_2;
      end else if (8'h74 == _T_9[7:0]) begin
        image_116 <= io_pixelVal_in_1;
      end else if (8'h74 == _T_5[7:0]) begin
        image_116 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_117 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h75 == _T_27[7:0]) begin
        image_117 <= io_pixelVal_in_7;
      end else if (8'h75 == _T_24[7:0]) begin
        image_117 <= io_pixelVal_in_6;
      end else if (8'h75 == _T_21[7:0]) begin
        image_117 <= io_pixelVal_in_5;
      end else if (8'h75 == _T_18[7:0]) begin
        image_117 <= io_pixelVal_in_4;
      end else if (8'h75 == _T_15[7:0]) begin
        image_117 <= io_pixelVal_in_3;
      end else if (8'h75 == _T_12[7:0]) begin
        image_117 <= io_pixelVal_in_2;
      end else if (8'h75 == _T_9[7:0]) begin
        image_117 <= io_pixelVal_in_1;
      end else if (8'h75 == _T_5[7:0]) begin
        image_117 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_118 <= 4'h4;
    end else if (io_valid_in) begin
      if (8'h76 == _T_27[7:0]) begin
        image_118 <= io_pixelVal_in_7;
      end else if (8'h76 == _T_24[7:0]) begin
        image_118 <= io_pixelVal_in_6;
      end else if (8'h76 == _T_21[7:0]) begin
        image_118 <= io_pixelVal_in_5;
      end else if (8'h76 == _T_18[7:0]) begin
        image_118 <= io_pixelVal_in_4;
      end else if (8'h76 == _T_15[7:0]) begin
        image_118 <= io_pixelVal_in_3;
      end else if (8'h76 == _T_12[7:0]) begin
        image_118 <= io_pixelVal_in_2;
      end else if (8'h76 == _T_9[7:0]) begin
        image_118 <= io_pixelVal_in_1;
      end else if (8'h76 == _T_5[7:0]) begin
        image_118 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_119 <= 4'h3;
    end else if (io_valid_in) begin
      if (8'h77 == _T_27[7:0]) begin
        image_119 <= io_pixelVal_in_7;
      end else if (8'h77 == _T_24[7:0]) begin
        image_119 <= io_pixelVal_in_6;
      end else if (8'h77 == _T_21[7:0]) begin
        image_119 <= io_pixelVal_in_5;
      end else if (8'h77 == _T_18[7:0]) begin
        image_119 <= io_pixelVal_in_4;
      end else if (8'h77 == _T_15[7:0]) begin
        image_119 <= io_pixelVal_in_3;
      end else if (8'h77 == _T_12[7:0]) begin
        image_119 <= io_pixelVal_in_2;
      end else if (8'h77 == _T_9[7:0]) begin
        image_119 <= io_pixelVal_in_1;
      end else if (8'h77 == _T_5[7:0]) begin
        image_119 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_120 <= 4'h4;
    end else if (io_valid_in) begin
      if (8'h78 == _T_27[7:0]) begin
        image_120 <= io_pixelVal_in_7;
      end else if (8'h78 == _T_24[7:0]) begin
        image_120 <= io_pixelVal_in_6;
      end else if (8'h78 == _T_21[7:0]) begin
        image_120 <= io_pixelVal_in_5;
      end else if (8'h78 == _T_18[7:0]) begin
        image_120 <= io_pixelVal_in_4;
      end else if (8'h78 == _T_15[7:0]) begin
        image_120 <= io_pixelVal_in_3;
      end else if (8'h78 == _T_12[7:0]) begin
        image_120 <= io_pixelVal_in_2;
      end else if (8'h78 == _T_9[7:0]) begin
        image_120 <= io_pixelVal_in_1;
      end else if (8'h78 == _T_5[7:0]) begin
        image_120 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_121 <= 4'h4;
    end else if (io_valid_in) begin
      if (8'h79 == _T_27[7:0]) begin
        image_121 <= io_pixelVal_in_7;
      end else if (8'h79 == _T_24[7:0]) begin
        image_121 <= io_pixelVal_in_6;
      end else if (8'h79 == _T_21[7:0]) begin
        image_121 <= io_pixelVal_in_5;
      end else if (8'h79 == _T_18[7:0]) begin
        image_121 <= io_pixelVal_in_4;
      end else if (8'h79 == _T_15[7:0]) begin
        image_121 <= io_pixelVal_in_3;
      end else if (8'h79 == _T_12[7:0]) begin
        image_121 <= io_pixelVal_in_2;
      end else if (8'h79 == _T_9[7:0]) begin
        image_121 <= io_pixelVal_in_1;
      end else if (8'h79 == _T_5[7:0]) begin
        image_121 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_122 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h7a == _T_27[7:0]) begin
        image_122 <= io_pixelVal_in_7;
      end else if (8'h7a == _T_24[7:0]) begin
        image_122 <= io_pixelVal_in_6;
      end else if (8'h7a == _T_21[7:0]) begin
        image_122 <= io_pixelVal_in_5;
      end else if (8'h7a == _T_18[7:0]) begin
        image_122 <= io_pixelVal_in_4;
      end else if (8'h7a == _T_15[7:0]) begin
        image_122 <= io_pixelVal_in_3;
      end else if (8'h7a == _T_12[7:0]) begin
        image_122 <= io_pixelVal_in_2;
      end else if (8'h7a == _T_9[7:0]) begin
        image_122 <= io_pixelVal_in_1;
      end else if (8'h7a == _T_5[7:0]) begin
        image_122 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_123 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h7b == _T_27[7:0]) begin
        image_123 <= io_pixelVal_in_7;
      end else if (8'h7b == _T_24[7:0]) begin
        image_123 <= io_pixelVal_in_6;
      end else if (8'h7b == _T_21[7:0]) begin
        image_123 <= io_pixelVal_in_5;
      end else if (8'h7b == _T_18[7:0]) begin
        image_123 <= io_pixelVal_in_4;
      end else if (8'h7b == _T_15[7:0]) begin
        image_123 <= io_pixelVal_in_3;
      end else if (8'h7b == _T_12[7:0]) begin
        image_123 <= io_pixelVal_in_2;
      end else if (8'h7b == _T_9[7:0]) begin
        image_123 <= io_pixelVal_in_1;
      end else if (8'h7b == _T_5[7:0]) begin
        image_123 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_124 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h7c == _T_27[7:0]) begin
        image_124 <= io_pixelVal_in_7;
      end else if (8'h7c == _T_24[7:0]) begin
        image_124 <= io_pixelVal_in_6;
      end else if (8'h7c == _T_21[7:0]) begin
        image_124 <= io_pixelVal_in_5;
      end else if (8'h7c == _T_18[7:0]) begin
        image_124 <= io_pixelVal_in_4;
      end else if (8'h7c == _T_15[7:0]) begin
        image_124 <= io_pixelVal_in_3;
      end else if (8'h7c == _T_12[7:0]) begin
        image_124 <= io_pixelVal_in_2;
      end else if (8'h7c == _T_9[7:0]) begin
        image_124 <= io_pixelVal_in_1;
      end else if (8'h7c == _T_5[7:0]) begin
        image_124 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_125 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h7d == _T_27[7:0]) begin
        image_125 <= io_pixelVal_in_7;
      end else if (8'h7d == _T_24[7:0]) begin
        image_125 <= io_pixelVal_in_6;
      end else if (8'h7d == _T_21[7:0]) begin
        image_125 <= io_pixelVal_in_5;
      end else if (8'h7d == _T_18[7:0]) begin
        image_125 <= io_pixelVal_in_4;
      end else if (8'h7d == _T_15[7:0]) begin
        image_125 <= io_pixelVal_in_3;
      end else if (8'h7d == _T_12[7:0]) begin
        image_125 <= io_pixelVal_in_2;
      end else if (8'h7d == _T_9[7:0]) begin
        image_125 <= io_pixelVal_in_1;
      end else if (8'h7d == _T_5[7:0]) begin
        image_125 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_126 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h7e == _T_27[7:0]) begin
        image_126 <= io_pixelVal_in_7;
      end else if (8'h7e == _T_24[7:0]) begin
        image_126 <= io_pixelVal_in_6;
      end else if (8'h7e == _T_21[7:0]) begin
        image_126 <= io_pixelVal_in_5;
      end else if (8'h7e == _T_18[7:0]) begin
        image_126 <= io_pixelVal_in_4;
      end else if (8'h7e == _T_15[7:0]) begin
        image_126 <= io_pixelVal_in_3;
      end else if (8'h7e == _T_12[7:0]) begin
        image_126 <= io_pixelVal_in_2;
      end else if (8'h7e == _T_9[7:0]) begin
        image_126 <= io_pixelVal_in_1;
      end else if (8'h7e == _T_5[7:0]) begin
        image_126 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_127 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7f == _T_27[7:0]) begin
        image_127 <= io_pixelVal_in_7;
      end else if (8'h7f == _T_24[7:0]) begin
        image_127 <= io_pixelVal_in_6;
      end else if (8'h7f == _T_21[7:0]) begin
        image_127 <= io_pixelVal_in_5;
      end else if (8'h7f == _T_18[7:0]) begin
        image_127 <= io_pixelVal_in_4;
      end else if (8'h7f == _T_15[7:0]) begin
        image_127 <= io_pixelVal_in_3;
      end else if (8'h7f == _T_12[7:0]) begin
        image_127 <= io_pixelVal_in_2;
      end else if (8'h7f == _T_9[7:0]) begin
        image_127 <= io_pixelVal_in_1;
      end else if (8'h7f == _T_5[7:0]) begin
        image_127 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_128 <= 4'h4;
    end else if (io_valid_in) begin
      if (8'h80 == _T_27[7:0]) begin
        image_128 <= io_pixelVal_in_7;
      end else if (8'h80 == _T_24[7:0]) begin
        image_128 <= io_pixelVal_in_6;
      end else if (8'h80 == _T_21[7:0]) begin
        image_128 <= io_pixelVal_in_5;
      end else if (8'h80 == _T_18[7:0]) begin
        image_128 <= io_pixelVal_in_4;
      end else if (8'h80 == _T_15[7:0]) begin
        image_128 <= io_pixelVal_in_3;
      end else if (8'h80 == _T_12[7:0]) begin
        image_128 <= io_pixelVal_in_2;
      end else if (8'h80 == _T_9[7:0]) begin
        image_128 <= io_pixelVal_in_1;
      end else if (8'h80 == _T_5[7:0]) begin
        image_128 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_129 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h81 == _T_27[7:0]) begin
        image_129 <= io_pixelVal_in_7;
      end else if (8'h81 == _T_24[7:0]) begin
        image_129 <= io_pixelVal_in_6;
      end else if (8'h81 == _T_21[7:0]) begin
        image_129 <= io_pixelVal_in_5;
      end else if (8'h81 == _T_18[7:0]) begin
        image_129 <= io_pixelVal_in_4;
      end else if (8'h81 == _T_15[7:0]) begin
        image_129 <= io_pixelVal_in_3;
      end else if (8'h81 == _T_12[7:0]) begin
        image_129 <= io_pixelVal_in_2;
      end else if (8'h81 == _T_9[7:0]) begin
        image_129 <= io_pixelVal_in_1;
      end else if (8'h81 == _T_5[7:0]) begin
        image_129 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_130 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h82 == _T_27[7:0]) begin
        image_130 <= io_pixelVal_in_7;
      end else if (8'h82 == _T_24[7:0]) begin
        image_130 <= io_pixelVal_in_6;
      end else if (8'h82 == _T_21[7:0]) begin
        image_130 <= io_pixelVal_in_5;
      end else if (8'h82 == _T_18[7:0]) begin
        image_130 <= io_pixelVal_in_4;
      end else if (8'h82 == _T_15[7:0]) begin
        image_130 <= io_pixelVal_in_3;
      end else if (8'h82 == _T_12[7:0]) begin
        image_130 <= io_pixelVal_in_2;
      end else if (8'h82 == _T_9[7:0]) begin
        image_130 <= io_pixelVal_in_1;
      end else if (8'h82 == _T_5[7:0]) begin
        image_130 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_131 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h83 == _T_27[7:0]) begin
        image_131 <= io_pixelVal_in_7;
      end else if (8'h83 == _T_24[7:0]) begin
        image_131 <= io_pixelVal_in_6;
      end else if (8'h83 == _T_21[7:0]) begin
        image_131 <= io_pixelVal_in_5;
      end else if (8'h83 == _T_18[7:0]) begin
        image_131 <= io_pixelVal_in_4;
      end else if (8'h83 == _T_15[7:0]) begin
        image_131 <= io_pixelVal_in_3;
      end else if (8'h83 == _T_12[7:0]) begin
        image_131 <= io_pixelVal_in_2;
      end else if (8'h83 == _T_9[7:0]) begin
        image_131 <= io_pixelVal_in_1;
      end else if (8'h83 == _T_5[7:0]) begin
        image_131 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_132 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h84 == _T_27[7:0]) begin
        image_132 <= io_pixelVal_in_7;
      end else if (8'h84 == _T_24[7:0]) begin
        image_132 <= io_pixelVal_in_6;
      end else if (8'h84 == _T_21[7:0]) begin
        image_132 <= io_pixelVal_in_5;
      end else if (8'h84 == _T_18[7:0]) begin
        image_132 <= io_pixelVal_in_4;
      end else if (8'h84 == _T_15[7:0]) begin
        image_132 <= io_pixelVal_in_3;
      end else if (8'h84 == _T_12[7:0]) begin
        image_132 <= io_pixelVal_in_2;
      end else if (8'h84 == _T_9[7:0]) begin
        image_132 <= io_pixelVal_in_1;
      end else if (8'h84 == _T_5[7:0]) begin
        image_132 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_133 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h85 == _T_27[7:0]) begin
        image_133 <= io_pixelVal_in_7;
      end else if (8'h85 == _T_24[7:0]) begin
        image_133 <= io_pixelVal_in_6;
      end else if (8'h85 == _T_21[7:0]) begin
        image_133 <= io_pixelVal_in_5;
      end else if (8'h85 == _T_18[7:0]) begin
        image_133 <= io_pixelVal_in_4;
      end else if (8'h85 == _T_15[7:0]) begin
        image_133 <= io_pixelVal_in_3;
      end else if (8'h85 == _T_12[7:0]) begin
        image_133 <= io_pixelVal_in_2;
      end else if (8'h85 == _T_9[7:0]) begin
        image_133 <= io_pixelVal_in_1;
      end else if (8'h85 == _T_5[7:0]) begin
        image_133 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_134 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h86 == _T_27[7:0]) begin
        image_134 <= io_pixelVal_in_7;
      end else if (8'h86 == _T_24[7:0]) begin
        image_134 <= io_pixelVal_in_6;
      end else if (8'h86 == _T_21[7:0]) begin
        image_134 <= io_pixelVal_in_5;
      end else if (8'h86 == _T_18[7:0]) begin
        image_134 <= io_pixelVal_in_4;
      end else if (8'h86 == _T_15[7:0]) begin
        image_134 <= io_pixelVal_in_3;
      end else if (8'h86 == _T_12[7:0]) begin
        image_134 <= io_pixelVal_in_2;
      end else if (8'h86 == _T_9[7:0]) begin
        image_134 <= io_pixelVal_in_1;
      end else if (8'h86 == _T_5[7:0]) begin
        image_134 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_135 <= 4'h4;
    end else if (io_valid_in) begin
      if (8'h87 == _T_27[7:0]) begin
        image_135 <= io_pixelVal_in_7;
      end else if (8'h87 == _T_24[7:0]) begin
        image_135 <= io_pixelVal_in_6;
      end else if (8'h87 == _T_21[7:0]) begin
        image_135 <= io_pixelVal_in_5;
      end else if (8'h87 == _T_18[7:0]) begin
        image_135 <= io_pixelVal_in_4;
      end else if (8'h87 == _T_15[7:0]) begin
        image_135 <= io_pixelVal_in_3;
      end else if (8'h87 == _T_12[7:0]) begin
        image_135 <= io_pixelVal_in_2;
      end else if (8'h87 == _T_9[7:0]) begin
        image_135 <= io_pixelVal_in_1;
      end else if (8'h87 == _T_5[7:0]) begin
        image_135 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_136 <= 4'h4;
    end else if (io_valid_in) begin
      if (8'h88 == _T_27[7:0]) begin
        image_136 <= io_pixelVal_in_7;
      end else if (8'h88 == _T_24[7:0]) begin
        image_136 <= io_pixelVal_in_6;
      end else if (8'h88 == _T_21[7:0]) begin
        image_136 <= io_pixelVal_in_5;
      end else if (8'h88 == _T_18[7:0]) begin
        image_136 <= io_pixelVal_in_4;
      end else if (8'h88 == _T_15[7:0]) begin
        image_136 <= io_pixelVal_in_3;
      end else if (8'h88 == _T_12[7:0]) begin
        image_136 <= io_pixelVal_in_2;
      end else if (8'h88 == _T_9[7:0]) begin
        image_136 <= io_pixelVal_in_1;
      end else if (8'h88 == _T_5[7:0]) begin
        image_136 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_137 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h89 == _T_27[7:0]) begin
        image_137 <= io_pixelVal_in_7;
      end else if (8'h89 == _T_24[7:0]) begin
        image_137 <= io_pixelVal_in_6;
      end else if (8'h89 == _T_21[7:0]) begin
        image_137 <= io_pixelVal_in_5;
      end else if (8'h89 == _T_18[7:0]) begin
        image_137 <= io_pixelVal_in_4;
      end else if (8'h89 == _T_15[7:0]) begin
        image_137 <= io_pixelVal_in_3;
      end else if (8'h89 == _T_12[7:0]) begin
        image_137 <= io_pixelVal_in_2;
      end else if (8'h89 == _T_9[7:0]) begin
        image_137 <= io_pixelVal_in_1;
      end else if (8'h89 == _T_5[7:0]) begin
        image_137 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_138 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h8a == _T_27[7:0]) begin
        image_138 <= io_pixelVal_in_7;
      end else if (8'h8a == _T_24[7:0]) begin
        image_138 <= io_pixelVal_in_6;
      end else if (8'h8a == _T_21[7:0]) begin
        image_138 <= io_pixelVal_in_5;
      end else if (8'h8a == _T_18[7:0]) begin
        image_138 <= io_pixelVal_in_4;
      end else if (8'h8a == _T_15[7:0]) begin
        image_138 <= io_pixelVal_in_3;
      end else if (8'h8a == _T_12[7:0]) begin
        image_138 <= io_pixelVal_in_2;
      end else if (8'h8a == _T_9[7:0]) begin
        image_138 <= io_pixelVal_in_1;
      end else if (8'h8a == _T_5[7:0]) begin
        image_138 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_139 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h8b == _T_27[7:0]) begin
        image_139 <= io_pixelVal_in_7;
      end else if (8'h8b == _T_24[7:0]) begin
        image_139 <= io_pixelVal_in_6;
      end else if (8'h8b == _T_21[7:0]) begin
        image_139 <= io_pixelVal_in_5;
      end else if (8'h8b == _T_18[7:0]) begin
        image_139 <= io_pixelVal_in_4;
      end else if (8'h8b == _T_15[7:0]) begin
        image_139 <= io_pixelVal_in_3;
      end else if (8'h8b == _T_12[7:0]) begin
        image_139 <= io_pixelVal_in_2;
      end else if (8'h8b == _T_9[7:0]) begin
        image_139 <= io_pixelVal_in_1;
      end else if (8'h8b == _T_5[7:0]) begin
        image_139 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_140 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h8c == _T_27[7:0]) begin
        image_140 <= io_pixelVal_in_7;
      end else if (8'h8c == _T_24[7:0]) begin
        image_140 <= io_pixelVal_in_6;
      end else if (8'h8c == _T_21[7:0]) begin
        image_140 <= io_pixelVal_in_5;
      end else if (8'h8c == _T_18[7:0]) begin
        image_140 <= io_pixelVal_in_4;
      end else if (8'h8c == _T_15[7:0]) begin
        image_140 <= io_pixelVal_in_3;
      end else if (8'h8c == _T_12[7:0]) begin
        image_140 <= io_pixelVal_in_2;
      end else if (8'h8c == _T_9[7:0]) begin
        image_140 <= io_pixelVal_in_1;
      end else if (8'h8c == _T_5[7:0]) begin
        image_140 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_141 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h8d == _T_27[7:0]) begin
        image_141 <= io_pixelVal_in_7;
      end else if (8'h8d == _T_24[7:0]) begin
        image_141 <= io_pixelVal_in_6;
      end else if (8'h8d == _T_21[7:0]) begin
        image_141 <= io_pixelVal_in_5;
      end else if (8'h8d == _T_18[7:0]) begin
        image_141 <= io_pixelVal_in_4;
      end else if (8'h8d == _T_15[7:0]) begin
        image_141 <= io_pixelVal_in_3;
      end else if (8'h8d == _T_12[7:0]) begin
        image_141 <= io_pixelVal_in_2;
      end else if (8'h8d == _T_9[7:0]) begin
        image_141 <= io_pixelVal_in_1;
      end else if (8'h8d == _T_5[7:0]) begin
        image_141 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_142 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h8e == _T_27[7:0]) begin
        image_142 <= io_pixelVal_in_7;
      end else if (8'h8e == _T_24[7:0]) begin
        image_142 <= io_pixelVal_in_6;
      end else if (8'h8e == _T_21[7:0]) begin
        image_142 <= io_pixelVal_in_5;
      end else if (8'h8e == _T_18[7:0]) begin
        image_142 <= io_pixelVal_in_4;
      end else if (8'h8e == _T_15[7:0]) begin
        image_142 <= io_pixelVal_in_3;
      end else if (8'h8e == _T_12[7:0]) begin
        image_142 <= io_pixelVal_in_2;
      end else if (8'h8e == _T_9[7:0]) begin
        image_142 <= io_pixelVal_in_1;
      end else if (8'h8e == _T_5[7:0]) begin
        image_142 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_143 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8f == _T_27[7:0]) begin
        image_143 <= io_pixelVal_in_7;
      end else if (8'h8f == _T_24[7:0]) begin
        image_143 <= io_pixelVal_in_6;
      end else if (8'h8f == _T_21[7:0]) begin
        image_143 <= io_pixelVal_in_5;
      end else if (8'h8f == _T_18[7:0]) begin
        image_143 <= io_pixelVal_in_4;
      end else if (8'h8f == _T_15[7:0]) begin
        image_143 <= io_pixelVal_in_3;
      end else if (8'h8f == _T_12[7:0]) begin
        image_143 <= io_pixelVal_in_2;
      end else if (8'h8f == _T_9[7:0]) begin
        image_143 <= io_pixelVal_in_1;
      end else if (8'h8f == _T_5[7:0]) begin
        image_143 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_144 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h90 == _T_27[7:0]) begin
        image_144 <= io_pixelVal_in_7;
      end else if (8'h90 == _T_24[7:0]) begin
        image_144 <= io_pixelVal_in_6;
      end else if (8'h90 == _T_21[7:0]) begin
        image_144 <= io_pixelVal_in_5;
      end else if (8'h90 == _T_18[7:0]) begin
        image_144 <= io_pixelVal_in_4;
      end else if (8'h90 == _T_15[7:0]) begin
        image_144 <= io_pixelVal_in_3;
      end else if (8'h90 == _T_12[7:0]) begin
        image_144 <= io_pixelVal_in_2;
      end else if (8'h90 == _T_9[7:0]) begin
        image_144 <= io_pixelVal_in_1;
      end else if (8'h90 == _T_5[7:0]) begin
        image_144 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_145 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h91 == _T_27[7:0]) begin
        image_145 <= io_pixelVal_in_7;
      end else if (8'h91 == _T_24[7:0]) begin
        image_145 <= io_pixelVal_in_6;
      end else if (8'h91 == _T_21[7:0]) begin
        image_145 <= io_pixelVal_in_5;
      end else if (8'h91 == _T_18[7:0]) begin
        image_145 <= io_pixelVal_in_4;
      end else if (8'h91 == _T_15[7:0]) begin
        image_145 <= io_pixelVal_in_3;
      end else if (8'h91 == _T_12[7:0]) begin
        image_145 <= io_pixelVal_in_2;
      end else if (8'h91 == _T_9[7:0]) begin
        image_145 <= io_pixelVal_in_1;
      end else if (8'h91 == _T_5[7:0]) begin
        image_145 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_146 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h92 == _T_27[7:0]) begin
        image_146 <= io_pixelVal_in_7;
      end else if (8'h92 == _T_24[7:0]) begin
        image_146 <= io_pixelVal_in_6;
      end else if (8'h92 == _T_21[7:0]) begin
        image_146 <= io_pixelVal_in_5;
      end else if (8'h92 == _T_18[7:0]) begin
        image_146 <= io_pixelVal_in_4;
      end else if (8'h92 == _T_15[7:0]) begin
        image_146 <= io_pixelVal_in_3;
      end else if (8'h92 == _T_12[7:0]) begin
        image_146 <= io_pixelVal_in_2;
      end else if (8'h92 == _T_9[7:0]) begin
        image_146 <= io_pixelVal_in_1;
      end else if (8'h92 == _T_5[7:0]) begin
        image_146 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_147 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h93 == _T_27[7:0]) begin
        image_147 <= io_pixelVal_in_7;
      end else if (8'h93 == _T_24[7:0]) begin
        image_147 <= io_pixelVal_in_6;
      end else if (8'h93 == _T_21[7:0]) begin
        image_147 <= io_pixelVal_in_5;
      end else if (8'h93 == _T_18[7:0]) begin
        image_147 <= io_pixelVal_in_4;
      end else if (8'h93 == _T_15[7:0]) begin
        image_147 <= io_pixelVal_in_3;
      end else if (8'h93 == _T_12[7:0]) begin
        image_147 <= io_pixelVal_in_2;
      end else if (8'h93 == _T_9[7:0]) begin
        image_147 <= io_pixelVal_in_1;
      end else if (8'h93 == _T_5[7:0]) begin
        image_147 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_148 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h94 == _T_27[7:0]) begin
        image_148 <= io_pixelVal_in_7;
      end else if (8'h94 == _T_24[7:0]) begin
        image_148 <= io_pixelVal_in_6;
      end else if (8'h94 == _T_21[7:0]) begin
        image_148 <= io_pixelVal_in_5;
      end else if (8'h94 == _T_18[7:0]) begin
        image_148 <= io_pixelVal_in_4;
      end else if (8'h94 == _T_15[7:0]) begin
        image_148 <= io_pixelVal_in_3;
      end else if (8'h94 == _T_12[7:0]) begin
        image_148 <= io_pixelVal_in_2;
      end else if (8'h94 == _T_9[7:0]) begin
        image_148 <= io_pixelVal_in_1;
      end else if (8'h94 == _T_5[7:0]) begin
        image_148 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_149 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h95 == _T_27[7:0]) begin
        image_149 <= io_pixelVal_in_7;
      end else if (8'h95 == _T_24[7:0]) begin
        image_149 <= io_pixelVal_in_6;
      end else if (8'h95 == _T_21[7:0]) begin
        image_149 <= io_pixelVal_in_5;
      end else if (8'h95 == _T_18[7:0]) begin
        image_149 <= io_pixelVal_in_4;
      end else if (8'h95 == _T_15[7:0]) begin
        image_149 <= io_pixelVal_in_3;
      end else if (8'h95 == _T_12[7:0]) begin
        image_149 <= io_pixelVal_in_2;
      end else if (8'h95 == _T_9[7:0]) begin
        image_149 <= io_pixelVal_in_1;
      end else if (8'h95 == _T_5[7:0]) begin
        image_149 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_150 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h96 == _T_27[7:0]) begin
        image_150 <= io_pixelVal_in_7;
      end else if (8'h96 == _T_24[7:0]) begin
        image_150 <= io_pixelVal_in_6;
      end else if (8'h96 == _T_21[7:0]) begin
        image_150 <= io_pixelVal_in_5;
      end else if (8'h96 == _T_18[7:0]) begin
        image_150 <= io_pixelVal_in_4;
      end else if (8'h96 == _T_15[7:0]) begin
        image_150 <= io_pixelVal_in_3;
      end else if (8'h96 == _T_12[7:0]) begin
        image_150 <= io_pixelVal_in_2;
      end else if (8'h96 == _T_9[7:0]) begin
        image_150 <= io_pixelVal_in_1;
      end else if (8'h96 == _T_5[7:0]) begin
        image_150 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_151 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h97 == _T_27[7:0]) begin
        image_151 <= io_pixelVal_in_7;
      end else if (8'h97 == _T_24[7:0]) begin
        image_151 <= io_pixelVal_in_6;
      end else if (8'h97 == _T_21[7:0]) begin
        image_151 <= io_pixelVal_in_5;
      end else if (8'h97 == _T_18[7:0]) begin
        image_151 <= io_pixelVal_in_4;
      end else if (8'h97 == _T_15[7:0]) begin
        image_151 <= io_pixelVal_in_3;
      end else if (8'h97 == _T_12[7:0]) begin
        image_151 <= io_pixelVal_in_2;
      end else if (8'h97 == _T_9[7:0]) begin
        image_151 <= io_pixelVal_in_1;
      end else if (8'h97 == _T_5[7:0]) begin
        image_151 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_152 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h98 == _T_27[7:0]) begin
        image_152 <= io_pixelVal_in_7;
      end else if (8'h98 == _T_24[7:0]) begin
        image_152 <= io_pixelVal_in_6;
      end else if (8'h98 == _T_21[7:0]) begin
        image_152 <= io_pixelVal_in_5;
      end else if (8'h98 == _T_18[7:0]) begin
        image_152 <= io_pixelVal_in_4;
      end else if (8'h98 == _T_15[7:0]) begin
        image_152 <= io_pixelVal_in_3;
      end else if (8'h98 == _T_12[7:0]) begin
        image_152 <= io_pixelVal_in_2;
      end else if (8'h98 == _T_9[7:0]) begin
        image_152 <= io_pixelVal_in_1;
      end else if (8'h98 == _T_5[7:0]) begin
        image_152 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_153 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h99 == _T_27[7:0]) begin
        image_153 <= io_pixelVal_in_7;
      end else if (8'h99 == _T_24[7:0]) begin
        image_153 <= io_pixelVal_in_6;
      end else if (8'h99 == _T_21[7:0]) begin
        image_153 <= io_pixelVal_in_5;
      end else if (8'h99 == _T_18[7:0]) begin
        image_153 <= io_pixelVal_in_4;
      end else if (8'h99 == _T_15[7:0]) begin
        image_153 <= io_pixelVal_in_3;
      end else if (8'h99 == _T_12[7:0]) begin
        image_153 <= io_pixelVal_in_2;
      end else if (8'h99 == _T_9[7:0]) begin
        image_153 <= io_pixelVal_in_1;
      end else if (8'h99 == _T_5[7:0]) begin
        image_153 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_154 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h9a == _T_27[7:0]) begin
        image_154 <= io_pixelVal_in_7;
      end else if (8'h9a == _T_24[7:0]) begin
        image_154 <= io_pixelVal_in_6;
      end else if (8'h9a == _T_21[7:0]) begin
        image_154 <= io_pixelVal_in_5;
      end else if (8'h9a == _T_18[7:0]) begin
        image_154 <= io_pixelVal_in_4;
      end else if (8'h9a == _T_15[7:0]) begin
        image_154 <= io_pixelVal_in_3;
      end else if (8'h9a == _T_12[7:0]) begin
        image_154 <= io_pixelVal_in_2;
      end else if (8'h9a == _T_9[7:0]) begin
        image_154 <= io_pixelVal_in_1;
      end else if (8'h9a == _T_5[7:0]) begin
        image_154 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_155 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h9b == _T_27[7:0]) begin
        image_155 <= io_pixelVal_in_7;
      end else if (8'h9b == _T_24[7:0]) begin
        image_155 <= io_pixelVal_in_6;
      end else if (8'h9b == _T_21[7:0]) begin
        image_155 <= io_pixelVal_in_5;
      end else if (8'h9b == _T_18[7:0]) begin
        image_155 <= io_pixelVal_in_4;
      end else if (8'h9b == _T_15[7:0]) begin
        image_155 <= io_pixelVal_in_3;
      end else if (8'h9b == _T_12[7:0]) begin
        image_155 <= io_pixelVal_in_2;
      end else if (8'h9b == _T_9[7:0]) begin
        image_155 <= io_pixelVal_in_1;
      end else if (8'h9b == _T_5[7:0]) begin
        image_155 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_156 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'h9c == _T_27[7:0]) begin
        image_156 <= io_pixelVal_in_7;
      end else if (8'h9c == _T_24[7:0]) begin
        image_156 <= io_pixelVal_in_6;
      end else if (8'h9c == _T_21[7:0]) begin
        image_156 <= io_pixelVal_in_5;
      end else if (8'h9c == _T_18[7:0]) begin
        image_156 <= io_pixelVal_in_4;
      end else if (8'h9c == _T_15[7:0]) begin
        image_156 <= io_pixelVal_in_3;
      end else if (8'h9c == _T_12[7:0]) begin
        image_156 <= io_pixelVal_in_2;
      end else if (8'h9c == _T_9[7:0]) begin
        image_156 <= io_pixelVal_in_1;
      end else if (8'h9c == _T_5[7:0]) begin
        image_156 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_157 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h9d == _T_27[7:0]) begin
        image_157 <= io_pixelVal_in_7;
      end else if (8'h9d == _T_24[7:0]) begin
        image_157 <= io_pixelVal_in_6;
      end else if (8'h9d == _T_21[7:0]) begin
        image_157 <= io_pixelVal_in_5;
      end else if (8'h9d == _T_18[7:0]) begin
        image_157 <= io_pixelVal_in_4;
      end else if (8'h9d == _T_15[7:0]) begin
        image_157 <= io_pixelVal_in_3;
      end else if (8'h9d == _T_12[7:0]) begin
        image_157 <= io_pixelVal_in_2;
      end else if (8'h9d == _T_9[7:0]) begin
        image_157 <= io_pixelVal_in_1;
      end else if (8'h9d == _T_5[7:0]) begin
        image_157 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_158 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'h9e == _T_27[7:0]) begin
        image_158 <= io_pixelVal_in_7;
      end else if (8'h9e == _T_24[7:0]) begin
        image_158 <= io_pixelVal_in_6;
      end else if (8'h9e == _T_21[7:0]) begin
        image_158 <= io_pixelVal_in_5;
      end else if (8'h9e == _T_18[7:0]) begin
        image_158 <= io_pixelVal_in_4;
      end else if (8'h9e == _T_15[7:0]) begin
        image_158 <= io_pixelVal_in_3;
      end else if (8'h9e == _T_12[7:0]) begin
        image_158 <= io_pixelVal_in_2;
      end else if (8'h9e == _T_9[7:0]) begin
        image_158 <= io_pixelVal_in_1;
      end else if (8'h9e == _T_5[7:0]) begin
        image_158 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_159 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9f == _T_27[7:0]) begin
        image_159 <= io_pixelVal_in_7;
      end else if (8'h9f == _T_24[7:0]) begin
        image_159 <= io_pixelVal_in_6;
      end else if (8'h9f == _T_21[7:0]) begin
        image_159 <= io_pixelVal_in_5;
      end else if (8'h9f == _T_18[7:0]) begin
        image_159 <= io_pixelVal_in_4;
      end else if (8'h9f == _T_15[7:0]) begin
        image_159 <= io_pixelVal_in_3;
      end else if (8'h9f == _T_12[7:0]) begin
        image_159 <= io_pixelVal_in_2;
      end else if (8'h9f == _T_9[7:0]) begin
        image_159 <= io_pixelVal_in_1;
      end else if (8'h9f == _T_5[7:0]) begin
        image_159 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_160 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha0 == _T_27[7:0]) begin
        image_160 <= io_pixelVal_in_7;
      end else if (8'ha0 == _T_24[7:0]) begin
        image_160 <= io_pixelVal_in_6;
      end else if (8'ha0 == _T_21[7:0]) begin
        image_160 <= io_pixelVal_in_5;
      end else if (8'ha0 == _T_18[7:0]) begin
        image_160 <= io_pixelVal_in_4;
      end else if (8'ha0 == _T_15[7:0]) begin
        image_160 <= io_pixelVal_in_3;
      end else if (8'ha0 == _T_12[7:0]) begin
        image_160 <= io_pixelVal_in_2;
      end else if (8'ha0 == _T_9[7:0]) begin
        image_160 <= io_pixelVal_in_1;
      end else if (8'ha0 == _T_5[7:0]) begin
        image_160 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_161 <= 4'h4;
    end else if (io_valid_in) begin
      if (8'ha1 == _T_27[7:0]) begin
        image_161 <= io_pixelVal_in_7;
      end else if (8'ha1 == _T_24[7:0]) begin
        image_161 <= io_pixelVal_in_6;
      end else if (8'ha1 == _T_21[7:0]) begin
        image_161 <= io_pixelVal_in_5;
      end else if (8'ha1 == _T_18[7:0]) begin
        image_161 <= io_pixelVal_in_4;
      end else if (8'ha1 == _T_15[7:0]) begin
        image_161 <= io_pixelVal_in_3;
      end else if (8'ha1 == _T_12[7:0]) begin
        image_161 <= io_pixelVal_in_2;
      end else if (8'ha1 == _T_9[7:0]) begin
        image_161 <= io_pixelVal_in_1;
      end else if (8'ha1 == _T_5[7:0]) begin
        image_161 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_162 <= 4'h4;
    end else if (io_valid_in) begin
      if (8'ha2 == _T_27[7:0]) begin
        image_162 <= io_pixelVal_in_7;
      end else if (8'ha2 == _T_24[7:0]) begin
        image_162 <= io_pixelVal_in_6;
      end else if (8'ha2 == _T_21[7:0]) begin
        image_162 <= io_pixelVal_in_5;
      end else if (8'ha2 == _T_18[7:0]) begin
        image_162 <= io_pixelVal_in_4;
      end else if (8'ha2 == _T_15[7:0]) begin
        image_162 <= io_pixelVal_in_3;
      end else if (8'ha2 == _T_12[7:0]) begin
        image_162 <= io_pixelVal_in_2;
      end else if (8'ha2 == _T_9[7:0]) begin
        image_162 <= io_pixelVal_in_1;
      end else if (8'ha2 == _T_5[7:0]) begin
        image_162 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_163 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'ha3 == _T_27[7:0]) begin
        image_163 <= io_pixelVal_in_7;
      end else if (8'ha3 == _T_24[7:0]) begin
        image_163 <= io_pixelVal_in_6;
      end else if (8'ha3 == _T_21[7:0]) begin
        image_163 <= io_pixelVal_in_5;
      end else if (8'ha3 == _T_18[7:0]) begin
        image_163 <= io_pixelVal_in_4;
      end else if (8'ha3 == _T_15[7:0]) begin
        image_163 <= io_pixelVal_in_3;
      end else if (8'ha3 == _T_12[7:0]) begin
        image_163 <= io_pixelVal_in_2;
      end else if (8'ha3 == _T_9[7:0]) begin
        image_163 <= io_pixelVal_in_1;
      end else if (8'ha3 == _T_5[7:0]) begin
        image_163 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_164 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'ha4 == _T_27[7:0]) begin
        image_164 <= io_pixelVal_in_7;
      end else if (8'ha4 == _T_24[7:0]) begin
        image_164 <= io_pixelVal_in_6;
      end else if (8'ha4 == _T_21[7:0]) begin
        image_164 <= io_pixelVal_in_5;
      end else if (8'ha4 == _T_18[7:0]) begin
        image_164 <= io_pixelVal_in_4;
      end else if (8'ha4 == _T_15[7:0]) begin
        image_164 <= io_pixelVal_in_3;
      end else if (8'ha4 == _T_12[7:0]) begin
        image_164 <= io_pixelVal_in_2;
      end else if (8'ha4 == _T_9[7:0]) begin
        image_164 <= io_pixelVal_in_1;
      end else if (8'ha4 == _T_5[7:0]) begin
        image_164 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_165 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'ha5 == _T_27[7:0]) begin
        image_165 <= io_pixelVal_in_7;
      end else if (8'ha5 == _T_24[7:0]) begin
        image_165 <= io_pixelVal_in_6;
      end else if (8'ha5 == _T_21[7:0]) begin
        image_165 <= io_pixelVal_in_5;
      end else if (8'ha5 == _T_18[7:0]) begin
        image_165 <= io_pixelVal_in_4;
      end else if (8'ha5 == _T_15[7:0]) begin
        image_165 <= io_pixelVal_in_3;
      end else if (8'ha5 == _T_12[7:0]) begin
        image_165 <= io_pixelVal_in_2;
      end else if (8'ha5 == _T_9[7:0]) begin
        image_165 <= io_pixelVal_in_1;
      end else if (8'ha5 == _T_5[7:0]) begin
        image_165 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_166 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'ha6 == _T_27[7:0]) begin
        image_166 <= io_pixelVal_in_7;
      end else if (8'ha6 == _T_24[7:0]) begin
        image_166 <= io_pixelVal_in_6;
      end else if (8'ha6 == _T_21[7:0]) begin
        image_166 <= io_pixelVal_in_5;
      end else if (8'ha6 == _T_18[7:0]) begin
        image_166 <= io_pixelVal_in_4;
      end else if (8'ha6 == _T_15[7:0]) begin
        image_166 <= io_pixelVal_in_3;
      end else if (8'ha6 == _T_12[7:0]) begin
        image_166 <= io_pixelVal_in_2;
      end else if (8'ha6 == _T_9[7:0]) begin
        image_166 <= io_pixelVal_in_1;
      end else if (8'ha6 == _T_5[7:0]) begin
        image_166 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_167 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'ha7 == _T_27[7:0]) begin
        image_167 <= io_pixelVal_in_7;
      end else if (8'ha7 == _T_24[7:0]) begin
        image_167 <= io_pixelVal_in_6;
      end else if (8'ha7 == _T_21[7:0]) begin
        image_167 <= io_pixelVal_in_5;
      end else if (8'ha7 == _T_18[7:0]) begin
        image_167 <= io_pixelVal_in_4;
      end else if (8'ha7 == _T_15[7:0]) begin
        image_167 <= io_pixelVal_in_3;
      end else if (8'ha7 == _T_12[7:0]) begin
        image_167 <= io_pixelVal_in_2;
      end else if (8'ha7 == _T_9[7:0]) begin
        image_167 <= io_pixelVal_in_1;
      end else if (8'ha7 == _T_5[7:0]) begin
        image_167 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_168 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'ha8 == _T_27[7:0]) begin
        image_168 <= io_pixelVal_in_7;
      end else if (8'ha8 == _T_24[7:0]) begin
        image_168 <= io_pixelVal_in_6;
      end else if (8'ha8 == _T_21[7:0]) begin
        image_168 <= io_pixelVal_in_5;
      end else if (8'ha8 == _T_18[7:0]) begin
        image_168 <= io_pixelVal_in_4;
      end else if (8'ha8 == _T_15[7:0]) begin
        image_168 <= io_pixelVal_in_3;
      end else if (8'ha8 == _T_12[7:0]) begin
        image_168 <= io_pixelVal_in_2;
      end else if (8'ha8 == _T_9[7:0]) begin
        image_168 <= io_pixelVal_in_1;
      end else if (8'ha8 == _T_5[7:0]) begin
        image_168 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_169 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'ha9 == _T_27[7:0]) begin
        image_169 <= io_pixelVal_in_7;
      end else if (8'ha9 == _T_24[7:0]) begin
        image_169 <= io_pixelVal_in_6;
      end else if (8'ha9 == _T_21[7:0]) begin
        image_169 <= io_pixelVal_in_5;
      end else if (8'ha9 == _T_18[7:0]) begin
        image_169 <= io_pixelVal_in_4;
      end else if (8'ha9 == _T_15[7:0]) begin
        image_169 <= io_pixelVal_in_3;
      end else if (8'ha9 == _T_12[7:0]) begin
        image_169 <= io_pixelVal_in_2;
      end else if (8'ha9 == _T_9[7:0]) begin
        image_169 <= io_pixelVal_in_1;
      end else if (8'ha9 == _T_5[7:0]) begin
        image_169 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_170 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'haa == _T_27[7:0]) begin
        image_170 <= io_pixelVal_in_7;
      end else if (8'haa == _T_24[7:0]) begin
        image_170 <= io_pixelVal_in_6;
      end else if (8'haa == _T_21[7:0]) begin
        image_170 <= io_pixelVal_in_5;
      end else if (8'haa == _T_18[7:0]) begin
        image_170 <= io_pixelVal_in_4;
      end else if (8'haa == _T_15[7:0]) begin
        image_170 <= io_pixelVal_in_3;
      end else if (8'haa == _T_12[7:0]) begin
        image_170 <= io_pixelVal_in_2;
      end else if (8'haa == _T_9[7:0]) begin
        image_170 <= io_pixelVal_in_1;
      end else if (8'haa == _T_5[7:0]) begin
        image_170 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_171 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'hab == _T_27[7:0]) begin
        image_171 <= io_pixelVal_in_7;
      end else if (8'hab == _T_24[7:0]) begin
        image_171 <= io_pixelVal_in_6;
      end else if (8'hab == _T_21[7:0]) begin
        image_171 <= io_pixelVal_in_5;
      end else if (8'hab == _T_18[7:0]) begin
        image_171 <= io_pixelVal_in_4;
      end else if (8'hab == _T_15[7:0]) begin
        image_171 <= io_pixelVal_in_3;
      end else if (8'hab == _T_12[7:0]) begin
        image_171 <= io_pixelVal_in_2;
      end else if (8'hab == _T_9[7:0]) begin
        image_171 <= io_pixelVal_in_1;
      end else if (8'hab == _T_5[7:0]) begin
        image_171 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_172 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'hac == _T_27[7:0]) begin
        image_172 <= io_pixelVal_in_7;
      end else if (8'hac == _T_24[7:0]) begin
        image_172 <= io_pixelVal_in_6;
      end else if (8'hac == _T_21[7:0]) begin
        image_172 <= io_pixelVal_in_5;
      end else if (8'hac == _T_18[7:0]) begin
        image_172 <= io_pixelVal_in_4;
      end else if (8'hac == _T_15[7:0]) begin
        image_172 <= io_pixelVal_in_3;
      end else if (8'hac == _T_12[7:0]) begin
        image_172 <= io_pixelVal_in_2;
      end else if (8'hac == _T_9[7:0]) begin
        image_172 <= io_pixelVal_in_1;
      end else if (8'hac == _T_5[7:0]) begin
        image_172 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_173 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'had == _T_27[7:0]) begin
        image_173 <= io_pixelVal_in_7;
      end else if (8'had == _T_24[7:0]) begin
        image_173 <= io_pixelVal_in_6;
      end else if (8'had == _T_21[7:0]) begin
        image_173 <= io_pixelVal_in_5;
      end else if (8'had == _T_18[7:0]) begin
        image_173 <= io_pixelVal_in_4;
      end else if (8'had == _T_15[7:0]) begin
        image_173 <= io_pixelVal_in_3;
      end else if (8'had == _T_12[7:0]) begin
        image_173 <= io_pixelVal_in_2;
      end else if (8'had == _T_9[7:0]) begin
        image_173 <= io_pixelVal_in_1;
      end else if (8'had == _T_5[7:0]) begin
        image_173 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_174 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'hae == _T_27[7:0]) begin
        image_174 <= io_pixelVal_in_7;
      end else if (8'hae == _T_24[7:0]) begin
        image_174 <= io_pixelVal_in_6;
      end else if (8'hae == _T_21[7:0]) begin
        image_174 <= io_pixelVal_in_5;
      end else if (8'hae == _T_18[7:0]) begin
        image_174 <= io_pixelVal_in_4;
      end else if (8'hae == _T_15[7:0]) begin
        image_174 <= io_pixelVal_in_3;
      end else if (8'hae == _T_12[7:0]) begin
        image_174 <= io_pixelVal_in_2;
      end else if (8'hae == _T_9[7:0]) begin
        image_174 <= io_pixelVal_in_1;
      end else if (8'hae == _T_5[7:0]) begin
        image_174 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_175 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'haf == _T_27[7:0]) begin
        image_175 <= io_pixelVal_in_7;
      end else if (8'haf == _T_24[7:0]) begin
        image_175 <= io_pixelVal_in_6;
      end else if (8'haf == _T_21[7:0]) begin
        image_175 <= io_pixelVal_in_5;
      end else if (8'haf == _T_18[7:0]) begin
        image_175 <= io_pixelVal_in_4;
      end else if (8'haf == _T_15[7:0]) begin
        image_175 <= io_pixelVal_in_3;
      end else if (8'haf == _T_12[7:0]) begin
        image_175 <= io_pixelVal_in_2;
      end else if (8'haf == _T_9[7:0]) begin
        image_175 <= io_pixelVal_in_1;
      end else if (8'haf == _T_5[7:0]) begin
        image_175 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_176 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb0 == _T_27[7:0]) begin
        image_176 <= io_pixelVal_in_7;
      end else if (8'hb0 == _T_24[7:0]) begin
        image_176 <= io_pixelVal_in_6;
      end else if (8'hb0 == _T_21[7:0]) begin
        image_176 <= io_pixelVal_in_5;
      end else if (8'hb0 == _T_18[7:0]) begin
        image_176 <= io_pixelVal_in_4;
      end else if (8'hb0 == _T_15[7:0]) begin
        image_176 <= io_pixelVal_in_3;
      end else if (8'hb0 == _T_12[7:0]) begin
        image_176 <= io_pixelVal_in_2;
      end else if (8'hb0 == _T_9[7:0]) begin
        image_176 <= io_pixelVal_in_1;
      end else if (8'hb0 == _T_5[7:0]) begin
        image_176 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_177 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb1 == _T_27[7:0]) begin
        image_177 <= io_pixelVal_in_7;
      end else if (8'hb1 == _T_24[7:0]) begin
        image_177 <= io_pixelVal_in_6;
      end else if (8'hb1 == _T_21[7:0]) begin
        image_177 <= io_pixelVal_in_5;
      end else if (8'hb1 == _T_18[7:0]) begin
        image_177 <= io_pixelVal_in_4;
      end else if (8'hb1 == _T_15[7:0]) begin
        image_177 <= io_pixelVal_in_3;
      end else if (8'hb1 == _T_12[7:0]) begin
        image_177 <= io_pixelVal_in_2;
      end else if (8'hb1 == _T_9[7:0]) begin
        image_177 <= io_pixelVal_in_1;
      end else if (8'hb1 == _T_5[7:0]) begin
        image_177 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_178 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb2 == _T_27[7:0]) begin
        image_178 <= io_pixelVal_in_7;
      end else if (8'hb2 == _T_24[7:0]) begin
        image_178 <= io_pixelVal_in_6;
      end else if (8'hb2 == _T_21[7:0]) begin
        image_178 <= io_pixelVal_in_5;
      end else if (8'hb2 == _T_18[7:0]) begin
        image_178 <= io_pixelVal_in_4;
      end else if (8'hb2 == _T_15[7:0]) begin
        image_178 <= io_pixelVal_in_3;
      end else if (8'hb2 == _T_12[7:0]) begin
        image_178 <= io_pixelVal_in_2;
      end else if (8'hb2 == _T_9[7:0]) begin
        image_178 <= io_pixelVal_in_1;
      end else if (8'hb2 == _T_5[7:0]) begin
        image_178 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_179 <= 4'h4;
    end else if (io_valid_in) begin
      if (8'hb3 == _T_27[7:0]) begin
        image_179 <= io_pixelVal_in_7;
      end else if (8'hb3 == _T_24[7:0]) begin
        image_179 <= io_pixelVal_in_6;
      end else if (8'hb3 == _T_21[7:0]) begin
        image_179 <= io_pixelVal_in_5;
      end else if (8'hb3 == _T_18[7:0]) begin
        image_179 <= io_pixelVal_in_4;
      end else if (8'hb3 == _T_15[7:0]) begin
        image_179 <= io_pixelVal_in_3;
      end else if (8'hb3 == _T_12[7:0]) begin
        image_179 <= io_pixelVal_in_2;
      end else if (8'hb3 == _T_9[7:0]) begin
        image_179 <= io_pixelVal_in_1;
      end else if (8'hb3 == _T_5[7:0]) begin
        image_179 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_180 <= 4'h4;
    end else if (io_valid_in) begin
      if (8'hb4 == _T_27[7:0]) begin
        image_180 <= io_pixelVal_in_7;
      end else if (8'hb4 == _T_24[7:0]) begin
        image_180 <= io_pixelVal_in_6;
      end else if (8'hb4 == _T_21[7:0]) begin
        image_180 <= io_pixelVal_in_5;
      end else if (8'hb4 == _T_18[7:0]) begin
        image_180 <= io_pixelVal_in_4;
      end else if (8'hb4 == _T_15[7:0]) begin
        image_180 <= io_pixelVal_in_3;
      end else if (8'hb4 == _T_12[7:0]) begin
        image_180 <= io_pixelVal_in_2;
      end else if (8'hb4 == _T_9[7:0]) begin
        image_180 <= io_pixelVal_in_1;
      end else if (8'hb4 == _T_5[7:0]) begin
        image_180 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_181 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'hb5 == _T_27[7:0]) begin
        image_181 <= io_pixelVal_in_7;
      end else if (8'hb5 == _T_24[7:0]) begin
        image_181 <= io_pixelVal_in_6;
      end else if (8'hb5 == _T_21[7:0]) begin
        image_181 <= io_pixelVal_in_5;
      end else if (8'hb5 == _T_18[7:0]) begin
        image_181 <= io_pixelVal_in_4;
      end else if (8'hb5 == _T_15[7:0]) begin
        image_181 <= io_pixelVal_in_3;
      end else if (8'hb5 == _T_12[7:0]) begin
        image_181 <= io_pixelVal_in_2;
      end else if (8'hb5 == _T_9[7:0]) begin
        image_181 <= io_pixelVal_in_1;
      end else if (8'hb5 == _T_5[7:0]) begin
        image_181 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_182 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'hb6 == _T_27[7:0]) begin
        image_182 <= io_pixelVal_in_7;
      end else if (8'hb6 == _T_24[7:0]) begin
        image_182 <= io_pixelVal_in_6;
      end else if (8'hb6 == _T_21[7:0]) begin
        image_182 <= io_pixelVal_in_5;
      end else if (8'hb6 == _T_18[7:0]) begin
        image_182 <= io_pixelVal_in_4;
      end else if (8'hb6 == _T_15[7:0]) begin
        image_182 <= io_pixelVal_in_3;
      end else if (8'hb6 == _T_12[7:0]) begin
        image_182 <= io_pixelVal_in_2;
      end else if (8'hb6 == _T_9[7:0]) begin
        image_182 <= io_pixelVal_in_1;
      end else if (8'hb6 == _T_5[7:0]) begin
        image_182 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_183 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'hb7 == _T_27[7:0]) begin
        image_183 <= io_pixelVal_in_7;
      end else if (8'hb7 == _T_24[7:0]) begin
        image_183 <= io_pixelVal_in_6;
      end else if (8'hb7 == _T_21[7:0]) begin
        image_183 <= io_pixelVal_in_5;
      end else if (8'hb7 == _T_18[7:0]) begin
        image_183 <= io_pixelVal_in_4;
      end else if (8'hb7 == _T_15[7:0]) begin
        image_183 <= io_pixelVal_in_3;
      end else if (8'hb7 == _T_12[7:0]) begin
        image_183 <= io_pixelVal_in_2;
      end else if (8'hb7 == _T_9[7:0]) begin
        image_183 <= io_pixelVal_in_1;
      end else if (8'hb7 == _T_5[7:0]) begin
        image_183 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_184 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'hb8 == _T_27[7:0]) begin
        image_184 <= io_pixelVal_in_7;
      end else if (8'hb8 == _T_24[7:0]) begin
        image_184 <= io_pixelVal_in_6;
      end else if (8'hb8 == _T_21[7:0]) begin
        image_184 <= io_pixelVal_in_5;
      end else if (8'hb8 == _T_18[7:0]) begin
        image_184 <= io_pixelVal_in_4;
      end else if (8'hb8 == _T_15[7:0]) begin
        image_184 <= io_pixelVal_in_3;
      end else if (8'hb8 == _T_12[7:0]) begin
        image_184 <= io_pixelVal_in_2;
      end else if (8'hb8 == _T_9[7:0]) begin
        image_184 <= io_pixelVal_in_1;
      end else if (8'hb8 == _T_5[7:0]) begin
        image_184 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_185 <= 4'h6;
    end else if (io_valid_in) begin
      if (8'hb9 == _T_27[7:0]) begin
        image_185 <= io_pixelVal_in_7;
      end else if (8'hb9 == _T_24[7:0]) begin
        image_185 <= io_pixelVal_in_6;
      end else if (8'hb9 == _T_21[7:0]) begin
        image_185 <= io_pixelVal_in_5;
      end else if (8'hb9 == _T_18[7:0]) begin
        image_185 <= io_pixelVal_in_4;
      end else if (8'hb9 == _T_15[7:0]) begin
        image_185 <= io_pixelVal_in_3;
      end else if (8'hb9 == _T_12[7:0]) begin
        image_185 <= io_pixelVal_in_2;
      end else if (8'hb9 == _T_9[7:0]) begin
        image_185 <= io_pixelVal_in_1;
      end else if (8'hb9 == _T_5[7:0]) begin
        image_185 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_186 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'hba == _T_27[7:0]) begin
        image_186 <= io_pixelVal_in_7;
      end else if (8'hba == _T_24[7:0]) begin
        image_186 <= io_pixelVal_in_6;
      end else if (8'hba == _T_21[7:0]) begin
        image_186 <= io_pixelVal_in_5;
      end else if (8'hba == _T_18[7:0]) begin
        image_186 <= io_pixelVal_in_4;
      end else if (8'hba == _T_15[7:0]) begin
        image_186 <= io_pixelVal_in_3;
      end else if (8'hba == _T_12[7:0]) begin
        image_186 <= io_pixelVal_in_2;
      end else if (8'hba == _T_9[7:0]) begin
        image_186 <= io_pixelVal_in_1;
      end else if (8'hba == _T_5[7:0]) begin
        image_186 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_187 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'hbb == _T_27[7:0]) begin
        image_187 <= io_pixelVal_in_7;
      end else if (8'hbb == _T_24[7:0]) begin
        image_187 <= io_pixelVal_in_6;
      end else if (8'hbb == _T_21[7:0]) begin
        image_187 <= io_pixelVal_in_5;
      end else if (8'hbb == _T_18[7:0]) begin
        image_187 <= io_pixelVal_in_4;
      end else if (8'hbb == _T_15[7:0]) begin
        image_187 <= io_pixelVal_in_3;
      end else if (8'hbb == _T_12[7:0]) begin
        image_187 <= io_pixelVal_in_2;
      end else if (8'hbb == _T_9[7:0]) begin
        image_187 <= io_pixelVal_in_1;
      end else if (8'hbb == _T_5[7:0]) begin
        image_187 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_188 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'hbc == _T_27[7:0]) begin
        image_188 <= io_pixelVal_in_7;
      end else if (8'hbc == _T_24[7:0]) begin
        image_188 <= io_pixelVal_in_6;
      end else if (8'hbc == _T_21[7:0]) begin
        image_188 <= io_pixelVal_in_5;
      end else if (8'hbc == _T_18[7:0]) begin
        image_188 <= io_pixelVal_in_4;
      end else if (8'hbc == _T_15[7:0]) begin
        image_188 <= io_pixelVal_in_3;
      end else if (8'hbc == _T_12[7:0]) begin
        image_188 <= io_pixelVal_in_2;
      end else if (8'hbc == _T_9[7:0]) begin
        image_188 <= io_pixelVal_in_1;
      end else if (8'hbc == _T_5[7:0]) begin
        image_188 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_189 <= 4'h5;
    end else if (io_valid_in) begin
      if (8'hbd == _T_27[7:0]) begin
        image_189 <= io_pixelVal_in_7;
      end else if (8'hbd == _T_24[7:0]) begin
        image_189 <= io_pixelVal_in_6;
      end else if (8'hbd == _T_21[7:0]) begin
        image_189 <= io_pixelVal_in_5;
      end else if (8'hbd == _T_18[7:0]) begin
        image_189 <= io_pixelVal_in_4;
      end else if (8'hbd == _T_15[7:0]) begin
        image_189 <= io_pixelVal_in_3;
      end else if (8'hbd == _T_12[7:0]) begin
        image_189 <= io_pixelVal_in_2;
      end else if (8'hbd == _T_9[7:0]) begin
        image_189 <= io_pixelVal_in_1;
      end else if (8'hbd == _T_5[7:0]) begin
        image_189 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_190 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbe == _T_27[7:0]) begin
        image_190 <= io_pixelVal_in_7;
      end else if (8'hbe == _T_24[7:0]) begin
        image_190 <= io_pixelVal_in_6;
      end else if (8'hbe == _T_21[7:0]) begin
        image_190 <= io_pixelVal_in_5;
      end else if (8'hbe == _T_18[7:0]) begin
        image_190 <= io_pixelVal_in_4;
      end else if (8'hbe == _T_15[7:0]) begin
        image_190 <= io_pixelVal_in_3;
      end else if (8'hbe == _T_12[7:0]) begin
        image_190 <= io_pixelVal_in_2;
      end else if (8'hbe == _T_9[7:0]) begin
        image_190 <= io_pixelVal_in_1;
      end else if (8'hbe == _T_5[7:0]) begin
        image_190 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      image_191 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbf == _T_27[7:0]) begin
        image_191 <= io_pixelVal_in_7;
      end else if (8'hbf == _T_24[7:0]) begin
        image_191 <= io_pixelVal_in_6;
      end else if (8'hbf == _T_21[7:0]) begin
        image_191 <= io_pixelVal_in_5;
      end else if (8'hbf == _T_18[7:0]) begin
        image_191 <= io_pixelVal_in_4;
      end else if (8'hbf == _T_15[7:0]) begin
        image_191 <= io_pixelVal_in_3;
      end else if (8'hbf == _T_12[7:0]) begin
        image_191 <= io_pixelVal_in_2;
      end else if (8'hbf == _T_9[7:0]) begin
        image_191 <= io_pixelVal_in_1;
      end else if (8'hbf == _T_5[7:0]) begin
        image_191 <= io_pixelVal_in_0;
      end
    end
    if (reset) begin
      pixelIndex <= 32'h0;
    end else if (io_valid_in) begin
      if (_T_32) begin
        pixelIndex <= 32'h0;
      end else begin
        pixelIndex <= _T_30;
      end
    end
  end
endmodule
