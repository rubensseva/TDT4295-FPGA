module DotProd(
  input        clock,
  input        reset,
  input  [7:0] io_dataInA,
  input  [7:0] io_dataInB,
  output [8:0] io_dataOut,
  output       io_outputValid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] countVal; // @[Counter.scala 29:33]
  wire  countReset = countVal == 4'h8; // @[Counter.scala 38:24]
  wire [3:0] _T_2 = countVal + 4'h1; // @[Counter.scala 39:22]
  reg [8:0] accumulator; // @[DotProd.scala 19:28]
  wire [15:0] product = $signed(io_dataInA) * $signed(io_dataInB); // @[DotProd.scala 20:35]
  wire [15:0] _GEN_5 = {{7{accumulator[8]}},accumulator}; // @[DotProd.scala 21:30]
  wire [15:0] _T_6 = $signed(_GEN_5) + $signed(product); // @[DotProd.scala 21:30]
  wire [15:0] _GEN_4 = countReset ? $signed(16'sh0) : $signed(_T_6); // @[DotProd.scala 25:20]
  assign io_dataOut = _T_6[8:0]; // @[DotProd.scala 23:14]
  assign io_outputValid = countVal == 4'h8; // @[DotProd.scala 26:20 DotProd.scala 29:20]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  countVal = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  accumulator = _RAND_1[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      countVal <= 4'h0;
    end else if (countReset) begin
      countVal <= 4'h0;
    end else begin
      countVal <= _T_2;
    end
    if (reset) begin
      accumulator <= 9'sh0;
    end else begin
      accumulator <= _GEN_4[8:0];
    end
  end
endmodule
module KernelConvolution(
  input        clock,
  input        reset,
  input  [4:0] io_kernelVal_in,
  input  [3:0] io_pixelVal_in_0,
  input  [3:0] io_pixelVal_in_1,
  input  [3:0] io_pixelVal_in_2,
  input  [3:0] io_pixelVal_in_3,
  input  [3:0] io_pixelVal_in_4,
  input  [3:0] io_pixelVal_in_5,
  input  [3:0] io_pixelVal_in_6,
  input  [3:0] io_pixelVal_in_7,
  output [8:0] io_pixelVal_out_0,
  output [8:0] io_pixelVal_out_1,
  output [8:0] io_pixelVal_out_2,
  output [8:0] io_pixelVal_out_3,
  output [8:0] io_pixelVal_out_4,
  output [8:0] io_pixelVal_out_5,
  output [8:0] io_pixelVal_out_6,
  output [8:0] io_pixelVal_out_7,
  output       io_valid_out
);
  wire  DotProd_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_1_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_1_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_1_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_1_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_1_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_1_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_2_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_2_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_2_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_2_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_2_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_2_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_3_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_3_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_3_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_3_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_3_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_3_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_4_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_4_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_4_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_4_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_4_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_4_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_5_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_5_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_5_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_5_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_5_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_5_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_6_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_6_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_6_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_6_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_6_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_6_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_7_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_7_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_7_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_7_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_7_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_7_io_outputValid; // @[KernelConvolution.scala 21:58]
  DotProd DotProd ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_clock),
    .reset(DotProd_reset),
    .io_dataInA(DotProd_io_dataInA),
    .io_dataInB(DotProd_io_dataInB),
    .io_dataOut(DotProd_io_dataOut),
    .io_outputValid(DotProd_io_outputValid)
  );
  DotProd DotProd_1 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_1_clock),
    .reset(DotProd_1_reset),
    .io_dataInA(DotProd_1_io_dataInA),
    .io_dataInB(DotProd_1_io_dataInB),
    .io_dataOut(DotProd_1_io_dataOut),
    .io_outputValid(DotProd_1_io_outputValid)
  );
  DotProd DotProd_2 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_2_clock),
    .reset(DotProd_2_reset),
    .io_dataInA(DotProd_2_io_dataInA),
    .io_dataInB(DotProd_2_io_dataInB),
    .io_dataOut(DotProd_2_io_dataOut),
    .io_outputValid(DotProd_2_io_outputValid)
  );
  DotProd DotProd_3 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_3_clock),
    .reset(DotProd_3_reset),
    .io_dataInA(DotProd_3_io_dataInA),
    .io_dataInB(DotProd_3_io_dataInB),
    .io_dataOut(DotProd_3_io_dataOut),
    .io_outputValid(DotProd_3_io_outputValid)
  );
  DotProd DotProd_4 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_4_clock),
    .reset(DotProd_4_reset),
    .io_dataInA(DotProd_4_io_dataInA),
    .io_dataInB(DotProd_4_io_dataInB),
    .io_dataOut(DotProd_4_io_dataOut),
    .io_outputValid(DotProd_4_io_outputValid)
  );
  DotProd DotProd_5 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_5_clock),
    .reset(DotProd_5_reset),
    .io_dataInA(DotProd_5_io_dataInA),
    .io_dataInB(DotProd_5_io_dataInB),
    .io_dataOut(DotProd_5_io_dataOut),
    .io_outputValid(DotProd_5_io_outputValid)
  );
  DotProd DotProd_6 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_6_clock),
    .reset(DotProd_6_reset),
    .io_dataInA(DotProd_6_io_dataInA),
    .io_dataInB(DotProd_6_io_dataInB),
    .io_dataOut(DotProd_6_io_dataOut),
    .io_outputValid(DotProd_6_io_outputValid)
  );
  DotProd DotProd_7 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_7_clock),
    .reset(DotProd_7_reset),
    .io_dataInA(DotProd_7_io_dataInA),
    .io_dataInB(DotProd_7_io_dataInB),
    .io_dataOut(DotProd_7_io_dataOut),
    .io_outputValid(DotProd_7_io_outputValid)
  );
  assign io_pixelVal_out_0 = DotProd_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_1 = DotProd_1_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_2 = DotProd_2_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_3 = DotProd_3_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_4 = DotProd_4_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_5 = DotProd_5_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_6 = DotProd_6_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_7 = DotProd_7_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_valid_out = DotProd_io_outputValid; // @[KernelConvolution.scala 35:30]
  assign DotProd_clock = clock;
  assign DotProd_reset = reset;
  assign DotProd_io_dataInA = {{4'd0}, io_pixelVal_in_0}; // @[KernelConvolution.scala 21:32]
  assign DotProd_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_1_clock = clock;
  assign DotProd_1_reset = reset;
  assign DotProd_1_io_dataInA = {{4'd0}, io_pixelVal_in_1}; // @[KernelConvolution.scala 21:32]
  assign DotProd_1_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_2_clock = clock;
  assign DotProd_2_reset = reset;
  assign DotProd_2_io_dataInA = {{4'd0}, io_pixelVal_in_2}; // @[KernelConvolution.scala 21:32]
  assign DotProd_2_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_3_clock = clock;
  assign DotProd_3_reset = reset;
  assign DotProd_3_io_dataInA = {{4'd0}, io_pixelVal_in_3}; // @[KernelConvolution.scala 21:32]
  assign DotProd_3_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_4_clock = clock;
  assign DotProd_4_reset = reset;
  assign DotProd_4_io_dataInA = {{4'd0}, io_pixelVal_in_4}; // @[KernelConvolution.scala 21:32]
  assign DotProd_4_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_5_clock = clock;
  assign DotProd_5_reset = reset;
  assign DotProd_5_io_dataInA = {{4'd0}, io_pixelVal_in_5}; // @[KernelConvolution.scala 21:32]
  assign DotProd_5_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_6_clock = clock;
  assign DotProd_6_reset = reset;
  assign DotProd_6_io_dataInA = {{4'd0}, io_pixelVal_in_6}; // @[KernelConvolution.scala 21:32]
  assign DotProd_6_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_7_clock = clock;
  assign DotProd_7_reset = reset;
  assign DotProd_7_io_dataInA = {{4'd0}, io_pixelVal_in_7}; // @[KernelConvolution.scala 21:32]
  assign DotProd_7_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
endmodule
module Filter(
  input        clock,
  input        reset,
  input  [5:0] io_SPI_filterIndex,
  input        io_SPI_distort,
  output [3:0] io_pixelVal_out_0_0,
  output [3:0] io_pixelVal_out_0_1,
  output [3:0] io_pixelVal_out_0_2,
  output [3:0] io_pixelVal_out_0_3,
  output [3:0] io_pixelVal_out_0_4,
  output [3:0] io_pixelVal_out_0_5,
  output [3:0] io_pixelVal_out_0_6,
  output [3:0] io_pixelVal_out_0_7,
  output [3:0] io_pixelVal_out_1_0,
  output [3:0] io_pixelVal_out_1_1,
  output [3:0] io_pixelVal_out_1_2,
  output [3:0] io_pixelVal_out_1_3,
  output [3:0] io_pixelVal_out_1_4,
  output [3:0] io_pixelVal_out_1_5,
  output [3:0] io_pixelVal_out_1_6,
  output [3:0] io_pixelVal_out_1_7,
  output [3:0] io_pixelVal_out_2_0,
  output [3:0] io_pixelVal_out_2_1,
  output [3:0] io_pixelVal_out_2_2,
  output [3:0] io_pixelVal_out_2_3,
  output [3:0] io_pixelVal_out_2_4,
  output [3:0] io_pixelVal_out_2_5,
  output [3:0] io_pixelVal_out_2_6,
  output [3:0] io_pixelVal_out_2_7,
  output       io_valid_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  KernelConvolution_clock; // @[Filter.scala 142:36]
  wire  KernelConvolution_reset; // @[Filter.scala 142:36]
  wire [4:0] KernelConvolution_io_kernelVal_in; // @[Filter.scala 142:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_0; // @[Filter.scala 142:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_1; // @[Filter.scala 142:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_2; // @[Filter.scala 142:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_3; // @[Filter.scala 142:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_4; // @[Filter.scala 142:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_5; // @[Filter.scala 142:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_6; // @[Filter.scala 142:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_7; // @[Filter.scala 142:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_0; // @[Filter.scala 142:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_1; // @[Filter.scala 142:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_2; // @[Filter.scala 142:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_3; // @[Filter.scala 142:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_4; // @[Filter.scala 142:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_5; // @[Filter.scala 142:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_6; // @[Filter.scala 142:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_7; // @[Filter.scala 142:36]
  wire  KernelConvolution_io_valid_out; // @[Filter.scala 142:36]
  wire  KernelConvolution_1_clock; // @[Filter.scala 143:36]
  wire  KernelConvolution_1_reset; // @[Filter.scala 143:36]
  wire [4:0] KernelConvolution_1_io_kernelVal_in; // @[Filter.scala 143:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_0; // @[Filter.scala 143:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_1; // @[Filter.scala 143:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_2; // @[Filter.scala 143:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_3; // @[Filter.scala 143:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_4; // @[Filter.scala 143:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_5; // @[Filter.scala 143:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_6; // @[Filter.scala 143:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_7; // @[Filter.scala 143:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_0; // @[Filter.scala 143:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_1; // @[Filter.scala 143:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_2; // @[Filter.scala 143:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_3; // @[Filter.scala 143:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_4; // @[Filter.scala 143:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_5; // @[Filter.scala 143:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_6; // @[Filter.scala 143:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_7; // @[Filter.scala 143:36]
  wire  KernelConvolution_1_io_valid_out; // @[Filter.scala 143:36]
  wire  KernelConvolution_2_clock; // @[Filter.scala 144:36]
  wire  KernelConvolution_2_reset; // @[Filter.scala 144:36]
  wire [4:0] KernelConvolution_2_io_kernelVal_in; // @[Filter.scala 144:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_0; // @[Filter.scala 144:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_1; // @[Filter.scala 144:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_2; // @[Filter.scala 144:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_3; // @[Filter.scala 144:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_4; // @[Filter.scala 144:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_5; // @[Filter.scala 144:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_6; // @[Filter.scala 144:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_7; // @[Filter.scala 144:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_0; // @[Filter.scala 144:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_1; // @[Filter.scala 144:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_2; // @[Filter.scala 144:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_3; // @[Filter.scala 144:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_4; // @[Filter.scala 144:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_5; // @[Filter.scala 144:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_6; // @[Filter.scala 144:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_7; // @[Filter.scala 144:36]
  wire  KernelConvolution_2_io_valid_out; // @[Filter.scala 144:36]
  reg [3:0] kernelCounter; // @[Counter.scala 29:33]
  wire  kernelCountReset = kernelCounter == 4'h8; // @[Counter.scala 38:24]
  wire [3:0] _T_14 = kernelCounter + 4'h1; // @[Counter.scala 39:22]
  wire  _GEN_9563 = 3'h0 == io_SPI_filterIndex[2:0]; // @[Filter.scala 150:41]
  wire  _GEN_9564 = 4'h4 == kernelCounter; // @[Filter.scala 150:41]
  wire [4:0] _GEN_7 = _GEN_9563 & _GEN_9564 ? $signed(5'sh1) : $signed(5'sh0); // @[Filter.scala 150:41]
  wire  _GEN_9566 = 4'h5 == kernelCounter; // @[Filter.scala 150:41]
  wire [4:0] _GEN_8 = _GEN_9563 & _GEN_9566 ? $signed(5'sh0) : $signed(_GEN_7); // @[Filter.scala 150:41]
  wire  _GEN_9568 = 4'h6 == kernelCounter; // @[Filter.scala 150:41]
  wire [4:0] _GEN_9 = _GEN_9563 & _GEN_9568 ? $signed(5'sh0) : $signed(_GEN_8); // @[Filter.scala 150:41]
  wire  _GEN_9570 = 4'h7 == kernelCounter; // @[Filter.scala 150:41]
  wire [4:0] _GEN_10 = _GEN_9563 & _GEN_9570 ? $signed(5'sh0) : $signed(_GEN_9); // @[Filter.scala 150:41]
  wire  _GEN_9572 = 4'h8 == kernelCounter; // @[Filter.scala 150:41]
  wire [4:0] _GEN_11 = _GEN_9563 & _GEN_9572 ? $signed(5'sh0) : $signed(_GEN_10); // @[Filter.scala 150:41]
  wire  _GEN_9573 = 3'h1 == io_SPI_filterIndex[2:0]; // @[Filter.scala 150:41]
  wire  _GEN_9574 = 4'h0 == kernelCounter; // @[Filter.scala 150:41]
  wire [4:0] _GEN_12 = _GEN_9573 & _GEN_9574 ? $signed(5'sh1) : $signed(_GEN_11); // @[Filter.scala 150:41]
  wire  _GEN_9576 = 4'h1 == kernelCounter; // @[Filter.scala 150:41]
  wire [4:0] _GEN_13 = _GEN_9573 & _GEN_9576 ? $signed(5'sh1) : $signed(_GEN_12); // @[Filter.scala 150:41]
  wire  _GEN_9578 = 4'h2 == kernelCounter; // @[Filter.scala 150:41]
  wire [4:0] _GEN_14 = _GEN_9573 & _GEN_9578 ? $signed(5'sh1) : $signed(_GEN_13); // @[Filter.scala 150:41]
  wire  _GEN_9580 = 4'h3 == kernelCounter; // @[Filter.scala 150:41]
  wire [4:0] _GEN_15 = _GEN_9573 & _GEN_9580 ? $signed(5'sh1) : $signed(_GEN_14); // @[Filter.scala 150:41]
  wire [4:0] _GEN_16 = _GEN_9573 & _GEN_9564 ? $signed(5'sh1) : $signed(_GEN_15); // @[Filter.scala 150:41]
  wire [4:0] _GEN_17 = _GEN_9573 & _GEN_9566 ? $signed(5'sh1) : $signed(_GEN_16); // @[Filter.scala 150:41]
  wire [4:0] _GEN_18 = _GEN_9573 & _GEN_9568 ? $signed(5'sh1) : $signed(_GEN_17); // @[Filter.scala 150:41]
  wire [4:0] _GEN_19 = _GEN_9573 & _GEN_9570 ? $signed(5'sh1) : $signed(_GEN_18); // @[Filter.scala 150:41]
  wire [4:0] _GEN_20 = _GEN_9573 & _GEN_9572 ? $signed(5'sh1) : $signed(_GEN_19); // @[Filter.scala 150:41]
  wire  _GEN_9591 = 3'h2 == io_SPI_filterIndex[2:0]; // @[Filter.scala 150:41]
  wire [4:0] _GEN_21 = _GEN_9591 & _GEN_9574 ? $signed(5'sh1) : $signed(_GEN_20); // @[Filter.scala 150:41]
  wire [4:0] _GEN_22 = _GEN_9591 & _GEN_9576 ? $signed(5'sh2) : $signed(_GEN_21); // @[Filter.scala 150:41]
  wire [4:0] _GEN_23 = _GEN_9591 & _GEN_9578 ? $signed(5'sh1) : $signed(_GEN_22); // @[Filter.scala 150:41]
  wire [4:0] _GEN_24 = _GEN_9591 & _GEN_9580 ? $signed(5'sh2) : $signed(_GEN_23); // @[Filter.scala 150:41]
  wire [4:0] _GEN_25 = _GEN_9591 & _GEN_9564 ? $signed(5'sh4) : $signed(_GEN_24); // @[Filter.scala 150:41]
  wire [4:0] _GEN_26 = _GEN_9591 & _GEN_9566 ? $signed(5'sh2) : $signed(_GEN_25); // @[Filter.scala 150:41]
  wire [4:0] _GEN_27 = _GEN_9591 & _GEN_9568 ? $signed(5'sh1) : $signed(_GEN_26); // @[Filter.scala 150:41]
  wire [4:0] _GEN_28 = _GEN_9591 & _GEN_9570 ? $signed(5'sh2) : $signed(_GEN_27); // @[Filter.scala 150:41]
  wire [4:0] _GEN_29 = _GEN_9591 & _GEN_9572 ? $signed(5'sh1) : $signed(_GEN_28); // @[Filter.scala 150:41]
  wire  _GEN_9609 = 3'h3 == io_SPI_filterIndex[2:0]; // @[Filter.scala 150:41]
  wire [4:0] _GEN_30 = _GEN_9609 & _GEN_9574 ? $signed(5'sh0) : $signed(_GEN_29); // @[Filter.scala 150:41]
  wire [4:0] _GEN_31 = _GEN_9609 & _GEN_9576 ? $signed(-5'sh1) : $signed(_GEN_30); // @[Filter.scala 150:41]
  wire [4:0] _GEN_32 = _GEN_9609 & _GEN_9578 ? $signed(5'sh0) : $signed(_GEN_31); // @[Filter.scala 150:41]
  wire [4:0] _GEN_33 = _GEN_9609 & _GEN_9580 ? $signed(-5'sh1) : $signed(_GEN_32); // @[Filter.scala 150:41]
  wire [4:0] _GEN_34 = _GEN_9609 & _GEN_9564 ? $signed(5'sh4) : $signed(_GEN_33); // @[Filter.scala 150:41]
  wire [4:0] _GEN_35 = _GEN_9609 & _GEN_9566 ? $signed(-5'sh1) : $signed(_GEN_34); // @[Filter.scala 150:41]
  wire [4:0] _GEN_36 = _GEN_9609 & _GEN_9568 ? $signed(5'sh0) : $signed(_GEN_35); // @[Filter.scala 150:41]
  wire [4:0] _GEN_37 = _GEN_9609 & _GEN_9570 ? $signed(-5'sh1) : $signed(_GEN_36); // @[Filter.scala 150:41]
  wire [4:0] _GEN_38 = _GEN_9609 & _GEN_9572 ? $signed(5'sh0) : $signed(_GEN_37); // @[Filter.scala 150:41]
  wire  _GEN_9627 = 3'h4 == io_SPI_filterIndex[2:0]; // @[Filter.scala 150:41]
  wire [4:0] _GEN_39 = _GEN_9627 & _GEN_9574 ? $signed(-5'sh1) : $signed(_GEN_38); // @[Filter.scala 150:41]
  wire [4:0] _GEN_40 = _GEN_9627 & _GEN_9576 ? $signed(-5'sh1) : $signed(_GEN_39); // @[Filter.scala 150:41]
  wire [4:0] _GEN_41 = _GEN_9627 & _GEN_9578 ? $signed(-5'sh1) : $signed(_GEN_40); // @[Filter.scala 150:41]
  wire [4:0] _GEN_42 = _GEN_9627 & _GEN_9580 ? $signed(-5'sh1) : $signed(_GEN_41); // @[Filter.scala 150:41]
  wire [4:0] _GEN_43 = _GEN_9627 & _GEN_9564 ? $signed(5'sh8) : $signed(_GEN_42); // @[Filter.scala 150:41]
  wire [4:0] _GEN_44 = _GEN_9627 & _GEN_9566 ? $signed(-5'sh1) : $signed(_GEN_43); // @[Filter.scala 150:41]
  wire [4:0] _GEN_45 = _GEN_9627 & _GEN_9568 ? $signed(-5'sh1) : $signed(_GEN_44); // @[Filter.scala 150:41]
  wire [4:0] _GEN_46 = _GEN_9627 & _GEN_9570 ? $signed(-5'sh1) : $signed(_GEN_45); // @[Filter.scala 150:41]
  wire [4:0] _GEN_47 = _GEN_9627 & _GEN_9572 ? $signed(-5'sh1) : $signed(_GEN_46); // @[Filter.scala 150:41]
  wire  _GEN_9645 = 3'h5 == io_SPI_filterIndex[2:0]; // @[Filter.scala 150:41]
  wire [4:0] _GEN_48 = _GEN_9645 & _GEN_9574 ? $signed(5'sh0) : $signed(_GEN_47); // @[Filter.scala 150:41]
  wire [4:0] _GEN_49 = _GEN_9645 & _GEN_9576 ? $signed(-5'sh1) : $signed(_GEN_48); // @[Filter.scala 150:41]
  wire [4:0] _GEN_50 = _GEN_9645 & _GEN_9578 ? $signed(5'sh0) : $signed(_GEN_49); // @[Filter.scala 150:41]
  wire [4:0] _GEN_51 = _GEN_9645 & _GEN_9580 ? $signed(-5'sh1) : $signed(_GEN_50); // @[Filter.scala 150:41]
  wire [4:0] _GEN_52 = _GEN_9645 & _GEN_9564 ? $signed(5'sh5) : $signed(_GEN_51); // @[Filter.scala 150:41]
  wire [4:0] _GEN_53 = _GEN_9645 & _GEN_9566 ? $signed(-5'sh1) : $signed(_GEN_52); // @[Filter.scala 150:41]
  wire [4:0] _GEN_54 = _GEN_9645 & _GEN_9568 ? $signed(5'sh0) : $signed(_GEN_53); // @[Filter.scala 150:41]
  wire [4:0] _GEN_55 = _GEN_9645 & _GEN_9570 ? $signed(-5'sh1) : $signed(_GEN_54); // @[Filter.scala 150:41]
  reg [1:0] imageCounterX; // @[Counter.scala 29:33]
  wire  imageCounterXReset = imageCounterX == 2'h2; // @[Counter.scala 38:24]
  wire [1:0] _T_20 = imageCounterX + 2'h1; // @[Counter.scala 39:22]
  reg [1:0] imageCounterY; // @[Counter.scala 29:33]
  wire  _T_21 = imageCounterY == 2'h2; // @[Counter.scala 38:24]
  wire [1:0] _T_23 = imageCounterY + 2'h1; // @[Counter.scala 39:22]
  reg [31:0] pixelIndex; // @[Filter.scala 155:31]
  wire [32:0] _T_24 = {{1'd0}, pixelIndex}; // @[Filter.scala 158:31]
  wire [31:0] _GEN_0 = _T_24[31:0] % 32'h10; // @[Filter.scala 158:38]
  wire [4:0] _T_26 = _GEN_0[4:0]; // @[Filter.scala 158:38]
  wire [4:0] _GEN_9863 = {{3'd0}, imageCounterX}; // @[Filter.scala 158:53]
  wire [4:0] _T_28 = _T_26 + _GEN_9863; // @[Filter.scala 158:53]
  wire [4:0] _T_30 = _T_28 - 5'h1; // @[Filter.scala 158:69]
  wire [31:0] _T_33 = _T_24[31:0] / 32'h10; // @[Filter.scala 159:38]
  wire [31:0] _GEN_9864 = {{30'd0}, imageCounterY}; // @[Filter.scala 159:53]
  wire [31:0] _T_35 = _T_33 + _GEN_9864; // @[Filter.scala 159:53]
  wire [31:0] _T_37 = _T_35 - 32'h1; // @[Filter.scala 159:69]
  wire [36:0] _T_38 = _T_37 * 32'h10; // @[Filter.scala 160:42]
  wire [36:0] _GEN_9865 = {{32'd0}, _T_30}; // @[Filter.scala 160:57]
  wire [36:0] _T_40 = _T_38 + _GEN_9865; // @[Filter.scala 160:57]
  wire [3:0] _GEN_179 = 8'h8 == _T_40[7:0] ? 4'h0 : 4'hf; // @[Filter.scala 160:62]
  wire [3:0] _GEN_180 = 8'h9 == _T_40[7:0] ? 4'h0 : _GEN_179; // @[Filter.scala 160:62]
  wire [3:0] _GEN_181 = 8'ha == _T_40[7:0] ? 4'h0 : _GEN_180; // @[Filter.scala 160:62]
  wire [3:0] _GEN_182 = 8'hb == _T_40[7:0] ? 4'h0 : _GEN_181; // @[Filter.scala 160:62]
  wire [3:0] _GEN_183 = 8'hc == _T_40[7:0] ? 4'h0 : _GEN_182; // @[Filter.scala 160:62]
  wire [3:0] _GEN_184 = 8'hd == _T_40[7:0] ? 4'h0 : _GEN_183; // @[Filter.scala 160:62]
  wire [3:0] _GEN_185 = 8'he == _T_40[7:0] ? 4'h0 : _GEN_184; // @[Filter.scala 160:62]
  wire [3:0] _GEN_186 = 8'hf == _T_40[7:0] ? 4'h0 : _GEN_185; // @[Filter.scala 160:62]
  wire [3:0] _GEN_187 = 8'h10 == _T_40[7:0] ? 4'hf : _GEN_186; // @[Filter.scala 160:62]
  wire [3:0] _GEN_188 = 8'h11 == _T_40[7:0] ? 4'hf : _GEN_187; // @[Filter.scala 160:62]
  wire [3:0] _GEN_189 = 8'h12 == _T_40[7:0] ? 4'hf : _GEN_188; // @[Filter.scala 160:62]
  wire [3:0] _GEN_190 = 8'h13 == _T_40[7:0] ? 4'hf : _GEN_189; // @[Filter.scala 160:62]
  wire [3:0] _GEN_191 = 8'h14 == _T_40[7:0] ? 4'hf : _GEN_190; // @[Filter.scala 160:62]
  wire [3:0] _GEN_192 = 8'h15 == _T_40[7:0] ? 4'hf : _GEN_191; // @[Filter.scala 160:62]
  wire [3:0] _GEN_193 = 8'h16 == _T_40[7:0] ? 4'hf : _GEN_192; // @[Filter.scala 160:62]
  wire [3:0] _GEN_194 = 8'h17 == _T_40[7:0] ? 4'hf : _GEN_193; // @[Filter.scala 160:62]
  wire [3:0] _GEN_195 = 8'h18 == _T_40[7:0] ? 4'h0 : _GEN_194; // @[Filter.scala 160:62]
  wire [3:0] _GEN_196 = 8'h19 == _T_40[7:0] ? 4'h0 : _GEN_195; // @[Filter.scala 160:62]
  wire [3:0] _GEN_197 = 8'h1a == _T_40[7:0] ? 4'h0 : _GEN_196; // @[Filter.scala 160:62]
  wire [3:0] _GEN_198 = 8'h1b == _T_40[7:0] ? 4'h0 : _GEN_197; // @[Filter.scala 160:62]
  wire [3:0] _GEN_199 = 8'h1c == _T_40[7:0] ? 4'h0 : _GEN_198; // @[Filter.scala 160:62]
  wire [3:0] _GEN_200 = 8'h1d == _T_40[7:0] ? 4'h0 : _GEN_199; // @[Filter.scala 160:62]
  wire [3:0] _GEN_201 = 8'h1e == _T_40[7:0] ? 4'h0 : _GEN_200; // @[Filter.scala 160:62]
  wire [3:0] _GEN_202 = 8'h1f == _T_40[7:0] ? 4'h0 : _GEN_201; // @[Filter.scala 160:62]
  wire [3:0] _GEN_203 = 8'h20 == _T_40[7:0] ? 4'hf : _GEN_202; // @[Filter.scala 160:62]
  wire [3:0] _GEN_204 = 8'h21 == _T_40[7:0] ? 4'hf : _GEN_203; // @[Filter.scala 160:62]
  wire [3:0] _GEN_205 = 8'h22 == _T_40[7:0] ? 4'hf : _GEN_204; // @[Filter.scala 160:62]
  wire [3:0] _GEN_206 = 8'h23 == _T_40[7:0] ? 4'hf : _GEN_205; // @[Filter.scala 160:62]
  wire [3:0] _GEN_207 = 8'h24 == _T_40[7:0] ? 4'hf : _GEN_206; // @[Filter.scala 160:62]
  wire [3:0] _GEN_208 = 8'h25 == _T_40[7:0] ? 4'hf : _GEN_207; // @[Filter.scala 160:62]
  wire [3:0] _GEN_209 = 8'h26 == _T_40[7:0] ? 4'hf : _GEN_208; // @[Filter.scala 160:62]
  wire [3:0] _GEN_210 = 8'h27 == _T_40[7:0] ? 4'hf : _GEN_209; // @[Filter.scala 160:62]
  wire [3:0] _GEN_211 = 8'h28 == _T_40[7:0] ? 4'h0 : _GEN_210; // @[Filter.scala 160:62]
  wire [3:0] _GEN_212 = 8'h29 == _T_40[7:0] ? 4'h0 : _GEN_211; // @[Filter.scala 160:62]
  wire [3:0] _GEN_213 = 8'h2a == _T_40[7:0] ? 4'h0 : _GEN_212; // @[Filter.scala 160:62]
  wire [3:0] _GEN_214 = 8'h2b == _T_40[7:0] ? 4'h0 : _GEN_213; // @[Filter.scala 160:62]
  wire [3:0] _GEN_215 = 8'h2c == _T_40[7:0] ? 4'h0 : _GEN_214; // @[Filter.scala 160:62]
  wire [3:0] _GEN_216 = 8'h2d == _T_40[7:0] ? 4'h0 : _GEN_215; // @[Filter.scala 160:62]
  wire [3:0] _GEN_217 = 8'h2e == _T_40[7:0] ? 4'h0 : _GEN_216; // @[Filter.scala 160:62]
  wire [3:0] _GEN_218 = 8'h2f == _T_40[7:0] ? 4'h0 : _GEN_217; // @[Filter.scala 160:62]
  wire [3:0] _GEN_219 = 8'h30 == _T_40[7:0] ? 4'hf : _GEN_218; // @[Filter.scala 160:62]
  wire [3:0] _GEN_220 = 8'h31 == _T_40[7:0] ? 4'hf : _GEN_219; // @[Filter.scala 160:62]
  wire [3:0] _GEN_221 = 8'h32 == _T_40[7:0] ? 4'hf : _GEN_220; // @[Filter.scala 160:62]
  wire [3:0] _GEN_222 = 8'h33 == _T_40[7:0] ? 4'hf : _GEN_221; // @[Filter.scala 160:62]
  wire [3:0] _GEN_223 = 8'h34 == _T_40[7:0] ? 4'hf : _GEN_222; // @[Filter.scala 160:62]
  wire [3:0] _GEN_224 = 8'h35 == _T_40[7:0] ? 4'hf : _GEN_223; // @[Filter.scala 160:62]
  wire [3:0] _GEN_225 = 8'h36 == _T_40[7:0] ? 4'hf : _GEN_224; // @[Filter.scala 160:62]
  wire [3:0] _GEN_226 = 8'h37 == _T_40[7:0] ? 4'hf : _GEN_225; // @[Filter.scala 160:62]
  wire [3:0] _GEN_227 = 8'h38 == _T_40[7:0] ? 4'h0 : _GEN_226; // @[Filter.scala 160:62]
  wire [3:0] _GEN_228 = 8'h39 == _T_40[7:0] ? 4'h0 : _GEN_227; // @[Filter.scala 160:62]
  wire [3:0] _GEN_229 = 8'h3a == _T_40[7:0] ? 4'h0 : _GEN_228; // @[Filter.scala 160:62]
  wire [3:0] _GEN_230 = 8'h3b == _T_40[7:0] ? 4'h0 : _GEN_229; // @[Filter.scala 160:62]
  wire [3:0] _GEN_231 = 8'h3c == _T_40[7:0] ? 4'h0 : _GEN_230; // @[Filter.scala 160:62]
  wire [3:0] _GEN_232 = 8'h3d == _T_40[7:0] ? 4'h0 : _GEN_231; // @[Filter.scala 160:62]
  wire [3:0] _GEN_233 = 8'h3e == _T_40[7:0] ? 4'h0 : _GEN_232; // @[Filter.scala 160:62]
  wire [3:0] _GEN_234 = 8'h3f == _T_40[7:0] ? 4'h0 : _GEN_233; // @[Filter.scala 160:62]
  wire [3:0] _GEN_235 = 8'h40 == _T_40[7:0] ? 4'hf : _GEN_234; // @[Filter.scala 160:62]
  wire [3:0] _GEN_236 = 8'h41 == _T_40[7:0] ? 4'hf : _GEN_235; // @[Filter.scala 160:62]
  wire [3:0] _GEN_237 = 8'h42 == _T_40[7:0] ? 4'hf : _GEN_236; // @[Filter.scala 160:62]
  wire [3:0] _GEN_238 = 8'h43 == _T_40[7:0] ? 4'hf : _GEN_237; // @[Filter.scala 160:62]
  wire [3:0] _GEN_239 = 8'h44 == _T_40[7:0] ? 4'hf : _GEN_238; // @[Filter.scala 160:62]
  wire [3:0] _GEN_240 = 8'h45 == _T_40[7:0] ? 4'hf : _GEN_239; // @[Filter.scala 160:62]
  wire [3:0] _GEN_241 = 8'h46 == _T_40[7:0] ? 4'hf : _GEN_240; // @[Filter.scala 160:62]
  wire [3:0] _GEN_242 = 8'h47 == _T_40[7:0] ? 4'hf : _GEN_241; // @[Filter.scala 160:62]
  wire [3:0] _GEN_243 = 8'h48 == _T_40[7:0] ? 4'h0 : _GEN_242; // @[Filter.scala 160:62]
  wire [3:0] _GEN_244 = 8'h49 == _T_40[7:0] ? 4'h0 : _GEN_243; // @[Filter.scala 160:62]
  wire [3:0] _GEN_245 = 8'h4a == _T_40[7:0] ? 4'h0 : _GEN_244; // @[Filter.scala 160:62]
  wire [3:0] _GEN_246 = 8'h4b == _T_40[7:0] ? 4'h0 : _GEN_245; // @[Filter.scala 160:62]
  wire [3:0] _GEN_247 = 8'h4c == _T_40[7:0] ? 4'h0 : _GEN_246; // @[Filter.scala 160:62]
  wire [3:0] _GEN_248 = 8'h4d == _T_40[7:0] ? 4'h0 : _GEN_247; // @[Filter.scala 160:62]
  wire [3:0] _GEN_249 = 8'h4e == _T_40[7:0] ? 4'h0 : _GEN_248; // @[Filter.scala 160:62]
  wire [3:0] _GEN_250 = 8'h4f == _T_40[7:0] ? 4'h0 : _GEN_249; // @[Filter.scala 160:62]
  wire [3:0] _GEN_251 = 8'h50 == _T_40[7:0] ? 4'hf : _GEN_250; // @[Filter.scala 160:62]
  wire [3:0] _GEN_252 = 8'h51 == _T_40[7:0] ? 4'hf : _GEN_251; // @[Filter.scala 160:62]
  wire [3:0] _GEN_253 = 8'h52 == _T_40[7:0] ? 4'hf : _GEN_252; // @[Filter.scala 160:62]
  wire [3:0] _GEN_254 = 8'h53 == _T_40[7:0] ? 4'hf : _GEN_253; // @[Filter.scala 160:62]
  wire [3:0] _GEN_255 = 8'h54 == _T_40[7:0] ? 4'hf : _GEN_254; // @[Filter.scala 160:62]
  wire [3:0] _GEN_256 = 8'h55 == _T_40[7:0] ? 4'hf : _GEN_255; // @[Filter.scala 160:62]
  wire [3:0] _GEN_257 = 8'h56 == _T_40[7:0] ? 4'hf : _GEN_256; // @[Filter.scala 160:62]
  wire [3:0] _GEN_258 = 8'h57 == _T_40[7:0] ? 4'hf : _GEN_257; // @[Filter.scala 160:62]
  wire [3:0] _GEN_259 = 8'h58 == _T_40[7:0] ? 4'h0 : _GEN_258; // @[Filter.scala 160:62]
  wire [3:0] _GEN_260 = 8'h59 == _T_40[7:0] ? 4'h0 : _GEN_259; // @[Filter.scala 160:62]
  wire [3:0] _GEN_261 = 8'h5a == _T_40[7:0] ? 4'h0 : _GEN_260; // @[Filter.scala 160:62]
  wire [3:0] _GEN_262 = 8'h5b == _T_40[7:0] ? 4'h0 : _GEN_261; // @[Filter.scala 160:62]
  wire [3:0] _GEN_263 = 8'h5c == _T_40[7:0] ? 4'h0 : _GEN_262; // @[Filter.scala 160:62]
  wire [3:0] _GEN_264 = 8'h5d == _T_40[7:0] ? 4'h0 : _GEN_263; // @[Filter.scala 160:62]
  wire [3:0] _GEN_265 = 8'h5e == _T_40[7:0] ? 4'h0 : _GEN_264; // @[Filter.scala 160:62]
  wire [3:0] _GEN_266 = 8'h5f == _T_40[7:0] ? 4'h0 : _GEN_265; // @[Filter.scala 160:62]
  wire [3:0] _GEN_267 = 8'h60 == _T_40[7:0] ? 4'h0 : _GEN_266; // @[Filter.scala 160:62]
  wire [3:0] _GEN_268 = 8'h61 == _T_40[7:0] ? 4'h0 : _GEN_267; // @[Filter.scala 160:62]
  wire [3:0] _GEN_269 = 8'h62 == _T_40[7:0] ? 4'h0 : _GEN_268; // @[Filter.scala 160:62]
  wire [3:0] _GEN_270 = 8'h63 == _T_40[7:0] ? 4'h0 : _GEN_269; // @[Filter.scala 160:62]
  wire [3:0] _GEN_271 = 8'h64 == _T_40[7:0] ? 4'h0 : _GEN_270; // @[Filter.scala 160:62]
  wire [3:0] _GEN_272 = 8'h65 == _T_40[7:0] ? 4'h0 : _GEN_271; // @[Filter.scala 160:62]
  wire [3:0] _GEN_273 = 8'h66 == _T_40[7:0] ? 4'h0 : _GEN_272; // @[Filter.scala 160:62]
  wire [3:0] _GEN_274 = 8'h67 == _T_40[7:0] ? 4'h0 : _GEN_273; // @[Filter.scala 160:62]
  wire [3:0] _GEN_275 = 8'h68 == _T_40[7:0] ? 4'hf : _GEN_274; // @[Filter.scala 160:62]
  wire [3:0] _GEN_276 = 8'h69 == _T_40[7:0] ? 4'hf : _GEN_275; // @[Filter.scala 160:62]
  wire [3:0] _GEN_277 = 8'h6a == _T_40[7:0] ? 4'hf : _GEN_276; // @[Filter.scala 160:62]
  wire [3:0] _GEN_278 = 8'h6b == _T_40[7:0] ? 4'hf : _GEN_277; // @[Filter.scala 160:62]
  wire [3:0] _GEN_279 = 8'h6c == _T_40[7:0] ? 4'hf : _GEN_278; // @[Filter.scala 160:62]
  wire [3:0] _GEN_280 = 8'h6d == _T_40[7:0] ? 4'hf : _GEN_279; // @[Filter.scala 160:62]
  wire [3:0] _GEN_281 = 8'h6e == _T_40[7:0] ? 4'hf : _GEN_280; // @[Filter.scala 160:62]
  wire [3:0] _GEN_282 = 8'h6f == _T_40[7:0] ? 4'hf : _GEN_281; // @[Filter.scala 160:62]
  wire [3:0] _GEN_283 = 8'h70 == _T_40[7:0] ? 4'h0 : _GEN_282; // @[Filter.scala 160:62]
  wire [3:0] _GEN_284 = 8'h71 == _T_40[7:0] ? 4'h0 : _GEN_283; // @[Filter.scala 160:62]
  wire [3:0] _GEN_285 = 8'h72 == _T_40[7:0] ? 4'h0 : _GEN_284; // @[Filter.scala 160:62]
  wire [3:0] _GEN_286 = 8'h73 == _T_40[7:0] ? 4'h0 : _GEN_285; // @[Filter.scala 160:62]
  wire [3:0] _GEN_287 = 8'h74 == _T_40[7:0] ? 4'h0 : _GEN_286; // @[Filter.scala 160:62]
  wire [3:0] _GEN_288 = 8'h75 == _T_40[7:0] ? 4'h0 : _GEN_287; // @[Filter.scala 160:62]
  wire [3:0] _GEN_289 = 8'h76 == _T_40[7:0] ? 4'h0 : _GEN_288; // @[Filter.scala 160:62]
  wire [3:0] _GEN_290 = 8'h77 == _T_40[7:0] ? 4'h0 : _GEN_289; // @[Filter.scala 160:62]
  wire [3:0] _GEN_291 = 8'h78 == _T_40[7:0] ? 4'hf : _GEN_290; // @[Filter.scala 160:62]
  wire [3:0] _GEN_292 = 8'h79 == _T_40[7:0] ? 4'hf : _GEN_291; // @[Filter.scala 160:62]
  wire [3:0] _GEN_293 = 8'h7a == _T_40[7:0] ? 4'hf : _GEN_292; // @[Filter.scala 160:62]
  wire [3:0] _GEN_294 = 8'h7b == _T_40[7:0] ? 4'hf : _GEN_293; // @[Filter.scala 160:62]
  wire [3:0] _GEN_295 = 8'h7c == _T_40[7:0] ? 4'hf : _GEN_294; // @[Filter.scala 160:62]
  wire [3:0] _GEN_296 = 8'h7d == _T_40[7:0] ? 4'hf : _GEN_295; // @[Filter.scala 160:62]
  wire [3:0] _GEN_297 = 8'h7e == _T_40[7:0] ? 4'hf : _GEN_296; // @[Filter.scala 160:62]
  wire [3:0] _GEN_298 = 8'h7f == _T_40[7:0] ? 4'hf : _GEN_297; // @[Filter.scala 160:62]
  wire [3:0] _GEN_299 = 8'h80 == _T_40[7:0] ? 4'h0 : _GEN_298; // @[Filter.scala 160:62]
  wire [3:0] _GEN_300 = 8'h81 == _T_40[7:0] ? 4'h0 : _GEN_299; // @[Filter.scala 160:62]
  wire [3:0] _GEN_301 = 8'h82 == _T_40[7:0] ? 4'h0 : _GEN_300; // @[Filter.scala 160:62]
  wire [3:0] _GEN_302 = 8'h83 == _T_40[7:0] ? 4'h0 : _GEN_301; // @[Filter.scala 160:62]
  wire [3:0] _GEN_303 = 8'h84 == _T_40[7:0] ? 4'h0 : _GEN_302; // @[Filter.scala 160:62]
  wire [3:0] _GEN_304 = 8'h85 == _T_40[7:0] ? 4'h0 : _GEN_303; // @[Filter.scala 160:62]
  wire [3:0] _GEN_305 = 8'h86 == _T_40[7:0] ? 4'h0 : _GEN_304; // @[Filter.scala 160:62]
  wire [3:0] _GEN_306 = 8'h87 == _T_40[7:0] ? 4'h0 : _GEN_305; // @[Filter.scala 160:62]
  wire [3:0] _GEN_307 = 8'h88 == _T_40[7:0] ? 4'hf : _GEN_306; // @[Filter.scala 160:62]
  wire [3:0] _GEN_308 = 8'h89 == _T_40[7:0] ? 4'hf : _GEN_307; // @[Filter.scala 160:62]
  wire [3:0] _GEN_309 = 8'h8a == _T_40[7:0] ? 4'hf : _GEN_308; // @[Filter.scala 160:62]
  wire [3:0] _GEN_310 = 8'h8b == _T_40[7:0] ? 4'hf : _GEN_309; // @[Filter.scala 160:62]
  wire [3:0] _GEN_311 = 8'h8c == _T_40[7:0] ? 4'hf : _GEN_310; // @[Filter.scala 160:62]
  wire [3:0] _GEN_312 = 8'h8d == _T_40[7:0] ? 4'hf : _GEN_311; // @[Filter.scala 160:62]
  wire [3:0] _GEN_313 = 8'h8e == _T_40[7:0] ? 4'hf : _GEN_312; // @[Filter.scala 160:62]
  wire [3:0] _GEN_314 = 8'h8f == _T_40[7:0] ? 4'hf : _GEN_313; // @[Filter.scala 160:62]
  wire [3:0] _GEN_315 = 8'h90 == _T_40[7:0] ? 4'h0 : _GEN_314; // @[Filter.scala 160:62]
  wire [3:0] _GEN_316 = 8'h91 == _T_40[7:0] ? 4'h0 : _GEN_315; // @[Filter.scala 160:62]
  wire [3:0] _GEN_317 = 8'h92 == _T_40[7:0] ? 4'h0 : _GEN_316; // @[Filter.scala 160:62]
  wire [3:0] _GEN_318 = 8'h93 == _T_40[7:0] ? 4'h0 : _GEN_317; // @[Filter.scala 160:62]
  wire [3:0] _GEN_319 = 8'h94 == _T_40[7:0] ? 4'h0 : _GEN_318; // @[Filter.scala 160:62]
  wire [3:0] _GEN_320 = 8'h95 == _T_40[7:0] ? 4'h0 : _GEN_319; // @[Filter.scala 160:62]
  wire [3:0] _GEN_321 = 8'h96 == _T_40[7:0] ? 4'h0 : _GEN_320; // @[Filter.scala 160:62]
  wire [3:0] _GEN_322 = 8'h97 == _T_40[7:0] ? 4'h0 : _GEN_321; // @[Filter.scala 160:62]
  wire [3:0] _GEN_323 = 8'h98 == _T_40[7:0] ? 4'hf : _GEN_322; // @[Filter.scala 160:62]
  wire [3:0] _GEN_324 = 8'h99 == _T_40[7:0] ? 4'hf : _GEN_323; // @[Filter.scala 160:62]
  wire [3:0] _GEN_325 = 8'h9a == _T_40[7:0] ? 4'hf : _GEN_324; // @[Filter.scala 160:62]
  wire [3:0] _GEN_326 = 8'h9b == _T_40[7:0] ? 4'hf : _GEN_325; // @[Filter.scala 160:62]
  wire [3:0] _GEN_327 = 8'h9c == _T_40[7:0] ? 4'hf : _GEN_326; // @[Filter.scala 160:62]
  wire [3:0] _GEN_328 = 8'h9d == _T_40[7:0] ? 4'hf : _GEN_327; // @[Filter.scala 160:62]
  wire [3:0] _GEN_329 = 8'h9e == _T_40[7:0] ? 4'hf : _GEN_328; // @[Filter.scala 160:62]
  wire [3:0] _GEN_330 = 8'h9f == _T_40[7:0] ? 4'hf : _GEN_329; // @[Filter.scala 160:62]
  wire [3:0] _GEN_331 = 8'ha0 == _T_40[7:0] ? 4'h0 : _GEN_330; // @[Filter.scala 160:62]
  wire [3:0] _GEN_332 = 8'ha1 == _T_40[7:0] ? 4'h0 : _GEN_331; // @[Filter.scala 160:62]
  wire [3:0] _GEN_333 = 8'ha2 == _T_40[7:0] ? 4'h0 : _GEN_332; // @[Filter.scala 160:62]
  wire [3:0] _GEN_334 = 8'ha3 == _T_40[7:0] ? 4'h0 : _GEN_333; // @[Filter.scala 160:62]
  wire [3:0] _GEN_335 = 8'ha4 == _T_40[7:0] ? 4'h0 : _GEN_334; // @[Filter.scala 160:62]
  wire [3:0] _GEN_336 = 8'ha5 == _T_40[7:0] ? 4'h0 : _GEN_335; // @[Filter.scala 160:62]
  wire [3:0] _GEN_337 = 8'ha6 == _T_40[7:0] ? 4'h0 : _GEN_336; // @[Filter.scala 160:62]
  wire [3:0] _GEN_338 = 8'ha7 == _T_40[7:0] ? 4'h0 : _GEN_337; // @[Filter.scala 160:62]
  wire [3:0] _GEN_339 = 8'ha8 == _T_40[7:0] ? 4'hf : _GEN_338; // @[Filter.scala 160:62]
  wire [3:0] _GEN_340 = 8'ha9 == _T_40[7:0] ? 4'hf : _GEN_339; // @[Filter.scala 160:62]
  wire [3:0] _GEN_341 = 8'haa == _T_40[7:0] ? 4'hf : _GEN_340; // @[Filter.scala 160:62]
  wire [3:0] _GEN_342 = 8'hab == _T_40[7:0] ? 4'hf : _GEN_341; // @[Filter.scala 160:62]
  wire [3:0] _GEN_343 = 8'hac == _T_40[7:0] ? 4'hf : _GEN_342; // @[Filter.scala 160:62]
  wire [3:0] _GEN_344 = 8'had == _T_40[7:0] ? 4'hf : _GEN_343; // @[Filter.scala 160:62]
  wire [3:0] _GEN_345 = 8'hae == _T_40[7:0] ? 4'hf : _GEN_344; // @[Filter.scala 160:62]
  wire [3:0] _GEN_346 = 8'haf == _T_40[7:0] ? 4'hf : _GEN_345; // @[Filter.scala 160:62]
  wire [3:0] _GEN_347 = 8'hb0 == _T_40[7:0] ? 4'h0 : _GEN_346; // @[Filter.scala 160:62]
  wire [3:0] _GEN_348 = 8'hb1 == _T_40[7:0] ? 4'h0 : _GEN_347; // @[Filter.scala 160:62]
  wire [3:0] _GEN_349 = 8'hb2 == _T_40[7:0] ? 4'h0 : _GEN_348; // @[Filter.scala 160:62]
  wire [3:0] _GEN_350 = 8'hb3 == _T_40[7:0] ? 4'h0 : _GEN_349; // @[Filter.scala 160:62]
  wire [3:0] _GEN_351 = 8'hb4 == _T_40[7:0] ? 4'h0 : _GEN_350; // @[Filter.scala 160:62]
  wire [3:0] _GEN_352 = 8'hb5 == _T_40[7:0] ? 4'h0 : _GEN_351; // @[Filter.scala 160:62]
  wire [3:0] _GEN_353 = 8'hb6 == _T_40[7:0] ? 4'h0 : _GEN_352; // @[Filter.scala 160:62]
  wire [3:0] _GEN_354 = 8'hb7 == _T_40[7:0] ? 4'h0 : _GEN_353; // @[Filter.scala 160:62]
  wire [3:0] _GEN_355 = 8'hb8 == _T_40[7:0] ? 4'hf : _GEN_354; // @[Filter.scala 160:62]
  wire [3:0] _GEN_356 = 8'hb9 == _T_40[7:0] ? 4'hf : _GEN_355; // @[Filter.scala 160:62]
  wire [3:0] _GEN_357 = 8'hba == _T_40[7:0] ? 4'hf : _GEN_356; // @[Filter.scala 160:62]
  wire [3:0] _GEN_358 = 8'hbb == _T_40[7:0] ? 4'hf : _GEN_357; // @[Filter.scala 160:62]
  wire [3:0] _GEN_359 = 8'hbc == _T_40[7:0] ? 4'hf : _GEN_358; // @[Filter.scala 160:62]
  wire [3:0] _GEN_360 = 8'hbd == _T_40[7:0] ? 4'hf : _GEN_359; // @[Filter.scala 160:62]
  wire [3:0] _GEN_361 = 8'hbe == _T_40[7:0] ? 4'hf : _GEN_360; // @[Filter.scala 160:62]
  wire [3:0] _GEN_362 = 8'hbf == _T_40[7:0] ? 4'hf : _GEN_361; // @[Filter.scala 160:62]
  wire [4:0] _GEN_9866 = {{1'd0}, _GEN_362}; // @[Filter.scala 160:62]
  wire [8:0] _T_42 = _GEN_9866 * 5'h14; // @[Filter.scala 160:62]
  wire [3:0] _GEN_459 = 8'h60 == _T_40[7:0] ? 4'hf : 4'h0; // @[Filter.scala 160:102]
  wire [3:0] _GEN_460 = 8'h61 == _T_40[7:0] ? 4'hf : _GEN_459; // @[Filter.scala 160:102]
  wire [3:0] _GEN_461 = 8'h62 == _T_40[7:0] ? 4'hf : _GEN_460; // @[Filter.scala 160:102]
  wire [3:0] _GEN_462 = 8'h63 == _T_40[7:0] ? 4'hf : _GEN_461; // @[Filter.scala 160:102]
  wire [3:0] _GEN_463 = 8'h64 == _T_40[7:0] ? 4'hf : _GEN_462; // @[Filter.scala 160:102]
  wire [3:0] _GEN_464 = 8'h65 == _T_40[7:0] ? 4'hf : _GEN_463; // @[Filter.scala 160:102]
  wire [3:0] _GEN_465 = 8'h66 == _T_40[7:0] ? 4'hf : _GEN_464; // @[Filter.scala 160:102]
  wire [3:0] _GEN_466 = 8'h67 == _T_40[7:0] ? 4'hf : _GEN_465; // @[Filter.scala 160:102]
  wire [3:0] _GEN_467 = 8'h68 == _T_40[7:0] ? 4'hf : _GEN_466; // @[Filter.scala 160:102]
  wire [3:0] _GEN_468 = 8'h69 == _T_40[7:0] ? 4'hf : _GEN_467; // @[Filter.scala 160:102]
  wire [3:0] _GEN_469 = 8'h6a == _T_40[7:0] ? 4'hf : _GEN_468; // @[Filter.scala 160:102]
  wire [3:0] _GEN_470 = 8'h6b == _T_40[7:0] ? 4'hf : _GEN_469; // @[Filter.scala 160:102]
  wire [3:0] _GEN_471 = 8'h6c == _T_40[7:0] ? 4'hf : _GEN_470; // @[Filter.scala 160:102]
  wire [3:0] _GEN_472 = 8'h6d == _T_40[7:0] ? 4'hf : _GEN_471; // @[Filter.scala 160:102]
  wire [3:0] _GEN_473 = 8'h6e == _T_40[7:0] ? 4'hf : _GEN_472; // @[Filter.scala 160:102]
  wire [3:0] _GEN_474 = 8'h6f == _T_40[7:0] ? 4'hf : _GEN_473; // @[Filter.scala 160:102]
  wire [3:0] _GEN_475 = 8'h70 == _T_40[7:0] ? 4'hf : _GEN_474; // @[Filter.scala 160:102]
  wire [3:0] _GEN_476 = 8'h71 == _T_40[7:0] ? 4'hf : _GEN_475; // @[Filter.scala 160:102]
  wire [3:0] _GEN_477 = 8'h72 == _T_40[7:0] ? 4'hf : _GEN_476; // @[Filter.scala 160:102]
  wire [3:0] _GEN_478 = 8'h73 == _T_40[7:0] ? 4'hf : _GEN_477; // @[Filter.scala 160:102]
  wire [3:0] _GEN_479 = 8'h74 == _T_40[7:0] ? 4'hf : _GEN_478; // @[Filter.scala 160:102]
  wire [3:0] _GEN_480 = 8'h75 == _T_40[7:0] ? 4'hf : _GEN_479; // @[Filter.scala 160:102]
  wire [3:0] _GEN_481 = 8'h76 == _T_40[7:0] ? 4'hf : _GEN_480; // @[Filter.scala 160:102]
  wire [3:0] _GEN_482 = 8'h77 == _T_40[7:0] ? 4'hf : _GEN_481; // @[Filter.scala 160:102]
  wire [3:0] _GEN_483 = 8'h78 == _T_40[7:0] ? 4'hf : _GEN_482; // @[Filter.scala 160:102]
  wire [3:0] _GEN_484 = 8'h79 == _T_40[7:0] ? 4'hf : _GEN_483; // @[Filter.scala 160:102]
  wire [3:0] _GEN_485 = 8'h7a == _T_40[7:0] ? 4'hf : _GEN_484; // @[Filter.scala 160:102]
  wire [3:0] _GEN_486 = 8'h7b == _T_40[7:0] ? 4'hf : _GEN_485; // @[Filter.scala 160:102]
  wire [3:0] _GEN_487 = 8'h7c == _T_40[7:0] ? 4'hf : _GEN_486; // @[Filter.scala 160:102]
  wire [3:0] _GEN_488 = 8'h7d == _T_40[7:0] ? 4'hf : _GEN_487; // @[Filter.scala 160:102]
  wire [3:0] _GEN_489 = 8'h7e == _T_40[7:0] ? 4'hf : _GEN_488; // @[Filter.scala 160:102]
  wire [3:0] _GEN_490 = 8'h7f == _T_40[7:0] ? 4'hf : _GEN_489; // @[Filter.scala 160:102]
  wire [3:0] _GEN_491 = 8'h80 == _T_40[7:0] ? 4'hf : _GEN_490; // @[Filter.scala 160:102]
  wire [3:0] _GEN_492 = 8'h81 == _T_40[7:0] ? 4'hf : _GEN_491; // @[Filter.scala 160:102]
  wire [3:0] _GEN_493 = 8'h82 == _T_40[7:0] ? 4'hf : _GEN_492; // @[Filter.scala 160:102]
  wire [3:0] _GEN_494 = 8'h83 == _T_40[7:0] ? 4'hf : _GEN_493; // @[Filter.scala 160:102]
  wire [3:0] _GEN_495 = 8'h84 == _T_40[7:0] ? 4'hf : _GEN_494; // @[Filter.scala 160:102]
  wire [3:0] _GEN_496 = 8'h85 == _T_40[7:0] ? 4'hf : _GEN_495; // @[Filter.scala 160:102]
  wire [3:0] _GEN_497 = 8'h86 == _T_40[7:0] ? 4'hf : _GEN_496; // @[Filter.scala 160:102]
  wire [3:0] _GEN_498 = 8'h87 == _T_40[7:0] ? 4'hf : _GEN_497; // @[Filter.scala 160:102]
  wire [3:0] _GEN_499 = 8'h88 == _T_40[7:0] ? 4'hf : _GEN_498; // @[Filter.scala 160:102]
  wire [3:0] _GEN_500 = 8'h89 == _T_40[7:0] ? 4'hf : _GEN_499; // @[Filter.scala 160:102]
  wire [3:0] _GEN_501 = 8'h8a == _T_40[7:0] ? 4'hf : _GEN_500; // @[Filter.scala 160:102]
  wire [3:0] _GEN_502 = 8'h8b == _T_40[7:0] ? 4'hf : _GEN_501; // @[Filter.scala 160:102]
  wire [3:0] _GEN_503 = 8'h8c == _T_40[7:0] ? 4'hf : _GEN_502; // @[Filter.scala 160:102]
  wire [3:0] _GEN_504 = 8'h8d == _T_40[7:0] ? 4'hf : _GEN_503; // @[Filter.scala 160:102]
  wire [3:0] _GEN_505 = 8'h8e == _T_40[7:0] ? 4'hf : _GEN_504; // @[Filter.scala 160:102]
  wire [3:0] _GEN_506 = 8'h8f == _T_40[7:0] ? 4'hf : _GEN_505; // @[Filter.scala 160:102]
  wire [3:0] _GEN_507 = 8'h90 == _T_40[7:0] ? 4'hf : _GEN_506; // @[Filter.scala 160:102]
  wire [3:0] _GEN_508 = 8'h91 == _T_40[7:0] ? 4'hf : _GEN_507; // @[Filter.scala 160:102]
  wire [3:0] _GEN_509 = 8'h92 == _T_40[7:0] ? 4'hf : _GEN_508; // @[Filter.scala 160:102]
  wire [3:0] _GEN_510 = 8'h93 == _T_40[7:0] ? 4'hf : _GEN_509; // @[Filter.scala 160:102]
  wire [3:0] _GEN_511 = 8'h94 == _T_40[7:0] ? 4'hf : _GEN_510; // @[Filter.scala 160:102]
  wire [3:0] _GEN_512 = 8'h95 == _T_40[7:0] ? 4'hf : _GEN_511; // @[Filter.scala 160:102]
  wire [3:0] _GEN_513 = 8'h96 == _T_40[7:0] ? 4'hf : _GEN_512; // @[Filter.scala 160:102]
  wire [3:0] _GEN_514 = 8'h97 == _T_40[7:0] ? 4'hf : _GEN_513; // @[Filter.scala 160:102]
  wire [3:0] _GEN_515 = 8'h98 == _T_40[7:0] ? 4'hf : _GEN_514; // @[Filter.scala 160:102]
  wire [3:0] _GEN_516 = 8'h99 == _T_40[7:0] ? 4'hf : _GEN_515; // @[Filter.scala 160:102]
  wire [3:0] _GEN_517 = 8'h9a == _T_40[7:0] ? 4'hf : _GEN_516; // @[Filter.scala 160:102]
  wire [3:0] _GEN_518 = 8'h9b == _T_40[7:0] ? 4'hf : _GEN_517; // @[Filter.scala 160:102]
  wire [3:0] _GEN_519 = 8'h9c == _T_40[7:0] ? 4'hf : _GEN_518; // @[Filter.scala 160:102]
  wire [3:0] _GEN_520 = 8'h9d == _T_40[7:0] ? 4'hf : _GEN_519; // @[Filter.scala 160:102]
  wire [3:0] _GEN_521 = 8'h9e == _T_40[7:0] ? 4'hf : _GEN_520; // @[Filter.scala 160:102]
  wire [3:0] _GEN_522 = 8'h9f == _T_40[7:0] ? 4'hf : _GEN_521; // @[Filter.scala 160:102]
  wire [3:0] _GEN_523 = 8'ha0 == _T_40[7:0] ? 4'hf : _GEN_522; // @[Filter.scala 160:102]
  wire [3:0] _GEN_524 = 8'ha1 == _T_40[7:0] ? 4'hf : _GEN_523; // @[Filter.scala 160:102]
  wire [3:0] _GEN_525 = 8'ha2 == _T_40[7:0] ? 4'hf : _GEN_524; // @[Filter.scala 160:102]
  wire [3:0] _GEN_526 = 8'ha3 == _T_40[7:0] ? 4'hf : _GEN_525; // @[Filter.scala 160:102]
  wire [3:0] _GEN_527 = 8'ha4 == _T_40[7:0] ? 4'hf : _GEN_526; // @[Filter.scala 160:102]
  wire [3:0] _GEN_528 = 8'ha5 == _T_40[7:0] ? 4'hf : _GEN_527; // @[Filter.scala 160:102]
  wire [3:0] _GEN_529 = 8'ha6 == _T_40[7:0] ? 4'hf : _GEN_528; // @[Filter.scala 160:102]
  wire [3:0] _GEN_530 = 8'ha7 == _T_40[7:0] ? 4'hf : _GEN_529; // @[Filter.scala 160:102]
  wire [3:0] _GEN_531 = 8'ha8 == _T_40[7:0] ? 4'hf : _GEN_530; // @[Filter.scala 160:102]
  wire [3:0] _GEN_532 = 8'ha9 == _T_40[7:0] ? 4'hf : _GEN_531; // @[Filter.scala 160:102]
  wire [3:0] _GEN_533 = 8'haa == _T_40[7:0] ? 4'hf : _GEN_532; // @[Filter.scala 160:102]
  wire [3:0] _GEN_534 = 8'hab == _T_40[7:0] ? 4'hf : _GEN_533; // @[Filter.scala 160:102]
  wire [3:0] _GEN_535 = 8'hac == _T_40[7:0] ? 4'hf : _GEN_534; // @[Filter.scala 160:102]
  wire [3:0] _GEN_536 = 8'had == _T_40[7:0] ? 4'hf : _GEN_535; // @[Filter.scala 160:102]
  wire [3:0] _GEN_537 = 8'hae == _T_40[7:0] ? 4'hf : _GEN_536; // @[Filter.scala 160:102]
  wire [3:0] _GEN_538 = 8'haf == _T_40[7:0] ? 4'hf : _GEN_537; // @[Filter.scala 160:102]
  wire [3:0] _GEN_539 = 8'hb0 == _T_40[7:0] ? 4'hf : _GEN_538; // @[Filter.scala 160:102]
  wire [3:0] _GEN_540 = 8'hb1 == _T_40[7:0] ? 4'hf : _GEN_539; // @[Filter.scala 160:102]
  wire [3:0] _GEN_541 = 8'hb2 == _T_40[7:0] ? 4'hf : _GEN_540; // @[Filter.scala 160:102]
  wire [3:0] _GEN_542 = 8'hb3 == _T_40[7:0] ? 4'hf : _GEN_541; // @[Filter.scala 160:102]
  wire [3:0] _GEN_543 = 8'hb4 == _T_40[7:0] ? 4'hf : _GEN_542; // @[Filter.scala 160:102]
  wire [3:0] _GEN_544 = 8'hb5 == _T_40[7:0] ? 4'hf : _GEN_543; // @[Filter.scala 160:102]
  wire [3:0] _GEN_545 = 8'hb6 == _T_40[7:0] ? 4'hf : _GEN_544; // @[Filter.scala 160:102]
  wire [3:0] _GEN_546 = 8'hb7 == _T_40[7:0] ? 4'hf : _GEN_545; // @[Filter.scala 160:102]
  wire [3:0] _GEN_547 = 8'hb8 == _T_40[7:0] ? 4'hf : _GEN_546; // @[Filter.scala 160:102]
  wire [3:0] _GEN_548 = 8'hb9 == _T_40[7:0] ? 4'hf : _GEN_547; // @[Filter.scala 160:102]
  wire [3:0] _GEN_549 = 8'hba == _T_40[7:0] ? 4'hf : _GEN_548; // @[Filter.scala 160:102]
  wire [3:0] _GEN_550 = 8'hbb == _T_40[7:0] ? 4'hf : _GEN_549; // @[Filter.scala 160:102]
  wire [3:0] _GEN_551 = 8'hbc == _T_40[7:0] ? 4'hf : _GEN_550; // @[Filter.scala 160:102]
  wire [3:0] _GEN_552 = 8'hbd == _T_40[7:0] ? 4'hf : _GEN_551; // @[Filter.scala 160:102]
  wire [3:0] _GEN_553 = 8'hbe == _T_40[7:0] ? 4'hf : _GEN_552; // @[Filter.scala 160:102]
  wire [3:0] _GEN_554 = 8'hbf == _T_40[7:0] ? 4'hf : _GEN_553; // @[Filter.scala 160:102]
  wire [6:0] _GEN_9868 = {{3'd0}, _GEN_554}; // @[Filter.scala 160:102]
  wire [10:0] _T_47 = _GEN_9868 * 7'h46; // @[Filter.scala 160:102]
  wire [10:0] _GEN_9869 = {{2'd0}, _T_42}; // @[Filter.scala 160:69]
  wire [10:0] _T_49 = _GEN_9869 + _T_47; // @[Filter.scala 160:69]
  wire [3:0] _GEN_563 = 8'h8 == _T_40[7:0] ? 4'hf : 4'h0; // @[Filter.scala 160:142]
  wire [3:0] _GEN_564 = 8'h9 == _T_40[7:0] ? 4'hf : _GEN_563; // @[Filter.scala 160:142]
  wire [3:0] _GEN_565 = 8'ha == _T_40[7:0] ? 4'hf : _GEN_564; // @[Filter.scala 160:142]
  wire [3:0] _GEN_566 = 8'hb == _T_40[7:0] ? 4'hf : _GEN_565; // @[Filter.scala 160:142]
  wire [3:0] _GEN_567 = 8'hc == _T_40[7:0] ? 4'hf : _GEN_566; // @[Filter.scala 160:142]
  wire [3:0] _GEN_568 = 8'hd == _T_40[7:0] ? 4'hf : _GEN_567; // @[Filter.scala 160:142]
  wire [3:0] _GEN_569 = 8'he == _T_40[7:0] ? 4'hf : _GEN_568; // @[Filter.scala 160:142]
  wire [3:0] _GEN_570 = 8'hf == _T_40[7:0] ? 4'hf : _GEN_569; // @[Filter.scala 160:142]
  wire [3:0] _GEN_571 = 8'h10 == _T_40[7:0] ? 4'h0 : _GEN_570; // @[Filter.scala 160:142]
  wire [3:0] _GEN_572 = 8'h11 == _T_40[7:0] ? 4'h0 : _GEN_571; // @[Filter.scala 160:142]
  wire [3:0] _GEN_573 = 8'h12 == _T_40[7:0] ? 4'h0 : _GEN_572; // @[Filter.scala 160:142]
  wire [3:0] _GEN_574 = 8'h13 == _T_40[7:0] ? 4'h0 : _GEN_573; // @[Filter.scala 160:142]
  wire [3:0] _GEN_575 = 8'h14 == _T_40[7:0] ? 4'h0 : _GEN_574; // @[Filter.scala 160:142]
  wire [3:0] _GEN_576 = 8'h15 == _T_40[7:0] ? 4'h0 : _GEN_575; // @[Filter.scala 160:142]
  wire [3:0] _GEN_577 = 8'h16 == _T_40[7:0] ? 4'h0 : _GEN_576; // @[Filter.scala 160:142]
  wire [3:0] _GEN_578 = 8'h17 == _T_40[7:0] ? 4'h0 : _GEN_577; // @[Filter.scala 160:142]
  wire [3:0] _GEN_579 = 8'h18 == _T_40[7:0] ? 4'hf : _GEN_578; // @[Filter.scala 160:142]
  wire [3:0] _GEN_580 = 8'h19 == _T_40[7:0] ? 4'hf : _GEN_579; // @[Filter.scala 160:142]
  wire [3:0] _GEN_581 = 8'h1a == _T_40[7:0] ? 4'hf : _GEN_580; // @[Filter.scala 160:142]
  wire [3:0] _GEN_582 = 8'h1b == _T_40[7:0] ? 4'hf : _GEN_581; // @[Filter.scala 160:142]
  wire [3:0] _GEN_583 = 8'h1c == _T_40[7:0] ? 4'hf : _GEN_582; // @[Filter.scala 160:142]
  wire [3:0] _GEN_584 = 8'h1d == _T_40[7:0] ? 4'hf : _GEN_583; // @[Filter.scala 160:142]
  wire [3:0] _GEN_585 = 8'h1e == _T_40[7:0] ? 4'hf : _GEN_584; // @[Filter.scala 160:142]
  wire [3:0] _GEN_586 = 8'h1f == _T_40[7:0] ? 4'hf : _GEN_585; // @[Filter.scala 160:142]
  wire [3:0] _GEN_587 = 8'h20 == _T_40[7:0] ? 4'h0 : _GEN_586; // @[Filter.scala 160:142]
  wire [3:0] _GEN_588 = 8'h21 == _T_40[7:0] ? 4'h0 : _GEN_587; // @[Filter.scala 160:142]
  wire [3:0] _GEN_589 = 8'h22 == _T_40[7:0] ? 4'h0 : _GEN_588; // @[Filter.scala 160:142]
  wire [3:0] _GEN_590 = 8'h23 == _T_40[7:0] ? 4'h0 : _GEN_589; // @[Filter.scala 160:142]
  wire [3:0] _GEN_591 = 8'h24 == _T_40[7:0] ? 4'h0 : _GEN_590; // @[Filter.scala 160:142]
  wire [3:0] _GEN_592 = 8'h25 == _T_40[7:0] ? 4'h0 : _GEN_591; // @[Filter.scala 160:142]
  wire [3:0] _GEN_593 = 8'h26 == _T_40[7:0] ? 4'h0 : _GEN_592; // @[Filter.scala 160:142]
  wire [3:0] _GEN_594 = 8'h27 == _T_40[7:0] ? 4'h0 : _GEN_593; // @[Filter.scala 160:142]
  wire [3:0] _GEN_595 = 8'h28 == _T_40[7:0] ? 4'hf : _GEN_594; // @[Filter.scala 160:142]
  wire [3:0] _GEN_596 = 8'h29 == _T_40[7:0] ? 4'hf : _GEN_595; // @[Filter.scala 160:142]
  wire [3:0] _GEN_597 = 8'h2a == _T_40[7:0] ? 4'hf : _GEN_596; // @[Filter.scala 160:142]
  wire [3:0] _GEN_598 = 8'h2b == _T_40[7:0] ? 4'hf : _GEN_597; // @[Filter.scala 160:142]
  wire [3:0] _GEN_599 = 8'h2c == _T_40[7:0] ? 4'hf : _GEN_598; // @[Filter.scala 160:142]
  wire [3:0] _GEN_600 = 8'h2d == _T_40[7:0] ? 4'hf : _GEN_599; // @[Filter.scala 160:142]
  wire [3:0] _GEN_601 = 8'h2e == _T_40[7:0] ? 4'hf : _GEN_600; // @[Filter.scala 160:142]
  wire [3:0] _GEN_602 = 8'h2f == _T_40[7:0] ? 4'hf : _GEN_601; // @[Filter.scala 160:142]
  wire [3:0] _GEN_603 = 8'h30 == _T_40[7:0] ? 4'h0 : _GEN_602; // @[Filter.scala 160:142]
  wire [3:0] _GEN_604 = 8'h31 == _T_40[7:0] ? 4'h0 : _GEN_603; // @[Filter.scala 160:142]
  wire [3:0] _GEN_605 = 8'h32 == _T_40[7:0] ? 4'h0 : _GEN_604; // @[Filter.scala 160:142]
  wire [3:0] _GEN_606 = 8'h33 == _T_40[7:0] ? 4'h0 : _GEN_605; // @[Filter.scala 160:142]
  wire [3:0] _GEN_607 = 8'h34 == _T_40[7:0] ? 4'h0 : _GEN_606; // @[Filter.scala 160:142]
  wire [3:0] _GEN_608 = 8'h35 == _T_40[7:0] ? 4'h0 : _GEN_607; // @[Filter.scala 160:142]
  wire [3:0] _GEN_609 = 8'h36 == _T_40[7:0] ? 4'h0 : _GEN_608; // @[Filter.scala 160:142]
  wire [3:0] _GEN_610 = 8'h37 == _T_40[7:0] ? 4'h0 : _GEN_609; // @[Filter.scala 160:142]
  wire [3:0] _GEN_611 = 8'h38 == _T_40[7:0] ? 4'hf : _GEN_610; // @[Filter.scala 160:142]
  wire [3:0] _GEN_612 = 8'h39 == _T_40[7:0] ? 4'hf : _GEN_611; // @[Filter.scala 160:142]
  wire [3:0] _GEN_613 = 8'h3a == _T_40[7:0] ? 4'hf : _GEN_612; // @[Filter.scala 160:142]
  wire [3:0] _GEN_614 = 8'h3b == _T_40[7:0] ? 4'hf : _GEN_613; // @[Filter.scala 160:142]
  wire [3:0] _GEN_615 = 8'h3c == _T_40[7:0] ? 4'hf : _GEN_614; // @[Filter.scala 160:142]
  wire [3:0] _GEN_616 = 8'h3d == _T_40[7:0] ? 4'hf : _GEN_615; // @[Filter.scala 160:142]
  wire [3:0] _GEN_617 = 8'h3e == _T_40[7:0] ? 4'hf : _GEN_616; // @[Filter.scala 160:142]
  wire [3:0] _GEN_618 = 8'h3f == _T_40[7:0] ? 4'hf : _GEN_617; // @[Filter.scala 160:142]
  wire [3:0] _GEN_619 = 8'h40 == _T_40[7:0] ? 4'h0 : _GEN_618; // @[Filter.scala 160:142]
  wire [3:0] _GEN_620 = 8'h41 == _T_40[7:0] ? 4'h0 : _GEN_619; // @[Filter.scala 160:142]
  wire [3:0] _GEN_621 = 8'h42 == _T_40[7:0] ? 4'h0 : _GEN_620; // @[Filter.scala 160:142]
  wire [3:0] _GEN_622 = 8'h43 == _T_40[7:0] ? 4'h0 : _GEN_621; // @[Filter.scala 160:142]
  wire [3:0] _GEN_623 = 8'h44 == _T_40[7:0] ? 4'h0 : _GEN_622; // @[Filter.scala 160:142]
  wire [3:0] _GEN_624 = 8'h45 == _T_40[7:0] ? 4'h0 : _GEN_623; // @[Filter.scala 160:142]
  wire [3:0] _GEN_625 = 8'h46 == _T_40[7:0] ? 4'h0 : _GEN_624; // @[Filter.scala 160:142]
  wire [3:0] _GEN_626 = 8'h47 == _T_40[7:0] ? 4'h0 : _GEN_625; // @[Filter.scala 160:142]
  wire [3:0] _GEN_627 = 8'h48 == _T_40[7:0] ? 4'hf : _GEN_626; // @[Filter.scala 160:142]
  wire [3:0] _GEN_628 = 8'h49 == _T_40[7:0] ? 4'hf : _GEN_627; // @[Filter.scala 160:142]
  wire [3:0] _GEN_629 = 8'h4a == _T_40[7:0] ? 4'hf : _GEN_628; // @[Filter.scala 160:142]
  wire [3:0] _GEN_630 = 8'h4b == _T_40[7:0] ? 4'hf : _GEN_629; // @[Filter.scala 160:142]
  wire [3:0] _GEN_631 = 8'h4c == _T_40[7:0] ? 4'hf : _GEN_630; // @[Filter.scala 160:142]
  wire [3:0] _GEN_632 = 8'h4d == _T_40[7:0] ? 4'hf : _GEN_631; // @[Filter.scala 160:142]
  wire [3:0] _GEN_633 = 8'h4e == _T_40[7:0] ? 4'hf : _GEN_632; // @[Filter.scala 160:142]
  wire [3:0] _GEN_634 = 8'h4f == _T_40[7:0] ? 4'hf : _GEN_633; // @[Filter.scala 160:142]
  wire [3:0] _GEN_635 = 8'h50 == _T_40[7:0] ? 4'h0 : _GEN_634; // @[Filter.scala 160:142]
  wire [3:0] _GEN_636 = 8'h51 == _T_40[7:0] ? 4'h0 : _GEN_635; // @[Filter.scala 160:142]
  wire [3:0] _GEN_637 = 8'h52 == _T_40[7:0] ? 4'h0 : _GEN_636; // @[Filter.scala 160:142]
  wire [3:0] _GEN_638 = 8'h53 == _T_40[7:0] ? 4'h0 : _GEN_637; // @[Filter.scala 160:142]
  wire [3:0] _GEN_639 = 8'h54 == _T_40[7:0] ? 4'h0 : _GEN_638; // @[Filter.scala 160:142]
  wire [3:0] _GEN_640 = 8'h55 == _T_40[7:0] ? 4'h0 : _GEN_639; // @[Filter.scala 160:142]
  wire [3:0] _GEN_641 = 8'h56 == _T_40[7:0] ? 4'h0 : _GEN_640; // @[Filter.scala 160:142]
  wire [3:0] _GEN_642 = 8'h57 == _T_40[7:0] ? 4'h0 : _GEN_641; // @[Filter.scala 160:142]
  wire [3:0] _GEN_643 = 8'h58 == _T_40[7:0] ? 4'hf : _GEN_642; // @[Filter.scala 160:142]
  wire [3:0] _GEN_644 = 8'h59 == _T_40[7:0] ? 4'hf : _GEN_643; // @[Filter.scala 160:142]
  wire [3:0] _GEN_645 = 8'h5a == _T_40[7:0] ? 4'hf : _GEN_644; // @[Filter.scala 160:142]
  wire [3:0] _GEN_646 = 8'h5b == _T_40[7:0] ? 4'hf : _GEN_645; // @[Filter.scala 160:142]
  wire [3:0] _GEN_647 = 8'h5c == _T_40[7:0] ? 4'hf : _GEN_646; // @[Filter.scala 160:142]
  wire [3:0] _GEN_648 = 8'h5d == _T_40[7:0] ? 4'hf : _GEN_647; // @[Filter.scala 160:142]
  wire [3:0] _GEN_649 = 8'h5e == _T_40[7:0] ? 4'hf : _GEN_648; // @[Filter.scala 160:142]
  wire [3:0] _GEN_650 = 8'h5f == _T_40[7:0] ? 4'hf : _GEN_649; // @[Filter.scala 160:142]
  wire [3:0] _GEN_651 = 8'h60 == _T_40[7:0] ? 4'h0 : _GEN_650; // @[Filter.scala 160:142]
  wire [3:0] _GEN_652 = 8'h61 == _T_40[7:0] ? 4'h0 : _GEN_651; // @[Filter.scala 160:142]
  wire [3:0] _GEN_653 = 8'h62 == _T_40[7:0] ? 4'h0 : _GEN_652; // @[Filter.scala 160:142]
  wire [3:0] _GEN_654 = 8'h63 == _T_40[7:0] ? 4'h0 : _GEN_653; // @[Filter.scala 160:142]
  wire [3:0] _GEN_655 = 8'h64 == _T_40[7:0] ? 4'h0 : _GEN_654; // @[Filter.scala 160:142]
  wire [3:0] _GEN_656 = 8'h65 == _T_40[7:0] ? 4'h0 : _GEN_655; // @[Filter.scala 160:142]
  wire [3:0] _GEN_657 = 8'h66 == _T_40[7:0] ? 4'h0 : _GEN_656; // @[Filter.scala 160:142]
  wire [3:0] _GEN_658 = 8'h67 == _T_40[7:0] ? 4'h0 : _GEN_657; // @[Filter.scala 160:142]
  wire [3:0] _GEN_659 = 8'h68 == _T_40[7:0] ? 4'hf : _GEN_658; // @[Filter.scala 160:142]
  wire [3:0] _GEN_660 = 8'h69 == _T_40[7:0] ? 4'hf : _GEN_659; // @[Filter.scala 160:142]
  wire [3:0] _GEN_661 = 8'h6a == _T_40[7:0] ? 4'hf : _GEN_660; // @[Filter.scala 160:142]
  wire [3:0] _GEN_662 = 8'h6b == _T_40[7:0] ? 4'hf : _GEN_661; // @[Filter.scala 160:142]
  wire [3:0] _GEN_663 = 8'h6c == _T_40[7:0] ? 4'hf : _GEN_662; // @[Filter.scala 160:142]
  wire [3:0] _GEN_664 = 8'h6d == _T_40[7:0] ? 4'hf : _GEN_663; // @[Filter.scala 160:142]
  wire [3:0] _GEN_665 = 8'h6e == _T_40[7:0] ? 4'hf : _GEN_664; // @[Filter.scala 160:142]
  wire [3:0] _GEN_666 = 8'h6f == _T_40[7:0] ? 4'hf : _GEN_665; // @[Filter.scala 160:142]
  wire [3:0] _GEN_667 = 8'h70 == _T_40[7:0] ? 4'h0 : _GEN_666; // @[Filter.scala 160:142]
  wire [3:0] _GEN_668 = 8'h71 == _T_40[7:0] ? 4'h0 : _GEN_667; // @[Filter.scala 160:142]
  wire [3:0] _GEN_669 = 8'h72 == _T_40[7:0] ? 4'h0 : _GEN_668; // @[Filter.scala 160:142]
  wire [3:0] _GEN_670 = 8'h73 == _T_40[7:0] ? 4'h0 : _GEN_669; // @[Filter.scala 160:142]
  wire [3:0] _GEN_671 = 8'h74 == _T_40[7:0] ? 4'h0 : _GEN_670; // @[Filter.scala 160:142]
  wire [3:0] _GEN_672 = 8'h75 == _T_40[7:0] ? 4'h0 : _GEN_671; // @[Filter.scala 160:142]
  wire [3:0] _GEN_673 = 8'h76 == _T_40[7:0] ? 4'h0 : _GEN_672; // @[Filter.scala 160:142]
  wire [3:0] _GEN_674 = 8'h77 == _T_40[7:0] ? 4'h0 : _GEN_673; // @[Filter.scala 160:142]
  wire [3:0] _GEN_675 = 8'h78 == _T_40[7:0] ? 4'hf : _GEN_674; // @[Filter.scala 160:142]
  wire [3:0] _GEN_676 = 8'h79 == _T_40[7:0] ? 4'hf : _GEN_675; // @[Filter.scala 160:142]
  wire [3:0] _GEN_677 = 8'h7a == _T_40[7:0] ? 4'hf : _GEN_676; // @[Filter.scala 160:142]
  wire [3:0] _GEN_678 = 8'h7b == _T_40[7:0] ? 4'hf : _GEN_677; // @[Filter.scala 160:142]
  wire [3:0] _GEN_679 = 8'h7c == _T_40[7:0] ? 4'hf : _GEN_678; // @[Filter.scala 160:142]
  wire [3:0] _GEN_680 = 8'h7d == _T_40[7:0] ? 4'hf : _GEN_679; // @[Filter.scala 160:142]
  wire [3:0] _GEN_681 = 8'h7e == _T_40[7:0] ? 4'hf : _GEN_680; // @[Filter.scala 160:142]
  wire [3:0] _GEN_682 = 8'h7f == _T_40[7:0] ? 4'hf : _GEN_681; // @[Filter.scala 160:142]
  wire [3:0] _GEN_683 = 8'h80 == _T_40[7:0] ? 4'h0 : _GEN_682; // @[Filter.scala 160:142]
  wire [3:0] _GEN_684 = 8'h81 == _T_40[7:0] ? 4'h0 : _GEN_683; // @[Filter.scala 160:142]
  wire [3:0] _GEN_685 = 8'h82 == _T_40[7:0] ? 4'h0 : _GEN_684; // @[Filter.scala 160:142]
  wire [3:0] _GEN_686 = 8'h83 == _T_40[7:0] ? 4'h0 : _GEN_685; // @[Filter.scala 160:142]
  wire [3:0] _GEN_687 = 8'h84 == _T_40[7:0] ? 4'h0 : _GEN_686; // @[Filter.scala 160:142]
  wire [3:0] _GEN_688 = 8'h85 == _T_40[7:0] ? 4'h0 : _GEN_687; // @[Filter.scala 160:142]
  wire [3:0] _GEN_689 = 8'h86 == _T_40[7:0] ? 4'h0 : _GEN_688; // @[Filter.scala 160:142]
  wire [3:0] _GEN_690 = 8'h87 == _T_40[7:0] ? 4'h0 : _GEN_689; // @[Filter.scala 160:142]
  wire [3:0] _GEN_691 = 8'h88 == _T_40[7:0] ? 4'hf : _GEN_690; // @[Filter.scala 160:142]
  wire [3:0] _GEN_692 = 8'h89 == _T_40[7:0] ? 4'hf : _GEN_691; // @[Filter.scala 160:142]
  wire [3:0] _GEN_693 = 8'h8a == _T_40[7:0] ? 4'hf : _GEN_692; // @[Filter.scala 160:142]
  wire [3:0] _GEN_694 = 8'h8b == _T_40[7:0] ? 4'hf : _GEN_693; // @[Filter.scala 160:142]
  wire [3:0] _GEN_695 = 8'h8c == _T_40[7:0] ? 4'hf : _GEN_694; // @[Filter.scala 160:142]
  wire [3:0] _GEN_696 = 8'h8d == _T_40[7:0] ? 4'hf : _GEN_695; // @[Filter.scala 160:142]
  wire [3:0] _GEN_697 = 8'h8e == _T_40[7:0] ? 4'hf : _GEN_696; // @[Filter.scala 160:142]
  wire [3:0] _GEN_698 = 8'h8f == _T_40[7:0] ? 4'hf : _GEN_697; // @[Filter.scala 160:142]
  wire [3:0] _GEN_699 = 8'h90 == _T_40[7:0] ? 4'h0 : _GEN_698; // @[Filter.scala 160:142]
  wire [3:0] _GEN_700 = 8'h91 == _T_40[7:0] ? 4'h0 : _GEN_699; // @[Filter.scala 160:142]
  wire [3:0] _GEN_701 = 8'h92 == _T_40[7:0] ? 4'h0 : _GEN_700; // @[Filter.scala 160:142]
  wire [3:0] _GEN_702 = 8'h93 == _T_40[7:0] ? 4'h0 : _GEN_701; // @[Filter.scala 160:142]
  wire [3:0] _GEN_703 = 8'h94 == _T_40[7:0] ? 4'h0 : _GEN_702; // @[Filter.scala 160:142]
  wire [3:0] _GEN_704 = 8'h95 == _T_40[7:0] ? 4'h0 : _GEN_703; // @[Filter.scala 160:142]
  wire [3:0] _GEN_705 = 8'h96 == _T_40[7:0] ? 4'h0 : _GEN_704; // @[Filter.scala 160:142]
  wire [3:0] _GEN_706 = 8'h97 == _T_40[7:0] ? 4'h0 : _GEN_705; // @[Filter.scala 160:142]
  wire [3:0] _GEN_707 = 8'h98 == _T_40[7:0] ? 4'hf : _GEN_706; // @[Filter.scala 160:142]
  wire [3:0] _GEN_708 = 8'h99 == _T_40[7:0] ? 4'hf : _GEN_707; // @[Filter.scala 160:142]
  wire [3:0] _GEN_709 = 8'h9a == _T_40[7:0] ? 4'hf : _GEN_708; // @[Filter.scala 160:142]
  wire [3:0] _GEN_710 = 8'h9b == _T_40[7:0] ? 4'hf : _GEN_709; // @[Filter.scala 160:142]
  wire [3:0] _GEN_711 = 8'h9c == _T_40[7:0] ? 4'hf : _GEN_710; // @[Filter.scala 160:142]
  wire [3:0] _GEN_712 = 8'h9d == _T_40[7:0] ? 4'hf : _GEN_711; // @[Filter.scala 160:142]
  wire [3:0] _GEN_713 = 8'h9e == _T_40[7:0] ? 4'hf : _GEN_712; // @[Filter.scala 160:142]
  wire [3:0] _GEN_714 = 8'h9f == _T_40[7:0] ? 4'hf : _GEN_713; // @[Filter.scala 160:142]
  wire [3:0] _GEN_715 = 8'ha0 == _T_40[7:0] ? 4'h0 : _GEN_714; // @[Filter.scala 160:142]
  wire [3:0] _GEN_716 = 8'ha1 == _T_40[7:0] ? 4'h0 : _GEN_715; // @[Filter.scala 160:142]
  wire [3:0] _GEN_717 = 8'ha2 == _T_40[7:0] ? 4'h0 : _GEN_716; // @[Filter.scala 160:142]
  wire [3:0] _GEN_718 = 8'ha3 == _T_40[7:0] ? 4'h0 : _GEN_717; // @[Filter.scala 160:142]
  wire [3:0] _GEN_719 = 8'ha4 == _T_40[7:0] ? 4'h0 : _GEN_718; // @[Filter.scala 160:142]
  wire [3:0] _GEN_720 = 8'ha5 == _T_40[7:0] ? 4'h0 : _GEN_719; // @[Filter.scala 160:142]
  wire [3:0] _GEN_721 = 8'ha6 == _T_40[7:0] ? 4'h0 : _GEN_720; // @[Filter.scala 160:142]
  wire [3:0] _GEN_722 = 8'ha7 == _T_40[7:0] ? 4'h0 : _GEN_721; // @[Filter.scala 160:142]
  wire [3:0] _GEN_723 = 8'ha8 == _T_40[7:0] ? 4'hf : _GEN_722; // @[Filter.scala 160:142]
  wire [3:0] _GEN_724 = 8'ha9 == _T_40[7:0] ? 4'hf : _GEN_723; // @[Filter.scala 160:142]
  wire [3:0] _GEN_725 = 8'haa == _T_40[7:0] ? 4'hf : _GEN_724; // @[Filter.scala 160:142]
  wire [3:0] _GEN_726 = 8'hab == _T_40[7:0] ? 4'hf : _GEN_725; // @[Filter.scala 160:142]
  wire [3:0] _GEN_727 = 8'hac == _T_40[7:0] ? 4'hf : _GEN_726; // @[Filter.scala 160:142]
  wire [3:0] _GEN_728 = 8'had == _T_40[7:0] ? 4'hf : _GEN_727; // @[Filter.scala 160:142]
  wire [3:0] _GEN_729 = 8'hae == _T_40[7:0] ? 4'hf : _GEN_728; // @[Filter.scala 160:142]
  wire [3:0] _GEN_730 = 8'haf == _T_40[7:0] ? 4'hf : _GEN_729; // @[Filter.scala 160:142]
  wire [3:0] _GEN_731 = 8'hb0 == _T_40[7:0] ? 4'h0 : _GEN_730; // @[Filter.scala 160:142]
  wire [3:0] _GEN_732 = 8'hb1 == _T_40[7:0] ? 4'h0 : _GEN_731; // @[Filter.scala 160:142]
  wire [3:0] _GEN_733 = 8'hb2 == _T_40[7:0] ? 4'h0 : _GEN_732; // @[Filter.scala 160:142]
  wire [3:0] _GEN_734 = 8'hb3 == _T_40[7:0] ? 4'h0 : _GEN_733; // @[Filter.scala 160:142]
  wire [3:0] _GEN_735 = 8'hb4 == _T_40[7:0] ? 4'h0 : _GEN_734; // @[Filter.scala 160:142]
  wire [3:0] _GEN_736 = 8'hb5 == _T_40[7:0] ? 4'h0 : _GEN_735; // @[Filter.scala 160:142]
  wire [3:0] _GEN_737 = 8'hb6 == _T_40[7:0] ? 4'h0 : _GEN_736; // @[Filter.scala 160:142]
  wire [3:0] _GEN_738 = 8'hb7 == _T_40[7:0] ? 4'h0 : _GEN_737; // @[Filter.scala 160:142]
  wire [3:0] _GEN_739 = 8'hb8 == _T_40[7:0] ? 4'hf : _GEN_738; // @[Filter.scala 160:142]
  wire [3:0] _GEN_740 = 8'hb9 == _T_40[7:0] ? 4'hf : _GEN_739; // @[Filter.scala 160:142]
  wire [3:0] _GEN_741 = 8'hba == _T_40[7:0] ? 4'hf : _GEN_740; // @[Filter.scala 160:142]
  wire [3:0] _GEN_742 = 8'hbb == _T_40[7:0] ? 4'hf : _GEN_741; // @[Filter.scala 160:142]
  wire [3:0] _GEN_743 = 8'hbc == _T_40[7:0] ? 4'hf : _GEN_742; // @[Filter.scala 160:142]
  wire [3:0] _GEN_744 = 8'hbd == _T_40[7:0] ? 4'hf : _GEN_743; // @[Filter.scala 160:142]
  wire [3:0] _GEN_745 = 8'hbe == _T_40[7:0] ? 4'hf : _GEN_744; // @[Filter.scala 160:142]
  wire [3:0] _GEN_746 = 8'hbf == _T_40[7:0] ? 4'hf : _GEN_745; // @[Filter.scala 160:142]
  wire [7:0] _T_54 = _GEN_746 * 4'ha; // @[Filter.scala 160:142]
  wire [10:0] _GEN_9871 = {{3'd0}, _T_54}; // @[Filter.scala 160:109]
  wire [10:0] _T_56 = _T_49 + _GEN_9871; // @[Filter.scala 160:109]
  wire [10:0] _T_57 = _T_56 / 11'h64; // @[Filter.scala 160:150]
  wire  _T_59 = _T_30 >= 5'h10; // @[Filter.scala 163:31]
  wire  _T_63 = _T_37 >= 32'hc; // @[Filter.scala 163:63]
  wire  _T_64 = _T_59 | _T_63; // @[Filter.scala 163:58]
  wire [10:0] _GEN_939 = io_SPI_distort ? _T_57 : {{7'd0}, _GEN_362}; // @[Filter.scala 165:35]
  wire [10:0] _GEN_940 = _T_64 ? 11'h0 : _GEN_939; // @[Filter.scala 163:80]
  wire [10:0] _GEN_1133 = io_SPI_distort ? _T_57 : {{7'd0}, _GEN_554}; // @[Filter.scala 165:35]
  wire [10:0] _GEN_1134 = _T_64 ? 11'h0 : _GEN_1133; // @[Filter.scala 163:80]
  wire [10:0] _GEN_1327 = io_SPI_distort ? _T_57 : {{7'd0}, _GEN_746}; // @[Filter.scala 165:35]
  wire [10:0] _GEN_1328 = _T_64 ? 11'h0 : _GEN_1327; // @[Filter.scala 163:80]
  wire [31:0] _T_92 = pixelIndex + 32'h1; // @[Filter.scala 158:31]
  wire [31:0] _GEN_1 = _T_92 % 32'h10; // @[Filter.scala 158:38]
  wire [4:0] _T_93 = _GEN_1[4:0]; // @[Filter.scala 158:38]
  wire [4:0] _T_95 = _T_93 + _GEN_9863; // @[Filter.scala 158:53]
  wire [4:0] _T_97 = _T_95 - 5'h1; // @[Filter.scala 158:69]
  wire [31:0] _T_100 = _T_92 / 32'h10; // @[Filter.scala 159:38]
  wire [31:0] _T_102 = _T_100 + _GEN_9864; // @[Filter.scala 159:53]
  wire [31:0] _T_104 = _T_102 - 32'h1; // @[Filter.scala 159:69]
  wire [36:0] _T_105 = _T_104 * 32'h10; // @[Filter.scala 160:42]
  wire [36:0] _GEN_9877 = {{32'd0}, _T_97}; // @[Filter.scala 160:57]
  wire [36:0] _T_107 = _T_105 + _GEN_9877; // @[Filter.scala 160:57]
  wire [3:0] _GEN_1337 = 8'h8 == _T_107[7:0] ? 4'h0 : 4'hf; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1338 = 8'h9 == _T_107[7:0] ? 4'h0 : _GEN_1337; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1339 = 8'ha == _T_107[7:0] ? 4'h0 : _GEN_1338; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1340 = 8'hb == _T_107[7:0] ? 4'h0 : _GEN_1339; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1341 = 8'hc == _T_107[7:0] ? 4'h0 : _GEN_1340; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1342 = 8'hd == _T_107[7:0] ? 4'h0 : _GEN_1341; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1343 = 8'he == _T_107[7:0] ? 4'h0 : _GEN_1342; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1344 = 8'hf == _T_107[7:0] ? 4'h0 : _GEN_1343; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1345 = 8'h10 == _T_107[7:0] ? 4'hf : _GEN_1344; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1346 = 8'h11 == _T_107[7:0] ? 4'hf : _GEN_1345; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1347 = 8'h12 == _T_107[7:0] ? 4'hf : _GEN_1346; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1348 = 8'h13 == _T_107[7:0] ? 4'hf : _GEN_1347; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1349 = 8'h14 == _T_107[7:0] ? 4'hf : _GEN_1348; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1350 = 8'h15 == _T_107[7:0] ? 4'hf : _GEN_1349; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1351 = 8'h16 == _T_107[7:0] ? 4'hf : _GEN_1350; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1352 = 8'h17 == _T_107[7:0] ? 4'hf : _GEN_1351; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1353 = 8'h18 == _T_107[7:0] ? 4'h0 : _GEN_1352; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1354 = 8'h19 == _T_107[7:0] ? 4'h0 : _GEN_1353; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1355 = 8'h1a == _T_107[7:0] ? 4'h0 : _GEN_1354; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1356 = 8'h1b == _T_107[7:0] ? 4'h0 : _GEN_1355; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1357 = 8'h1c == _T_107[7:0] ? 4'h0 : _GEN_1356; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1358 = 8'h1d == _T_107[7:0] ? 4'h0 : _GEN_1357; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1359 = 8'h1e == _T_107[7:0] ? 4'h0 : _GEN_1358; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1360 = 8'h1f == _T_107[7:0] ? 4'h0 : _GEN_1359; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1361 = 8'h20 == _T_107[7:0] ? 4'hf : _GEN_1360; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1362 = 8'h21 == _T_107[7:0] ? 4'hf : _GEN_1361; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1363 = 8'h22 == _T_107[7:0] ? 4'hf : _GEN_1362; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1364 = 8'h23 == _T_107[7:0] ? 4'hf : _GEN_1363; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1365 = 8'h24 == _T_107[7:0] ? 4'hf : _GEN_1364; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1366 = 8'h25 == _T_107[7:0] ? 4'hf : _GEN_1365; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1367 = 8'h26 == _T_107[7:0] ? 4'hf : _GEN_1366; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1368 = 8'h27 == _T_107[7:0] ? 4'hf : _GEN_1367; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1369 = 8'h28 == _T_107[7:0] ? 4'h0 : _GEN_1368; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1370 = 8'h29 == _T_107[7:0] ? 4'h0 : _GEN_1369; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1371 = 8'h2a == _T_107[7:0] ? 4'h0 : _GEN_1370; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1372 = 8'h2b == _T_107[7:0] ? 4'h0 : _GEN_1371; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1373 = 8'h2c == _T_107[7:0] ? 4'h0 : _GEN_1372; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1374 = 8'h2d == _T_107[7:0] ? 4'h0 : _GEN_1373; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1375 = 8'h2e == _T_107[7:0] ? 4'h0 : _GEN_1374; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1376 = 8'h2f == _T_107[7:0] ? 4'h0 : _GEN_1375; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1377 = 8'h30 == _T_107[7:0] ? 4'hf : _GEN_1376; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1378 = 8'h31 == _T_107[7:0] ? 4'hf : _GEN_1377; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1379 = 8'h32 == _T_107[7:0] ? 4'hf : _GEN_1378; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1380 = 8'h33 == _T_107[7:0] ? 4'hf : _GEN_1379; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1381 = 8'h34 == _T_107[7:0] ? 4'hf : _GEN_1380; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1382 = 8'h35 == _T_107[7:0] ? 4'hf : _GEN_1381; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1383 = 8'h36 == _T_107[7:0] ? 4'hf : _GEN_1382; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1384 = 8'h37 == _T_107[7:0] ? 4'hf : _GEN_1383; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1385 = 8'h38 == _T_107[7:0] ? 4'h0 : _GEN_1384; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1386 = 8'h39 == _T_107[7:0] ? 4'h0 : _GEN_1385; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1387 = 8'h3a == _T_107[7:0] ? 4'h0 : _GEN_1386; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1388 = 8'h3b == _T_107[7:0] ? 4'h0 : _GEN_1387; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1389 = 8'h3c == _T_107[7:0] ? 4'h0 : _GEN_1388; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1390 = 8'h3d == _T_107[7:0] ? 4'h0 : _GEN_1389; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1391 = 8'h3e == _T_107[7:0] ? 4'h0 : _GEN_1390; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1392 = 8'h3f == _T_107[7:0] ? 4'h0 : _GEN_1391; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1393 = 8'h40 == _T_107[7:0] ? 4'hf : _GEN_1392; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1394 = 8'h41 == _T_107[7:0] ? 4'hf : _GEN_1393; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1395 = 8'h42 == _T_107[7:0] ? 4'hf : _GEN_1394; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1396 = 8'h43 == _T_107[7:0] ? 4'hf : _GEN_1395; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1397 = 8'h44 == _T_107[7:0] ? 4'hf : _GEN_1396; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1398 = 8'h45 == _T_107[7:0] ? 4'hf : _GEN_1397; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1399 = 8'h46 == _T_107[7:0] ? 4'hf : _GEN_1398; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1400 = 8'h47 == _T_107[7:0] ? 4'hf : _GEN_1399; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1401 = 8'h48 == _T_107[7:0] ? 4'h0 : _GEN_1400; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1402 = 8'h49 == _T_107[7:0] ? 4'h0 : _GEN_1401; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1403 = 8'h4a == _T_107[7:0] ? 4'h0 : _GEN_1402; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1404 = 8'h4b == _T_107[7:0] ? 4'h0 : _GEN_1403; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1405 = 8'h4c == _T_107[7:0] ? 4'h0 : _GEN_1404; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1406 = 8'h4d == _T_107[7:0] ? 4'h0 : _GEN_1405; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1407 = 8'h4e == _T_107[7:0] ? 4'h0 : _GEN_1406; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1408 = 8'h4f == _T_107[7:0] ? 4'h0 : _GEN_1407; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1409 = 8'h50 == _T_107[7:0] ? 4'hf : _GEN_1408; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1410 = 8'h51 == _T_107[7:0] ? 4'hf : _GEN_1409; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1411 = 8'h52 == _T_107[7:0] ? 4'hf : _GEN_1410; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1412 = 8'h53 == _T_107[7:0] ? 4'hf : _GEN_1411; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1413 = 8'h54 == _T_107[7:0] ? 4'hf : _GEN_1412; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1414 = 8'h55 == _T_107[7:0] ? 4'hf : _GEN_1413; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1415 = 8'h56 == _T_107[7:0] ? 4'hf : _GEN_1414; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1416 = 8'h57 == _T_107[7:0] ? 4'hf : _GEN_1415; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1417 = 8'h58 == _T_107[7:0] ? 4'h0 : _GEN_1416; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1418 = 8'h59 == _T_107[7:0] ? 4'h0 : _GEN_1417; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1419 = 8'h5a == _T_107[7:0] ? 4'h0 : _GEN_1418; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1420 = 8'h5b == _T_107[7:0] ? 4'h0 : _GEN_1419; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1421 = 8'h5c == _T_107[7:0] ? 4'h0 : _GEN_1420; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1422 = 8'h5d == _T_107[7:0] ? 4'h0 : _GEN_1421; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1423 = 8'h5e == _T_107[7:0] ? 4'h0 : _GEN_1422; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1424 = 8'h5f == _T_107[7:0] ? 4'h0 : _GEN_1423; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1425 = 8'h60 == _T_107[7:0] ? 4'h0 : _GEN_1424; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1426 = 8'h61 == _T_107[7:0] ? 4'h0 : _GEN_1425; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1427 = 8'h62 == _T_107[7:0] ? 4'h0 : _GEN_1426; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1428 = 8'h63 == _T_107[7:0] ? 4'h0 : _GEN_1427; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1429 = 8'h64 == _T_107[7:0] ? 4'h0 : _GEN_1428; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1430 = 8'h65 == _T_107[7:0] ? 4'h0 : _GEN_1429; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1431 = 8'h66 == _T_107[7:0] ? 4'h0 : _GEN_1430; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1432 = 8'h67 == _T_107[7:0] ? 4'h0 : _GEN_1431; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1433 = 8'h68 == _T_107[7:0] ? 4'hf : _GEN_1432; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1434 = 8'h69 == _T_107[7:0] ? 4'hf : _GEN_1433; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1435 = 8'h6a == _T_107[7:0] ? 4'hf : _GEN_1434; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1436 = 8'h6b == _T_107[7:0] ? 4'hf : _GEN_1435; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1437 = 8'h6c == _T_107[7:0] ? 4'hf : _GEN_1436; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1438 = 8'h6d == _T_107[7:0] ? 4'hf : _GEN_1437; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1439 = 8'h6e == _T_107[7:0] ? 4'hf : _GEN_1438; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1440 = 8'h6f == _T_107[7:0] ? 4'hf : _GEN_1439; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1441 = 8'h70 == _T_107[7:0] ? 4'h0 : _GEN_1440; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1442 = 8'h71 == _T_107[7:0] ? 4'h0 : _GEN_1441; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1443 = 8'h72 == _T_107[7:0] ? 4'h0 : _GEN_1442; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1444 = 8'h73 == _T_107[7:0] ? 4'h0 : _GEN_1443; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1445 = 8'h74 == _T_107[7:0] ? 4'h0 : _GEN_1444; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1446 = 8'h75 == _T_107[7:0] ? 4'h0 : _GEN_1445; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1447 = 8'h76 == _T_107[7:0] ? 4'h0 : _GEN_1446; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1448 = 8'h77 == _T_107[7:0] ? 4'h0 : _GEN_1447; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1449 = 8'h78 == _T_107[7:0] ? 4'hf : _GEN_1448; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1450 = 8'h79 == _T_107[7:0] ? 4'hf : _GEN_1449; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1451 = 8'h7a == _T_107[7:0] ? 4'hf : _GEN_1450; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1452 = 8'h7b == _T_107[7:0] ? 4'hf : _GEN_1451; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1453 = 8'h7c == _T_107[7:0] ? 4'hf : _GEN_1452; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1454 = 8'h7d == _T_107[7:0] ? 4'hf : _GEN_1453; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1455 = 8'h7e == _T_107[7:0] ? 4'hf : _GEN_1454; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1456 = 8'h7f == _T_107[7:0] ? 4'hf : _GEN_1455; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1457 = 8'h80 == _T_107[7:0] ? 4'h0 : _GEN_1456; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1458 = 8'h81 == _T_107[7:0] ? 4'h0 : _GEN_1457; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1459 = 8'h82 == _T_107[7:0] ? 4'h0 : _GEN_1458; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1460 = 8'h83 == _T_107[7:0] ? 4'h0 : _GEN_1459; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1461 = 8'h84 == _T_107[7:0] ? 4'h0 : _GEN_1460; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1462 = 8'h85 == _T_107[7:0] ? 4'h0 : _GEN_1461; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1463 = 8'h86 == _T_107[7:0] ? 4'h0 : _GEN_1462; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1464 = 8'h87 == _T_107[7:0] ? 4'h0 : _GEN_1463; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1465 = 8'h88 == _T_107[7:0] ? 4'hf : _GEN_1464; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1466 = 8'h89 == _T_107[7:0] ? 4'hf : _GEN_1465; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1467 = 8'h8a == _T_107[7:0] ? 4'hf : _GEN_1466; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1468 = 8'h8b == _T_107[7:0] ? 4'hf : _GEN_1467; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1469 = 8'h8c == _T_107[7:0] ? 4'hf : _GEN_1468; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1470 = 8'h8d == _T_107[7:0] ? 4'hf : _GEN_1469; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1471 = 8'h8e == _T_107[7:0] ? 4'hf : _GEN_1470; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1472 = 8'h8f == _T_107[7:0] ? 4'hf : _GEN_1471; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1473 = 8'h90 == _T_107[7:0] ? 4'h0 : _GEN_1472; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1474 = 8'h91 == _T_107[7:0] ? 4'h0 : _GEN_1473; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1475 = 8'h92 == _T_107[7:0] ? 4'h0 : _GEN_1474; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1476 = 8'h93 == _T_107[7:0] ? 4'h0 : _GEN_1475; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1477 = 8'h94 == _T_107[7:0] ? 4'h0 : _GEN_1476; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1478 = 8'h95 == _T_107[7:0] ? 4'h0 : _GEN_1477; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1479 = 8'h96 == _T_107[7:0] ? 4'h0 : _GEN_1478; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1480 = 8'h97 == _T_107[7:0] ? 4'h0 : _GEN_1479; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1481 = 8'h98 == _T_107[7:0] ? 4'hf : _GEN_1480; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1482 = 8'h99 == _T_107[7:0] ? 4'hf : _GEN_1481; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1483 = 8'h9a == _T_107[7:0] ? 4'hf : _GEN_1482; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1484 = 8'h9b == _T_107[7:0] ? 4'hf : _GEN_1483; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1485 = 8'h9c == _T_107[7:0] ? 4'hf : _GEN_1484; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1486 = 8'h9d == _T_107[7:0] ? 4'hf : _GEN_1485; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1487 = 8'h9e == _T_107[7:0] ? 4'hf : _GEN_1486; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1488 = 8'h9f == _T_107[7:0] ? 4'hf : _GEN_1487; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1489 = 8'ha0 == _T_107[7:0] ? 4'h0 : _GEN_1488; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1490 = 8'ha1 == _T_107[7:0] ? 4'h0 : _GEN_1489; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1491 = 8'ha2 == _T_107[7:0] ? 4'h0 : _GEN_1490; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1492 = 8'ha3 == _T_107[7:0] ? 4'h0 : _GEN_1491; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1493 = 8'ha4 == _T_107[7:0] ? 4'h0 : _GEN_1492; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1494 = 8'ha5 == _T_107[7:0] ? 4'h0 : _GEN_1493; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1495 = 8'ha6 == _T_107[7:0] ? 4'h0 : _GEN_1494; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1496 = 8'ha7 == _T_107[7:0] ? 4'h0 : _GEN_1495; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1497 = 8'ha8 == _T_107[7:0] ? 4'hf : _GEN_1496; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1498 = 8'ha9 == _T_107[7:0] ? 4'hf : _GEN_1497; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1499 = 8'haa == _T_107[7:0] ? 4'hf : _GEN_1498; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1500 = 8'hab == _T_107[7:0] ? 4'hf : _GEN_1499; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1501 = 8'hac == _T_107[7:0] ? 4'hf : _GEN_1500; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1502 = 8'had == _T_107[7:0] ? 4'hf : _GEN_1501; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1503 = 8'hae == _T_107[7:0] ? 4'hf : _GEN_1502; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1504 = 8'haf == _T_107[7:0] ? 4'hf : _GEN_1503; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1505 = 8'hb0 == _T_107[7:0] ? 4'h0 : _GEN_1504; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1506 = 8'hb1 == _T_107[7:0] ? 4'h0 : _GEN_1505; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1507 = 8'hb2 == _T_107[7:0] ? 4'h0 : _GEN_1506; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1508 = 8'hb3 == _T_107[7:0] ? 4'h0 : _GEN_1507; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1509 = 8'hb4 == _T_107[7:0] ? 4'h0 : _GEN_1508; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1510 = 8'hb5 == _T_107[7:0] ? 4'h0 : _GEN_1509; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1511 = 8'hb6 == _T_107[7:0] ? 4'h0 : _GEN_1510; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1512 = 8'hb7 == _T_107[7:0] ? 4'h0 : _GEN_1511; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1513 = 8'hb8 == _T_107[7:0] ? 4'hf : _GEN_1512; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1514 = 8'hb9 == _T_107[7:0] ? 4'hf : _GEN_1513; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1515 = 8'hba == _T_107[7:0] ? 4'hf : _GEN_1514; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1516 = 8'hbb == _T_107[7:0] ? 4'hf : _GEN_1515; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1517 = 8'hbc == _T_107[7:0] ? 4'hf : _GEN_1516; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1518 = 8'hbd == _T_107[7:0] ? 4'hf : _GEN_1517; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1519 = 8'hbe == _T_107[7:0] ? 4'hf : _GEN_1518; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1520 = 8'hbf == _T_107[7:0] ? 4'hf : _GEN_1519; // @[Filter.scala 160:62]
  wire [4:0] _GEN_9878 = {{1'd0}, _GEN_1520}; // @[Filter.scala 160:62]
  wire [8:0] _T_109 = _GEN_9878 * 5'h14; // @[Filter.scala 160:62]
  wire [3:0] _GEN_1617 = 8'h60 == _T_107[7:0] ? 4'hf : 4'h0; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1618 = 8'h61 == _T_107[7:0] ? 4'hf : _GEN_1617; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1619 = 8'h62 == _T_107[7:0] ? 4'hf : _GEN_1618; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1620 = 8'h63 == _T_107[7:0] ? 4'hf : _GEN_1619; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1621 = 8'h64 == _T_107[7:0] ? 4'hf : _GEN_1620; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1622 = 8'h65 == _T_107[7:0] ? 4'hf : _GEN_1621; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1623 = 8'h66 == _T_107[7:0] ? 4'hf : _GEN_1622; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1624 = 8'h67 == _T_107[7:0] ? 4'hf : _GEN_1623; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1625 = 8'h68 == _T_107[7:0] ? 4'hf : _GEN_1624; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1626 = 8'h69 == _T_107[7:0] ? 4'hf : _GEN_1625; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1627 = 8'h6a == _T_107[7:0] ? 4'hf : _GEN_1626; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1628 = 8'h6b == _T_107[7:0] ? 4'hf : _GEN_1627; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1629 = 8'h6c == _T_107[7:0] ? 4'hf : _GEN_1628; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1630 = 8'h6d == _T_107[7:0] ? 4'hf : _GEN_1629; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1631 = 8'h6e == _T_107[7:0] ? 4'hf : _GEN_1630; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1632 = 8'h6f == _T_107[7:0] ? 4'hf : _GEN_1631; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1633 = 8'h70 == _T_107[7:0] ? 4'hf : _GEN_1632; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1634 = 8'h71 == _T_107[7:0] ? 4'hf : _GEN_1633; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1635 = 8'h72 == _T_107[7:0] ? 4'hf : _GEN_1634; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1636 = 8'h73 == _T_107[7:0] ? 4'hf : _GEN_1635; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1637 = 8'h74 == _T_107[7:0] ? 4'hf : _GEN_1636; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1638 = 8'h75 == _T_107[7:0] ? 4'hf : _GEN_1637; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1639 = 8'h76 == _T_107[7:0] ? 4'hf : _GEN_1638; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1640 = 8'h77 == _T_107[7:0] ? 4'hf : _GEN_1639; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1641 = 8'h78 == _T_107[7:0] ? 4'hf : _GEN_1640; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1642 = 8'h79 == _T_107[7:0] ? 4'hf : _GEN_1641; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1643 = 8'h7a == _T_107[7:0] ? 4'hf : _GEN_1642; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1644 = 8'h7b == _T_107[7:0] ? 4'hf : _GEN_1643; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1645 = 8'h7c == _T_107[7:0] ? 4'hf : _GEN_1644; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1646 = 8'h7d == _T_107[7:0] ? 4'hf : _GEN_1645; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1647 = 8'h7e == _T_107[7:0] ? 4'hf : _GEN_1646; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1648 = 8'h7f == _T_107[7:0] ? 4'hf : _GEN_1647; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1649 = 8'h80 == _T_107[7:0] ? 4'hf : _GEN_1648; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1650 = 8'h81 == _T_107[7:0] ? 4'hf : _GEN_1649; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1651 = 8'h82 == _T_107[7:0] ? 4'hf : _GEN_1650; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1652 = 8'h83 == _T_107[7:0] ? 4'hf : _GEN_1651; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1653 = 8'h84 == _T_107[7:0] ? 4'hf : _GEN_1652; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1654 = 8'h85 == _T_107[7:0] ? 4'hf : _GEN_1653; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1655 = 8'h86 == _T_107[7:0] ? 4'hf : _GEN_1654; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1656 = 8'h87 == _T_107[7:0] ? 4'hf : _GEN_1655; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1657 = 8'h88 == _T_107[7:0] ? 4'hf : _GEN_1656; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1658 = 8'h89 == _T_107[7:0] ? 4'hf : _GEN_1657; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1659 = 8'h8a == _T_107[7:0] ? 4'hf : _GEN_1658; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1660 = 8'h8b == _T_107[7:0] ? 4'hf : _GEN_1659; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1661 = 8'h8c == _T_107[7:0] ? 4'hf : _GEN_1660; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1662 = 8'h8d == _T_107[7:0] ? 4'hf : _GEN_1661; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1663 = 8'h8e == _T_107[7:0] ? 4'hf : _GEN_1662; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1664 = 8'h8f == _T_107[7:0] ? 4'hf : _GEN_1663; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1665 = 8'h90 == _T_107[7:0] ? 4'hf : _GEN_1664; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1666 = 8'h91 == _T_107[7:0] ? 4'hf : _GEN_1665; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1667 = 8'h92 == _T_107[7:0] ? 4'hf : _GEN_1666; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1668 = 8'h93 == _T_107[7:0] ? 4'hf : _GEN_1667; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1669 = 8'h94 == _T_107[7:0] ? 4'hf : _GEN_1668; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1670 = 8'h95 == _T_107[7:0] ? 4'hf : _GEN_1669; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1671 = 8'h96 == _T_107[7:0] ? 4'hf : _GEN_1670; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1672 = 8'h97 == _T_107[7:0] ? 4'hf : _GEN_1671; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1673 = 8'h98 == _T_107[7:0] ? 4'hf : _GEN_1672; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1674 = 8'h99 == _T_107[7:0] ? 4'hf : _GEN_1673; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1675 = 8'h9a == _T_107[7:0] ? 4'hf : _GEN_1674; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1676 = 8'h9b == _T_107[7:0] ? 4'hf : _GEN_1675; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1677 = 8'h9c == _T_107[7:0] ? 4'hf : _GEN_1676; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1678 = 8'h9d == _T_107[7:0] ? 4'hf : _GEN_1677; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1679 = 8'h9e == _T_107[7:0] ? 4'hf : _GEN_1678; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1680 = 8'h9f == _T_107[7:0] ? 4'hf : _GEN_1679; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1681 = 8'ha0 == _T_107[7:0] ? 4'hf : _GEN_1680; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1682 = 8'ha1 == _T_107[7:0] ? 4'hf : _GEN_1681; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1683 = 8'ha2 == _T_107[7:0] ? 4'hf : _GEN_1682; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1684 = 8'ha3 == _T_107[7:0] ? 4'hf : _GEN_1683; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1685 = 8'ha4 == _T_107[7:0] ? 4'hf : _GEN_1684; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1686 = 8'ha5 == _T_107[7:0] ? 4'hf : _GEN_1685; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1687 = 8'ha6 == _T_107[7:0] ? 4'hf : _GEN_1686; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1688 = 8'ha7 == _T_107[7:0] ? 4'hf : _GEN_1687; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1689 = 8'ha8 == _T_107[7:0] ? 4'hf : _GEN_1688; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1690 = 8'ha9 == _T_107[7:0] ? 4'hf : _GEN_1689; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1691 = 8'haa == _T_107[7:0] ? 4'hf : _GEN_1690; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1692 = 8'hab == _T_107[7:0] ? 4'hf : _GEN_1691; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1693 = 8'hac == _T_107[7:0] ? 4'hf : _GEN_1692; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1694 = 8'had == _T_107[7:0] ? 4'hf : _GEN_1693; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1695 = 8'hae == _T_107[7:0] ? 4'hf : _GEN_1694; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1696 = 8'haf == _T_107[7:0] ? 4'hf : _GEN_1695; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1697 = 8'hb0 == _T_107[7:0] ? 4'hf : _GEN_1696; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1698 = 8'hb1 == _T_107[7:0] ? 4'hf : _GEN_1697; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1699 = 8'hb2 == _T_107[7:0] ? 4'hf : _GEN_1698; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1700 = 8'hb3 == _T_107[7:0] ? 4'hf : _GEN_1699; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1701 = 8'hb4 == _T_107[7:0] ? 4'hf : _GEN_1700; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1702 = 8'hb5 == _T_107[7:0] ? 4'hf : _GEN_1701; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1703 = 8'hb6 == _T_107[7:0] ? 4'hf : _GEN_1702; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1704 = 8'hb7 == _T_107[7:0] ? 4'hf : _GEN_1703; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1705 = 8'hb8 == _T_107[7:0] ? 4'hf : _GEN_1704; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1706 = 8'hb9 == _T_107[7:0] ? 4'hf : _GEN_1705; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1707 = 8'hba == _T_107[7:0] ? 4'hf : _GEN_1706; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1708 = 8'hbb == _T_107[7:0] ? 4'hf : _GEN_1707; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1709 = 8'hbc == _T_107[7:0] ? 4'hf : _GEN_1708; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1710 = 8'hbd == _T_107[7:0] ? 4'hf : _GEN_1709; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1711 = 8'hbe == _T_107[7:0] ? 4'hf : _GEN_1710; // @[Filter.scala 160:102]
  wire [3:0] _GEN_1712 = 8'hbf == _T_107[7:0] ? 4'hf : _GEN_1711; // @[Filter.scala 160:102]
  wire [6:0] _GEN_9880 = {{3'd0}, _GEN_1712}; // @[Filter.scala 160:102]
  wire [10:0] _T_114 = _GEN_9880 * 7'h46; // @[Filter.scala 160:102]
  wire [10:0] _GEN_9881 = {{2'd0}, _T_109}; // @[Filter.scala 160:69]
  wire [10:0] _T_116 = _GEN_9881 + _T_114; // @[Filter.scala 160:69]
  wire [3:0] _GEN_1721 = 8'h8 == _T_107[7:0] ? 4'hf : 4'h0; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1722 = 8'h9 == _T_107[7:0] ? 4'hf : _GEN_1721; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1723 = 8'ha == _T_107[7:0] ? 4'hf : _GEN_1722; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1724 = 8'hb == _T_107[7:0] ? 4'hf : _GEN_1723; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1725 = 8'hc == _T_107[7:0] ? 4'hf : _GEN_1724; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1726 = 8'hd == _T_107[7:0] ? 4'hf : _GEN_1725; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1727 = 8'he == _T_107[7:0] ? 4'hf : _GEN_1726; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1728 = 8'hf == _T_107[7:0] ? 4'hf : _GEN_1727; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1729 = 8'h10 == _T_107[7:0] ? 4'h0 : _GEN_1728; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1730 = 8'h11 == _T_107[7:0] ? 4'h0 : _GEN_1729; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1731 = 8'h12 == _T_107[7:0] ? 4'h0 : _GEN_1730; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1732 = 8'h13 == _T_107[7:0] ? 4'h0 : _GEN_1731; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1733 = 8'h14 == _T_107[7:0] ? 4'h0 : _GEN_1732; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1734 = 8'h15 == _T_107[7:0] ? 4'h0 : _GEN_1733; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1735 = 8'h16 == _T_107[7:0] ? 4'h0 : _GEN_1734; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1736 = 8'h17 == _T_107[7:0] ? 4'h0 : _GEN_1735; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1737 = 8'h18 == _T_107[7:0] ? 4'hf : _GEN_1736; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1738 = 8'h19 == _T_107[7:0] ? 4'hf : _GEN_1737; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1739 = 8'h1a == _T_107[7:0] ? 4'hf : _GEN_1738; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1740 = 8'h1b == _T_107[7:0] ? 4'hf : _GEN_1739; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1741 = 8'h1c == _T_107[7:0] ? 4'hf : _GEN_1740; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1742 = 8'h1d == _T_107[7:0] ? 4'hf : _GEN_1741; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1743 = 8'h1e == _T_107[7:0] ? 4'hf : _GEN_1742; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1744 = 8'h1f == _T_107[7:0] ? 4'hf : _GEN_1743; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1745 = 8'h20 == _T_107[7:0] ? 4'h0 : _GEN_1744; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1746 = 8'h21 == _T_107[7:0] ? 4'h0 : _GEN_1745; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1747 = 8'h22 == _T_107[7:0] ? 4'h0 : _GEN_1746; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1748 = 8'h23 == _T_107[7:0] ? 4'h0 : _GEN_1747; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1749 = 8'h24 == _T_107[7:0] ? 4'h0 : _GEN_1748; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1750 = 8'h25 == _T_107[7:0] ? 4'h0 : _GEN_1749; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1751 = 8'h26 == _T_107[7:0] ? 4'h0 : _GEN_1750; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1752 = 8'h27 == _T_107[7:0] ? 4'h0 : _GEN_1751; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1753 = 8'h28 == _T_107[7:0] ? 4'hf : _GEN_1752; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1754 = 8'h29 == _T_107[7:0] ? 4'hf : _GEN_1753; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1755 = 8'h2a == _T_107[7:0] ? 4'hf : _GEN_1754; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1756 = 8'h2b == _T_107[7:0] ? 4'hf : _GEN_1755; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1757 = 8'h2c == _T_107[7:0] ? 4'hf : _GEN_1756; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1758 = 8'h2d == _T_107[7:0] ? 4'hf : _GEN_1757; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1759 = 8'h2e == _T_107[7:0] ? 4'hf : _GEN_1758; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1760 = 8'h2f == _T_107[7:0] ? 4'hf : _GEN_1759; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1761 = 8'h30 == _T_107[7:0] ? 4'h0 : _GEN_1760; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1762 = 8'h31 == _T_107[7:0] ? 4'h0 : _GEN_1761; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1763 = 8'h32 == _T_107[7:0] ? 4'h0 : _GEN_1762; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1764 = 8'h33 == _T_107[7:0] ? 4'h0 : _GEN_1763; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1765 = 8'h34 == _T_107[7:0] ? 4'h0 : _GEN_1764; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1766 = 8'h35 == _T_107[7:0] ? 4'h0 : _GEN_1765; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1767 = 8'h36 == _T_107[7:0] ? 4'h0 : _GEN_1766; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1768 = 8'h37 == _T_107[7:0] ? 4'h0 : _GEN_1767; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1769 = 8'h38 == _T_107[7:0] ? 4'hf : _GEN_1768; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1770 = 8'h39 == _T_107[7:0] ? 4'hf : _GEN_1769; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1771 = 8'h3a == _T_107[7:0] ? 4'hf : _GEN_1770; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1772 = 8'h3b == _T_107[7:0] ? 4'hf : _GEN_1771; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1773 = 8'h3c == _T_107[7:0] ? 4'hf : _GEN_1772; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1774 = 8'h3d == _T_107[7:0] ? 4'hf : _GEN_1773; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1775 = 8'h3e == _T_107[7:0] ? 4'hf : _GEN_1774; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1776 = 8'h3f == _T_107[7:0] ? 4'hf : _GEN_1775; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1777 = 8'h40 == _T_107[7:0] ? 4'h0 : _GEN_1776; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1778 = 8'h41 == _T_107[7:0] ? 4'h0 : _GEN_1777; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1779 = 8'h42 == _T_107[7:0] ? 4'h0 : _GEN_1778; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1780 = 8'h43 == _T_107[7:0] ? 4'h0 : _GEN_1779; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1781 = 8'h44 == _T_107[7:0] ? 4'h0 : _GEN_1780; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1782 = 8'h45 == _T_107[7:0] ? 4'h0 : _GEN_1781; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1783 = 8'h46 == _T_107[7:0] ? 4'h0 : _GEN_1782; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1784 = 8'h47 == _T_107[7:0] ? 4'h0 : _GEN_1783; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1785 = 8'h48 == _T_107[7:0] ? 4'hf : _GEN_1784; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1786 = 8'h49 == _T_107[7:0] ? 4'hf : _GEN_1785; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1787 = 8'h4a == _T_107[7:0] ? 4'hf : _GEN_1786; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1788 = 8'h4b == _T_107[7:0] ? 4'hf : _GEN_1787; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1789 = 8'h4c == _T_107[7:0] ? 4'hf : _GEN_1788; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1790 = 8'h4d == _T_107[7:0] ? 4'hf : _GEN_1789; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1791 = 8'h4e == _T_107[7:0] ? 4'hf : _GEN_1790; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1792 = 8'h4f == _T_107[7:0] ? 4'hf : _GEN_1791; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1793 = 8'h50 == _T_107[7:0] ? 4'h0 : _GEN_1792; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1794 = 8'h51 == _T_107[7:0] ? 4'h0 : _GEN_1793; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1795 = 8'h52 == _T_107[7:0] ? 4'h0 : _GEN_1794; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1796 = 8'h53 == _T_107[7:0] ? 4'h0 : _GEN_1795; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1797 = 8'h54 == _T_107[7:0] ? 4'h0 : _GEN_1796; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1798 = 8'h55 == _T_107[7:0] ? 4'h0 : _GEN_1797; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1799 = 8'h56 == _T_107[7:0] ? 4'h0 : _GEN_1798; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1800 = 8'h57 == _T_107[7:0] ? 4'h0 : _GEN_1799; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1801 = 8'h58 == _T_107[7:0] ? 4'hf : _GEN_1800; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1802 = 8'h59 == _T_107[7:0] ? 4'hf : _GEN_1801; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1803 = 8'h5a == _T_107[7:0] ? 4'hf : _GEN_1802; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1804 = 8'h5b == _T_107[7:0] ? 4'hf : _GEN_1803; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1805 = 8'h5c == _T_107[7:0] ? 4'hf : _GEN_1804; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1806 = 8'h5d == _T_107[7:0] ? 4'hf : _GEN_1805; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1807 = 8'h5e == _T_107[7:0] ? 4'hf : _GEN_1806; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1808 = 8'h5f == _T_107[7:0] ? 4'hf : _GEN_1807; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1809 = 8'h60 == _T_107[7:0] ? 4'h0 : _GEN_1808; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1810 = 8'h61 == _T_107[7:0] ? 4'h0 : _GEN_1809; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1811 = 8'h62 == _T_107[7:0] ? 4'h0 : _GEN_1810; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1812 = 8'h63 == _T_107[7:0] ? 4'h0 : _GEN_1811; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1813 = 8'h64 == _T_107[7:0] ? 4'h0 : _GEN_1812; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1814 = 8'h65 == _T_107[7:0] ? 4'h0 : _GEN_1813; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1815 = 8'h66 == _T_107[7:0] ? 4'h0 : _GEN_1814; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1816 = 8'h67 == _T_107[7:0] ? 4'h0 : _GEN_1815; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1817 = 8'h68 == _T_107[7:0] ? 4'hf : _GEN_1816; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1818 = 8'h69 == _T_107[7:0] ? 4'hf : _GEN_1817; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1819 = 8'h6a == _T_107[7:0] ? 4'hf : _GEN_1818; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1820 = 8'h6b == _T_107[7:0] ? 4'hf : _GEN_1819; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1821 = 8'h6c == _T_107[7:0] ? 4'hf : _GEN_1820; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1822 = 8'h6d == _T_107[7:0] ? 4'hf : _GEN_1821; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1823 = 8'h6e == _T_107[7:0] ? 4'hf : _GEN_1822; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1824 = 8'h6f == _T_107[7:0] ? 4'hf : _GEN_1823; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1825 = 8'h70 == _T_107[7:0] ? 4'h0 : _GEN_1824; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1826 = 8'h71 == _T_107[7:0] ? 4'h0 : _GEN_1825; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1827 = 8'h72 == _T_107[7:0] ? 4'h0 : _GEN_1826; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1828 = 8'h73 == _T_107[7:0] ? 4'h0 : _GEN_1827; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1829 = 8'h74 == _T_107[7:0] ? 4'h0 : _GEN_1828; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1830 = 8'h75 == _T_107[7:0] ? 4'h0 : _GEN_1829; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1831 = 8'h76 == _T_107[7:0] ? 4'h0 : _GEN_1830; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1832 = 8'h77 == _T_107[7:0] ? 4'h0 : _GEN_1831; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1833 = 8'h78 == _T_107[7:0] ? 4'hf : _GEN_1832; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1834 = 8'h79 == _T_107[7:0] ? 4'hf : _GEN_1833; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1835 = 8'h7a == _T_107[7:0] ? 4'hf : _GEN_1834; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1836 = 8'h7b == _T_107[7:0] ? 4'hf : _GEN_1835; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1837 = 8'h7c == _T_107[7:0] ? 4'hf : _GEN_1836; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1838 = 8'h7d == _T_107[7:0] ? 4'hf : _GEN_1837; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1839 = 8'h7e == _T_107[7:0] ? 4'hf : _GEN_1838; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1840 = 8'h7f == _T_107[7:0] ? 4'hf : _GEN_1839; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1841 = 8'h80 == _T_107[7:0] ? 4'h0 : _GEN_1840; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1842 = 8'h81 == _T_107[7:0] ? 4'h0 : _GEN_1841; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1843 = 8'h82 == _T_107[7:0] ? 4'h0 : _GEN_1842; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1844 = 8'h83 == _T_107[7:0] ? 4'h0 : _GEN_1843; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1845 = 8'h84 == _T_107[7:0] ? 4'h0 : _GEN_1844; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1846 = 8'h85 == _T_107[7:0] ? 4'h0 : _GEN_1845; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1847 = 8'h86 == _T_107[7:0] ? 4'h0 : _GEN_1846; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1848 = 8'h87 == _T_107[7:0] ? 4'h0 : _GEN_1847; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1849 = 8'h88 == _T_107[7:0] ? 4'hf : _GEN_1848; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1850 = 8'h89 == _T_107[7:0] ? 4'hf : _GEN_1849; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1851 = 8'h8a == _T_107[7:0] ? 4'hf : _GEN_1850; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1852 = 8'h8b == _T_107[7:0] ? 4'hf : _GEN_1851; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1853 = 8'h8c == _T_107[7:0] ? 4'hf : _GEN_1852; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1854 = 8'h8d == _T_107[7:0] ? 4'hf : _GEN_1853; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1855 = 8'h8e == _T_107[7:0] ? 4'hf : _GEN_1854; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1856 = 8'h8f == _T_107[7:0] ? 4'hf : _GEN_1855; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1857 = 8'h90 == _T_107[7:0] ? 4'h0 : _GEN_1856; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1858 = 8'h91 == _T_107[7:0] ? 4'h0 : _GEN_1857; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1859 = 8'h92 == _T_107[7:0] ? 4'h0 : _GEN_1858; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1860 = 8'h93 == _T_107[7:0] ? 4'h0 : _GEN_1859; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1861 = 8'h94 == _T_107[7:0] ? 4'h0 : _GEN_1860; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1862 = 8'h95 == _T_107[7:0] ? 4'h0 : _GEN_1861; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1863 = 8'h96 == _T_107[7:0] ? 4'h0 : _GEN_1862; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1864 = 8'h97 == _T_107[7:0] ? 4'h0 : _GEN_1863; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1865 = 8'h98 == _T_107[7:0] ? 4'hf : _GEN_1864; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1866 = 8'h99 == _T_107[7:0] ? 4'hf : _GEN_1865; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1867 = 8'h9a == _T_107[7:0] ? 4'hf : _GEN_1866; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1868 = 8'h9b == _T_107[7:0] ? 4'hf : _GEN_1867; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1869 = 8'h9c == _T_107[7:0] ? 4'hf : _GEN_1868; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1870 = 8'h9d == _T_107[7:0] ? 4'hf : _GEN_1869; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1871 = 8'h9e == _T_107[7:0] ? 4'hf : _GEN_1870; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1872 = 8'h9f == _T_107[7:0] ? 4'hf : _GEN_1871; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1873 = 8'ha0 == _T_107[7:0] ? 4'h0 : _GEN_1872; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1874 = 8'ha1 == _T_107[7:0] ? 4'h0 : _GEN_1873; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1875 = 8'ha2 == _T_107[7:0] ? 4'h0 : _GEN_1874; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1876 = 8'ha3 == _T_107[7:0] ? 4'h0 : _GEN_1875; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1877 = 8'ha4 == _T_107[7:0] ? 4'h0 : _GEN_1876; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1878 = 8'ha5 == _T_107[7:0] ? 4'h0 : _GEN_1877; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1879 = 8'ha6 == _T_107[7:0] ? 4'h0 : _GEN_1878; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1880 = 8'ha7 == _T_107[7:0] ? 4'h0 : _GEN_1879; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1881 = 8'ha8 == _T_107[7:0] ? 4'hf : _GEN_1880; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1882 = 8'ha9 == _T_107[7:0] ? 4'hf : _GEN_1881; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1883 = 8'haa == _T_107[7:0] ? 4'hf : _GEN_1882; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1884 = 8'hab == _T_107[7:0] ? 4'hf : _GEN_1883; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1885 = 8'hac == _T_107[7:0] ? 4'hf : _GEN_1884; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1886 = 8'had == _T_107[7:0] ? 4'hf : _GEN_1885; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1887 = 8'hae == _T_107[7:0] ? 4'hf : _GEN_1886; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1888 = 8'haf == _T_107[7:0] ? 4'hf : _GEN_1887; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1889 = 8'hb0 == _T_107[7:0] ? 4'h0 : _GEN_1888; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1890 = 8'hb1 == _T_107[7:0] ? 4'h0 : _GEN_1889; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1891 = 8'hb2 == _T_107[7:0] ? 4'h0 : _GEN_1890; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1892 = 8'hb3 == _T_107[7:0] ? 4'h0 : _GEN_1891; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1893 = 8'hb4 == _T_107[7:0] ? 4'h0 : _GEN_1892; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1894 = 8'hb5 == _T_107[7:0] ? 4'h0 : _GEN_1893; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1895 = 8'hb6 == _T_107[7:0] ? 4'h0 : _GEN_1894; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1896 = 8'hb7 == _T_107[7:0] ? 4'h0 : _GEN_1895; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1897 = 8'hb8 == _T_107[7:0] ? 4'hf : _GEN_1896; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1898 = 8'hb9 == _T_107[7:0] ? 4'hf : _GEN_1897; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1899 = 8'hba == _T_107[7:0] ? 4'hf : _GEN_1898; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1900 = 8'hbb == _T_107[7:0] ? 4'hf : _GEN_1899; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1901 = 8'hbc == _T_107[7:0] ? 4'hf : _GEN_1900; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1902 = 8'hbd == _T_107[7:0] ? 4'hf : _GEN_1901; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1903 = 8'hbe == _T_107[7:0] ? 4'hf : _GEN_1902; // @[Filter.scala 160:142]
  wire [3:0] _GEN_1904 = 8'hbf == _T_107[7:0] ? 4'hf : _GEN_1903; // @[Filter.scala 160:142]
  wire [7:0] _T_121 = _GEN_1904 * 4'ha; // @[Filter.scala 160:142]
  wire [10:0] _GEN_9883 = {{3'd0}, _T_121}; // @[Filter.scala 160:109]
  wire [10:0] _T_123 = _T_116 + _GEN_9883; // @[Filter.scala 160:109]
  wire [10:0] _T_124 = _T_123 / 11'h64; // @[Filter.scala 160:150]
  wire  _T_126 = _T_97 >= 5'h10; // @[Filter.scala 163:31]
  wire  _T_130 = _T_104 >= 32'hc; // @[Filter.scala 163:63]
  wire  _T_131 = _T_126 | _T_130; // @[Filter.scala 163:58]
  wire [10:0] _GEN_2097 = io_SPI_distort ? _T_124 : {{7'd0}, _GEN_1520}; // @[Filter.scala 165:35]
  wire [10:0] _GEN_2098 = _T_131 ? 11'h0 : _GEN_2097; // @[Filter.scala 163:80]
  wire [10:0] _GEN_2291 = io_SPI_distort ? _T_124 : {{7'd0}, _GEN_1712}; // @[Filter.scala 165:35]
  wire [10:0] _GEN_2292 = _T_131 ? 11'h0 : _GEN_2291; // @[Filter.scala 163:80]
  wire [10:0] _GEN_2485 = io_SPI_distort ? _T_124 : {{7'd0}, _GEN_1904}; // @[Filter.scala 165:35]
  wire [10:0] _GEN_2486 = _T_131 ? 11'h0 : _GEN_2485; // @[Filter.scala 163:80]
  wire [31:0] _T_159 = pixelIndex + 32'h2; // @[Filter.scala 158:31]
  wire [31:0] _GEN_2 = _T_159 % 32'h10; // @[Filter.scala 158:38]
  wire [4:0] _T_160 = _GEN_2[4:0]; // @[Filter.scala 158:38]
  wire [4:0] _T_162 = _T_160 + _GEN_9863; // @[Filter.scala 158:53]
  wire [4:0] _T_164 = _T_162 - 5'h1; // @[Filter.scala 158:69]
  wire [31:0] _T_167 = _T_159 / 32'h10; // @[Filter.scala 159:38]
  wire [31:0] _T_169 = _T_167 + _GEN_9864; // @[Filter.scala 159:53]
  wire [31:0] _T_171 = _T_169 - 32'h1; // @[Filter.scala 159:69]
  wire [36:0] _T_172 = _T_171 * 32'h10; // @[Filter.scala 160:42]
  wire [36:0] _GEN_9889 = {{32'd0}, _T_164}; // @[Filter.scala 160:57]
  wire [36:0] _T_174 = _T_172 + _GEN_9889; // @[Filter.scala 160:57]
  wire [3:0] _GEN_2495 = 8'h8 == _T_174[7:0] ? 4'h0 : 4'hf; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2496 = 8'h9 == _T_174[7:0] ? 4'h0 : _GEN_2495; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2497 = 8'ha == _T_174[7:0] ? 4'h0 : _GEN_2496; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2498 = 8'hb == _T_174[7:0] ? 4'h0 : _GEN_2497; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2499 = 8'hc == _T_174[7:0] ? 4'h0 : _GEN_2498; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2500 = 8'hd == _T_174[7:0] ? 4'h0 : _GEN_2499; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2501 = 8'he == _T_174[7:0] ? 4'h0 : _GEN_2500; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2502 = 8'hf == _T_174[7:0] ? 4'h0 : _GEN_2501; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2503 = 8'h10 == _T_174[7:0] ? 4'hf : _GEN_2502; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2504 = 8'h11 == _T_174[7:0] ? 4'hf : _GEN_2503; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2505 = 8'h12 == _T_174[7:0] ? 4'hf : _GEN_2504; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2506 = 8'h13 == _T_174[7:0] ? 4'hf : _GEN_2505; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2507 = 8'h14 == _T_174[7:0] ? 4'hf : _GEN_2506; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2508 = 8'h15 == _T_174[7:0] ? 4'hf : _GEN_2507; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2509 = 8'h16 == _T_174[7:0] ? 4'hf : _GEN_2508; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2510 = 8'h17 == _T_174[7:0] ? 4'hf : _GEN_2509; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2511 = 8'h18 == _T_174[7:0] ? 4'h0 : _GEN_2510; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2512 = 8'h19 == _T_174[7:0] ? 4'h0 : _GEN_2511; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2513 = 8'h1a == _T_174[7:0] ? 4'h0 : _GEN_2512; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2514 = 8'h1b == _T_174[7:0] ? 4'h0 : _GEN_2513; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2515 = 8'h1c == _T_174[7:0] ? 4'h0 : _GEN_2514; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2516 = 8'h1d == _T_174[7:0] ? 4'h0 : _GEN_2515; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2517 = 8'h1e == _T_174[7:0] ? 4'h0 : _GEN_2516; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2518 = 8'h1f == _T_174[7:0] ? 4'h0 : _GEN_2517; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2519 = 8'h20 == _T_174[7:0] ? 4'hf : _GEN_2518; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2520 = 8'h21 == _T_174[7:0] ? 4'hf : _GEN_2519; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2521 = 8'h22 == _T_174[7:0] ? 4'hf : _GEN_2520; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2522 = 8'h23 == _T_174[7:0] ? 4'hf : _GEN_2521; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2523 = 8'h24 == _T_174[7:0] ? 4'hf : _GEN_2522; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2524 = 8'h25 == _T_174[7:0] ? 4'hf : _GEN_2523; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2525 = 8'h26 == _T_174[7:0] ? 4'hf : _GEN_2524; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2526 = 8'h27 == _T_174[7:0] ? 4'hf : _GEN_2525; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2527 = 8'h28 == _T_174[7:0] ? 4'h0 : _GEN_2526; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2528 = 8'h29 == _T_174[7:0] ? 4'h0 : _GEN_2527; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2529 = 8'h2a == _T_174[7:0] ? 4'h0 : _GEN_2528; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2530 = 8'h2b == _T_174[7:0] ? 4'h0 : _GEN_2529; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2531 = 8'h2c == _T_174[7:0] ? 4'h0 : _GEN_2530; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2532 = 8'h2d == _T_174[7:0] ? 4'h0 : _GEN_2531; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2533 = 8'h2e == _T_174[7:0] ? 4'h0 : _GEN_2532; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2534 = 8'h2f == _T_174[7:0] ? 4'h0 : _GEN_2533; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2535 = 8'h30 == _T_174[7:0] ? 4'hf : _GEN_2534; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2536 = 8'h31 == _T_174[7:0] ? 4'hf : _GEN_2535; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2537 = 8'h32 == _T_174[7:0] ? 4'hf : _GEN_2536; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2538 = 8'h33 == _T_174[7:0] ? 4'hf : _GEN_2537; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2539 = 8'h34 == _T_174[7:0] ? 4'hf : _GEN_2538; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2540 = 8'h35 == _T_174[7:0] ? 4'hf : _GEN_2539; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2541 = 8'h36 == _T_174[7:0] ? 4'hf : _GEN_2540; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2542 = 8'h37 == _T_174[7:0] ? 4'hf : _GEN_2541; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2543 = 8'h38 == _T_174[7:0] ? 4'h0 : _GEN_2542; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2544 = 8'h39 == _T_174[7:0] ? 4'h0 : _GEN_2543; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2545 = 8'h3a == _T_174[7:0] ? 4'h0 : _GEN_2544; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2546 = 8'h3b == _T_174[7:0] ? 4'h0 : _GEN_2545; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2547 = 8'h3c == _T_174[7:0] ? 4'h0 : _GEN_2546; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2548 = 8'h3d == _T_174[7:0] ? 4'h0 : _GEN_2547; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2549 = 8'h3e == _T_174[7:0] ? 4'h0 : _GEN_2548; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2550 = 8'h3f == _T_174[7:0] ? 4'h0 : _GEN_2549; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2551 = 8'h40 == _T_174[7:0] ? 4'hf : _GEN_2550; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2552 = 8'h41 == _T_174[7:0] ? 4'hf : _GEN_2551; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2553 = 8'h42 == _T_174[7:0] ? 4'hf : _GEN_2552; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2554 = 8'h43 == _T_174[7:0] ? 4'hf : _GEN_2553; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2555 = 8'h44 == _T_174[7:0] ? 4'hf : _GEN_2554; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2556 = 8'h45 == _T_174[7:0] ? 4'hf : _GEN_2555; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2557 = 8'h46 == _T_174[7:0] ? 4'hf : _GEN_2556; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2558 = 8'h47 == _T_174[7:0] ? 4'hf : _GEN_2557; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2559 = 8'h48 == _T_174[7:0] ? 4'h0 : _GEN_2558; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2560 = 8'h49 == _T_174[7:0] ? 4'h0 : _GEN_2559; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2561 = 8'h4a == _T_174[7:0] ? 4'h0 : _GEN_2560; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2562 = 8'h4b == _T_174[7:0] ? 4'h0 : _GEN_2561; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2563 = 8'h4c == _T_174[7:0] ? 4'h0 : _GEN_2562; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2564 = 8'h4d == _T_174[7:0] ? 4'h0 : _GEN_2563; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2565 = 8'h4e == _T_174[7:0] ? 4'h0 : _GEN_2564; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2566 = 8'h4f == _T_174[7:0] ? 4'h0 : _GEN_2565; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2567 = 8'h50 == _T_174[7:0] ? 4'hf : _GEN_2566; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2568 = 8'h51 == _T_174[7:0] ? 4'hf : _GEN_2567; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2569 = 8'h52 == _T_174[7:0] ? 4'hf : _GEN_2568; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2570 = 8'h53 == _T_174[7:0] ? 4'hf : _GEN_2569; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2571 = 8'h54 == _T_174[7:0] ? 4'hf : _GEN_2570; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2572 = 8'h55 == _T_174[7:0] ? 4'hf : _GEN_2571; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2573 = 8'h56 == _T_174[7:0] ? 4'hf : _GEN_2572; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2574 = 8'h57 == _T_174[7:0] ? 4'hf : _GEN_2573; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2575 = 8'h58 == _T_174[7:0] ? 4'h0 : _GEN_2574; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2576 = 8'h59 == _T_174[7:0] ? 4'h0 : _GEN_2575; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2577 = 8'h5a == _T_174[7:0] ? 4'h0 : _GEN_2576; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2578 = 8'h5b == _T_174[7:0] ? 4'h0 : _GEN_2577; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2579 = 8'h5c == _T_174[7:0] ? 4'h0 : _GEN_2578; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2580 = 8'h5d == _T_174[7:0] ? 4'h0 : _GEN_2579; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2581 = 8'h5e == _T_174[7:0] ? 4'h0 : _GEN_2580; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2582 = 8'h5f == _T_174[7:0] ? 4'h0 : _GEN_2581; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2583 = 8'h60 == _T_174[7:0] ? 4'h0 : _GEN_2582; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2584 = 8'h61 == _T_174[7:0] ? 4'h0 : _GEN_2583; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2585 = 8'h62 == _T_174[7:0] ? 4'h0 : _GEN_2584; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2586 = 8'h63 == _T_174[7:0] ? 4'h0 : _GEN_2585; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2587 = 8'h64 == _T_174[7:0] ? 4'h0 : _GEN_2586; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2588 = 8'h65 == _T_174[7:0] ? 4'h0 : _GEN_2587; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2589 = 8'h66 == _T_174[7:0] ? 4'h0 : _GEN_2588; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2590 = 8'h67 == _T_174[7:0] ? 4'h0 : _GEN_2589; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2591 = 8'h68 == _T_174[7:0] ? 4'hf : _GEN_2590; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2592 = 8'h69 == _T_174[7:0] ? 4'hf : _GEN_2591; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2593 = 8'h6a == _T_174[7:0] ? 4'hf : _GEN_2592; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2594 = 8'h6b == _T_174[7:0] ? 4'hf : _GEN_2593; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2595 = 8'h6c == _T_174[7:0] ? 4'hf : _GEN_2594; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2596 = 8'h6d == _T_174[7:0] ? 4'hf : _GEN_2595; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2597 = 8'h6e == _T_174[7:0] ? 4'hf : _GEN_2596; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2598 = 8'h6f == _T_174[7:0] ? 4'hf : _GEN_2597; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2599 = 8'h70 == _T_174[7:0] ? 4'h0 : _GEN_2598; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2600 = 8'h71 == _T_174[7:0] ? 4'h0 : _GEN_2599; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2601 = 8'h72 == _T_174[7:0] ? 4'h0 : _GEN_2600; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2602 = 8'h73 == _T_174[7:0] ? 4'h0 : _GEN_2601; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2603 = 8'h74 == _T_174[7:0] ? 4'h0 : _GEN_2602; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2604 = 8'h75 == _T_174[7:0] ? 4'h0 : _GEN_2603; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2605 = 8'h76 == _T_174[7:0] ? 4'h0 : _GEN_2604; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2606 = 8'h77 == _T_174[7:0] ? 4'h0 : _GEN_2605; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2607 = 8'h78 == _T_174[7:0] ? 4'hf : _GEN_2606; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2608 = 8'h79 == _T_174[7:0] ? 4'hf : _GEN_2607; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2609 = 8'h7a == _T_174[7:0] ? 4'hf : _GEN_2608; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2610 = 8'h7b == _T_174[7:0] ? 4'hf : _GEN_2609; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2611 = 8'h7c == _T_174[7:0] ? 4'hf : _GEN_2610; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2612 = 8'h7d == _T_174[7:0] ? 4'hf : _GEN_2611; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2613 = 8'h7e == _T_174[7:0] ? 4'hf : _GEN_2612; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2614 = 8'h7f == _T_174[7:0] ? 4'hf : _GEN_2613; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2615 = 8'h80 == _T_174[7:0] ? 4'h0 : _GEN_2614; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2616 = 8'h81 == _T_174[7:0] ? 4'h0 : _GEN_2615; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2617 = 8'h82 == _T_174[7:0] ? 4'h0 : _GEN_2616; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2618 = 8'h83 == _T_174[7:0] ? 4'h0 : _GEN_2617; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2619 = 8'h84 == _T_174[7:0] ? 4'h0 : _GEN_2618; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2620 = 8'h85 == _T_174[7:0] ? 4'h0 : _GEN_2619; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2621 = 8'h86 == _T_174[7:0] ? 4'h0 : _GEN_2620; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2622 = 8'h87 == _T_174[7:0] ? 4'h0 : _GEN_2621; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2623 = 8'h88 == _T_174[7:0] ? 4'hf : _GEN_2622; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2624 = 8'h89 == _T_174[7:0] ? 4'hf : _GEN_2623; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2625 = 8'h8a == _T_174[7:0] ? 4'hf : _GEN_2624; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2626 = 8'h8b == _T_174[7:0] ? 4'hf : _GEN_2625; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2627 = 8'h8c == _T_174[7:0] ? 4'hf : _GEN_2626; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2628 = 8'h8d == _T_174[7:0] ? 4'hf : _GEN_2627; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2629 = 8'h8e == _T_174[7:0] ? 4'hf : _GEN_2628; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2630 = 8'h8f == _T_174[7:0] ? 4'hf : _GEN_2629; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2631 = 8'h90 == _T_174[7:0] ? 4'h0 : _GEN_2630; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2632 = 8'h91 == _T_174[7:0] ? 4'h0 : _GEN_2631; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2633 = 8'h92 == _T_174[7:0] ? 4'h0 : _GEN_2632; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2634 = 8'h93 == _T_174[7:0] ? 4'h0 : _GEN_2633; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2635 = 8'h94 == _T_174[7:0] ? 4'h0 : _GEN_2634; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2636 = 8'h95 == _T_174[7:0] ? 4'h0 : _GEN_2635; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2637 = 8'h96 == _T_174[7:0] ? 4'h0 : _GEN_2636; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2638 = 8'h97 == _T_174[7:0] ? 4'h0 : _GEN_2637; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2639 = 8'h98 == _T_174[7:0] ? 4'hf : _GEN_2638; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2640 = 8'h99 == _T_174[7:0] ? 4'hf : _GEN_2639; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2641 = 8'h9a == _T_174[7:0] ? 4'hf : _GEN_2640; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2642 = 8'h9b == _T_174[7:0] ? 4'hf : _GEN_2641; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2643 = 8'h9c == _T_174[7:0] ? 4'hf : _GEN_2642; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2644 = 8'h9d == _T_174[7:0] ? 4'hf : _GEN_2643; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2645 = 8'h9e == _T_174[7:0] ? 4'hf : _GEN_2644; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2646 = 8'h9f == _T_174[7:0] ? 4'hf : _GEN_2645; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2647 = 8'ha0 == _T_174[7:0] ? 4'h0 : _GEN_2646; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2648 = 8'ha1 == _T_174[7:0] ? 4'h0 : _GEN_2647; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2649 = 8'ha2 == _T_174[7:0] ? 4'h0 : _GEN_2648; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2650 = 8'ha3 == _T_174[7:0] ? 4'h0 : _GEN_2649; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2651 = 8'ha4 == _T_174[7:0] ? 4'h0 : _GEN_2650; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2652 = 8'ha5 == _T_174[7:0] ? 4'h0 : _GEN_2651; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2653 = 8'ha6 == _T_174[7:0] ? 4'h0 : _GEN_2652; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2654 = 8'ha7 == _T_174[7:0] ? 4'h0 : _GEN_2653; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2655 = 8'ha8 == _T_174[7:0] ? 4'hf : _GEN_2654; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2656 = 8'ha9 == _T_174[7:0] ? 4'hf : _GEN_2655; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2657 = 8'haa == _T_174[7:0] ? 4'hf : _GEN_2656; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2658 = 8'hab == _T_174[7:0] ? 4'hf : _GEN_2657; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2659 = 8'hac == _T_174[7:0] ? 4'hf : _GEN_2658; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2660 = 8'had == _T_174[7:0] ? 4'hf : _GEN_2659; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2661 = 8'hae == _T_174[7:0] ? 4'hf : _GEN_2660; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2662 = 8'haf == _T_174[7:0] ? 4'hf : _GEN_2661; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2663 = 8'hb0 == _T_174[7:0] ? 4'h0 : _GEN_2662; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2664 = 8'hb1 == _T_174[7:0] ? 4'h0 : _GEN_2663; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2665 = 8'hb2 == _T_174[7:0] ? 4'h0 : _GEN_2664; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2666 = 8'hb3 == _T_174[7:0] ? 4'h0 : _GEN_2665; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2667 = 8'hb4 == _T_174[7:0] ? 4'h0 : _GEN_2666; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2668 = 8'hb5 == _T_174[7:0] ? 4'h0 : _GEN_2667; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2669 = 8'hb6 == _T_174[7:0] ? 4'h0 : _GEN_2668; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2670 = 8'hb7 == _T_174[7:0] ? 4'h0 : _GEN_2669; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2671 = 8'hb8 == _T_174[7:0] ? 4'hf : _GEN_2670; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2672 = 8'hb9 == _T_174[7:0] ? 4'hf : _GEN_2671; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2673 = 8'hba == _T_174[7:0] ? 4'hf : _GEN_2672; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2674 = 8'hbb == _T_174[7:0] ? 4'hf : _GEN_2673; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2675 = 8'hbc == _T_174[7:0] ? 4'hf : _GEN_2674; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2676 = 8'hbd == _T_174[7:0] ? 4'hf : _GEN_2675; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2677 = 8'hbe == _T_174[7:0] ? 4'hf : _GEN_2676; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2678 = 8'hbf == _T_174[7:0] ? 4'hf : _GEN_2677; // @[Filter.scala 160:62]
  wire [4:0] _GEN_9890 = {{1'd0}, _GEN_2678}; // @[Filter.scala 160:62]
  wire [8:0] _T_176 = _GEN_9890 * 5'h14; // @[Filter.scala 160:62]
  wire [3:0] _GEN_2775 = 8'h60 == _T_174[7:0] ? 4'hf : 4'h0; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2776 = 8'h61 == _T_174[7:0] ? 4'hf : _GEN_2775; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2777 = 8'h62 == _T_174[7:0] ? 4'hf : _GEN_2776; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2778 = 8'h63 == _T_174[7:0] ? 4'hf : _GEN_2777; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2779 = 8'h64 == _T_174[7:0] ? 4'hf : _GEN_2778; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2780 = 8'h65 == _T_174[7:0] ? 4'hf : _GEN_2779; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2781 = 8'h66 == _T_174[7:0] ? 4'hf : _GEN_2780; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2782 = 8'h67 == _T_174[7:0] ? 4'hf : _GEN_2781; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2783 = 8'h68 == _T_174[7:0] ? 4'hf : _GEN_2782; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2784 = 8'h69 == _T_174[7:0] ? 4'hf : _GEN_2783; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2785 = 8'h6a == _T_174[7:0] ? 4'hf : _GEN_2784; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2786 = 8'h6b == _T_174[7:0] ? 4'hf : _GEN_2785; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2787 = 8'h6c == _T_174[7:0] ? 4'hf : _GEN_2786; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2788 = 8'h6d == _T_174[7:0] ? 4'hf : _GEN_2787; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2789 = 8'h6e == _T_174[7:0] ? 4'hf : _GEN_2788; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2790 = 8'h6f == _T_174[7:0] ? 4'hf : _GEN_2789; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2791 = 8'h70 == _T_174[7:0] ? 4'hf : _GEN_2790; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2792 = 8'h71 == _T_174[7:0] ? 4'hf : _GEN_2791; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2793 = 8'h72 == _T_174[7:0] ? 4'hf : _GEN_2792; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2794 = 8'h73 == _T_174[7:0] ? 4'hf : _GEN_2793; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2795 = 8'h74 == _T_174[7:0] ? 4'hf : _GEN_2794; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2796 = 8'h75 == _T_174[7:0] ? 4'hf : _GEN_2795; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2797 = 8'h76 == _T_174[7:0] ? 4'hf : _GEN_2796; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2798 = 8'h77 == _T_174[7:0] ? 4'hf : _GEN_2797; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2799 = 8'h78 == _T_174[7:0] ? 4'hf : _GEN_2798; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2800 = 8'h79 == _T_174[7:0] ? 4'hf : _GEN_2799; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2801 = 8'h7a == _T_174[7:0] ? 4'hf : _GEN_2800; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2802 = 8'h7b == _T_174[7:0] ? 4'hf : _GEN_2801; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2803 = 8'h7c == _T_174[7:0] ? 4'hf : _GEN_2802; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2804 = 8'h7d == _T_174[7:0] ? 4'hf : _GEN_2803; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2805 = 8'h7e == _T_174[7:0] ? 4'hf : _GEN_2804; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2806 = 8'h7f == _T_174[7:0] ? 4'hf : _GEN_2805; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2807 = 8'h80 == _T_174[7:0] ? 4'hf : _GEN_2806; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2808 = 8'h81 == _T_174[7:0] ? 4'hf : _GEN_2807; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2809 = 8'h82 == _T_174[7:0] ? 4'hf : _GEN_2808; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2810 = 8'h83 == _T_174[7:0] ? 4'hf : _GEN_2809; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2811 = 8'h84 == _T_174[7:0] ? 4'hf : _GEN_2810; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2812 = 8'h85 == _T_174[7:0] ? 4'hf : _GEN_2811; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2813 = 8'h86 == _T_174[7:0] ? 4'hf : _GEN_2812; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2814 = 8'h87 == _T_174[7:0] ? 4'hf : _GEN_2813; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2815 = 8'h88 == _T_174[7:0] ? 4'hf : _GEN_2814; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2816 = 8'h89 == _T_174[7:0] ? 4'hf : _GEN_2815; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2817 = 8'h8a == _T_174[7:0] ? 4'hf : _GEN_2816; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2818 = 8'h8b == _T_174[7:0] ? 4'hf : _GEN_2817; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2819 = 8'h8c == _T_174[7:0] ? 4'hf : _GEN_2818; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2820 = 8'h8d == _T_174[7:0] ? 4'hf : _GEN_2819; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2821 = 8'h8e == _T_174[7:0] ? 4'hf : _GEN_2820; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2822 = 8'h8f == _T_174[7:0] ? 4'hf : _GEN_2821; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2823 = 8'h90 == _T_174[7:0] ? 4'hf : _GEN_2822; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2824 = 8'h91 == _T_174[7:0] ? 4'hf : _GEN_2823; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2825 = 8'h92 == _T_174[7:0] ? 4'hf : _GEN_2824; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2826 = 8'h93 == _T_174[7:0] ? 4'hf : _GEN_2825; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2827 = 8'h94 == _T_174[7:0] ? 4'hf : _GEN_2826; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2828 = 8'h95 == _T_174[7:0] ? 4'hf : _GEN_2827; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2829 = 8'h96 == _T_174[7:0] ? 4'hf : _GEN_2828; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2830 = 8'h97 == _T_174[7:0] ? 4'hf : _GEN_2829; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2831 = 8'h98 == _T_174[7:0] ? 4'hf : _GEN_2830; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2832 = 8'h99 == _T_174[7:0] ? 4'hf : _GEN_2831; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2833 = 8'h9a == _T_174[7:0] ? 4'hf : _GEN_2832; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2834 = 8'h9b == _T_174[7:0] ? 4'hf : _GEN_2833; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2835 = 8'h9c == _T_174[7:0] ? 4'hf : _GEN_2834; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2836 = 8'h9d == _T_174[7:0] ? 4'hf : _GEN_2835; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2837 = 8'h9e == _T_174[7:0] ? 4'hf : _GEN_2836; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2838 = 8'h9f == _T_174[7:0] ? 4'hf : _GEN_2837; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2839 = 8'ha0 == _T_174[7:0] ? 4'hf : _GEN_2838; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2840 = 8'ha1 == _T_174[7:0] ? 4'hf : _GEN_2839; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2841 = 8'ha2 == _T_174[7:0] ? 4'hf : _GEN_2840; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2842 = 8'ha3 == _T_174[7:0] ? 4'hf : _GEN_2841; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2843 = 8'ha4 == _T_174[7:0] ? 4'hf : _GEN_2842; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2844 = 8'ha5 == _T_174[7:0] ? 4'hf : _GEN_2843; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2845 = 8'ha6 == _T_174[7:0] ? 4'hf : _GEN_2844; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2846 = 8'ha7 == _T_174[7:0] ? 4'hf : _GEN_2845; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2847 = 8'ha8 == _T_174[7:0] ? 4'hf : _GEN_2846; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2848 = 8'ha9 == _T_174[7:0] ? 4'hf : _GEN_2847; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2849 = 8'haa == _T_174[7:0] ? 4'hf : _GEN_2848; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2850 = 8'hab == _T_174[7:0] ? 4'hf : _GEN_2849; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2851 = 8'hac == _T_174[7:0] ? 4'hf : _GEN_2850; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2852 = 8'had == _T_174[7:0] ? 4'hf : _GEN_2851; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2853 = 8'hae == _T_174[7:0] ? 4'hf : _GEN_2852; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2854 = 8'haf == _T_174[7:0] ? 4'hf : _GEN_2853; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2855 = 8'hb0 == _T_174[7:0] ? 4'hf : _GEN_2854; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2856 = 8'hb1 == _T_174[7:0] ? 4'hf : _GEN_2855; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2857 = 8'hb2 == _T_174[7:0] ? 4'hf : _GEN_2856; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2858 = 8'hb3 == _T_174[7:0] ? 4'hf : _GEN_2857; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2859 = 8'hb4 == _T_174[7:0] ? 4'hf : _GEN_2858; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2860 = 8'hb5 == _T_174[7:0] ? 4'hf : _GEN_2859; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2861 = 8'hb6 == _T_174[7:0] ? 4'hf : _GEN_2860; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2862 = 8'hb7 == _T_174[7:0] ? 4'hf : _GEN_2861; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2863 = 8'hb8 == _T_174[7:0] ? 4'hf : _GEN_2862; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2864 = 8'hb9 == _T_174[7:0] ? 4'hf : _GEN_2863; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2865 = 8'hba == _T_174[7:0] ? 4'hf : _GEN_2864; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2866 = 8'hbb == _T_174[7:0] ? 4'hf : _GEN_2865; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2867 = 8'hbc == _T_174[7:0] ? 4'hf : _GEN_2866; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2868 = 8'hbd == _T_174[7:0] ? 4'hf : _GEN_2867; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2869 = 8'hbe == _T_174[7:0] ? 4'hf : _GEN_2868; // @[Filter.scala 160:102]
  wire [3:0] _GEN_2870 = 8'hbf == _T_174[7:0] ? 4'hf : _GEN_2869; // @[Filter.scala 160:102]
  wire [6:0] _GEN_9892 = {{3'd0}, _GEN_2870}; // @[Filter.scala 160:102]
  wire [10:0] _T_181 = _GEN_9892 * 7'h46; // @[Filter.scala 160:102]
  wire [10:0] _GEN_9893 = {{2'd0}, _T_176}; // @[Filter.scala 160:69]
  wire [10:0] _T_183 = _GEN_9893 + _T_181; // @[Filter.scala 160:69]
  wire [3:0] _GEN_2879 = 8'h8 == _T_174[7:0] ? 4'hf : 4'h0; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2880 = 8'h9 == _T_174[7:0] ? 4'hf : _GEN_2879; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2881 = 8'ha == _T_174[7:0] ? 4'hf : _GEN_2880; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2882 = 8'hb == _T_174[7:0] ? 4'hf : _GEN_2881; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2883 = 8'hc == _T_174[7:0] ? 4'hf : _GEN_2882; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2884 = 8'hd == _T_174[7:0] ? 4'hf : _GEN_2883; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2885 = 8'he == _T_174[7:0] ? 4'hf : _GEN_2884; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2886 = 8'hf == _T_174[7:0] ? 4'hf : _GEN_2885; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2887 = 8'h10 == _T_174[7:0] ? 4'h0 : _GEN_2886; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2888 = 8'h11 == _T_174[7:0] ? 4'h0 : _GEN_2887; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2889 = 8'h12 == _T_174[7:0] ? 4'h0 : _GEN_2888; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2890 = 8'h13 == _T_174[7:0] ? 4'h0 : _GEN_2889; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2891 = 8'h14 == _T_174[7:0] ? 4'h0 : _GEN_2890; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2892 = 8'h15 == _T_174[7:0] ? 4'h0 : _GEN_2891; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2893 = 8'h16 == _T_174[7:0] ? 4'h0 : _GEN_2892; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2894 = 8'h17 == _T_174[7:0] ? 4'h0 : _GEN_2893; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2895 = 8'h18 == _T_174[7:0] ? 4'hf : _GEN_2894; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2896 = 8'h19 == _T_174[7:0] ? 4'hf : _GEN_2895; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2897 = 8'h1a == _T_174[7:0] ? 4'hf : _GEN_2896; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2898 = 8'h1b == _T_174[7:0] ? 4'hf : _GEN_2897; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2899 = 8'h1c == _T_174[7:0] ? 4'hf : _GEN_2898; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2900 = 8'h1d == _T_174[7:0] ? 4'hf : _GEN_2899; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2901 = 8'h1e == _T_174[7:0] ? 4'hf : _GEN_2900; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2902 = 8'h1f == _T_174[7:0] ? 4'hf : _GEN_2901; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2903 = 8'h20 == _T_174[7:0] ? 4'h0 : _GEN_2902; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2904 = 8'h21 == _T_174[7:0] ? 4'h0 : _GEN_2903; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2905 = 8'h22 == _T_174[7:0] ? 4'h0 : _GEN_2904; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2906 = 8'h23 == _T_174[7:0] ? 4'h0 : _GEN_2905; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2907 = 8'h24 == _T_174[7:0] ? 4'h0 : _GEN_2906; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2908 = 8'h25 == _T_174[7:0] ? 4'h0 : _GEN_2907; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2909 = 8'h26 == _T_174[7:0] ? 4'h0 : _GEN_2908; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2910 = 8'h27 == _T_174[7:0] ? 4'h0 : _GEN_2909; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2911 = 8'h28 == _T_174[7:0] ? 4'hf : _GEN_2910; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2912 = 8'h29 == _T_174[7:0] ? 4'hf : _GEN_2911; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2913 = 8'h2a == _T_174[7:0] ? 4'hf : _GEN_2912; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2914 = 8'h2b == _T_174[7:0] ? 4'hf : _GEN_2913; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2915 = 8'h2c == _T_174[7:0] ? 4'hf : _GEN_2914; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2916 = 8'h2d == _T_174[7:0] ? 4'hf : _GEN_2915; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2917 = 8'h2e == _T_174[7:0] ? 4'hf : _GEN_2916; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2918 = 8'h2f == _T_174[7:0] ? 4'hf : _GEN_2917; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2919 = 8'h30 == _T_174[7:0] ? 4'h0 : _GEN_2918; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2920 = 8'h31 == _T_174[7:0] ? 4'h0 : _GEN_2919; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2921 = 8'h32 == _T_174[7:0] ? 4'h0 : _GEN_2920; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2922 = 8'h33 == _T_174[7:0] ? 4'h0 : _GEN_2921; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2923 = 8'h34 == _T_174[7:0] ? 4'h0 : _GEN_2922; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2924 = 8'h35 == _T_174[7:0] ? 4'h0 : _GEN_2923; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2925 = 8'h36 == _T_174[7:0] ? 4'h0 : _GEN_2924; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2926 = 8'h37 == _T_174[7:0] ? 4'h0 : _GEN_2925; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2927 = 8'h38 == _T_174[7:0] ? 4'hf : _GEN_2926; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2928 = 8'h39 == _T_174[7:0] ? 4'hf : _GEN_2927; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2929 = 8'h3a == _T_174[7:0] ? 4'hf : _GEN_2928; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2930 = 8'h3b == _T_174[7:0] ? 4'hf : _GEN_2929; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2931 = 8'h3c == _T_174[7:0] ? 4'hf : _GEN_2930; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2932 = 8'h3d == _T_174[7:0] ? 4'hf : _GEN_2931; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2933 = 8'h3e == _T_174[7:0] ? 4'hf : _GEN_2932; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2934 = 8'h3f == _T_174[7:0] ? 4'hf : _GEN_2933; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2935 = 8'h40 == _T_174[7:0] ? 4'h0 : _GEN_2934; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2936 = 8'h41 == _T_174[7:0] ? 4'h0 : _GEN_2935; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2937 = 8'h42 == _T_174[7:0] ? 4'h0 : _GEN_2936; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2938 = 8'h43 == _T_174[7:0] ? 4'h0 : _GEN_2937; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2939 = 8'h44 == _T_174[7:0] ? 4'h0 : _GEN_2938; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2940 = 8'h45 == _T_174[7:0] ? 4'h0 : _GEN_2939; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2941 = 8'h46 == _T_174[7:0] ? 4'h0 : _GEN_2940; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2942 = 8'h47 == _T_174[7:0] ? 4'h0 : _GEN_2941; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2943 = 8'h48 == _T_174[7:0] ? 4'hf : _GEN_2942; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2944 = 8'h49 == _T_174[7:0] ? 4'hf : _GEN_2943; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2945 = 8'h4a == _T_174[7:0] ? 4'hf : _GEN_2944; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2946 = 8'h4b == _T_174[7:0] ? 4'hf : _GEN_2945; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2947 = 8'h4c == _T_174[7:0] ? 4'hf : _GEN_2946; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2948 = 8'h4d == _T_174[7:0] ? 4'hf : _GEN_2947; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2949 = 8'h4e == _T_174[7:0] ? 4'hf : _GEN_2948; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2950 = 8'h4f == _T_174[7:0] ? 4'hf : _GEN_2949; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2951 = 8'h50 == _T_174[7:0] ? 4'h0 : _GEN_2950; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2952 = 8'h51 == _T_174[7:0] ? 4'h0 : _GEN_2951; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2953 = 8'h52 == _T_174[7:0] ? 4'h0 : _GEN_2952; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2954 = 8'h53 == _T_174[7:0] ? 4'h0 : _GEN_2953; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2955 = 8'h54 == _T_174[7:0] ? 4'h0 : _GEN_2954; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2956 = 8'h55 == _T_174[7:0] ? 4'h0 : _GEN_2955; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2957 = 8'h56 == _T_174[7:0] ? 4'h0 : _GEN_2956; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2958 = 8'h57 == _T_174[7:0] ? 4'h0 : _GEN_2957; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2959 = 8'h58 == _T_174[7:0] ? 4'hf : _GEN_2958; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2960 = 8'h59 == _T_174[7:0] ? 4'hf : _GEN_2959; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2961 = 8'h5a == _T_174[7:0] ? 4'hf : _GEN_2960; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2962 = 8'h5b == _T_174[7:0] ? 4'hf : _GEN_2961; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2963 = 8'h5c == _T_174[7:0] ? 4'hf : _GEN_2962; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2964 = 8'h5d == _T_174[7:0] ? 4'hf : _GEN_2963; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2965 = 8'h5e == _T_174[7:0] ? 4'hf : _GEN_2964; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2966 = 8'h5f == _T_174[7:0] ? 4'hf : _GEN_2965; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2967 = 8'h60 == _T_174[7:0] ? 4'h0 : _GEN_2966; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2968 = 8'h61 == _T_174[7:0] ? 4'h0 : _GEN_2967; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2969 = 8'h62 == _T_174[7:0] ? 4'h0 : _GEN_2968; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2970 = 8'h63 == _T_174[7:0] ? 4'h0 : _GEN_2969; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2971 = 8'h64 == _T_174[7:0] ? 4'h0 : _GEN_2970; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2972 = 8'h65 == _T_174[7:0] ? 4'h0 : _GEN_2971; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2973 = 8'h66 == _T_174[7:0] ? 4'h0 : _GEN_2972; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2974 = 8'h67 == _T_174[7:0] ? 4'h0 : _GEN_2973; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2975 = 8'h68 == _T_174[7:0] ? 4'hf : _GEN_2974; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2976 = 8'h69 == _T_174[7:0] ? 4'hf : _GEN_2975; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2977 = 8'h6a == _T_174[7:0] ? 4'hf : _GEN_2976; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2978 = 8'h6b == _T_174[7:0] ? 4'hf : _GEN_2977; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2979 = 8'h6c == _T_174[7:0] ? 4'hf : _GEN_2978; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2980 = 8'h6d == _T_174[7:0] ? 4'hf : _GEN_2979; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2981 = 8'h6e == _T_174[7:0] ? 4'hf : _GEN_2980; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2982 = 8'h6f == _T_174[7:0] ? 4'hf : _GEN_2981; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2983 = 8'h70 == _T_174[7:0] ? 4'h0 : _GEN_2982; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2984 = 8'h71 == _T_174[7:0] ? 4'h0 : _GEN_2983; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2985 = 8'h72 == _T_174[7:0] ? 4'h0 : _GEN_2984; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2986 = 8'h73 == _T_174[7:0] ? 4'h0 : _GEN_2985; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2987 = 8'h74 == _T_174[7:0] ? 4'h0 : _GEN_2986; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2988 = 8'h75 == _T_174[7:0] ? 4'h0 : _GEN_2987; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2989 = 8'h76 == _T_174[7:0] ? 4'h0 : _GEN_2988; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2990 = 8'h77 == _T_174[7:0] ? 4'h0 : _GEN_2989; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2991 = 8'h78 == _T_174[7:0] ? 4'hf : _GEN_2990; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2992 = 8'h79 == _T_174[7:0] ? 4'hf : _GEN_2991; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2993 = 8'h7a == _T_174[7:0] ? 4'hf : _GEN_2992; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2994 = 8'h7b == _T_174[7:0] ? 4'hf : _GEN_2993; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2995 = 8'h7c == _T_174[7:0] ? 4'hf : _GEN_2994; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2996 = 8'h7d == _T_174[7:0] ? 4'hf : _GEN_2995; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2997 = 8'h7e == _T_174[7:0] ? 4'hf : _GEN_2996; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2998 = 8'h7f == _T_174[7:0] ? 4'hf : _GEN_2997; // @[Filter.scala 160:142]
  wire [3:0] _GEN_2999 = 8'h80 == _T_174[7:0] ? 4'h0 : _GEN_2998; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3000 = 8'h81 == _T_174[7:0] ? 4'h0 : _GEN_2999; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3001 = 8'h82 == _T_174[7:0] ? 4'h0 : _GEN_3000; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3002 = 8'h83 == _T_174[7:0] ? 4'h0 : _GEN_3001; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3003 = 8'h84 == _T_174[7:0] ? 4'h0 : _GEN_3002; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3004 = 8'h85 == _T_174[7:0] ? 4'h0 : _GEN_3003; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3005 = 8'h86 == _T_174[7:0] ? 4'h0 : _GEN_3004; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3006 = 8'h87 == _T_174[7:0] ? 4'h0 : _GEN_3005; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3007 = 8'h88 == _T_174[7:0] ? 4'hf : _GEN_3006; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3008 = 8'h89 == _T_174[7:0] ? 4'hf : _GEN_3007; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3009 = 8'h8a == _T_174[7:0] ? 4'hf : _GEN_3008; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3010 = 8'h8b == _T_174[7:0] ? 4'hf : _GEN_3009; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3011 = 8'h8c == _T_174[7:0] ? 4'hf : _GEN_3010; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3012 = 8'h8d == _T_174[7:0] ? 4'hf : _GEN_3011; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3013 = 8'h8e == _T_174[7:0] ? 4'hf : _GEN_3012; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3014 = 8'h8f == _T_174[7:0] ? 4'hf : _GEN_3013; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3015 = 8'h90 == _T_174[7:0] ? 4'h0 : _GEN_3014; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3016 = 8'h91 == _T_174[7:0] ? 4'h0 : _GEN_3015; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3017 = 8'h92 == _T_174[7:0] ? 4'h0 : _GEN_3016; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3018 = 8'h93 == _T_174[7:0] ? 4'h0 : _GEN_3017; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3019 = 8'h94 == _T_174[7:0] ? 4'h0 : _GEN_3018; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3020 = 8'h95 == _T_174[7:0] ? 4'h0 : _GEN_3019; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3021 = 8'h96 == _T_174[7:0] ? 4'h0 : _GEN_3020; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3022 = 8'h97 == _T_174[7:0] ? 4'h0 : _GEN_3021; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3023 = 8'h98 == _T_174[7:0] ? 4'hf : _GEN_3022; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3024 = 8'h99 == _T_174[7:0] ? 4'hf : _GEN_3023; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3025 = 8'h9a == _T_174[7:0] ? 4'hf : _GEN_3024; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3026 = 8'h9b == _T_174[7:0] ? 4'hf : _GEN_3025; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3027 = 8'h9c == _T_174[7:0] ? 4'hf : _GEN_3026; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3028 = 8'h9d == _T_174[7:0] ? 4'hf : _GEN_3027; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3029 = 8'h9e == _T_174[7:0] ? 4'hf : _GEN_3028; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3030 = 8'h9f == _T_174[7:0] ? 4'hf : _GEN_3029; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3031 = 8'ha0 == _T_174[7:0] ? 4'h0 : _GEN_3030; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3032 = 8'ha1 == _T_174[7:0] ? 4'h0 : _GEN_3031; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3033 = 8'ha2 == _T_174[7:0] ? 4'h0 : _GEN_3032; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3034 = 8'ha3 == _T_174[7:0] ? 4'h0 : _GEN_3033; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3035 = 8'ha4 == _T_174[7:0] ? 4'h0 : _GEN_3034; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3036 = 8'ha5 == _T_174[7:0] ? 4'h0 : _GEN_3035; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3037 = 8'ha6 == _T_174[7:0] ? 4'h0 : _GEN_3036; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3038 = 8'ha7 == _T_174[7:0] ? 4'h0 : _GEN_3037; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3039 = 8'ha8 == _T_174[7:0] ? 4'hf : _GEN_3038; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3040 = 8'ha9 == _T_174[7:0] ? 4'hf : _GEN_3039; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3041 = 8'haa == _T_174[7:0] ? 4'hf : _GEN_3040; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3042 = 8'hab == _T_174[7:0] ? 4'hf : _GEN_3041; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3043 = 8'hac == _T_174[7:0] ? 4'hf : _GEN_3042; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3044 = 8'had == _T_174[7:0] ? 4'hf : _GEN_3043; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3045 = 8'hae == _T_174[7:0] ? 4'hf : _GEN_3044; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3046 = 8'haf == _T_174[7:0] ? 4'hf : _GEN_3045; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3047 = 8'hb0 == _T_174[7:0] ? 4'h0 : _GEN_3046; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3048 = 8'hb1 == _T_174[7:0] ? 4'h0 : _GEN_3047; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3049 = 8'hb2 == _T_174[7:0] ? 4'h0 : _GEN_3048; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3050 = 8'hb3 == _T_174[7:0] ? 4'h0 : _GEN_3049; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3051 = 8'hb4 == _T_174[7:0] ? 4'h0 : _GEN_3050; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3052 = 8'hb5 == _T_174[7:0] ? 4'h0 : _GEN_3051; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3053 = 8'hb6 == _T_174[7:0] ? 4'h0 : _GEN_3052; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3054 = 8'hb7 == _T_174[7:0] ? 4'h0 : _GEN_3053; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3055 = 8'hb8 == _T_174[7:0] ? 4'hf : _GEN_3054; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3056 = 8'hb9 == _T_174[7:0] ? 4'hf : _GEN_3055; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3057 = 8'hba == _T_174[7:0] ? 4'hf : _GEN_3056; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3058 = 8'hbb == _T_174[7:0] ? 4'hf : _GEN_3057; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3059 = 8'hbc == _T_174[7:0] ? 4'hf : _GEN_3058; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3060 = 8'hbd == _T_174[7:0] ? 4'hf : _GEN_3059; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3061 = 8'hbe == _T_174[7:0] ? 4'hf : _GEN_3060; // @[Filter.scala 160:142]
  wire [3:0] _GEN_3062 = 8'hbf == _T_174[7:0] ? 4'hf : _GEN_3061; // @[Filter.scala 160:142]
  wire [7:0] _T_188 = _GEN_3062 * 4'ha; // @[Filter.scala 160:142]
  wire [10:0] _GEN_9895 = {{3'd0}, _T_188}; // @[Filter.scala 160:109]
  wire [10:0] _T_190 = _T_183 + _GEN_9895; // @[Filter.scala 160:109]
  wire [10:0] _T_191 = _T_190 / 11'h64; // @[Filter.scala 160:150]
  wire  _T_193 = _T_164 >= 5'h10; // @[Filter.scala 163:31]
  wire  _T_197 = _T_171 >= 32'hc; // @[Filter.scala 163:63]
  wire  _T_198 = _T_193 | _T_197; // @[Filter.scala 163:58]
  wire [10:0] _GEN_3255 = io_SPI_distort ? _T_191 : {{7'd0}, _GEN_2678}; // @[Filter.scala 165:35]
  wire [10:0] _GEN_3256 = _T_198 ? 11'h0 : _GEN_3255; // @[Filter.scala 163:80]
  wire [10:0] _GEN_3449 = io_SPI_distort ? _T_191 : {{7'd0}, _GEN_2870}; // @[Filter.scala 165:35]
  wire [10:0] _GEN_3450 = _T_198 ? 11'h0 : _GEN_3449; // @[Filter.scala 163:80]
  wire [10:0] _GEN_3643 = io_SPI_distort ? _T_191 : {{7'd0}, _GEN_3062}; // @[Filter.scala 165:35]
  wire [10:0] _GEN_3644 = _T_198 ? 11'h0 : _GEN_3643; // @[Filter.scala 163:80]
  wire [31:0] _T_226 = pixelIndex + 32'h3; // @[Filter.scala 158:31]
  wire [31:0] _GEN_3 = _T_226 % 32'h10; // @[Filter.scala 158:38]
  wire [4:0] _T_227 = _GEN_3[4:0]; // @[Filter.scala 158:38]
  wire [4:0] _T_229 = _T_227 + _GEN_9863; // @[Filter.scala 158:53]
  wire [4:0] _T_231 = _T_229 - 5'h1; // @[Filter.scala 158:69]
  wire [31:0] _T_234 = _T_226 / 32'h10; // @[Filter.scala 159:38]
  wire [31:0] _T_236 = _T_234 + _GEN_9864; // @[Filter.scala 159:53]
  wire [31:0] _T_238 = _T_236 - 32'h1; // @[Filter.scala 159:69]
  wire [36:0] _T_239 = _T_238 * 32'h10; // @[Filter.scala 160:42]
  wire [36:0] _GEN_9901 = {{32'd0}, _T_231}; // @[Filter.scala 160:57]
  wire [36:0] _T_241 = _T_239 + _GEN_9901; // @[Filter.scala 160:57]
  wire [3:0] _GEN_3653 = 8'h8 == _T_241[7:0] ? 4'h0 : 4'hf; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3654 = 8'h9 == _T_241[7:0] ? 4'h0 : _GEN_3653; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3655 = 8'ha == _T_241[7:0] ? 4'h0 : _GEN_3654; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3656 = 8'hb == _T_241[7:0] ? 4'h0 : _GEN_3655; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3657 = 8'hc == _T_241[7:0] ? 4'h0 : _GEN_3656; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3658 = 8'hd == _T_241[7:0] ? 4'h0 : _GEN_3657; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3659 = 8'he == _T_241[7:0] ? 4'h0 : _GEN_3658; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3660 = 8'hf == _T_241[7:0] ? 4'h0 : _GEN_3659; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3661 = 8'h10 == _T_241[7:0] ? 4'hf : _GEN_3660; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3662 = 8'h11 == _T_241[7:0] ? 4'hf : _GEN_3661; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3663 = 8'h12 == _T_241[7:0] ? 4'hf : _GEN_3662; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3664 = 8'h13 == _T_241[7:0] ? 4'hf : _GEN_3663; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3665 = 8'h14 == _T_241[7:0] ? 4'hf : _GEN_3664; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3666 = 8'h15 == _T_241[7:0] ? 4'hf : _GEN_3665; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3667 = 8'h16 == _T_241[7:0] ? 4'hf : _GEN_3666; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3668 = 8'h17 == _T_241[7:0] ? 4'hf : _GEN_3667; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3669 = 8'h18 == _T_241[7:0] ? 4'h0 : _GEN_3668; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3670 = 8'h19 == _T_241[7:0] ? 4'h0 : _GEN_3669; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3671 = 8'h1a == _T_241[7:0] ? 4'h0 : _GEN_3670; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3672 = 8'h1b == _T_241[7:0] ? 4'h0 : _GEN_3671; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3673 = 8'h1c == _T_241[7:0] ? 4'h0 : _GEN_3672; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3674 = 8'h1d == _T_241[7:0] ? 4'h0 : _GEN_3673; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3675 = 8'h1e == _T_241[7:0] ? 4'h0 : _GEN_3674; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3676 = 8'h1f == _T_241[7:0] ? 4'h0 : _GEN_3675; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3677 = 8'h20 == _T_241[7:0] ? 4'hf : _GEN_3676; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3678 = 8'h21 == _T_241[7:0] ? 4'hf : _GEN_3677; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3679 = 8'h22 == _T_241[7:0] ? 4'hf : _GEN_3678; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3680 = 8'h23 == _T_241[7:0] ? 4'hf : _GEN_3679; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3681 = 8'h24 == _T_241[7:0] ? 4'hf : _GEN_3680; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3682 = 8'h25 == _T_241[7:0] ? 4'hf : _GEN_3681; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3683 = 8'h26 == _T_241[7:0] ? 4'hf : _GEN_3682; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3684 = 8'h27 == _T_241[7:0] ? 4'hf : _GEN_3683; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3685 = 8'h28 == _T_241[7:0] ? 4'h0 : _GEN_3684; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3686 = 8'h29 == _T_241[7:0] ? 4'h0 : _GEN_3685; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3687 = 8'h2a == _T_241[7:0] ? 4'h0 : _GEN_3686; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3688 = 8'h2b == _T_241[7:0] ? 4'h0 : _GEN_3687; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3689 = 8'h2c == _T_241[7:0] ? 4'h0 : _GEN_3688; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3690 = 8'h2d == _T_241[7:0] ? 4'h0 : _GEN_3689; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3691 = 8'h2e == _T_241[7:0] ? 4'h0 : _GEN_3690; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3692 = 8'h2f == _T_241[7:0] ? 4'h0 : _GEN_3691; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3693 = 8'h30 == _T_241[7:0] ? 4'hf : _GEN_3692; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3694 = 8'h31 == _T_241[7:0] ? 4'hf : _GEN_3693; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3695 = 8'h32 == _T_241[7:0] ? 4'hf : _GEN_3694; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3696 = 8'h33 == _T_241[7:0] ? 4'hf : _GEN_3695; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3697 = 8'h34 == _T_241[7:0] ? 4'hf : _GEN_3696; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3698 = 8'h35 == _T_241[7:0] ? 4'hf : _GEN_3697; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3699 = 8'h36 == _T_241[7:0] ? 4'hf : _GEN_3698; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3700 = 8'h37 == _T_241[7:0] ? 4'hf : _GEN_3699; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3701 = 8'h38 == _T_241[7:0] ? 4'h0 : _GEN_3700; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3702 = 8'h39 == _T_241[7:0] ? 4'h0 : _GEN_3701; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3703 = 8'h3a == _T_241[7:0] ? 4'h0 : _GEN_3702; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3704 = 8'h3b == _T_241[7:0] ? 4'h0 : _GEN_3703; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3705 = 8'h3c == _T_241[7:0] ? 4'h0 : _GEN_3704; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3706 = 8'h3d == _T_241[7:0] ? 4'h0 : _GEN_3705; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3707 = 8'h3e == _T_241[7:0] ? 4'h0 : _GEN_3706; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3708 = 8'h3f == _T_241[7:0] ? 4'h0 : _GEN_3707; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3709 = 8'h40 == _T_241[7:0] ? 4'hf : _GEN_3708; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3710 = 8'h41 == _T_241[7:0] ? 4'hf : _GEN_3709; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3711 = 8'h42 == _T_241[7:0] ? 4'hf : _GEN_3710; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3712 = 8'h43 == _T_241[7:0] ? 4'hf : _GEN_3711; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3713 = 8'h44 == _T_241[7:0] ? 4'hf : _GEN_3712; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3714 = 8'h45 == _T_241[7:0] ? 4'hf : _GEN_3713; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3715 = 8'h46 == _T_241[7:0] ? 4'hf : _GEN_3714; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3716 = 8'h47 == _T_241[7:0] ? 4'hf : _GEN_3715; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3717 = 8'h48 == _T_241[7:0] ? 4'h0 : _GEN_3716; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3718 = 8'h49 == _T_241[7:0] ? 4'h0 : _GEN_3717; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3719 = 8'h4a == _T_241[7:0] ? 4'h0 : _GEN_3718; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3720 = 8'h4b == _T_241[7:0] ? 4'h0 : _GEN_3719; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3721 = 8'h4c == _T_241[7:0] ? 4'h0 : _GEN_3720; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3722 = 8'h4d == _T_241[7:0] ? 4'h0 : _GEN_3721; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3723 = 8'h4e == _T_241[7:0] ? 4'h0 : _GEN_3722; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3724 = 8'h4f == _T_241[7:0] ? 4'h0 : _GEN_3723; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3725 = 8'h50 == _T_241[7:0] ? 4'hf : _GEN_3724; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3726 = 8'h51 == _T_241[7:0] ? 4'hf : _GEN_3725; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3727 = 8'h52 == _T_241[7:0] ? 4'hf : _GEN_3726; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3728 = 8'h53 == _T_241[7:0] ? 4'hf : _GEN_3727; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3729 = 8'h54 == _T_241[7:0] ? 4'hf : _GEN_3728; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3730 = 8'h55 == _T_241[7:0] ? 4'hf : _GEN_3729; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3731 = 8'h56 == _T_241[7:0] ? 4'hf : _GEN_3730; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3732 = 8'h57 == _T_241[7:0] ? 4'hf : _GEN_3731; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3733 = 8'h58 == _T_241[7:0] ? 4'h0 : _GEN_3732; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3734 = 8'h59 == _T_241[7:0] ? 4'h0 : _GEN_3733; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3735 = 8'h5a == _T_241[7:0] ? 4'h0 : _GEN_3734; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3736 = 8'h5b == _T_241[7:0] ? 4'h0 : _GEN_3735; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3737 = 8'h5c == _T_241[7:0] ? 4'h0 : _GEN_3736; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3738 = 8'h5d == _T_241[7:0] ? 4'h0 : _GEN_3737; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3739 = 8'h5e == _T_241[7:0] ? 4'h0 : _GEN_3738; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3740 = 8'h5f == _T_241[7:0] ? 4'h0 : _GEN_3739; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3741 = 8'h60 == _T_241[7:0] ? 4'h0 : _GEN_3740; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3742 = 8'h61 == _T_241[7:0] ? 4'h0 : _GEN_3741; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3743 = 8'h62 == _T_241[7:0] ? 4'h0 : _GEN_3742; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3744 = 8'h63 == _T_241[7:0] ? 4'h0 : _GEN_3743; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3745 = 8'h64 == _T_241[7:0] ? 4'h0 : _GEN_3744; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3746 = 8'h65 == _T_241[7:0] ? 4'h0 : _GEN_3745; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3747 = 8'h66 == _T_241[7:0] ? 4'h0 : _GEN_3746; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3748 = 8'h67 == _T_241[7:0] ? 4'h0 : _GEN_3747; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3749 = 8'h68 == _T_241[7:0] ? 4'hf : _GEN_3748; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3750 = 8'h69 == _T_241[7:0] ? 4'hf : _GEN_3749; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3751 = 8'h6a == _T_241[7:0] ? 4'hf : _GEN_3750; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3752 = 8'h6b == _T_241[7:0] ? 4'hf : _GEN_3751; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3753 = 8'h6c == _T_241[7:0] ? 4'hf : _GEN_3752; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3754 = 8'h6d == _T_241[7:0] ? 4'hf : _GEN_3753; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3755 = 8'h6e == _T_241[7:0] ? 4'hf : _GEN_3754; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3756 = 8'h6f == _T_241[7:0] ? 4'hf : _GEN_3755; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3757 = 8'h70 == _T_241[7:0] ? 4'h0 : _GEN_3756; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3758 = 8'h71 == _T_241[7:0] ? 4'h0 : _GEN_3757; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3759 = 8'h72 == _T_241[7:0] ? 4'h0 : _GEN_3758; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3760 = 8'h73 == _T_241[7:0] ? 4'h0 : _GEN_3759; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3761 = 8'h74 == _T_241[7:0] ? 4'h0 : _GEN_3760; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3762 = 8'h75 == _T_241[7:0] ? 4'h0 : _GEN_3761; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3763 = 8'h76 == _T_241[7:0] ? 4'h0 : _GEN_3762; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3764 = 8'h77 == _T_241[7:0] ? 4'h0 : _GEN_3763; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3765 = 8'h78 == _T_241[7:0] ? 4'hf : _GEN_3764; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3766 = 8'h79 == _T_241[7:0] ? 4'hf : _GEN_3765; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3767 = 8'h7a == _T_241[7:0] ? 4'hf : _GEN_3766; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3768 = 8'h7b == _T_241[7:0] ? 4'hf : _GEN_3767; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3769 = 8'h7c == _T_241[7:0] ? 4'hf : _GEN_3768; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3770 = 8'h7d == _T_241[7:0] ? 4'hf : _GEN_3769; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3771 = 8'h7e == _T_241[7:0] ? 4'hf : _GEN_3770; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3772 = 8'h7f == _T_241[7:0] ? 4'hf : _GEN_3771; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3773 = 8'h80 == _T_241[7:0] ? 4'h0 : _GEN_3772; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3774 = 8'h81 == _T_241[7:0] ? 4'h0 : _GEN_3773; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3775 = 8'h82 == _T_241[7:0] ? 4'h0 : _GEN_3774; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3776 = 8'h83 == _T_241[7:0] ? 4'h0 : _GEN_3775; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3777 = 8'h84 == _T_241[7:0] ? 4'h0 : _GEN_3776; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3778 = 8'h85 == _T_241[7:0] ? 4'h0 : _GEN_3777; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3779 = 8'h86 == _T_241[7:0] ? 4'h0 : _GEN_3778; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3780 = 8'h87 == _T_241[7:0] ? 4'h0 : _GEN_3779; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3781 = 8'h88 == _T_241[7:0] ? 4'hf : _GEN_3780; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3782 = 8'h89 == _T_241[7:0] ? 4'hf : _GEN_3781; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3783 = 8'h8a == _T_241[7:0] ? 4'hf : _GEN_3782; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3784 = 8'h8b == _T_241[7:0] ? 4'hf : _GEN_3783; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3785 = 8'h8c == _T_241[7:0] ? 4'hf : _GEN_3784; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3786 = 8'h8d == _T_241[7:0] ? 4'hf : _GEN_3785; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3787 = 8'h8e == _T_241[7:0] ? 4'hf : _GEN_3786; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3788 = 8'h8f == _T_241[7:0] ? 4'hf : _GEN_3787; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3789 = 8'h90 == _T_241[7:0] ? 4'h0 : _GEN_3788; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3790 = 8'h91 == _T_241[7:0] ? 4'h0 : _GEN_3789; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3791 = 8'h92 == _T_241[7:0] ? 4'h0 : _GEN_3790; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3792 = 8'h93 == _T_241[7:0] ? 4'h0 : _GEN_3791; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3793 = 8'h94 == _T_241[7:0] ? 4'h0 : _GEN_3792; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3794 = 8'h95 == _T_241[7:0] ? 4'h0 : _GEN_3793; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3795 = 8'h96 == _T_241[7:0] ? 4'h0 : _GEN_3794; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3796 = 8'h97 == _T_241[7:0] ? 4'h0 : _GEN_3795; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3797 = 8'h98 == _T_241[7:0] ? 4'hf : _GEN_3796; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3798 = 8'h99 == _T_241[7:0] ? 4'hf : _GEN_3797; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3799 = 8'h9a == _T_241[7:0] ? 4'hf : _GEN_3798; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3800 = 8'h9b == _T_241[7:0] ? 4'hf : _GEN_3799; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3801 = 8'h9c == _T_241[7:0] ? 4'hf : _GEN_3800; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3802 = 8'h9d == _T_241[7:0] ? 4'hf : _GEN_3801; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3803 = 8'h9e == _T_241[7:0] ? 4'hf : _GEN_3802; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3804 = 8'h9f == _T_241[7:0] ? 4'hf : _GEN_3803; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3805 = 8'ha0 == _T_241[7:0] ? 4'h0 : _GEN_3804; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3806 = 8'ha1 == _T_241[7:0] ? 4'h0 : _GEN_3805; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3807 = 8'ha2 == _T_241[7:0] ? 4'h0 : _GEN_3806; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3808 = 8'ha3 == _T_241[7:0] ? 4'h0 : _GEN_3807; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3809 = 8'ha4 == _T_241[7:0] ? 4'h0 : _GEN_3808; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3810 = 8'ha5 == _T_241[7:0] ? 4'h0 : _GEN_3809; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3811 = 8'ha6 == _T_241[7:0] ? 4'h0 : _GEN_3810; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3812 = 8'ha7 == _T_241[7:0] ? 4'h0 : _GEN_3811; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3813 = 8'ha8 == _T_241[7:0] ? 4'hf : _GEN_3812; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3814 = 8'ha9 == _T_241[7:0] ? 4'hf : _GEN_3813; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3815 = 8'haa == _T_241[7:0] ? 4'hf : _GEN_3814; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3816 = 8'hab == _T_241[7:0] ? 4'hf : _GEN_3815; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3817 = 8'hac == _T_241[7:0] ? 4'hf : _GEN_3816; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3818 = 8'had == _T_241[7:0] ? 4'hf : _GEN_3817; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3819 = 8'hae == _T_241[7:0] ? 4'hf : _GEN_3818; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3820 = 8'haf == _T_241[7:0] ? 4'hf : _GEN_3819; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3821 = 8'hb0 == _T_241[7:0] ? 4'h0 : _GEN_3820; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3822 = 8'hb1 == _T_241[7:0] ? 4'h0 : _GEN_3821; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3823 = 8'hb2 == _T_241[7:0] ? 4'h0 : _GEN_3822; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3824 = 8'hb3 == _T_241[7:0] ? 4'h0 : _GEN_3823; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3825 = 8'hb4 == _T_241[7:0] ? 4'h0 : _GEN_3824; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3826 = 8'hb5 == _T_241[7:0] ? 4'h0 : _GEN_3825; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3827 = 8'hb6 == _T_241[7:0] ? 4'h0 : _GEN_3826; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3828 = 8'hb7 == _T_241[7:0] ? 4'h0 : _GEN_3827; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3829 = 8'hb8 == _T_241[7:0] ? 4'hf : _GEN_3828; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3830 = 8'hb9 == _T_241[7:0] ? 4'hf : _GEN_3829; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3831 = 8'hba == _T_241[7:0] ? 4'hf : _GEN_3830; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3832 = 8'hbb == _T_241[7:0] ? 4'hf : _GEN_3831; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3833 = 8'hbc == _T_241[7:0] ? 4'hf : _GEN_3832; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3834 = 8'hbd == _T_241[7:0] ? 4'hf : _GEN_3833; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3835 = 8'hbe == _T_241[7:0] ? 4'hf : _GEN_3834; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3836 = 8'hbf == _T_241[7:0] ? 4'hf : _GEN_3835; // @[Filter.scala 160:62]
  wire [4:0] _GEN_9902 = {{1'd0}, _GEN_3836}; // @[Filter.scala 160:62]
  wire [8:0] _T_243 = _GEN_9902 * 5'h14; // @[Filter.scala 160:62]
  wire [3:0] _GEN_3933 = 8'h60 == _T_241[7:0] ? 4'hf : 4'h0; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3934 = 8'h61 == _T_241[7:0] ? 4'hf : _GEN_3933; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3935 = 8'h62 == _T_241[7:0] ? 4'hf : _GEN_3934; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3936 = 8'h63 == _T_241[7:0] ? 4'hf : _GEN_3935; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3937 = 8'h64 == _T_241[7:0] ? 4'hf : _GEN_3936; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3938 = 8'h65 == _T_241[7:0] ? 4'hf : _GEN_3937; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3939 = 8'h66 == _T_241[7:0] ? 4'hf : _GEN_3938; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3940 = 8'h67 == _T_241[7:0] ? 4'hf : _GEN_3939; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3941 = 8'h68 == _T_241[7:0] ? 4'hf : _GEN_3940; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3942 = 8'h69 == _T_241[7:0] ? 4'hf : _GEN_3941; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3943 = 8'h6a == _T_241[7:0] ? 4'hf : _GEN_3942; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3944 = 8'h6b == _T_241[7:0] ? 4'hf : _GEN_3943; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3945 = 8'h6c == _T_241[7:0] ? 4'hf : _GEN_3944; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3946 = 8'h6d == _T_241[7:0] ? 4'hf : _GEN_3945; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3947 = 8'h6e == _T_241[7:0] ? 4'hf : _GEN_3946; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3948 = 8'h6f == _T_241[7:0] ? 4'hf : _GEN_3947; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3949 = 8'h70 == _T_241[7:0] ? 4'hf : _GEN_3948; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3950 = 8'h71 == _T_241[7:0] ? 4'hf : _GEN_3949; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3951 = 8'h72 == _T_241[7:0] ? 4'hf : _GEN_3950; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3952 = 8'h73 == _T_241[7:0] ? 4'hf : _GEN_3951; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3953 = 8'h74 == _T_241[7:0] ? 4'hf : _GEN_3952; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3954 = 8'h75 == _T_241[7:0] ? 4'hf : _GEN_3953; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3955 = 8'h76 == _T_241[7:0] ? 4'hf : _GEN_3954; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3956 = 8'h77 == _T_241[7:0] ? 4'hf : _GEN_3955; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3957 = 8'h78 == _T_241[7:0] ? 4'hf : _GEN_3956; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3958 = 8'h79 == _T_241[7:0] ? 4'hf : _GEN_3957; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3959 = 8'h7a == _T_241[7:0] ? 4'hf : _GEN_3958; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3960 = 8'h7b == _T_241[7:0] ? 4'hf : _GEN_3959; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3961 = 8'h7c == _T_241[7:0] ? 4'hf : _GEN_3960; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3962 = 8'h7d == _T_241[7:0] ? 4'hf : _GEN_3961; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3963 = 8'h7e == _T_241[7:0] ? 4'hf : _GEN_3962; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3964 = 8'h7f == _T_241[7:0] ? 4'hf : _GEN_3963; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3965 = 8'h80 == _T_241[7:0] ? 4'hf : _GEN_3964; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3966 = 8'h81 == _T_241[7:0] ? 4'hf : _GEN_3965; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3967 = 8'h82 == _T_241[7:0] ? 4'hf : _GEN_3966; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3968 = 8'h83 == _T_241[7:0] ? 4'hf : _GEN_3967; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3969 = 8'h84 == _T_241[7:0] ? 4'hf : _GEN_3968; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3970 = 8'h85 == _T_241[7:0] ? 4'hf : _GEN_3969; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3971 = 8'h86 == _T_241[7:0] ? 4'hf : _GEN_3970; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3972 = 8'h87 == _T_241[7:0] ? 4'hf : _GEN_3971; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3973 = 8'h88 == _T_241[7:0] ? 4'hf : _GEN_3972; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3974 = 8'h89 == _T_241[7:0] ? 4'hf : _GEN_3973; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3975 = 8'h8a == _T_241[7:0] ? 4'hf : _GEN_3974; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3976 = 8'h8b == _T_241[7:0] ? 4'hf : _GEN_3975; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3977 = 8'h8c == _T_241[7:0] ? 4'hf : _GEN_3976; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3978 = 8'h8d == _T_241[7:0] ? 4'hf : _GEN_3977; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3979 = 8'h8e == _T_241[7:0] ? 4'hf : _GEN_3978; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3980 = 8'h8f == _T_241[7:0] ? 4'hf : _GEN_3979; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3981 = 8'h90 == _T_241[7:0] ? 4'hf : _GEN_3980; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3982 = 8'h91 == _T_241[7:0] ? 4'hf : _GEN_3981; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3983 = 8'h92 == _T_241[7:0] ? 4'hf : _GEN_3982; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3984 = 8'h93 == _T_241[7:0] ? 4'hf : _GEN_3983; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3985 = 8'h94 == _T_241[7:0] ? 4'hf : _GEN_3984; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3986 = 8'h95 == _T_241[7:0] ? 4'hf : _GEN_3985; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3987 = 8'h96 == _T_241[7:0] ? 4'hf : _GEN_3986; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3988 = 8'h97 == _T_241[7:0] ? 4'hf : _GEN_3987; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3989 = 8'h98 == _T_241[7:0] ? 4'hf : _GEN_3988; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3990 = 8'h99 == _T_241[7:0] ? 4'hf : _GEN_3989; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3991 = 8'h9a == _T_241[7:0] ? 4'hf : _GEN_3990; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3992 = 8'h9b == _T_241[7:0] ? 4'hf : _GEN_3991; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3993 = 8'h9c == _T_241[7:0] ? 4'hf : _GEN_3992; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3994 = 8'h9d == _T_241[7:0] ? 4'hf : _GEN_3993; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3995 = 8'h9e == _T_241[7:0] ? 4'hf : _GEN_3994; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3996 = 8'h9f == _T_241[7:0] ? 4'hf : _GEN_3995; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3997 = 8'ha0 == _T_241[7:0] ? 4'hf : _GEN_3996; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3998 = 8'ha1 == _T_241[7:0] ? 4'hf : _GEN_3997; // @[Filter.scala 160:102]
  wire [3:0] _GEN_3999 = 8'ha2 == _T_241[7:0] ? 4'hf : _GEN_3998; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4000 = 8'ha3 == _T_241[7:0] ? 4'hf : _GEN_3999; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4001 = 8'ha4 == _T_241[7:0] ? 4'hf : _GEN_4000; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4002 = 8'ha5 == _T_241[7:0] ? 4'hf : _GEN_4001; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4003 = 8'ha6 == _T_241[7:0] ? 4'hf : _GEN_4002; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4004 = 8'ha7 == _T_241[7:0] ? 4'hf : _GEN_4003; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4005 = 8'ha8 == _T_241[7:0] ? 4'hf : _GEN_4004; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4006 = 8'ha9 == _T_241[7:0] ? 4'hf : _GEN_4005; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4007 = 8'haa == _T_241[7:0] ? 4'hf : _GEN_4006; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4008 = 8'hab == _T_241[7:0] ? 4'hf : _GEN_4007; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4009 = 8'hac == _T_241[7:0] ? 4'hf : _GEN_4008; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4010 = 8'had == _T_241[7:0] ? 4'hf : _GEN_4009; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4011 = 8'hae == _T_241[7:0] ? 4'hf : _GEN_4010; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4012 = 8'haf == _T_241[7:0] ? 4'hf : _GEN_4011; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4013 = 8'hb0 == _T_241[7:0] ? 4'hf : _GEN_4012; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4014 = 8'hb1 == _T_241[7:0] ? 4'hf : _GEN_4013; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4015 = 8'hb2 == _T_241[7:0] ? 4'hf : _GEN_4014; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4016 = 8'hb3 == _T_241[7:0] ? 4'hf : _GEN_4015; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4017 = 8'hb4 == _T_241[7:0] ? 4'hf : _GEN_4016; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4018 = 8'hb5 == _T_241[7:0] ? 4'hf : _GEN_4017; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4019 = 8'hb6 == _T_241[7:0] ? 4'hf : _GEN_4018; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4020 = 8'hb7 == _T_241[7:0] ? 4'hf : _GEN_4019; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4021 = 8'hb8 == _T_241[7:0] ? 4'hf : _GEN_4020; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4022 = 8'hb9 == _T_241[7:0] ? 4'hf : _GEN_4021; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4023 = 8'hba == _T_241[7:0] ? 4'hf : _GEN_4022; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4024 = 8'hbb == _T_241[7:0] ? 4'hf : _GEN_4023; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4025 = 8'hbc == _T_241[7:0] ? 4'hf : _GEN_4024; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4026 = 8'hbd == _T_241[7:0] ? 4'hf : _GEN_4025; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4027 = 8'hbe == _T_241[7:0] ? 4'hf : _GEN_4026; // @[Filter.scala 160:102]
  wire [3:0] _GEN_4028 = 8'hbf == _T_241[7:0] ? 4'hf : _GEN_4027; // @[Filter.scala 160:102]
  wire [6:0] _GEN_9904 = {{3'd0}, _GEN_4028}; // @[Filter.scala 160:102]
  wire [10:0] _T_248 = _GEN_9904 * 7'h46; // @[Filter.scala 160:102]
  wire [10:0] _GEN_9905 = {{2'd0}, _T_243}; // @[Filter.scala 160:69]
  wire [10:0] _T_250 = _GEN_9905 + _T_248; // @[Filter.scala 160:69]
  wire [3:0] _GEN_4037 = 8'h8 == _T_241[7:0] ? 4'hf : 4'h0; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4038 = 8'h9 == _T_241[7:0] ? 4'hf : _GEN_4037; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4039 = 8'ha == _T_241[7:0] ? 4'hf : _GEN_4038; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4040 = 8'hb == _T_241[7:0] ? 4'hf : _GEN_4039; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4041 = 8'hc == _T_241[7:0] ? 4'hf : _GEN_4040; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4042 = 8'hd == _T_241[7:0] ? 4'hf : _GEN_4041; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4043 = 8'he == _T_241[7:0] ? 4'hf : _GEN_4042; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4044 = 8'hf == _T_241[7:0] ? 4'hf : _GEN_4043; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4045 = 8'h10 == _T_241[7:0] ? 4'h0 : _GEN_4044; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4046 = 8'h11 == _T_241[7:0] ? 4'h0 : _GEN_4045; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4047 = 8'h12 == _T_241[7:0] ? 4'h0 : _GEN_4046; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4048 = 8'h13 == _T_241[7:0] ? 4'h0 : _GEN_4047; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4049 = 8'h14 == _T_241[7:0] ? 4'h0 : _GEN_4048; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4050 = 8'h15 == _T_241[7:0] ? 4'h0 : _GEN_4049; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4051 = 8'h16 == _T_241[7:0] ? 4'h0 : _GEN_4050; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4052 = 8'h17 == _T_241[7:0] ? 4'h0 : _GEN_4051; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4053 = 8'h18 == _T_241[7:0] ? 4'hf : _GEN_4052; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4054 = 8'h19 == _T_241[7:0] ? 4'hf : _GEN_4053; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4055 = 8'h1a == _T_241[7:0] ? 4'hf : _GEN_4054; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4056 = 8'h1b == _T_241[7:0] ? 4'hf : _GEN_4055; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4057 = 8'h1c == _T_241[7:0] ? 4'hf : _GEN_4056; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4058 = 8'h1d == _T_241[7:0] ? 4'hf : _GEN_4057; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4059 = 8'h1e == _T_241[7:0] ? 4'hf : _GEN_4058; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4060 = 8'h1f == _T_241[7:0] ? 4'hf : _GEN_4059; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4061 = 8'h20 == _T_241[7:0] ? 4'h0 : _GEN_4060; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4062 = 8'h21 == _T_241[7:0] ? 4'h0 : _GEN_4061; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4063 = 8'h22 == _T_241[7:0] ? 4'h0 : _GEN_4062; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4064 = 8'h23 == _T_241[7:0] ? 4'h0 : _GEN_4063; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4065 = 8'h24 == _T_241[7:0] ? 4'h0 : _GEN_4064; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4066 = 8'h25 == _T_241[7:0] ? 4'h0 : _GEN_4065; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4067 = 8'h26 == _T_241[7:0] ? 4'h0 : _GEN_4066; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4068 = 8'h27 == _T_241[7:0] ? 4'h0 : _GEN_4067; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4069 = 8'h28 == _T_241[7:0] ? 4'hf : _GEN_4068; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4070 = 8'h29 == _T_241[7:0] ? 4'hf : _GEN_4069; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4071 = 8'h2a == _T_241[7:0] ? 4'hf : _GEN_4070; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4072 = 8'h2b == _T_241[7:0] ? 4'hf : _GEN_4071; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4073 = 8'h2c == _T_241[7:0] ? 4'hf : _GEN_4072; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4074 = 8'h2d == _T_241[7:0] ? 4'hf : _GEN_4073; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4075 = 8'h2e == _T_241[7:0] ? 4'hf : _GEN_4074; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4076 = 8'h2f == _T_241[7:0] ? 4'hf : _GEN_4075; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4077 = 8'h30 == _T_241[7:0] ? 4'h0 : _GEN_4076; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4078 = 8'h31 == _T_241[7:0] ? 4'h0 : _GEN_4077; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4079 = 8'h32 == _T_241[7:0] ? 4'h0 : _GEN_4078; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4080 = 8'h33 == _T_241[7:0] ? 4'h0 : _GEN_4079; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4081 = 8'h34 == _T_241[7:0] ? 4'h0 : _GEN_4080; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4082 = 8'h35 == _T_241[7:0] ? 4'h0 : _GEN_4081; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4083 = 8'h36 == _T_241[7:0] ? 4'h0 : _GEN_4082; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4084 = 8'h37 == _T_241[7:0] ? 4'h0 : _GEN_4083; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4085 = 8'h38 == _T_241[7:0] ? 4'hf : _GEN_4084; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4086 = 8'h39 == _T_241[7:0] ? 4'hf : _GEN_4085; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4087 = 8'h3a == _T_241[7:0] ? 4'hf : _GEN_4086; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4088 = 8'h3b == _T_241[7:0] ? 4'hf : _GEN_4087; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4089 = 8'h3c == _T_241[7:0] ? 4'hf : _GEN_4088; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4090 = 8'h3d == _T_241[7:0] ? 4'hf : _GEN_4089; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4091 = 8'h3e == _T_241[7:0] ? 4'hf : _GEN_4090; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4092 = 8'h3f == _T_241[7:0] ? 4'hf : _GEN_4091; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4093 = 8'h40 == _T_241[7:0] ? 4'h0 : _GEN_4092; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4094 = 8'h41 == _T_241[7:0] ? 4'h0 : _GEN_4093; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4095 = 8'h42 == _T_241[7:0] ? 4'h0 : _GEN_4094; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4096 = 8'h43 == _T_241[7:0] ? 4'h0 : _GEN_4095; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4097 = 8'h44 == _T_241[7:0] ? 4'h0 : _GEN_4096; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4098 = 8'h45 == _T_241[7:0] ? 4'h0 : _GEN_4097; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4099 = 8'h46 == _T_241[7:0] ? 4'h0 : _GEN_4098; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4100 = 8'h47 == _T_241[7:0] ? 4'h0 : _GEN_4099; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4101 = 8'h48 == _T_241[7:0] ? 4'hf : _GEN_4100; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4102 = 8'h49 == _T_241[7:0] ? 4'hf : _GEN_4101; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4103 = 8'h4a == _T_241[7:0] ? 4'hf : _GEN_4102; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4104 = 8'h4b == _T_241[7:0] ? 4'hf : _GEN_4103; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4105 = 8'h4c == _T_241[7:0] ? 4'hf : _GEN_4104; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4106 = 8'h4d == _T_241[7:0] ? 4'hf : _GEN_4105; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4107 = 8'h4e == _T_241[7:0] ? 4'hf : _GEN_4106; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4108 = 8'h4f == _T_241[7:0] ? 4'hf : _GEN_4107; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4109 = 8'h50 == _T_241[7:0] ? 4'h0 : _GEN_4108; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4110 = 8'h51 == _T_241[7:0] ? 4'h0 : _GEN_4109; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4111 = 8'h52 == _T_241[7:0] ? 4'h0 : _GEN_4110; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4112 = 8'h53 == _T_241[7:0] ? 4'h0 : _GEN_4111; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4113 = 8'h54 == _T_241[7:0] ? 4'h0 : _GEN_4112; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4114 = 8'h55 == _T_241[7:0] ? 4'h0 : _GEN_4113; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4115 = 8'h56 == _T_241[7:0] ? 4'h0 : _GEN_4114; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4116 = 8'h57 == _T_241[7:0] ? 4'h0 : _GEN_4115; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4117 = 8'h58 == _T_241[7:0] ? 4'hf : _GEN_4116; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4118 = 8'h59 == _T_241[7:0] ? 4'hf : _GEN_4117; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4119 = 8'h5a == _T_241[7:0] ? 4'hf : _GEN_4118; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4120 = 8'h5b == _T_241[7:0] ? 4'hf : _GEN_4119; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4121 = 8'h5c == _T_241[7:0] ? 4'hf : _GEN_4120; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4122 = 8'h5d == _T_241[7:0] ? 4'hf : _GEN_4121; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4123 = 8'h5e == _T_241[7:0] ? 4'hf : _GEN_4122; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4124 = 8'h5f == _T_241[7:0] ? 4'hf : _GEN_4123; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4125 = 8'h60 == _T_241[7:0] ? 4'h0 : _GEN_4124; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4126 = 8'h61 == _T_241[7:0] ? 4'h0 : _GEN_4125; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4127 = 8'h62 == _T_241[7:0] ? 4'h0 : _GEN_4126; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4128 = 8'h63 == _T_241[7:0] ? 4'h0 : _GEN_4127; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4129 = 8'h64 == _T_241[7:0] ? 4'h0 : _GEN_4128; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4130 = 8'h65 == _T_241[7:0] ? 4'h0 : _GEN_4129; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4131 = 8'h66 == _T_241[7:0] ? 4'h0 : _GEN_4130; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4132 = 8'h67 == _T_241[7:0] ? 4'h0 : _GEN_4131; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4133 = 8'h68 == _T_241[7:0] ? 4'hf : _GEN_4132; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4134 = 8'h69 == _T_241[7:0] ? 4'hf : _GEN_4133; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4135 = 8'h6a == _T_241[7:0] ? 4'hf : _GEN_4134; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4136 = 8'h6b == _T_241[7:0] ? 4'hf : _GEN_4135; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4137 = 8'h6c == _T_241[7:0] ? 4'hf : _GEN_4136; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4138 = 8'h6d == _T_241[7:0] ? 4'hf : _GEN_4137; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4139 = 8'h6e == _T_241[7:0] ? 4'hf : _GEN_4138; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4140 = 8'h6f == _T_241[7:0] ? 4'hf : _GEN_4139; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4141 = 8'h70 == _T_241[7:0] ? 4'h0 : _GEN_4140; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4142 = 8'h71 == _T_241[7:0] ? 4'h0 : _GEN_4141; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4143 = 8'h72 == _T_241[7:0] ? 4'h0 : _GEN_4142; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4144 = 8'h73 == _T_241[7:0] ? 4'h0 : _GEN_4143; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4145 = 8'h74 == _T_241[7:0] ? 4'h0 : _GEN_4144; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4146 = 8'h75 == _T_241[7:0] ? 4'h0 : _GEN_4145; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4147 = 8'h76 == _T_241[7:0] ? 4'h0 : _GEN_4146; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4148 = 8'h77 == _T_241[7:0] ? 4'h0 : _GEN_4147; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4149 = 8'h78 == _T_241[7:0] ? 4'hf : _GEN_4148; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4150 = 8'h79 == _T_241[7:0] ? 4'hf : _GEN_4149; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4151 = 8'h7a == _T_241[7:0] ? 4'hf : _GEN_4150; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4152 = 8'h7b == _T_241[7:0] ? 4'hf : _GEN_4151; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4153 = 8'h7c == _T_241[7:0] ? 4'hf : _GEN_4152; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4154 = 8'h7d == _T_241[7:0] ? 4'hf : _GEN_4153; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4155 = 8'h7e == _T_241[7:0] ? 4'hf : _GEN_4154; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4156 = 8'h7f == _T_241[7:0] ? 4'hf : _GEN_4155; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4157 = 8'h80 == _T_241[7:0] ? 4'h0 : _GEN_4156; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4158 = 8'h81 == _T_241[7:0] ? 4'h0 : _GEN_4157; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4159 = 8'h82 == _T_241[7:0] ? 4'h0 : _GEN_4158; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4160 = 8'h83 == _T_241[7:0] ? 4'h0 : _GEN_4159; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4161 = 8'h84 == _T_241[7:0] ? 4'h0 : _GEN_4160; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4162 = 8'h85 == _T_241[7:0] ? 4'h0 : _GEN_4161; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4163 = 8'h86 == _T_241[7:0] ? 4'h0 : _GEN_4162; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4164 = 8'h87 == _T_241[7:0] ? 4'h0 : _GEN_4163; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4165 = 8'h88 == _T_241[7:0] ? 4'hf : _GEN_4164; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4166 = 8'h89 == _T_241[7:0] ? 4'hf : _GEN_4165; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4167 = 8'h8a == _T_241[7:0] ? 4'hf : _GEN_4166; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4168 = 8'h8b == _T_241[7:0] ? 4'hf : _GEN_4167; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4169 = 8'h8c == _T_241[7:0] ? 4'hf : _GEN_4168; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4170 = 8'h8d == _T_241[7:0] ? 4'hf : _GEN_4169; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4171 = 8'h8e == _T_241[7:0] ? 4'hf : _GEN_4170; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4172 = 8'h8f == _T_241[7:0] ? 4'hf : _GEN_4171; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4173 = 8'h90 == _T_241[7:0] ? 4'h0 : _GEN_4172; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4174 = 8'h91 == _T_241[7:0] ? 4'h0 : _GEN_4173; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4175 = 8'h92 == _T_241[7:0] ? 4'h0 : _GEN_4174; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4176 = 8'h93 == _T_241[7:0] ? 4'h0 : _GEN_4175; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4177 = 8'h94 == _T_241[7:0] ? 4'h0 : _GEN_4176; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4178 = 8'h95 == _T_241[7:0] ? 4'h0 : _GEN_4177; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4179 = 8'h96 == _T_241[7:0] ? 4'h0 : _GEN_4178; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4180 = 8'h97 == _T_241[7:0] ? 4'h0 : _GEN_4179; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4181 = 8'h98 == _T_241[7:0] ? 4'hf : _GEN_4180; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4182 = 8'h99 == _T_241[7:0] ? 4'hf : _GEN_4181; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4183 = 8'h9a == _T_241[7:0] ? 4'hf : _GEN_4182; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4184 = 8'h9b == _T_241[7:0] ? 4'hf : _GEN_4183; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4185 = 8'h9c == _T_241[7:0] ? 4'hf : _GEN_4184; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4186 = 8'h9d == _T_241[7:0] ? 4'hf : _GEN_4185; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4187 = 8'h9e == _T_241[7:0] ? 4'hf : _GEN_4186; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4188 = 8'h9f == _T_241[7:0] ? 4'hf : _GEN_4187; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4189 = 8'ha0 == _T_241[7:0] ? 4'h0 : _GEN_4188; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4190 = 8'ha1 == _T_241[7:0] ? 4'h0 : _GEN_4189; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4191 = 8'ha2 == _T_241[7:0] ? 4'h0 : _GEN_4190; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4192 = 8'ha3 == _T_241[7:0] ? 4'h0 : _GEN_4191; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4193 = 8'ha4 == _T_241[7:0] ? 4'h0 : _GEN_4192; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4194 = 8'ha5 == _T_241[7:0] ? 4'h0 : _GEN_4193; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4195 = 8'ha6 == _T_241[7:0] ? 4'h0 : _GEN_4194; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4196 = 8'ha7 == _T_241[7:0] ? 4'h0 : _GEN_4195; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4197 = 8'ha8 == _T_241[7:0] ? 4'hf : _GEN_4196; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4198 = 8'ha9 == _T_241[7:0] ? 4'hf : _GEN_4197; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4199 = 8'haa == _T_241[7:0] ? 4'hf : _GEN_4198; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4200 = 8'hab == _T_241[7:0] ? 4'hf : _GEN_4199; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4201 = 8'hac == _T_241[7:0] ? 4'hf : _GEN_4200; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4202 = 8'had == _T_241[7:0] ? 4'hf : _GEN_4201; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4203 = 8'hae == _T_241[7:0] ? 4'hf : _GEN_4202; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4204 = 8'haf == _T_241[7:0] ? 4'hf : _GEN_4203; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4205 = 8'hb0 == _T_241[7:0] ? 4'h0 : _GEN_4204; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4206 = 8'hb1 == _T_241[7:0] ? 4'h0 : _GEN_4205; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4207 = 8'hb2 == _T_241[7:0] ? 4'h0 : _GEN_4206; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4208 = 8'hb3 == _T_241[7:0] ? 4'h0 : _GEN_4207; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4209 = 8'hb4 == _T_241[7:0] ? 4'h0 : _GEN_4208; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4210 = 8'hb5 == _T_241[7:0] ? 4'h0 : _GEN_4209; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4211 = 8'hb6 == _T_241[7:0] ? 4'h0 : _GEN_4210; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4212 = 8'hb7 == _T_241[7:0] ? 4'h0 : _GEN_4211; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4213 = 8'hb8 == _T_241[7:0] ? 4'hf : _GEN_4212; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4214 = 8'hb9 == _T_241[7:0] ? 4'hf : _GEN_4213; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4215 = 8'hba == _T_241[7:0] ? 4'hf : _GEN_4214; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4216 = 8'hbb == _T_241[7:0] ? 4'hf : _GEN_4215; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4217 = 8'hbc == _T_241[7:0] ? 4'hf : _GEN_4216; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4218 = 8'hbd == _T_241[7:0] ? 4'hf : _GEN_4217; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4219 = 8'hbe == _T_241[7:0] ? 4'hf : _GEN_4218; // @[Filter.scala 160:142]
  wire [3:0] _GEN_4220 = 8'hbf == _T_241[7:0] ? 4'hf : _GEN_4219; // @[Filter.scala 160:142]
  wire [7:0] _T_255 = _GEN_4220 * 4'ha; // @[Filter.scala 160:142]
  wire [10:0] _GEN_9907 = {{3'd0}, _T_255}; // @[Filter.scala 160:109]
  wire [10:0] _T_257 = _T_250 + _GEN_9907; // @[Filter.scala 160:109]
  wire [10:0] _T_258 = _T_257 / 11'h64; // @[Filter.scala 160:150]
  wire  _T_260 = _T_231 >= 5'h10; // @[Filter.scala 163:31]
  wire  _T_264 = _T_238 >= 32'hc; // @[Filter.scala 163:63]
  wire  _T_265 = _T_260 | _T_264; // @[Filter.scala 163:58]
  wire [10:0] _GEN_4413 = io_SPI_distort ? _T_258 : {{7'd0}, _GEN_3836}; // @[Filter.scala 165:35]
  wire [10:0] _GEN_4414 = _T_265 ? 11'h0 : _GEN_4413; // @[Filter.scala 163:80]
  wire [10:0] _GEN_4607 = io_SPI_distort ? _T_258 : {{7'd0}, _GEN_4028}; // @[Filter.scala 165:35]
  wire [10:0] _GEN_4608 = _T_265 ? 11'h0 : _GEN_4607; // @[Filter.scala 163:80]
  wire [10:0] _GEN_4801 = io_SPI_distort ? _T_258 : {{7'd0}, _GEN_4220}; // @[Filter.scala 165:35]
  wire [10:0] _GEN_4802 = _T_265 ? 11'h0 : _GEN_4801; // @[Filter.scala 163:80]
  wire [31:0] _T_293 = pixelIndex + 32'h4; // @[Filter.scala 158:31]
  wire [31:0] _GEN_4 = _T_293 % 32'h10; // @[Filter.scala 158:38]
  wire [4:0] _T_294 = _GEN_4[4:0]; // @[Filter.scala 158:38]
  wire [4:0] _T_296 = _T_294 + _GEN_9863; // @[Filter.scala 158:53]
  wire [4:0] _T_298 = _T_296 - 5'h1; // @[Filter.scala 158:69]
  wire [31:0] _T_301 = _T_293 / 32'h10; // @[Filter.scala 159:38]
  wire [31:0] _T_303 = _T_301 + _GEN_9864; // @[Filter.scala 159:53]
  wire [31:0] _T_305 = _T_303 - 32'h1; // @[Filter.scala 159:69]
  wire [36:0] _T_306 = _T_305 * 32'h10; // @[Filter.scala 160:42]
  wire [36:0] _GEN_9913 = {{32'd0}, _T_298}; // @[Filter.scala 160:57]
  wire [36:0] _T_308 = _T_306 + _GEN_9913; // @[Filter.scala 160:57]
  wire [3:0] _GEN_4811 = 8'h8 == _T_308[7:0] ? 4'h0 : 4'hf; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4812 = 8'h9 == _T_308[7:0] ? 4'h0 : _GEN_4811; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4813 = 8'ha == _T_308[7:0] ? 4'h0 : _GEN_4812; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4814 = 8'hb == _T_308[7:0] ? 4'h0 : _GEN_4813; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4815 = 8'hc == _T_308[7:0] ? 4'h0 : _GEN_4814; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4816 = 8'hd == _T_308[7:0] ? 4'h0 : _GEN_4815; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4817 = 8'he == _T_308[7:0] ? 4'h0 : _GEN_4816; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4818 = 8'hf == _T_308[7:0] ? 4'h0 : _GEN_4817; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4819 = 8'h10 == _T_308[7:0] ? 4'hf : _GEN_4818; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4820 = 8'h11 == _T_308[7:0] ? 4'hf : _GEN_4819; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4821 = 8'h12 == _T_308[7:0] ? 4'hf : _GEN_4820; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4822 = 8'h13 == _T_308[7:0] ? 4'hf : _GEN_4821; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4823 = 8'h14 == _T_308[7:0] ? 4'hf : _GEN_4822; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4824 = 8'h15 == _T_308[7:0] ? 4'hf : _GEN_4823; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4825 = 8'h16 == _T_308[7:0] ? 4'hf : _GEN_4824; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4826 = 8'h17 == _T_308[7:0] ? 4'hf : _GEN_4825; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4827 = 8'h18 == _T_308[7:0] ? 4'h0 : _GEN_4826; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4828 = 8'h19 == _T_308[7:0] ? 4'h0 : _GEN_4827; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4829 = 8'h1a == _T_308[7:0] ? 4'h0 : _GEN_4828; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4830 = 8'h1b == _T_308[7:0] ? 4'h0 : _GEN_4829; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4831 = 8'h1c == _T_308[7:0] ? 4'h0 : _GEN_4830; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4832 = 8'h1d == _T_308[7:0] ? 4'h0 : _GEN_4831; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4833 = 8'h1e == _T_308[7:0] ? 4'h0 : _GEN_4832; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4834 = 8'h1f == _T_308[7:0] ? 4'h0 : _GEN_4833; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4835 = 8'h20 == _T_308[7:0] ? 4'hf : _GEN_4834; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4836 = 8'h21 == _T_308[7:0] ? 4'hf : _GEN_4835; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4837 = 8'h22 == _T_308[7:0] ? 4'hf : _GEN_4836; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4838 = 8'h23 == _T_308[7:0] ? 4'hf : _GEN_4837; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4839 = 8'h24 == _T_308[7:0] ? 4'hf : _GEN_4838; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4840 = 8'h25 == _T_308[7:0] ? 4'hf : _GEN_4839; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4841 = 8'h26 == _T_308[7:0] ? 4'hf : _GEN_4840; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4842 = 8'h27 == _T_308[7:0] ? 4'hf : _GEN_4841; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4843 = 8'h28 == _T_308[7:0] ? 4'h0 : _GEN_4842; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4844 = 8'h29 == _T_308[7:0] ? 4'h0 : _GEN_4843; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4845 = 8'h2a == _T_308[7:0] ? 4'h0 : _GEN_4844; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4846 = 8'h2b == _T_308[7:0] ? 4'h0 : _GEN_4845; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4847 = 8'h2c == _T_308[7:0] ? 4'h0 : _GEN_4846; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4848 = 8'h2d == _T_308[7:0] ? 4'h0 : _GEN_4847; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4849 = 8'h2e == _T_308[7:0] ? 4'h0 : _GEN_4848; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4850 = 8'h2f == _T_308[7:0] ? 4'h0 : _GEN_4849; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4851 = 8'h30 == _T_308[7:0] ? 4'hf : _GEN_4850; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4852 = 8'h31 == _T_308[7:0] ? 4'hf : _GEN_4851; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4853 = 8'h32 == _T_308[7:0] ? 4'hf : _GEN_4852; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4854 = 8'h33 == _T_308[7:0] ? 4'hf : _GEN_4853; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4855 = 8'h34 == _T_308[7:0] ? 4'hf : _GEN_4854; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4856 = 8'h35 == _T_308[7:0] ? 4'hf : _GEN_4855; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4857 = 8'h36 == _T_308[7:0] ? 4'hf : _GEN_4856; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4858 = 8'h37 == _T_308[7:0] ? 4'hf : _GEN_4857; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4859 = 8'h38 == _T_308[7:0] ? 4'h0 : _GEN_4858; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4860 = 8'h39 == _T_308[7:0] ? 4'h0 : _GEN_4859; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4861 = 8'h3a == _T_308[7:0] ? 4'h0 : _GEN_4860; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4862 = 8'h3b == _T_308[7:0] ? 4'h0 : _GEN_4861; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4863 = 8'h3c == _T_308[7:0] ? 4'h0 : _GEN_4862; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4864 = 8'h3d == _T_308[7:0] ? 4'h0 : _GEN_4863; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4865 = 8'h3e == _T_308[7:0] ? 4'h0 : _GEN_4864; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4866 = 8'h3f == _T_308[7:0] ? 4'h0 : _GEN_4865; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4867 = 8'h40 == _T_308[7:0] ? 4'hf : _GEN_4866; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4868 = 8'h41 == _T_308[7:0] ? 4'hf : _GEN_4867; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4869 = 8'h42 == _T_308[7:0] ? 4'hf : _GEN_4868; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4870 = 8'h43 == _T_308[7:0] ? 4'hf : _GEN_4869; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4871 = 8'h44 == _T_308[7:0] ? 4'hf : _GEN_4870; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4872 = 8'h45 == _T_308[7:0] ? 4'hf : _GEN_4871; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4873 = 8'h46 == _T_308[7:0] ? 4'hf : _GEN_4872; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4874 = 8'h47 == _T_308[7:0] ? 4'hf : _GEN_4873; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4875 = 8'h48 == _T_308[7:0] ? 4'h0 : _GEN_4874; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4876 = 8'h49 == _T_308[7:0] ? 4'h0 : _GEN_4875; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4877 = 8'h4a == _T_308[7:0] ? 4'h0 : _GEN_4876; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4878 = 8'h4b == _T_308[7:0] ? 4'h0 : _GEN_4877; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4879 = 8'h4c == _T_308[7:0] ? 4'h0 : _GEN_4878; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4880 = 8'h4d == _T_308[7:0] ? 4'h0 : _GEN_4879; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4881 = 8'h4e == _T_308[7:0] ? 4'h0 : _GEN_4880; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4882 = 8'h4f == _T_308[7:0] ? 4'h0 : _GEN_4881; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4883 = 8'h50 == _T_308[7:0] ? 4'hf : _GEN_4882; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4884 = 8'h51 == _T_308[7:0] ? 4'hf : _GEN_4883; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4885 = 8'h52 == _T_308[7:0] ? 4'hf : _GEN_4884; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4886 = 8'h53 == _T_308[7:0] ? 4'hf : _GEN_4885; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4887 = 8'h54 == _T_308[7:0] ? 4'hf : _GEN_4886; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4888 = 8'h55 == _T_308[7:0] ? 4'hf : _GEN_4887; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4889 = 8'h56 == _T_308[7:0] ? 4'hf : _GEN_4888; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4890 = 8'h57 == _T_308[7:0] ? 4'hf : _GEN_4889; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4891 = 8'h58 == _T_308[7:0] ? 4'h0 : _GEN_4890; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4892 = 8'h59 == _T_308[7:0] ? 4'h0 : _GEN_4891; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4893 = 8'h5a == _T_308[7:0] ? 4'h0 : _GEN_4892; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4894 = 8'h5b == _T_308[7:0] ? 4'h0 : _GEN_4893; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4895 = 8'h5c == _T_308[7:0] ? 4'h0 : _GEN_4894; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4896 = 8'h5d == _T_308[7:0] ? 4'h0 : _GEN_4895; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4897 = 8'h5e == _T_308[7:0] ? 4'h0 : _GEN_4896; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4898 = 8'h5f == _T_308[7:0] ? 4'h0 : _GEN_4897; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4899 = 8'h60 == _T_308[7:0] ? 4'h0 : _GEN_4898; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4900 = 8'h61 == _T_308[7:0] ? 4'h0 : _GEN_4899; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4901 = 8'h62 == _T_308[7:0] ? 4'h0 : _GEN_4900; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4902 = 8'h63 == _T_308[7:0] ? 4'h0 : _GEN_4901; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4903 = 8'h64 == _T_308[7:0] ? 4'h0 : _GEN_4902; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4904 = 8'h65 == _T_308[7:0] ? 4'h0 : _GEN_4903; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4905 = 8'h66 == _T_308[7:0] ? 4'h0 : _GEN_4904; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4906 = 8'h67 == _T_308[7:0] ? 4'h0 : _GEN_4905; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4907 = 8'h68 == _T_308[7:0] ? 4'hf : _GEN_4906; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4908 = 8'h69 == _T_308[7:0] ? 4'hf : _GEN_4907; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4909 = 8'h6a == _T_308[7:0] ? 4'hf : _GEN_4908; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4910 = 8'h6b == _T_308[7:0] ? 4'hf : _GEN_4909; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4911 = 8'h6c == _T_308[7:0] ? 4'hf : _GEN_4910; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4912 = 8'h6d == _T_308[7:0] ? 4'hf : _GEN_4911; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4913 = 8'h6e == _T_308[7:0] ? 4'hf : _GEN_4912; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4914 = 8'h6f == _T_308[7:0] ? 4'hf : _GEN_4913; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4915 = 8'h70 == _T_308[7:0] ? 4'h0 : _GEN_4914; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4916 = 8'h71 == _T_308[7:0] ? 4'h0 : _GEN_4915; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4917 = 8'h72 == _T_308[7:0] ? 4'h0 : _GEN_4916; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4918 = 8'h73 == _T_308[7:0] ? 4'h0 : _GEN_4917; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4919 = 8'h74 == _T_308[7:0] ? 4'h0 : _GEN_4918; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4920 = 8'h75 == _T_308[7:0] ? 4'h0 : _GEN_4919; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4921 = 8'h76 == _T_308[7:0] ? 4'h0 : _GEN_4920; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4922 = 8'h77 == _T_308[7:0] ? 4'h0 : _GEN_4921; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4923 = 8'h78 == _T_308[7:0] ? 4'hf : _GEN_4922; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4924 = 8'h79 == _T_308[7:0] ? 4'hf : _GEN_4923; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4925 = 8'h7a == _T_308[7:0] ? 4'hf : _GEN_4924; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4926 = 8'h7b == _T_308[7:0] ? 4'hf : _GEN_4925; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4927 = 8'h7c == _T_308[7:0] ? 4'hf : _GEN_4926; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4928 = 8'h7d == _T_308[7:0] ? 4'hf : _GEN_4927; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4929 = 8'h7e == _T_308[7:0] ? 4'hf : _GEN_4928; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4930 = 8'h7f == _T_308[7:0] ? 4'hf : _GEN_4929; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4931 = 8'h80 == _T_308[7:0] ? 4'h0 : _GEN_4930; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4932 = 8'h81 == _T_308[7:0] ? 4'h0 : _GEN_4931; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4933 = 8'h82 == _T_308[7:0] ? 4'h0 : _GEN_4932; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4934 = 8'h83 == _T_308[7:0] ? 4'h0 : _GEN_4933; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4935 = 8'h84 == _T_308[7:0] ? 4'h0 : _GEN_4934; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4936 = 8'h85 == _T_308[7:0] ? 4'h0 : _GEN_4935; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4937 = 8'h86 == _T_308[7:0] ? 4'h0 : _GEN_4936; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4938 = 8'h87 == _T_308[7:0] ? 4'h0 : _GEN_4937; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4939 = 8'h88 == _T_308[7:0] ? 4'hf : _GEN_4938; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4940 = 8'h89 == _T_308[7:0] ? 4'hf : _GEN_4939; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4941 = 8'h8a == _T_308[7:0] ? 4'hf : _GEN_4940; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4942 = 8'h8b == _T_308[7:0] ? 4'hf : _GEN_4941; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4943 = 8'h8c == _T_308[7:0] ? 4'hf : _GEN_4942; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4944 = 8'h8d == _T_308[7:0] ? 4'hf : _GEN_4943; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4945 = 8'h8e == _T_308[7:0] ? 4'hf : _GEN_4944; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4946 = 8'h8f == _T_308[7:0] ? 4'hf : _GEN_4945; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4947 = 8'h90 == _T_308[7:0] ? 4'h0 : _GEN_4946; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4948 = 8'h91 == _T_308[7:0] ? 4'h0 : _GEN_4947; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4949 = 8'h92 == _T_308[7:0] ? 4'h0 : _GEN_4948; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4950 = 8'h93 == _T_308[7:0] ? 4'h0 : _GEN_4949; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4951 = 8'h94 == _T_308[7:0] ? 4'h0 : _GEN_4950; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4952 = 8'h95 == _T_308[7:0] ? 4'h0 : _GEN_4951; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4953 = 8'h96 == _T_308[7:0] ? 4'h0 : _GEN_4952; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4954 = 8'h97 == _T_308[7:0] ? 4'h0 : _GEN_4953; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4955 = 8'h98 == _T_308[7:0] ? 4'hf : _GEN_4954; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4956 = 8'h99 == _T_308[7:0] ? 4'hf : _GEN_4955; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4957 = 8'h9a == _T_308[7:0] ? 4'hf : _GEN_4956; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4958 = 8'h9b == _T_308[7:0] ? 4'hf : _GEN_4957; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4959 = 8'h9c == _T_308[7:0] ? 4'hf : _GEN_4958; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4960 = 8'h9d == _T_308[7:0] ? 4'hf : _GEN_4959; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4961 = 8'h9e == _T_308[7:0] ? 4'hf : _GEN_4960; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4962 = 8'h9f == _T_308[7:0] ? 4'hf : _GEN_4961; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4963 = 8'ha0 == _T_308[7:0] ? 4'h0 : _GEN_4962; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4964 = 8'ha1 == _T_308[7:0] ? 4'h0 : _GEN_4963; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4965 = 8'ha2 == _T_308[7:0] ? 4'h0 : _GEN_4964; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4966 = 8'ha3 == _T_308[7:0] ? 4'h0 : _GEN_4965; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4967 = 8'ha4 == _T_308[7:0] ? 4'h0 : _GEN_4966; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4968 = 8'ha5 == _T_308[7:0] ? 4'h0 : _GEN_4967; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4969 = 8'ha6 == _T_308[7:0] ? 4'h0 : _GEN_4968; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4970 = 8'ha7 == _T_308[7:0] ? 4'h0 : _GEN_4969; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4971 = 8'ha8 == _T_308[7:0] ? 4'hf : _GEN_4970; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4972 = 8'ha9 == _T_308[7:0] ? 4'hf : _GEN_4971; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4973 = 8'haa == _T_308[7:0] ? 4'hf : _GEN_4972; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4974 = 8'hab == _T_308[7:0] ? 4'hf : _GEN_4973; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4975 = 8'hac == _T_308[7:0] ? 4'hf : _GEN_4974; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4976 = 8'had == _T_308[7:0] ? 4'hf : _GEN_4975; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4977 = 8'hae == _T_308[7:0] ? 4'hf : _GEN_4976; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4978 = 8'haf == _T_308[7:0] ? 4'hf : _GEN_4977; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4979 = 8'hb0 == _T_308[7:0] ? 4'h0 : _GEN_4978; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4980 = 8'hb1 == _T_308[7:0] ? 4'h0 : _GEN_4979; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4981 = 8'hb2 == _T_308[7:0] ? 4'h0 : _GEN_4980; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4982 = 8'hb3 == _T_308[7:0] ? 4'h0 : _GEN_4981; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4983 = 8'hb4 == _T_308[7:0] ? 4'h0 : _GEN_4982; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4984 = 8'hb5 == _T_308[7:0] ? 4'h0 : _GEN_4983; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4985 = 8'hb6 == _T_308[7:0] ? 4'h0 : _GEN_4984; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4986 = 8'hb7 == _T_308[7:0] ? 4'h0 : _GEN_4985; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4987 = 8'hb8 == _T_308[7:0] ? 4'hf : _GEN_4986; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4988 = 8'hb9 == _T_308[7:0] ? 4'hf : _GEN_4987; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4989 = 8'hba == _T_308[7:0] ? 4'hf : _GEN_4988; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4990 = 8'hbb == _T_308[7:0] ? 4'hf : _GEN_4989; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4991 = 8'hbc == _T_308[7:0] ? 4'hf : _GEN_4990; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4992 = 8'hbd == _T_308[7:0] ? 4'hf : _GEN_4991; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4993 = 8'hbe == _T_308[7:0] ? 4'hf : _GEN_4992; // @[Filter.scala 160:62]
  wire [3:0] _GEN_4994 = 8'hbf == _T_308[7:0] ? 4'hf : _GEN_4993; // @[Filter.scala 160:62]
  wire [4:0] _GEN_9914 = {{1'd0}, _GEN_4994}; // @[Filter.scala 160:62]
  wire [8:0] _T_310 = _GEN_9914 * 5'h14; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5091 = 8'h60 == _T_308[7:0] ? 4'hf : 4'h0; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5092 = 8'h61 == _T_308[7:0] ? 4'hf : _GEN_5091; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5093 = 8'h62 == _T_308[7:0] ? 4'hf : _GEN_5092; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5094 = 8'h63 == _T_308[7:0] ? 4'hf : _GEN_5093; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5095 = 8'h64 == _T_308[7:0] ? 4'hf : _GEN_5094; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5096 = 8'h65 == _T_308[7:0] ? 4'hf : _GEN_5095; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5097 = 8'h66 == _T_308[7:0] ? 4'hf : _GEN_5096; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5098 = 8'h67 == _T_308[7:0] ? 4'hf : _GEN_5097; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5099 = 8'h68 == _T_308[7:0] ? 4'hf : _GEN_5098; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5100 = 8'h69 == _T_308[7:0] ? 4'hf : _GEN_5099; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5101 = 8'h6a == _T_308[7:0] ? 4'hf : _GEN_5100; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5102 = 8'h6b == _T_308[7:0] ? 4'hf : _GEN_5101; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5103 = 8'h6c == _T_308[7:0] ? 4'hf : _GEN_5102; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5104 = 8'h6d == _T_308[7:0] ? 4'hf : _GEN_5103; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5105 = 8'h6e == _T_308[7:0] ? 4'hf : _GEN_5104; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5106 = 8'h6f == _T_308[7:0] ? 4'hf : _GEN_5105; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5107 = 8'h70 == _T_308[7:0] ? 4'hf : _GEN_5106; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5108 = 8'h71 == _T_308[7:0] ? 4'hf : _GEN_5107; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5109 = 8'h72 == _T_308[7:0] ? 4'hf : _GEN_5108; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5110 = 8'h73 == _T_308[7:0] ? 4'hf : _GEN_5109; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5111 = 8'h74 == _T_308[7:0] ? 4'hf : _GEN_5110; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5112 = 8'h75 == _T_308[7:0] ? 4'hf : _GEN_5111; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5113 = 8'h76 == _T_308[7:0] ? 4'hf : _GEN_5112; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5114 = 8'h77 == _T_308[7:0] ? 4'hf : _GEN_5113; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5115 = 8'h78 == _T_308[7:0] ? 4'hf : _GEN_5114; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5116 = 8'h79 == _T_308[7:0] ? 4'hf : _GEN_5115; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5117 = 8'h7a == _T_308[7:0] ? 4'hf : _GEN_5116; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5118 = 8'h7b == _T_308[7:0] ? 4'hf : _GEN_5117; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5119 = 8'h7c == _T_308[7:0] ? 4'hf : _GEN_5118; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5120 = 8'h7d == _T_308[7:0] ? 4'hf : _GEN_5119; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5121 = 8'h7e == _T_308[7:0] ? 4'hf : _GEN_5120; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5122 = 8'h7f == _T_308[7:0] ? 4'hf : _GEN_5121; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5123 = 8'h80 == _T_308[7:0] ? 4'hf : _GEN_5122; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5124 = 8'h81 == _T_308[7:0] ? 4'hf : _GEN_5123; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5125 = 8'h82 == _T_308[7:0] ? 4'hf : _GEN_5124; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5126 = 8'h83 == _T_308[7:0] ? 4'hf : _GEN_5125; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5127 = 8'h84 == _T_308[7:0] ? 4'hf : _GEN_5126; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5128 = 8'h85 == _T_308[7:0] ? 4'hf : _GEN_5127; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5129 = 8'h86 == _T_308[7:0] ? 4'hf : _GEN_5128; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5130 = 8'h87 == _T_308[7:0] ? 4'hf : _GEN_5129; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5131 = 8'h88 == _T_308[7:0] ? 4'hf : _GEN_5130; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5132 = 8'h89 == _T_308[7:0] ? 4'hf : _GEN_5131; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5133 = 8'h8a == _T_308[7:0] ? 4'hf : _GEN_5132; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5134 = 8'h8b == _T_308[7:0] ? 4'hf : _GEN_5133; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5135 = 8'h8c == _T_308[7:0] ? 4'hf : _GEN_5134; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5136 = 8'h8d == _T_308[7:0] ? 4'hf : _GEN_5135; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5137 = 8'h8e == _T_308[7:0] ? 4'hf : _GEN_5136; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5138 = 8'h8f == _T_308[7:0] ? 4'hf : _GEN_5137; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5139 = 8'h90 == _T_308[7:0] ? 4'hf : _GEN_5138; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5140 = 8'h91 == _T_308[7:0] ? 4'hf : _GEN_5139; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5141 = 8'h92 == _T_308[7:0] ? 4'hf : _GEN_5140; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5142 = 8'h93 == _T_308[7:0] ? 4'hf : _GEN_5141; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5143 = 8'h94 == _T_308[7:0] ? 4'hf : _GEN_5142; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5144 = 8'h95 == _T_308[7:0] ? 4'hf : _GEN_5143; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5145 = 8'h96 == _T_308[7:0] ? 4'hf : _GEN_5144; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5146 = 8'h97 == _T_308[7:0] ? 4'hf : _GEN_5145; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5147 = 8'h98 == _T_308[7:0] ? 4'hf : _GEN_5146; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5148 = 8'h99 == _T_308[7:0] ? 4'hf : _GEN_5147; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5149 = 8'h9a == _T_308[7:0] ? 4'hf : _GEN_5148; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5150 = 8'h9b == _T_308[7:0] ? 4'hf : _GEN_5149; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5151 = 8'h9c == _T_308[7:0] ? 4'hf : _GEN_5150; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5152 = 8'h9d == _T_308[7:0] ? 4'hf : _GEN_5151; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5153 = 8'h9e == _T_308[7:0] ? 4'hf : _GEN_5152; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5154 = 8'h9f == _T_308[7:0] ? 4'hf : _GEN_5153; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5155 = 8'ha0 == _T_308[7:0] ? 4'hf : _GEN_5154; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5156 = 8'ha1 == _T_308[7:0] ? 4'hf : _GEN_5155; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5157 = 8'ha2 == _T_308[7:0] ? 4'hf : _GEN_5156; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5158 = 8'ha3 == _T_308[7:0] ? 4'hf : _GEN_5157; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5159 = 8'ha4 == _T_308[7:0] ? 4'hf : _GEN_5158; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5160 = 8'ha5 == _T_308[7:0] ? 4'hf : _GEN_5159; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5161 = 8'ha6 == _T_308[7:0] ? 4'hf : _GEN_5160; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5162 = 8'ha7 == _T_308[7:0] ? 4'hf : _GEN_5161; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5163 = 8'ha8 == _T_308[7:0] ? 4'hf : _GEN_5162; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5164 = 8'ha9 == _T_308[7:0] ? 4'hf : _GEN_5163; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5165 = 8'haa == _T_308[7:0] ? 4'hf : _GEN_5164; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5166 = 8'hab == _T_308[7:0] ? 4'hf : _GEN_5165; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5167 = 8'hac == _T_308[7:0] ? 4'hf : _GEN_5166; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5168 = 8'had == _T_308[7:0] ? 4'hf : _GEN_5167; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5169 = 8'hae == _T_308[7:0] ? 4'hf : _GEN_5168; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5170 = 8'haf == _T_308[7:0] ? 4'hf : _GEN_5169; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5171 = 8'hb0 == _T_308[7:0] ? 4'hf : _GEN_5170; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5172 = 8'hb1 == _T_308[7:0] ? 4'hf : _GEN_5171; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5173 = 8'hb2 == _T_308[7:0] ? 4'hf : _GEN_5172; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5174 = 8'hb3 == _T_308[7:0] ? 4'hf : _GEN_5173; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5175 = 8'hb4 == _T_308[7:0] ? 4'hf : _GEN_5174; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5176 = 8'hb5 == _T_308[7:0] ? 4'hf : _GEN_5175; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5177 = 8'hb6 == _T_308[7:0] ? 4'hf : _GEN_5176; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5178 = 8'hb7 == _T_308[7:0] ? 4'hf : _GEN_5177; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5179 = 8'hb8 == _T_308[7:0] ? 4'hf : _GEN_5178; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5180 = 8'hb9 == _T_308[7:0] ? 4'hf : _GEN_5179; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5181 = 8'hba == _T_308[7:0] ? 4'hf : _GEN_5180; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5182 = 8'hbb == _T_308[7:0] ? 4'hf : _GEN_5181; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5183 = 8'hbc == _T_308[7:0] ? 4'hf : _GEN_5182; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5184 = 8'hbd == _T_308[7:0] ? 4'hf : _GEN_5183; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5185 = 8'hbe == _T_308[7:0] ? 4'hf : _GEN_5184; // @[Filter.scala 160:102]
  wire [3:0] _GEN_5186 = 8'hbf == _T_308[7:0] ? 4'hf : _GEN_5185; // @[Filter.scala 160:102]
  wire [6:0] _GEN_9916 = {{3'd0}, _GEN_5186}; // @[Filter.scala 160:102]
  wire [10:0] _T_315 = _GEN_9916 * 7'h46; // @[Filter.scala 160:102]
  wire [10:0] _GEN_9917 = {{2'd0}, _T_310}; // @[Filter.scala 160:69]
  wire [10:0] _T_317 = _GEN_9917 + _T_315; // @[Filter.scala 160:69]
  wire [3:0] _GEN_5195 = 8'h8 == _T_308[7:0] ? 4'hf : 4'h0; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5196 = 8'h9 == _T_308[7:0] ? 4'hf : _GEN_5195; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5197 = 8'ha == _T_308[7:0] ? 4'hf : _GEN_5196; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5198 = 8'hb == _T_308[7:0] ? 4'hf : _GEN_5197; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5199 = 8'hc == _T_308[7:0] ? 4'hf : _GEN_5198; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5200 = 8'hd == _T_308[7:0] ? 4'hf : _GEN_5199; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5201 = 8'he == _T_308[7:0] ? 4'hf : _GEN_5200; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5202 = 8'hf == _T_308[7:0] ? 4'hf : _GEN_5201; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5203 = 8'h10 == _T_308[7:0] ? 4'h0 : _GEN_5202; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5204 = 8'h11 == _T_308[7:0] ? 4'h0 : _GEN_5203; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5205 = 8'h12 == _T_308[7:0] ? 4'h0 : _GEN_5204; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5206 = 8'h13 == _T_308[7:0] ? 4'h0 : _GEN_5205; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5207 = 8'h14 == _T_308[7:0] ? 4'h0 : _GEN_5206; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5208 = 8'h15 == _T_308[7:0] ? 4'h0 : _GEN_5207; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5209 = 8'h16 == _T_308[7:0] ? 4'h0 : _GEN_5208; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5210 = 8'h17 == _T_308[7:0] ? 4'h0 : _GEN_5209; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5211 = 8'h18 == _T_308[7:0] ? 4'hf : _GEN_5210; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5212 = 8'h19 == _T_308[7:0] ? 4'hf : _GEN_5211; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5213 = 8'h1a == _T_308[7:0] ? 4'hf : _GEN_5212; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5214 = 8'h1b == _T_308[7:0] ? 4'hf : _GEN_5213; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5215 = 8'h1c == _T_308[7:0] ? 4'hf : _GEN_5214; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5216 = 8'h1d == _T_308[7:0] ? 4'hf : _GEN_5215; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5217 = 8'h1e == _T_308[7:0] ? 4'hf : _GEN_5216; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5218 = 8'h1f == _T_308[7:0] ? 4'hf : _GEN_5217; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5219 = 8'h20 == _T_308[7:0] ? 4'h0 : _GEN_5218; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5220 = 8'h21 == _T_308[7:0] ? 4'h0 : _GEN_5219; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5221 = 8'h22 == _T_308[7:0] ? 4'h0 : _GEN_5220; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5222 = 8'h23 == _T_308[7:0] ? 4'h0 : _GEN_5221; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5223 = 8'h24 == _T_308[7:0] ? 4'h0 : _GEN_5222; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5224 = 8'h25 == _T_308[7:0] ? 4'h0 : _GEN_5223; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5225 = 8'h26 == _T_308[7:0] ? 4'h0 : _GEN_5224; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5226 = 8'h27 == _T_308[7:0] ? 4'h0 : _GEN_5225; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5227 = 8'h28 == _T_308[7:0] ? 4'hf : _GEN_5226; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5228 = 8'h29 == _T_308[7:0] ? 4'hf : _GEN_5227; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5229 = 8'h2a == _T_308[7:0] ? 4'hf : _GEN_5228; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5230 = 8'h2b == _T_308[7:0] ? 4'hf : _GEN_5229; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5231 = 8'h2c == _T_308[7:0] ? 4'hf : _GEN_5230; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5232 = 8'h2d == _T_308[7:0] ? 4'hf : _GEN_5231; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5233 = 8'h2e == _T_308[7:0] ? 4'hf : _GEN_5232; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5234 = 8'h2f == _T_308[7:0] ? 4'hf : _GEN_5233; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5235 = 8'h30 == _T_308[7:0] ? 4'h0 : _GEN_5234; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5236 = 8'h31 == _T_308[7:0] ? 4'h0 : _GEN_5235; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5237 = 8'h32 == _T_308[7:0] ? 4'h0 : _GEN_5236; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5238 = 8'h33 == _T_308[7:0] ? 4'h0 : _GEN_5237; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5239 = 8'h34 == _T_308[7:0] ? 4'h0 : _GEN_5238; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5240 = 8'h35 == _T_308[7:0] ? 4'h0 : _GEN_5239; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5241 = 8'h36 == _T_308[7:0] ? 4'h0 : _GEN_5240; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5242 = 8'h37 == _T_308[7:0] ? 4'h0 : _GEN_5241; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5243 = 8'h38 == _T_308[7:0] ? 4'hf : _GEN_5242; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5244 = 8'h39 == _T_308[7:0] ? 4'hf : _GEN_5243; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5245 = 8'h3a == _T_308[7:0] ? 4'hf : _GEN_5244; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5246 = 8'h3b == _T_308[7:0] ? 4'hf : _GEN_5245; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5247 = 8'h3c == _T_308[7:0] ? 4'hf : _GEN_5246; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5248 = 8'h3d == _T_308[7:0] ? 4'hf : _GEN_5247; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5249 = 8'h3e == _T_308[7:0] ? 4'hf : _GEN_5248; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5250 = 8'h3f == _T_308[7:0] ? 4'hf : _GEN_5249; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5251 = 8'h40 == _T_308[7:0] ? 4'h0 : _GEN_5250; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5252 = 8'h41 == _T_308[7:0] ? 4'h0 : _GEN_5251; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5253 = 8'h42 == _T_308[7:0] ? 4'h0 : _GEN_5252; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5254 = 8'h43 == _T_308[7:0] ? 4'h0 : _GEN_5253; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5255 = 8'h44 == _T_308[7:0] ? 4'h0 : _GEN_5254; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5256 = 8'h45 == _T_308[7:0] ? 4'h0 : _GEN_5255; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5257 = 8'h46 == _T_308[7:0] ? 4'h0 : _GEN_5256; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5258 = 8'h47 == _T_308[7:0] ? 4'h0 : _GEN_5257; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5259 = 8'h48 == _T_308[7:0] ? 4'hf : _GEN_5258; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5260 = 8'h49 == _T_308[7:0] ? 4'hf : _GEN_5259; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5261 = 8'h4a == _T_308[7:0] ? 4'hf : _GEN_5260; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5262 = 8'h4b == _T_308[7:0] ? 4'hf : _GEN_5261; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5263 = 8'h4c == _T_308[7:0] ? 4'hf : _GEN_5262; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5264 = 8'h4d == _T_308[7:0] ? 4'hf : _GEN_5263; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5265 = 8'h4e == _T_308[7:0] ? 4'hf : _GEN_5264; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5266 = 8'h4f == _T_308[7:0] ? 4'hf : _GEN_5265; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5267 = 8'h50 == _T_308[7:0] ? 4'h0 : _GEN_5266; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5268 = 8'h51 == _T_308[7:0] ? 4'h0 : _GEN_5267; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5269 = 8'h52 == _T_308[7:0] ? 4'h0 : _GEN_5268; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5270 = 8'h53 == _T_308[7:0] ? 4'h0 : _GEN_5269; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5271 = 8'h54 == _T_308[7:0] ? 4'h0 : _GEN_5270; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5272 = 8'h55 == _T_308[7:0] ? 4'h0 : _GEN_5271; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5273 = 8'h56 == _T_308[7:0] ? 4'h0 : _GEN_5272; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5274 = 8'h57 == _T_308[7:0] ? 4'h0 : _GEN_5273; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5275 = 8'h58 == _T_308[7:0] ? 4'hf : _GEN_5274; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5276 = 8'h59 == _T_308[7:0] ? 4'hf : _GEN_5275; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5277 = 8'h5a == _T_308[7:0] ? 4'hf : _GEN_5276; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5278 = 8'h5b == _T_308[7:0] ? 4'hf : _GEN_5277; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5279 = 8'h5c == _T_308[7:0] ? 4'hf : _GEN_5278; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5280 = 8'h5d == _T_308[7:0] ? 4'hf : _GEN_5279; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5281 = 8'h5e == _T_308[7:0] ? 4'hf : _GEN_5280; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5282 = 8'h5f == _T_308[7:0] ? 4'hf : _GEN_5281; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5283 = 8'h60 == _T_308[7:0] ? 4'h0 : _GEN_5282; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5284 = 8'h61 == _T_308[7:0] ? 4'h0 : _GEN_5283; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5285 = 8'h62 == _T_308[7:0] ? 4'h0 : _GEN_5284; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5286 = 8'h63 == _T_308[7:0] ? 4'h0 : _GEN_5285; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5287 = 8'h64 == _T_308[7:0] ? 4'h0 : _GEN_5286; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5288 = 8'h65 == _T_308[7:0] ? 4'h0 : _GEN_5287; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5289 = 8'h66 == _T_308[7:0] ? 4'h0 : _GEN_5288; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5290 = 8'h67 == _T_308[7:0] ? 4'h0 : _GEN_5289; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5291 = 8'h68 == _T_308[7:0] ? 4'hf : _GEN_5290; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5292 = 8'h69 == _T_308[7:0] ? 4'hf : _GEN_5291; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5293 = 8'h6a == _T_308[7:0] ? 4'hf : _GEN_5292; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5294 = 8'h6b == _T_308[7:0] ? 4'hf : _GEN_5293; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5295 = 8'h6c == _T_308[7:0] ? 4'hf : _GEN_5294; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5296 = 8'h6d == _T_308[7:0] ? 4'hf : _GEN_5295; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5297 = 8'h6e == _T_308[7:0] ? 4'hf : _GEN_5296; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5298 = 8'h6f == _T_308[7:0] ? 4'hf : _GEN_5297; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5299 = 8'h70 == _T_308[7:0] ? 4'h0 : _GEN_5298; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5300 = 8'h71 == _T_308[7:0] ? 4'h0 : _GEN_5299; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5301 = 8'h72 == _T_308[7:0] ? 4'h0 : _GEN_5300; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5302 = 8'h73 == _T_308[7:0] ? 4'h0 : _GEN_5301; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5303 = 8'h74 == _T_308[7:0] ? 4'h0 : _GEN_5302; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5304 = 8'h75 == _T_308[7:0] ? 4'h0 : _GEN_5303; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5305 = 8'h76 == _T_308[7:0] ? 4'h0 : _GEN_5304; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5306 = 8'h77 == _T_308[7:0] ? 4'h0 : _GEN_5305; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5307 = 8'h78 == _T_308[7:0] ? 4'hf : _GEN_5306; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5308 = 8'h79 == _T_308[7:0] ? 4'hf : _GEN_5307; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5309 = 8'h7a == _T_308[7:0] ? 4'hf : _GEN_5308; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5310 = 8'h7b == _T_308[7:0] ? 4'hf : _GEN_5309; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5311 = 8'h7c == _T_308[7:0] ? 4'hf : _GEN_5310; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5312 = 8'h7d == _T_308[7:0] ? 4'hf : _GEN_5311; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5313 = 8'h7e == _T_308[7:0] ? 4'hf : _GEN_5312; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5314 = 8'h7f == _T_308[7:0] ? 4'hf : _GEN_5313; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5315 = 8'h80 == _T_308[7:0] ? 4'h0 : _GEN_5314; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5316 = 8'h81 == _T_308[7:0] ? 4'h0 : _GEN_5315; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5317 = 8'h82 == _T_308[7:0] ? 4'h0 : _GEN_5316; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5318 = 8'h83 == _T_308[7:0] ? 4'h0 : _GEN_5317; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5319 = 8'h84 == _T_308[7:0] ? 4'h0 : _GEN_5318; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5320 = 8'h85 == _T_308[7:0] ? 4'h0 : _GEN_5319; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5321 = 8'h86 == _T_308[7:0] ? 4'h0 : _GEN_5320; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5322 = 8'h87 == _T_308[7:0] ? 4'h0 : _GEN_5321; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5323 = 8'h88 == _T_308[7:0] ? 4'hf : _GEN_5322; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5324 = 8'h89 == _T_308[7:0] ? 4'hf : _GEN_5323; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5325 = 8'h8a == _T_308[7:0] ? 4'hf : _GEN_5324; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5326 = 8'h8b == _T_308[7:0] ? 4'hf : _GEN_5325; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5327 = 8'h8c == _T_308[7:0] ? 4'hf : _GEN_5326; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5328 = 8'h8d == _T_308[7:0] ? 4'hf : _GEN_5327; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5329 = 8'h8e == _T_308[7:0] ? 4'hf : _GEN_5328; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5330 = 8'h8f == _T_308[7:0] ? 4'hf : _GEN_5329; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5331 = 8'h90 == _T_308[7:0] ? 4'h0 : _GEN_5330; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5332 = 8'h91 == _T_308[7:0] ? 4'h0 : _GEN_5331; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5333 = 8'h92 == _T_308[7:0] ? 4'h0 : _GEN_5332; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5334 = 8'h93 == _T_308[7:0] ? 4'h0 : _GEN_5333; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5335 = 8'h94 == _T_308[7:0] ? 4'h0 : _GEN_5334; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5336 = 8'h95 == _T_308[7:0] ? 4'h0 : _GEN_5335; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5337 = 8'h96 == _T_308[7:0] ? 4'h0 : _GEN_5336; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5338 = 8'h97 == _T_308[7:0] ? 4'h0 : _GEN_5337; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5339 = 8'h98 == _T_308[7:0] ? 4'hf : _GEN_5338; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5340 = 8'h99 == _T_308[7:0] ? 4'hf : _GEN_5339; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5341 = 8'h9a == _T_308[7:0] ? 4'hf : _GEN_5340; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5342 = 8'h9b == _T_308[7:0] ? 4'hf : _GEN_5341; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5343 = 8'h9c == _T_308[7:0] ? 4'hf : _GEN_5342; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5344 = 8'h9d == _T_308[7:0] ? 4'hf : _GEN_5343; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5345 = 8'h9e == _T_308[7:0] ? 4'hf : _GEN_5344; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5346 = 8'h9f == _T_308[7:0] ? 4'hf : _GEN_5345; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5347 = 8'ha0 == _T_308[7:0] ? 4'h0 : _GEN_5346; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5348 = 8'ha1 == _T_308[7:0] ? 4'h0 : _GEN_5347; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5349 = 8'ha2 == _T_308[7:0] ? 4'h0 : _GEN_5348; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5350 = 8'ha3 == _T_308[7:0] ? 4'h0 : _GEN_5349; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5351 = 8'ha4 == _T_308[7:0] ? 4'h0 : _GEN_5350; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5352 = 8'ha5 == _T_308[7:0] ? 4'h0 : _GEN_5351; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5353 = 8'ha6 == _T_308[7:0] ? 4'h0 : _GEN_5352; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5354 = 8'ha7 == _T_308[7:0] ? 4'h0 : _GEN_5353; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5355 = 8'ha8 == _T_308[7:0] ? 4'hf : _GEN_5354; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5356 = 8'ha9 == _T_308[7:0] ? 4'hf : _GEN_5355; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5357 = 8'haa == _T_308[7:0] ? 4'hf : _GEN_5356; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5358 = 8'hab == _T_308[7:0] ? 4'hf : _GEN_5357; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5359 = 8'hac == _T_308[7:0] ? 4'hf : _GEN_5358; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5360 = 8'had == _T_308[7:0] ? 4'hf : _GEN_5359; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5361 = 8'hae == _T_308[7:0] ? 4'hf : _GEN_5360; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5362 = 8'haf == _T_308[7:0] ? 4'hf : _GEN_5361; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5363 = 8'hb0 == _T_308[7:0] ? 4'h0 : _GEN_5362; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5364 = 8'hb1 == _T_308[7:0] ? 4'h0 : _GEN_5363; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5365 = 8'hb2 == _T_308[7:0] ? 4'h0 : _GEN_5364; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5366 = 8'hb3 == _T_308[7:0] ? 4'h0 : _GEN_5365; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5367 = 8'hb4 == _T_308[7:0] ? 4'h0 : _GEN_5366; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5368 = 8'hb5 == _T_308[7:0] ? 4'h0 : _GEN_5367; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5369 = 8'hb6 == _T_308[7:0] ? 4'h0 : _GEN_5368; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5370 = 8'hb7 == _T_308[7:0] ? 4'h0 : _GEN_5369; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5371 = 8'hb8 == _T_308[7:0] ? 4'hf : _GEN_5370; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5372 = 8'hb9 == _T_308[7:0] ? 4'hf : _GEN_5371; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5373 = 8'hba == _T_308[7:0] ? 4'hf : _GEN_5372; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5374 = 8'hbb == _T_308[7:0] ? 4'hf : _GEN_5373; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5375 = 8'hbc == _T_308[7:0] ? 4'hf : _GEN_5374; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5376 = 8'hbd == _T_308[7:0] ? 4'hf : _GEN_5375; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5377 = 8'hbe == _T_308[7:0] ? 4'hf : _GEN_5376; // @[Filter.scala 160:142]
  wire [3:0] _GEN_5378 = 8'hbf == _T_308[7:0] ? 4'hf : _GEN_5377; // @[Filter.scala 160:142]
  wire [7:0] _T_322 = _GEN_5378 * 4'ha; // @[Filter.scala 160:142]
  wire [10:0] _GEN_9919 = {{3'd0}, _T_322}; // @[Filter.scala 160:109]
  wire [10:0] _T_324 = _T_317 + _GEN_9919; // @[Filter.scala 160:109]
  wire [10:0] _T_325 = _T_324 / 11'h64; // @[Filter.scala 160:150]
  wire  _T_327 = _T_298 >= 5'h10; // @[Filter.scala 163:31]
  wire  _T_331 = _T_305 >= 32'hc; // @[Filter.scala 163:63]
  wire  _T_332 = _T_327 | _T_331; // @[Filter.scala 163:58]
  wire [10:0] _GEN_5571 = io_SPI_distort ? _T_325 : {{7'd0}, _GEN_4994}; // @[Filter.scala 165:35]
  wire [10:0] _GEN_5572 = _T_332 ? 11'h0 : _GEN_5571; // @[Filter.scala 163:80]
  wire [10:0] _GEN_5765 = io_SPI_distort ? _T_325 : {{7'd0}, _GEN_5186}; // @[Filter.scala 165:35]
  wire [10:0] _GEN_5766 = _T_332 ? 11'h0 : _GEN_5765; // @[Filter.scala 163:80]
  wire [10:0] _GEN_5959 = io_SPI_distort ? _T_325 : {{7'd0}, _GEN_5378}; // @[Filter.scala 165:35]
  wire [10:0] _GEN_5960 = _T_332 ? 11'h0 : _GEN_5959; // @[Filter.scala 163:80]
  wire [31:0] _T_360 = pixelIndex + 32'h5; // @[Filter.scala 158:31]
  wire [31:0] _GEN_5 = _T_360 % 32'h10; // @[Filter.scala 158:38]
  wire [4:0] _T_361 = _GEN_5[4:0]; // @[Filter.scala 158:38]
  wire [4:0] _T_363 = _T_361 + _GEN_9863; // @[Filter.scala 158:53]
  wire [4:0] _T_365 = _T_363 - 5'h1; // @[Filter.scala 158:69]
  wire [31:0] _T_368 = _T_360 / 32'h10; // @[Filter.scala 159:38]
  wire [31:0] _T_370 = _T_368 + _GEN_9864; // @[Filter.scala 159:53]
  wire [31:0] _T_372 = _T_370 - 32'h1; // @[Filter.scala 159:69]
  wire [36:0] _T_373 = _T_372 * 32'h10; // @[Filter.scala 160:42]
  wire [36:0] _GEN_9925 = {{32'd0}, _T_365}; // @[Filter.scala 160:57]
  wire [36:0] _T_375 = _T_373 + _GEN_9925; // @[Filter.scala 160:57]
  wire [3:0] _GEN_5969 = 8'h8 == _T_375[7:0] ? 4'h0 : 4'hf; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5970 = 8'h9 == _T_375[7:0] ? 4'h0 : _GEN_5969; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5971 = 8'ha == _T_375[7:0] ? 4'h0 : _GEN_5970; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5972 = 8'hb == _T_375[7:0] ? 4'h0 : _GEN_5971; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5973 = 8'hc == _T_375[7:0] ? 4'h0 : _GEN_5972; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5974 = 8'hd == _T_375[7:0] ? 4'h0 : _GEN_5973; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5975 = 8'he == _T_375[7:0] ? 4'h0 : _GEN_5974; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5976 = 8'hf == _T_375[7:0] ? 4'h0 : _GEN_5975; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5977 = 8'h10 == _T_375[7:0] ? 4'hf : _GEN_5976; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5978 = 8'h11 == _T_375[7:0] ? 4'hf : _GEN_5977; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5979 = 8'h12 == _T_375[7:0] ? 4'hf : _GEN_5978; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5980 = 8'h13 == _T_375[7:0] ? 4'hf : _GEN_5979; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5981 = 8'h14 == _T_375[7:0] ? 4'hf : _GEN_5980; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5982 = 8'h15 == _T_375[7:0] ? 4'hf : _GEN_5981; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5983 = 8'h16 == _T_375[7:0] ? 4'hf : _GEN_5982; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5984 = 8'h17 == _T_375[7:0] ? 4'hf : _GEN_5983; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5985 = 8'h18 == _T_375[7:0] ? 4'h0 : _GEN_5984; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5986 = 8'h19 == _T_375[7:0] ? 4'h0 : _GEN_5985; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5987 = 8'h1a == _T_375[7:0] ? 4'h0 : _GEN_5986; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5988 = 8'h1b == _T_375[7:0] ? 4'h0 : _GEN_5987; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5989 = 8'h1c == _T_375[7:0] ? 4'h0 : _GEN_5988; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5990 = 8'h1d == _T_375[7:0] ? 4'h0 : _GEN_5989; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5991 = 8'h1e == _T_375[7:0] ? 4'h0 : _GEN_5990; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5992 = 8'h1f == _T_375[7:0] ? 4'h0 : _GEN_5991; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5993 = 8'h20 == _T_375[7:0] ? 4'hf : _GEN_5992; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5994 = 8'h21 == _T_375[7:0] ? 4'hf : _GEN_5993; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5995 = 8'h22 == _T_375[7:0] ? 4'hf : _GEN_5994; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5996 = 8'h23 == _T_375[7:0] ? 4'hf : _GEN_5995; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5997 = 8'h24 == _T_375[7:0] ? 4'hf : _GEN_5996; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5998 = 8'h25 == _T_375[7:0] ? 4'hf : _GEN_5997; // @[Filter.scala 160:62]
  wire [3:0] _GEN_5999 = 8'h26 == _T_375[7:0] ? 4'hf : _GEN_5998; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6000 = 8'h27 == _T_375[7:0] ? 4'hf : _GEN_5999; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6001 = 8'h28 == _T_375[7:0] ? 4'h0 : _GEN_6000; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6002 = 8'h29 == _T_375[7:0] ? 4'h0 : _GEN_6001; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6003 = 8'h2a == _T_375[7:0] ? 4'h0 : _GEN_6002; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6004 = 8'h2b == _T_375[7:0] ? 4'h0 : _GEN_6003; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6005 = 8'h2c == _T_375[7:0] ? 4'h0 : _GEN_6004; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6006 = 8'h2d == _T_375[7:0] ? 4'h0 : _GEN_6005; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6007 = 8'h2e == _T_375[7:0] ? 4'h0 : _GEN_6006; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6008 = 8'h2f == _T_375[7:0] ? 4'h0 : _GEN_6007; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6009 = 8'h30 == _T_375[7:0] ? 4'hf : _GEN_6008; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6010 = 8'h31 == _T_375[7:0] ? 4'hf : _GEN_6009; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6011 = 8'h32 == _T_375[7:0] ? 4'hf : _GEN_6010; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6012 = 8'h33 == _T_375[7:0] ? 4'hf : _GEN_6011; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6013 = 8'h34 == _T_375[7:0] ? 4'hf : _GEN_6012; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6014 = 8'h35 == _T_375[7:0] ? 4'hf : _GEN_6013; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6015 = 8'h36 == _T_375[7:0] ? 4'hf : _GEN_6014; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6016 = 8'h37 == _T_375[7:0] ? 4'hf : _GEN_6015; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6017 = 8'h38 == _T_375[7:0] ? 4'h0 : _GEN_6016; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6018 = 8'h39 == _T_375[7:0] ? 4'h0 : _GEN_6017; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6019 = 8'h3a == _T_375[7:0] ? 4'h0 : _GEN_6018; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6020 = 8'h3b == _T_375[7:0] ? 4'h0 : _GEN_6019; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6021 = 8'h3c == _T_375[7:0] ? 4'h0 : _GEN_6020; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6022 = 8'h3d == _T_375[7:0] ? 4'h0 : _GEN_6021; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6023 = 8'h3e == _T_375[7:0] ? 4'h0 : _GEN_6022; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6024 = 8'h3f == _T_375[7:0] ? 4'h0 : _GEN_6023; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6025 = 8'h40 == _T_375[7:0] ? 4'hf : _GEN_6024; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6026 = 8'h41 == _T_375[7:0] ? 4'hf : _GEN_6025; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6027 = 8'h42 == _T_375[7:0] ? 4'hf : _GEN_6026; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6028 = 8'h43 == _T_375[7:0] ? 4'hf : _GEN_6027; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6029 = 8'h44 == _T_375[7:0] ? 4'hf : _GEN_6028; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6030 = 8'h45 == _T_375[7:0] ? 4'hf : _GEN_6029; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6031 = 8'h46 == _T_375[7:0] ? 4'hf : _GEN_6030; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6032 = 8'h47 == _T_375[7:0] ? 4'hf : _GEN_6031; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6033 = 8'h48 == _T_375[7:0] ? 4'h0 : _GEN_6032; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6034 = 8'h49 == _T_375[7:0] ? 4'h0 : _GEN_6033; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6035 = 8'h4a == _T_375[7:0] ? 4'h0 : _GEN_6034; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6036 = 8'h4b == _T_375[7:0] ? 4'h0 : _GEN_6035; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6037 = 8'h4c == _T_375[7:0] ? 4'h0 : _GEN_6036; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6038 = 8'h4d == _T_375[7:0] ? 4'h0 : _GEN_6037; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6039 = 8'h4e == _T_375[7:0] ? 4'h0 : _GEN_6038; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6040 = 8'h4f == _T_375[7:0] ? 4'h0 : _GEN_6039; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6041 = 8'h50 == _T_375[7:0] ? 4'hf : _GEN_6040; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6042 = 8'h51 == _T_375[7:0] ? 4'hf : _GEN_6041; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6043 = 8'h52 == _T_375[7:0] ? 4'hf : _GEN_6042; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6044 = 8'h53 == _T_375[7:0] ? 4'hf : _GEN_6043; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6045 = 8'h54 == _T_375[7:0] ? 4'hf : _GEN_6044; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6046 = 8'h55 == _T_375[7:0] ? 4'hf : _GEN_6045; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6047 = 8'h56 == _T_375[7:0] ? 4'hf : _GEN_6046; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6048 = 8'h57 == _T_375[7:0] ? 4'hf : _GEN_6047; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6049 = 8'h58 == _T_375[7:0] ? 4'h0 : _GEN_6048; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6050 = 8'h59 == _T_375[7:0] ? 4'h0 : _GEN_6049; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6051 = 8'h5a == _T_375[7:0] ? 4'h0 : _GEN_6050; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6052 = 8'h5b == _T_375[7:0] ? 4'h0 : _GEN_6051; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6053 = 8'h5c == _T_375[7:0] ? 4'h0 : _GEN_6052; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6054 = 8'h5d == _T_375[7:0] ? 4'h0 : _GEN_6053; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6055 = 8'h5e == _T_375[7:0] ? 4'h0 : _GEN_6054; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6056 = 8'h5f == _T_375[7:0] ? 4'h0 : _GEN_6055; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6057 = 8'h60 == _T_375[7:0] ? 4'h0 : _GEN_6056; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6058 = 8'h61 == _T_375[7:0] ? 4'h0 : _GEN_6057; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6059 = 8'h62 == _T_375[7:0] ? 4'h0 : _GEN_6058; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6060 = 8'h63 == _T_375[7:0] ? 4'h0 : _GEN_6059; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6061 = 8'h64 == _T_375[7:0] ? 4'h0 : _GEN_6060; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6062 = 8'h65 == _T_375[7:0] ? 4'h0 : _GEN_6061; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6063 = 8'h66 == _T_375[7:0] ? 4'h0 : _GEN_6062; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6064 = 8'h67 == _T_375[7:0] ? 4'h0 : _GEN_6063; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6065 = 8'h68 == _T_375[7:0] ? 4'hf : _GEN_6064; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6066 = 8'h69 == _T_375[7:0] ? 4'hf : _GEN_6065; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6067 = 8'h6a == _T_375[7:0] ? 4'hf : _GEN_6066; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6068 = 8'h6b == _T_375[7:0] ? 4'hf : _GEN_6067; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6069 = 8'h6c == _T_375[7:0] ? 4'hf : _GEN_6068; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6070 = 8'h6d == _T_375[7:0] ? 4'hf : _GEN_6069; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6071 = 8'h6e == _T_375[7:0] ? 4'hf : _GEN_6070; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6072 = 8'h6f == _T_375[7:0] ? 4'hf : _GEN_6071; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6073 = 8'h70 == _T_375[7:0] ? 4'h0 : _GEN_6072; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6074 = 8'h71 == _T_375[7:0] ? 4'h0 : _GEN_6073; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6075 = 8'h72 == _T_375[7:0] ? 4'h0 : _GEN_6074; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6076 = 8'h73 == _T_375[7:0] ? 4'h0 : _GEN_6075; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6077 = 8'h74 == _T_375[7:0] ? 4'h0 : _GEN_6076; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6078 = 8'h75 == _T_375[7:0] ? 4'h0 : _GEN_6077; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6079 = 8'h76 == _T_375[7:0] ? 4'h0 : _GEN_6078; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6080 = 8'h77 == _T_375[7:0] ? 4'h0 : _GEN_6079; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6081 = 8'h78 == _T_375[7:0] ? 4'hf : _GEN_6080; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6082 = 8'h79 == _T_375[7:0] ? 4'hf : _GEN_6081; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6083 = 8'h7a == _T_375[7:0] ? 4'hf : _GEN_6082; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6084 = 8'h7b == _T_375[7:0] ? 4'hf : _GEN_6083; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6085 = 8'h7c == _T_375[7:0] ? 4'hf : _GEN_6084; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6086 = 8'h7d == _T_375[7:0] ? 4'hf : _GEN_6085; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6087 = 8'h7e == _T_375[7:0] ? 4'hf : _GEN_6086; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6088 = 8'h7f == _T_375[7:0] ? 4'hf : _GEN_6087; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6089 = 8'h80 == _T_375[7:0] ? 4'h0 : _GEN_6088; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6090 = 8'h81 == _T_375[7:0] ? 4'h0 : _GEN_6089; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6091 = 8'h82 == _T_375[7:0] ? 4'h0 : _GEN_6090; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6092 = 8'h83 == _T_375[7:0] ? 4'h0 : _GEN_6091; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6093 = 8'h84 == _T_375[7:0] ? 4'h0 : _GEN_6092; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6094 = 8'h85 == _T_375[7:0] ? 4'h0 : _GEN_6093; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6095 = 8'h86 == _T_375[7:0] ? 4'h0 : _GEN_6094; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6096 = 8'h87 == _T_375[7:0] ? 4'h0 : _GEN_6095; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6097 = 8'h88 == _T_375[7:0] ? 4'hf : _GEN_6096; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6098 = 8'h89 == _T_375[7:0] ? 4'hf : _GEN_6097; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6099 = 8'h8a == _T_375[7:0] ? 4'hf : _GEN_6098; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6100 = 8'h8b == _T_375[7:0] ? 4'hf : _GEN_6099; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6101 = 8'h8c == _T_375[7:0] ? 4'hf : _GEN_6100; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6102 = 8'h8d == _T_375[7:0] ? 4'hf : _GEN_6101; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6103 = 8'h8e == _T_375[7:0] ? 4'hf : _GEN_6102; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6104 = 8'h8f == _T_375[7:0] ? 4'hf : _GEN_6103; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6105 = 8'h90 == _T_375[7:0] ? 4'h0 : _GEN_6104; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6106 = 8'h91 == _T_375[7:0] ? 4'h0 : _GEN_6105; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6107 = 8'h92 == _T_375[7:0] ? 4'h0 : _GEN_6106; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6108 = 8'h93 == _T_375[7:0] ? 4'h0 : _GEN_6107; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6109 = 8'h94 == _T_375[7:0] ? 4'h0 : _GEN_6108; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6110 = 8'h95 == _T_375[7:0] ? 4'h0 : _GEN_6109; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6111 = 8'h96 == _T_375[7:0] ? 4'h0 : _GEN_6110; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6112 = 8'h97 == _T_375[7:0] ? 4'h0 : _GEN_6111; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6113 = 8'h98 == _T_375[7:0] ? 4'hf : _GEN_6112; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6114 = 8'h99 == _T_375[7:0] ? 4'hf : _GEN_6113; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6115 = 8'h9a == _T_375[7:0] ? 4'hf : _GEN_6114; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6116 = 8'h9b == _T_375[7:0] ? 4'hf : _GEN_6115; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6117 = 8'h9c == _T_375[7:0] ? 4'hf : _GEN_6116; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6118 = 8'h9d == _T_375[7:0] ? 4'hf : _GEN_6117; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6119 = 8'h9e == _T_375[7:0] ? 4'hf : _GEN_6118; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6120 = 8'h9f == _T_375[7:0] ? 4'hf : _GEN_6119; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6121 = 8'ha0 == _T_375[7:0] ? 4'h0 : _GEN_6120; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6122 = 8'ha1 == _T_375[7:0] ? 4'h0 : _GEN_6121; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6123 = 8'ha2 == _T_375[7:0] ? 4'h0 : _GEN_6122; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6124 = 8'ha3 == _T_375[7:0] ? 4'h0 : _GEN_6123; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6125 = 8'ha4 == _T_375[7:0] ? 4'h0 : _GEN_6124; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6126 = 8'ha5 == _T_375[7:0] ? 4'h0 : _GEN_6125; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6127 = 8'ha6 == _T_375[7:0] ? 4'h0 : _GEN_6126; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6128 = 8'ha7 == _T_375[7:0] ? 4'h0 : _GEN_6127; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6129 = 8'ha8 == _T_375[7:0] ? 4'hf : _GEN_6128; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6130 = 8'ha9 == _T_375[7:0] ? 4'hf : _GEN_6129; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6131 = 8'haa == _T_375[7:0] ? 4'hf : _GEN_6130; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6132 = 8'hab == _T_375[7:0] ? 4'hf : _GEN_6131; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6133 = 8'hac == _T_375[7:0] ? 4'hf : _GEN_6132; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6134 = 8'had == _T_375[7:0] ? 4'hf : _GEN_6133; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6135 = 8'hae == _T_375[7:0] ? 4'hf : _GEN_6134; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6136 = 8'haf == _T_375[7:0] ? 4'hf : _GEN_6135; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6137 = 8'hb0 == _T_375[7:0] ? 4'h0 : _GEN_6136; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6138 = 8'hb1 == _T_375[7:0] ? 4'h0 : _GEN_6137; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6139 = 8'hb2 == _T_375[7:0] ? 4'h0 : _GEN_6138; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6140 = 8'hb3 == _T_375[7:0] ? 4'h0 : _GEN_6139; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6141 = 8'hb4 == _T_375[7:0] ? 4'h0 : _GEN_6140; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6142 = 8'hb5 == _T_375[7:0] ? 4'h0 : _GEN_6141; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6143 = 8'hb6 == _T_375[7:0] ? 4'h0 : _GEN_6142; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6144 = 8'hb7 == _T_375[7:0] ? 4'h0 : _GEN_6143; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6145 = 8'hb8 == _T_375[7:0] ? 4'hf : _GEN_6144; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6146 = 8'hb9 == _T_375[7:0] ? 4'hf : _GEN_6145; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6147 = 8'hba == _T_375[7:0] ? 4'hf : _GEN_6146; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6148 = 8'hbb == _T_375[7:0] ? 4'hf : _GEN_6147; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6149 = 8'hbc == _T_375[7:0] ? 4'hf : _GEN_6148; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6150 = 8'hbd == _T_375[7:0] ? 4'hf : _GEN_6149; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6151 = 8'hbe == _T_375[7:0] ? 4'hf : _GEN_6150; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6152 = 8'hbf == _T_375[7:0] ? 4'hf : _GEN_6151; // @[Filter.scala 160:62]
  wire [4:0] _GEN_9926 = {{1'd0}, _GEN_6152}; // @[Filter.scala 160:62]
  wire [8:0] _T_377 = _GEN_9926 * 5'h14; // @[Filter.scala 160:62]
  wire [3:0] _GEN_6249 = 8'h60 == _T_375[7:0] ? 4'hf : 4'h0; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6250 = 8'h61 == _T_375[7:0] ? 4'hf : _GEN_6249; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6251 = 8'h62 == _T_375[7:0] ? 4'hf : _GEN_6250; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6252 = 8'h63 == _T_375[7:0] ? 4'hf : _GEN_6251; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6253 = 8'h64 == _T_375[7:0] ? 4'hf : _GEN_6252; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6254 = 8'h65 == _T_375[7:0] ? 4'hf : _GEN_6253; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6255 = 8'h66 == _T_375[7:0] ? 4'hf : _GEN_6254; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6256 = 8'h67 == _T_375[7:0] ? 4'hf : _GEN_6255; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6257 = 8'h68 == _T_375[7:0] ? 4'hf : _GEN_6256; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6258 = 8'h69 == _T_375[7:0] ? 4'hf : _GEN_6257; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6259 = 8'h6a == _T_375[7:0] ? 4'hf : _GEN_6258; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6260 = 8'h6b == _T_375[7:0] ? 4'hf : _GEN_6259; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6261 = 8'h6c == _T_375[7:0] ? 4'hf : _GEN_6260; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6262 = 8'h6d == _T_375[7:0] ? 4'hf : _GEN_6261; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6263 = 8'h6e == _T_375[7:0] ? 4'hf : _GEN_6262; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6264 = 8'h6f == _T_375[7:0] ? 4'hf : _GEN_6263; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6265 = 8'h70 == _T_375[7:0] ? 4'hf : _GEN_6264; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6266 = 8'h71 == _T_375[7:0] ? 4'hf : _GEN_6265; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6267 = 8'h72 == _T_375[7:0] ? 4'hf : _GEN_6266; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6268 = 8'h73 == _T_375[7:0] ? 4'hf : _GEN_6267; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6269 = 8'h74 == _T_375[7:0] ? 4'hf : _GEN_6268; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6270 = 8'h75 == _T_375[7:0] ? 4'hf : _GEN_6269; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6271 = 8'h76 == _T_375[7:0] ? 4'hf : _GEN_6270; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6272 = 8'h77 == _T_375[7:0] ? 4'hf : _GEN_6271; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6273 = 8'h78 == _T_375[7:0] ? 4'hf : _GEN_6272; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6274 = 8'h79 == _T_375[7:0] ? 4'hf : _GEN_6273; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6275 = 8'h7a == _T_375[7:0] ? 4'hf : _GEN_6274; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6276 = 8'h7b == _T_375[7:0] ? 4'hf : _GEN_6275; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6277 = 8'h7c == _T_375[7:0] ? 4'hf : _GEN_6276; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6278 = 8'h7d == _T_375[7:0] ? 4'hf : _GEN_6277; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6279 = 8'h7e == _T_375[7:0] ? 4'hf : _GEN_6278; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6280 = 8'h7f == _T_375[7:0] ? 4'hf : _GEN_6279; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6281 = 8'h80 == _T_375[7:0] ? 4'hf : _GEN_6280; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6282 = 8'h81 == _T_375[7:0] ? 4'hf : _GEN_6281; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6283 = 8'h82 == _T_375[7:0] ? 4'hf : _GEN_6282; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6284 = 8'h83 == _T_375[7:0] ? 4'hf : _GEN_6283; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6285 = 8'h84 == _T_375[7:0] ? 4'hf : _GEN_6284; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6286 = 8'h85 == _T_375[7:0] ? 4'hf : _GEN_6285; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6287 = 8'h86 == _T_375[7:0] ? 4'hf : _GEN_6286; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6288 = 8'h87 == _T_375[7:0] ? 4'hf : _GEN_6287; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6289 = 8'h88 == _T_375[7:0] ? 4'hf : _GEN_6288; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6290 = 8'h89 == _T_375[7:0] ? 4'hf : _GEN_6289; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6291 = 8'h8a == _T_375[7:0] ? 4'hf : _GEN_6290; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6292 = 8'h8b == _T_375[7:0] ? 4'hf : _GEN_6291; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6293 = 8'h8c == _T_375[7:0] ? 4'hf : _GEN_6292; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6294 = 8'h8d == _T_375[7:0] ? 4'hf : _GEN_6293; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6295 = 8'h8e == _T_375[7:0] ? 4'hf : _GEN_6294; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6296 = 8'h8f == _T_375[7:0] ? 4'hf : _GEN_6295; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6297 = 8'h90 == _T_375[7:0] ? 4'hf : _GEN_6296; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6298 = 8'h91 == _T_375[7:0] ? 4'hf : _GEN_6297; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6299 = 8'h92 == _T_375[7:0] ? 4'hf : _GEN_6298; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6300 = 8'h93 == _T_375[7:0] ? 4'hf : _GEN_6299; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6301 = 8'h94 == _T_375[7:0] ? 4'hf : _GEN_6300; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6302 = 8'h95 == _T_375[7:0] ? 4'hf : _GEN_6301; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6303 = 8'h96 == _T_375[7:0] ? 4'hf : _GEN_6302; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6304 = 8'h97 == _T_375[7:0] ? 4'hf : _GEN_6303; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6305 = 8'h98 == _T_375[7:0] ? 4'hf : _GEN_6304; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6306 = 8'h99 == _T_375[7:0] ? 4'hf : _GEN_6305; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6307 = 8'h9a == _T_375[7:0] ? 4'hf : _GEN_6306; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6308 = 8'h9b == _T_375[7:0] ? 4'hf : _GEN_6307; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6309 = 8'h9c == _T_375[7:0] ? 4'hf : _GEN_6308; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6310 = 8'h9d == _T_375[7:0] ? 4'hf : _GEN_6309; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6311 = 8'h9e == _T_375[7:0] ? 4'hf : _GEN_6310; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6312 = 8'h9f == _T_375[7:0] ? 4'hf : _GEN_6311; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6313 = 8'ha0 == _T_375[7:0] ? 4'hf : _GEN_6312; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6314 = 8'ha1 == _T_375[7:0] ? 4'hf : _GEN_6313; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6315 = 8'ha2 == _T_375[7:0] ? 4'hf : _GEN_6314; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6316 = 8'ha3 == _T_375[7:0] ? 4'hf : _GEN_6315; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6317 = 8'ha4 == _T_375[7:0] ? 4'hf : _GEN_6316; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6318 = 8'ha5 == _T_375[7:0] ? 4'hf : _GEN_6317; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6319 = 8'ha6 == _T_375[7:0] ? 4'hf : _GEN_6318; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6320 = 8'ha7 == _T_375[7:0] ? 4'hf : _GEN_6319; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6321 = 8'ha8 == _T_375[7:0] ? 4'hf : _GEN_6320; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6322 = 8'ha9 == _T_375[7:0] ? 4'hf : _GEN_6321; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6323 = 8'haa == _T_375[7:0] ? 4'hf : _GEN_6322; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6324 = 8'hab == _T_375[7:0] ? 4'hf : _GEN_6323; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6325 = 8'hac == _T_375[7:0] ? 4'hf : _GEN_6324; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6326 = 8'had == _T_375[7:0] ? 4'hf : _GEN_6325; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6327 = 8'hae == _T_375[7:0] ? 4'hf : _GEN_6326; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6328 = 8'haf == _T_375[7:0] ? 4'hf : _GEN_6327; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6329 = 8'hb0 == _T_375[7:0] ? 4'hf : _GEN_6328; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6330 = 8'hb1 == _T_375[7:0] ? 4'hf : _GEN_6329; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6331 = 8'hb2 == _T_375[7:0] ? 4'hf : _GEN_6330; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6332 = 8'hb3 == _T_375[7:0] ? 4'hf : _GEN_6331; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6333 = 8'hb4 == _T_375[7:0] ? 4'hf : _GEN_6332; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6334 = 8'hb5 == _T_375[7:0] ? 4'hf : _GEN_6333; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6335 = 8'hb6 == _T_375[7:0] ? 4'hf : _GEN_6334; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6336 = 8'hb7 == _T_375[7:0] ? 4'hf : _GEN_6335; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6337 = 8'hb8 == _T_375[7:0] ? 4'hf : _GEN_6336; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6338 = 8'hb9 == _T_375[7:0] ? 4'hf : _GEN_6337; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6339 = 8'hba == _T_375[7:0] ? 4'hf : _GEN_6338; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6340 = 8'hbb == _T_375[7:0] ? 4'hf : _GEN_6339; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6341 = 8'hbc == _T_375[7:0] ? 4'hf : _GEN_6340; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6342 = 8'hbd == _T_375[7:0] ? 4'hf : _GEN_6341; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6343 = 8'hbe == _T_375[7:0] ? 4'hf : _GEN_6342; // @[Filter.scala 160:102]
  wire [3:0] _GEN_6344 = 8'hbf == _T_375[7:0] ? 4'hf : _GEN_6343; // @[Filter.scala 160:102]
  wire [6:0] _GEN_9928 = {{3'd0}, _GEN_6344}; // @[Filter.scala 160:102]
  wire [10:0] _T_382 = _GEN_9928 * 7'h46; // @[Filter.scala 160:102]
  wire [10:0] _GEN_9929 = {{2'd0}, _T_377}; // @[Filter.scala 160:69]
  wire [10:0] _T_384 = _GEN_9929 + _T_382; // @[Filter.scala 160:69]
  wire [3:0] _GEN_6353 = 8'h8 == _T_375[7:0] ? 4'hf : 4'h0; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6354 = 8'h9 == _T_375[7:0] ? 4'hf : _GEN_6353; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6355 = 8'ha == _T_375[7:0] ? 4'hf : _GEN_6354; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6356 = 8'hb == _T_375[7:0] ? 4'hf : _GEN_6355; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6357 = 8'hc == _T_375[7:0] ? 4'hf : _GEN_6356; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6358 = 8'hd == _T_375[7:0] ? 4'hf : _GEN_6357; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6359 = 8'he == _T_375[7:0] ? 4'hf : _GEN_6358; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6360 = 8'hf == _T_375[7:0] ? 4'hf : _GEN_6359; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6361 = 8'h10 == _T_375[7:0] ? 4'h0 : _GEN_6360; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6362 = 8'h11 == _T_375[7:0] ? 4'h0 : _GEN_6361; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6363 = 8'h12 == _T_375[7:0] ? 4'h0 : _GEN_6362; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6364 = 8'h13 == _T_375[7:0] ? 4'h0 : _GEN_6363; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6365 = 8'h14 == _T_375[7:0] ? 4'h0 : _GEN_6364; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6366 = 8'h15 == _T_375[7:0] ? 4'h0 : _GEN_6365; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6367 = 8'h16 == _T_375[7:0] ? 4'h0 : _GEN_6366; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6368 = 8'h17 == _T_375[7:0] ? 4'h0 : _GEN_6367; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6369 = 8'h18 == _T_375[7:0] ? 4'hf : _GEN_6368; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6370 = 8'h19 == _T_375[7:0] ? 4'hf : _GEN_6369; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6371 = 8'h1a == _T_375[7:0] ? 4'hf : _GEN_6370; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6372 = 8'h1b == _T_375[7:0] ? 4'hf : _GEN_6371; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6373 = 8'h1c == _T_375[7:0] ? 4'hf : _GEN_6372; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6374 = 8'h1d == _T_375[7:0] ? 4'hf : _GEN_6373; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6375 = 8'h1e == _T_375[7:0] ? 4'hf : _GEN_6374; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6376 = 8'h1f == _T_375[7:0] ? 4'hf : _GEN_6375; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6377 = 8'h20 == _T_375[7:0] ? 4'h0 : _GEN_6376; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6378 = 8'h21 == _T_375[7:0] ? 4'h0 : _GEN_6377; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6379 = 8'h22 == _T_375[7:0] ? 4'h0 : _GEN_6378; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6380 = 8'h23 == _T_375[7:0] ? 4'h0 : _GEN_6379; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6381 = 8'h24 == _T_375[7:0] ? 4'h0 : _GEN_6380; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6382 = 8'h25 == _T_375[7:0] ? 4'h0 : _GEN_6381; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6383 = 8'h26 == _T_375[7:0] ? 4'h0 : _GEN_6382; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6384 = 8'h27 == _T_375[7:0] ? 4'h0 : _GEN_6383; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6385 = 8'h28 == _T_375[7:0] ? 4'hf : _GEN_6384; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6386 = 8'h29 == _T_375[7:0] ? 4'hf : _GEN_6385; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6387 = 8'h2a == _T_375[7:0] ? 4'hf : _GEN_6386; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6388 = 8'h2b == _T_375[7:0] ? 4'hf : _GEN_6387; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6389 = 8'h2c == _T_375[7:0] ? 4'hf : _GEN_6388; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6390 = 8'h2d == _T_375[7:0] ? 4'hf : _GEN_6389; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6391 = 8'h2e == _T_375[7:0] ? 4'hf : _GEN_6390; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6392 = 8'h2f == _T_375[7:0] ? 4'hf : _GEN_6391; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6393 = 8'h30 == _T_375[7:0] ? 4'h0 : _GEN_6392; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6394 = 8'h31 == _T_375[7:0] ? 4'h0 : _GEN_6393; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6395 = 8'h32 == _T_375[7:0] ? 4'h0 : _GEN_6394; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6396 = 8'h33 == _T_375[7:0] ? 4'h0 : _GEN_6395; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6397 = 8'h34 == _T_375[7:0] ? 4'h0 : _GEN_6396; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6398 = 8'h35 == _T_375[7:0] ? 4'h0 : _GEN_6397; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6399 = 8'h36 == _T_375[7:0] ? 4'h0 : _GEN_6398; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6400 = 8'h37 == _T_375[7:0] ? 4'h0 : _GEN_6399; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6401 = 8'h38 == _T_375[7:0] ? 4'hf : _GEN_6400; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6402 = 8'h39 == _T_375[7:0] ? 4'hf : _GEN_6401; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6403 = 8'h3a == _T_375[7:0] ? 4'hf : _GEN_6402; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6404 = 8'h3b == _T_375[7:0] ? 4'hf : _GEN_6403; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6405 = 8'h3c == _T_375[7:0] ? 4'hf : _GEN_6404; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6406 = 8'h3d == _T_375[7:0] ? 4'hf : _GEN_6405; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6407 = 8'h3e == _T_375[7:0] ? 4'hf : _GEN_6406; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6408 = 8'h3f == _T_375[7:0] ? 4'hf : _GEN_6407; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6409 = 8'h40 == _T_375[7:0] ? 4'h0 : _GEN_6408; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6410 = 8'h41 == _T_375[7:0] ? 4'h0 : _GEN_6409; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6411 = 8'h42 == _T_375[7:0] ? 4'h0 : _GEN_6410; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6412 = 8'h43 == _T_375[7:0] ? 4'h0 : _GEN_6411; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6413 = 8'h44 == _T_375[7:0] ? 4'h0 : _GEN_6412; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6414 = 8'h45 == _T_375[7:0] ? 4'h0 : _GEN_6413; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6415 = 8'h46 == _T_375[7:0] ? 4'h0 : _GEN_6414; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6416 = 8'h47 == _T_375[7:0] ? 4'h0 : _GEN_6415; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6417 = 8'h48 == _T_375[7:0] ? 4'hf : _GEN_6416; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6418 = 8'h49 == _T_375[7:0] ? 4'hf : _GEN_6417; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6419 = 8'h4a == _T_375[7:0] ? 4'hf : _GEN_6418; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6420 = 8'h4b == _T_375[7:0] ? 4'hf : _GEN_6419; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6421 = 8'h4c == _T_375[7:0] ? 4'hf : _GEN_6420; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6422 = 8'h4d == _T_375[7:0] ? 4'hf : _GEN_6421; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6423 = 8'h4e == _T_375[7:0] ? 4'hf : _GEN_6422; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6424 = 8'h4f == _T_375[7:0] ? 4'hf : _GEN_6423; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6425 = 8'h50 == _T_375[7:0] ? 4'h0 : _GEN_6424; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6426 = 8'h51 == _T_375[7:0] ? 4'h0 : _GEN_6425; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6427 = 8'h52 == _T_375[7:0] ? 4'h0 : _GEN_6426; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6428 = 8'h53 == _T_375[7:0] ? 4'h0 : _GEN_6427; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6429 = 8'h54 == _T_375[7:0] ? 4'h0 : _GEN_6428; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6430 = 8'h55 == _T_375[7:0] ? 4'h0 : _GEN_6429; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6431 = 8'h56 == _T_375[7:0] ? 4'h0 : _GEN_6430; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6432 = 8'h57 == _T_375[7:0] ? 4'h0 : _GEN_6431; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6433 = 8'h58 == _T_375[7:0] ? 4'hf : _GEN_6432; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6434 = 8'h59 == _T_375[7:0] ? 4'hf : _GEN_6433; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6435 = 8'h5a == _T_375[7:0] ? 4'hf : _GEN_6434; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6436 = 8'h5b == _T_375[7:0] ? 4'hf : _GEN_6435; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6437 = 8'h5c == _T_375[7:0] ? 4'hf : _GEN_6436; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6438 = 8'h5d == _T_375[7:0] ? 4'hf : _GEN_6437; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6439 = 8'h5e == _T_375[7:0] ? 4'hf : _GEN_6438; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6440 = 8'h5f == _T_375[7:0] ? 4'hf : _GEN_6439; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6441 = 8'h60 == _T_375[7:0] ? 4'h0 : _GEN_6440; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6442 = 8'h61 == _T_375[7:0] ? 4'h0 : _GEN_6441; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6443 = 8'h62 == _T_375[7:0] ? 4'h0 : _GEN_6442; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6444 = 8'h63 == _T_375[7:0] ? 4'h0 : _GEN_6443; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6445 = 8'h64 == _T_375[7:0] ? 4'h0 : _GEN_6444; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6446 = 8'h65 == _T_375[7:0] ? 4'h0 : _GEN_6445; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6447 = 8'h66 == _T_375[7:0] ? 4'h0 : _GEN_6446; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6448 = 8'h67 == _T_375[7:0] ? 4'h0 : _GEN_6447; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6449 = 8'h68 == _T_375[7:0] ? 4'hf : _GEN_6448; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6450 = 8'h69 == _T_375[7:0] ? 4'hf : _GEN_6449; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6451 = 8'h6a == _T_375[7:0] ? 4'hf : _GEN_6450; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6452 = 8'h6b == _T_375[7:0] ? 4'hf : _GEN_6451; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6453 = 8'h6c == _T_375[7:0] ? 4'hf : _GEN_6452; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6454 = 8'h6d == _T_375[7:0] ? 4'hf : _GEN_6453; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6455 = 8'h6e == _T_375[7:0] ? 4'hf : _GEN_6454; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6456 = 8'h6f == _T_375[7:0] ? 4'hf : _GEN_6455; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6457 = 8'h70 == _T_375[7:0] ? 4'h0 : _GEN_6456; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6458 = 8'h71 == _T_375[7:0] ? 4'h0 : _GEN_6457; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6459 = 8'h72 == _T_375[7:0] ? 4'h0 : _GEN_6458; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6460 = 8'h73 == _T_375[7:0] ? 4'h0 : _GEN_6459; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6461 = 8'h74 == _T_375[7:0] ? 4'h0 : _GEN_6460; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6462 = 8'h75 == _T_375[7:0] ? 4'h0 : _GEN_6461; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6463 = 8'h76 == _T_375[7:0] ? 4'h0 : _GEN_6462; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6464 = 8'h77 == _T_375[7:0] ? 4'h0 : _GEN_6463; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6465 = 8'h78 == _T_375[7:0] ? 4'hf : _GEN_6464; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6466 = 8'h79 == _T_375[7:0] ? 4'hf : _GEN_6465; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6467 = 8'h7a == _T_375[7:0] ? 4'hf : _GEN_6466; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6468 = 8'h7b == _T_375[7:0] ? 4'hf : _GEN_6467; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6469 = 8'h7c == _T_375[7:0] ? 4'hf : _GEN_6468; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6470 = 8'h7d == _T_375[7:0] ? 4'hf : _GEN_6469; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6471 = 8'h7e == _T_375[7:0] ? 4'hf : _GEN_6470; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6472 = 8'h7f == _T_375[7:0] ? 4'hf : _GEN_6471; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6473 = 8'h80 == _T_375[7:0] ? 4'h0 : _GEN_6472; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6474 = 8'h81 == _T_375[7:0] ? 4'h0 : _GEN_6473; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6475 = 8'h82 == _T_375[7:0] ? 4'h0 : _GEN_6474; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6476 = 8'h83 == _T_375[7:0] ? 4'h0 : _GEN_6475; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6477 = 8'h84 == _T_375[7:0] ? 4'h0 : _GEN_6476; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6478 = 8'h85 == _T_375[7:0] ? 4'h0 : _GEN_6477; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6479 = 8'h86 == _T_375[7:0] ? 4'h0 : _GEN_6478; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6480 = 8'h87 == _T_375[7:0] ? 4'h0 : _GEN_6479; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6481 = 8'h88 == _T_375[7:0] ? 4'hf : _GEN_6480; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6482 = 8'h89 == _T_375[7:0] ? 4'hf : _GEN_6481; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6483 = 8'h8a == _T_375[7:0] ? 4'hf : _GEN_6482; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6484 = 8'h8b == _T_375[7:0] ? 4'hf : _GEN_6483; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6485 = 8'h8c == _T_375[7:0] ? 4'hf : _GEN_6484; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6486 = 8'h8d == _T_375[7:0] ? 4'hf : _GEN_6485; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6487 = 8'h8e == _T_375[7:0] ? 4'hf : _GEN_6486; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6488 = 8'h8f == _T_375[7:0] ? 4'hf : _GEN_6487; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6489 = 8'h90 == _T_375[7:0] ? 4'h0 : _GEN_6488; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6490 = 8'h91 == _T_375[7:0] ? 4'h0 : _GEN_6489; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6491 = 8'h92 == _T_375[7:0] ? 4'h0 : _GEN_6490; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6492 = 8'h93 == _T_375[7:0] ? 4'h0 : _GEN_6491; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6493 = 8'h94 == _T_375[7:0] ? 4'h0 : _GEN_6492; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6494 = 8'h95 == _T_375[7:0] ? 4'h0 : _GEN_6493; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6495 = 8'h96 == _T_375[7:0] ? 4'h0 : _GEN_6494; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6496 = 8'h97 == _T_375[7:0] ? 4'h0 : _GEN_6495; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6497 = 8'h98 == _T_375[7:0] ? 4'hf : _GEN_6496; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6498 = 8'h99 == _T_375[7:0] ? 4'hf : _GEN_6497; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6499 = 8'h9a == _T_375[7:0] ? 4'hf : _GEN_6498; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6500 = 8'h9b == _T_375[7:0] ? 4'hf : _GEN_6499; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6501 = 8'h9c == _T_375[7:0] ? 4'hf : _GEN_6500; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6502 = 8'h9d == _T_375[7:0] ? 4'hf : _GEN_6501; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6503 = 8'h9e == _T_375[7:0] ? 4'hf : _GEN_6502; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6504 = 8'h9f == _T_375[7:0] ? 4'hf : _GEN_6503; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6505 = 8'ha0 == _T_375[7:0] ? 4'h0 : _GEN_6504; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6506 = 8'ha1 == _T_375[7:0] ? 4'h0 : _GEN_6505; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6507 = 8'ha2 == _T_375[7:0] ? 4'h0 : _GEN_6506; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6508 = 8'ha3 == _T_375[7:0] ? 4'h0 : _GEN_6507; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6509 = 8'ha4 == _T_375[7:0] ? 4'h0 : _GEN_6508; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6510 = 8'ha5 == _T_375[7:0] ? 4'h0 : _GEN_6509; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6511 = 8'ha6 == _T_375[7:0] ? 4'h0 : _GEN_6510; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6512 = 8'ha7 == _T_375[7:0] ? 4'h0 : _GEN_6511; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6513 = 8'ha8 == _T_375[7:0] ? 4'hf : _GEN_6512; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6514 = 8'ha9 == _T_375[7:0] ? 4'hf : _GEN_6513; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6515 = 8'haa == _T_375[7:0] ? 4'hf : _GEN_6514; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6516 = 8'hab == _T_375[7:0] ? 4'hf : _GEN_6515; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6517 = 8'hac == _T_375[7:0] ? 4'hf : _GEN_6516; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6518 = 8'had == _T_375[7:0] ? 4'hf : _GEN_6517; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6519 = 8'hae == _T_375[7:0] ? 4'hf : _GEN_6518; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6520 = 8'haf == _T_375[7:0] ? 4'hf : _GEN_6519; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6521 = 8'hb0 == _T_375[7:0] ? 4'h0 : _GEN_6520; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6522 = 8'hb1 == _T_375[7:0] ? 4'h0 : _GEN_6521; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6523 = 8'hb2 == _T_375[7:0] ? 4'h0 : _GEN_6522; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6524 = 8'hb3 == _T_375[7:0] ? 4'h0 : _GEN_6523; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6525 = 8'hb4 == _T_375[7:0] ? 4'h0 : _GEN_6524; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6526 = 8'hb5 == _T_375[7:0] ? 4'h0 : _GEN_6525; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6527 = 8'hb6 == _T_375[7:0] ? 4'h0 : _GEN_6526; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6528 = 8'hb7 == _T_375[7:0] ? 4'h0 : _GEN_6527; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6529 = 8'hb8 == _T_375[7:0] ? 4'hf : _GEN_6528; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6530 = 8'hb9 == _T_375[7:0] ? 4'hf : _GEN_6529; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6531 = 8'hba == _T_375[7:0] ? 4'hf : _GEN_6530; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6532 = 8'hbb == _T_375[7:0] ? 4'hf : _GEN_6531; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6533 = 8'hbc == _T_375[7:0] ? 4'hf : _GEN_6532; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6534 = 8'hbd == _T_375[7:0] ? 4'hf : _GEN_6533; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6535 = 8'hbe == _T_375[7:0] ? 4'hf : _GEN_6534; // @[Filter.scala 160:142]
  wire [3:0] _GEN_6536 = 8'hbf == _T_375[7:0] ? 4'hf : _GEN_6535; // @[Filter.scala 160:142]
  wire [7:0] _T_389 = _GEN_6536 * 4'ha; // @[Filter.scala 160:142]
  wire [10:0] _GEN_9931 = {{3'd0}, _T_389}; // @[Filter.scala 160:109]
  wire [10:0] _T_391 = _T_384 + _GEN_9931; // @[Filter.scala 160:109]
  wire [10:0] _T_392 = _T_391 / 11'h64; // @[Filter.scala 160:150]
  wire  _T_394 = _T_365 >= 5'h10; // @[Filter.scala 163:31]
  wire  _T_398 = _T_372 >= 32'hc; // @[Filter.scala 163:63]
  wire  _T_399 = _T_394 | _T_398; // @[Filter.scala 163:58]
  wire [10:0] _GEN_6729 = io_SPI_distort ? _T_392 : {{7'd0}, _GEN_6152}; // @[Filter.scala 165:35]
  wire [10:0] _GEN_6730 = _T_399 ? 11'h0 : _GEN_6729; // @[Filter.scala 163:80]
  wire [10:0] _GEN_6923 = io_SPI_distort ? _T_392 : {{7'd0}, _GEN_6344}; // @[Filter.scala 165:35]
  wire [10:0] _GEN_6924 = _T_399 ? 11'h0 : _GEN_6923; // @[Filter.scala 163:80]
  wire [10:0] _GEN_7117 = io_SPI_distort ? _T_392 : {{7'd0}, _GEN_6536}; // @[Filter.scala 165:35]
  wire [10:0] _GEN_7118 = _T_399 ? 11'h0 : _GEN_7117; // @[Filter.scala 163:80]
  wire [31:0] _T_427 = pixelIndex + 32'h6; // @[Filter.scala 158:31]
  wire [31:0] _GEN_6 = _T_427 % 32'h10; // @[Filter.scala 158:38]
  wire [4:0] _T_428 = _GEN_6[4:0]; // @[Filter.scala 158:38]
  wire [4:0] _T_430 = _T_428 + _GEN_9863; // @[Filter.scala 158:53]
  wire [4:0] _T_432 = _T_430 - 5'h1; // @[Filter.scala 158:69]
  wire [31:0] _T_435 = _T_427 / 32'h10; // @[Filter.scala 159:38]
  wire [31:0] _T_437 = _T_435 + _GEN_9864; // @[Filter.scala 159:53]
  wire [31:0] _T_439 = _T_437 - 32'h1; // @[Filter.scala 159:69]
  wire [36:0] _T_440 = _T_439 * 32'h10; // @[Filter.scala 160:42]
  wire [36:0] _GEN_9937 = {{32'd0}, _T_432}; // @[Filter.scala 160:57]
  wire [36:0] _T_442 = _T_440 + _GEN_9937; // @[Filter.scala 160:57]
  wire [3:0] _GEN_7127 = 8'h8 == _T_442[7:0] ? 4'h0 : 4'hf; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7128 = 8'h9 == _T_442[7:0] ? 4'h0 : _GEN_7127; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7129 = 8'ha == _T_442[7:0] ? 4'h0 : _GEN_7128; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7130 = 8'hb == _T_442[7:0] ? 4'h0 : _GEN_7129; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7131 = 8'hc == _T_442[7:0] ? 4'h0 : _GEN_7130; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7132 = 8'hd == _T_442[7:0] ? 4'h0 : _GEN_7131; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7133 = 8'he == _T_442[7:0] ? 4'h0 : _GEN_7132; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7134 = 8'hf == _T_442[7:0] ? 4'h0 : _GEN_7133; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7135 = 8'h10 == _T_442[7:0] ? 4'hf : _GEN_7134; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7136 = 8'h11 == _T_442[7:0] ? 4'hf : _GEN_7135; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7137 = 8'h12 == _T_442[7:0] ? 4'hf : _GEN_7136; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7138 = 8'h13 == _T_442[7:0] ? 4'hf : _GEN_7137; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7139 = 8'h14 == _T_442[7:0] ? 4'hf : _GEN_7138; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7140 = 8'h15 == _T_442[7:0] ? 4'hf : _GEN_7139; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7141 = 8'h16 == _T_442[7:0] ? 4'hf : _GEN_7140; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7142 = 8'h17 == _T_442[7:0] ? 4'hf : _GEN_7141; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7143 = 8'h18 == _T_442[7:0] ? 4'h0 : _GEN_7142; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7144 = 8'h19 == _T_442[7:0] ? 4'h0 : _GEN_7143; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7145 = 8'h1a == _T_442[7:0] ? 4'h0 : _GEN_7144; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7146 = 8'h1b == _T_442[7:0] ? 4'h0 : _GEN_7145; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7147 = 8'h1c == _T_442[7:0] ? 4'h0 : _GEN_7146; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7148 = 8'h1d == _T_442[7:0] ? 4'h0 : _GEN_7147; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7149 = 8'h1e == _T_442[7:0] ? 4'h0 : _GEN_7148; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7150 = 8'h1f == _T_442[7:0] ? 4'h0 : _GEN_7149; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7151 = 8'h20 == _T_442[7:0] ? 4'hf : _GEN_7150; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7152 = 8'h21 == _T_442[7:0] ? 4'hf : _GEN_7151; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7153 = 8'h22 == _T_442[7:0] ? 4'hf : _GEN_7152; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7154 = 8'h23 == _T_442[7:0] ? 4'hf : _GEN_7153; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7155 = 8'h24 == _T_442[7:0] ? 4'hf : _GEN_7154; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7156 = 8'h25 == _T_442[7:0] ? 4'hf : _GEN_7155; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7157 = 8'h26 == _T_442[7:0] ? 4'hf : _GEN_7156; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7158 = 8'h27 == _T_442[7:0] ? 4'hf : _GEN_7157; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7159 = 8'h28 == _T_442[7:0] ? 4'h0 : _GEN_7158; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7160 = 8'h29 == _T_442[7:0] ? 4'h0 : _GEN_7159; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7161 = 8'h2a == _T_442[7:0] ? 4'h0 : _GEN_7160; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7162 = 8'h2b == _T_442[7:0] ? 4'h0 : _GEN_7161; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7163 = 8'h2c == _T_442[7:0] ? 4'h0 : _GEN_7162; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7164 = 8'h2d == _T_442[7:0] ? 4'h0 : _GEN_7163; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7165 = 8'h2e == _T_442[7:0] ? 4'h0 : _GEN_7164; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7166 = 8'h2f == _T_442[7:0] ? 4'h0 : _GEN_7165; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7167 = 8'h30 == _T_442[7:0] ? 4'hf : _GEN_7166; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7168 = 8'h31 == _T_442[7:0] ? 4'hf : _GEN_7167; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7169 = 8'h32 == _T_442[7:0] ? 4'hf : _GEN_7168; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7170 = 8'h33 == _T_442[7:0] ? 4'hf : _GEN_7169; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7171 = 8'h34 == _T_442[7:0] ? 4'hf : _GEN_7170; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7172 = 8'h35 == _T_442[7:0] ? 4'hf : _GEN_7171; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7173 = 8'h36 == _T_442[7:0] ? 4'hf : _GEN_7172; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7174 = 8'h37 == _T_442[7:0] ? 4'hf : _GEN_7173; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7175 = 8'h38 == _T_442[7:0] ? 4'h0 : _GEN_7174; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7176 = 8'h39 == _T_442[7:0] ? 4'h0 : _GEN_7175; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7177 = 8'h3a == _T_442[7:0] ? 4'h0 : _GEN_7176; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7178 = 8'h3b == _T_442[7:0] ? 4'h0 : _GEN_7177; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7179 = 8'h3c == _T_442[7:0] ? 4'h0 : _GEN_7178; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7180 = 8'h3d == _T_442[7:0] ? 4'h0 : _GEN_7179; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7181 = 8'h3e == _T_442[7:0] ? 4'h0 : _GEN_7180; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7182 = 8'h3f == _T_442[7:0] ? 4'h0 : _GEN_7181; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7183 = 8'h40 == _T_442[7:0] ? 4'hf : _GEN_7182; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7184 = 8'h41 == _T_442[7:0] ? 4'hf : _GEN_7183; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7185 = 8'h42 == _T_442[7:0] ? 4'hf : _GEN_7184; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7186 = 8'h43 == _T_442[7:0] ? 4'hf : _GEN_7185; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7187 = 8'h44 == _T_442[7:0] ? 4'hf : _GEN_7186; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7188 = 8'h45 == _T_442[7:0] ? 4'hf : _GEN_7187; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7189 = 8'h46 == _T_442[7:0] ? 4'hf : _GEN_7188; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7190 = 8'h47 == _T_442[7:0] ? 4'hf : _GEN_7189; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7191 = 8'h48 == _T_442[7:0] ? 4'h0 : _GEN_7190; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7192 = 8'h49 == _T_442[7:0] ? 4'h0 : _GEN_7191; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7193 = 8'h4a == _T_442[7:0] ? 4'h0 : _GEN_7192; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7194 = 8'h4b == _T_442[7:0] ? 4'h0 : _GEN_7193; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7195 = 8'h4c == _T_442[7:0] ? 4'h0 : _GEN_7194; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7196 = 8'h4d == _T_442[7:0] ? 4'h0 : _GEN_7195; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7197 = 8'h4e == _T_442[7:0] ? 4'h0 : _GEN_7196; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7198 = 8'h4f == _T_442[7:0] ? 4'h0 : _GEN_7197; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7199 = 8'h50 == _T_442[7:0] ? 4'hf : _GEN_7198; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7200 = 8'h51 == _T_442[7:0] ? 4'hf : _GEN_7199; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7201 = 8'h52 == _T_442[7:0] ? 4'hf : _GEN_7200; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7202 = 8'h53 == _T_442[7:0] ? 4'hf : _GEN_7201; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7203 = 8'h54 == _T_442[7:0] ? 4'hf : _GEN_7202; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7204 = 8'h55 == _T_442[7:0] ? 4'hf : _GEN_7203; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7205 = 8'h56 == _T_442[7:0] ? 4'hf : _GEN_7204; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7206 = 8'h57 == _T_442[7:0] ? 4'hf : _GEN_7205; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7207 = 8'h58 == _T_442[7:0] ? 4'h0 : _GEN_7206; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7208 = 8'h59 == _T_442[7:0] ? 4'h0 : _GEN_7207; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7209 = 8'h5a == _T_442[7:0] ? 4'h0 : _GEN_7208; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7210 = 8'h5b == _T_442[7:0] ? 4'h0 : _GEN_7209; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7211 = 8'h5c == _T_442[7:0] ? 4'h0 : _GEN_7210; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7212 = 8'h5d == _T_442[7:0] ? 4'h0 : _GEN_7211; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7213 = 8'h5e == _T_442[7:0] ? 4'h0 : _GEN_7212; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7214 = 8'h5f == _T_442[7:0] ? 4'h0 : _GEN_7213; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7215 = 8'h60 == _T_442[7:0] ? 4'h0 : _GEN_7214; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7216 = 8'h61 == _T_442[7:0] ? 4'h0 : _GEN_7215; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7217 = 8'h62 == _T_442[7:0] ? 4'h0 : _GEN_7216; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7218 = 8'h63 == _T_442[7:0] ? 4'h0 : _GEN_7217; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7219 = 8'h64 == _T_442[7:0] ? 4'h0 : _GEN_7218; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7220 = 8'h65 == _T_442[7:0] ? 4'h0 : _GEN_7219; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7221 = 8'h66 == _T_442[7:0] ? 4'h0 : _GEN_7220; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7222 = 8'h67 == _T_442[7:0] ? 4'h0 : _GEN_7221; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7223 = 8'h68 == _T_442[7:0] ? 4'hf : _GEN_7222; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7224 = 8'h69 == _T_442[7:0] ? 4'hf : _GEN_7223; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7225 = 8'h6a == _T_442[7:0] ? 4'hf : _GEN_7224; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7226 = 8'h6b == _T_442[7:0] ? 4'hf : _GEN_7225; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7227 = 8'h6c == _T_442[7:0] ? 4'hf : _GEN_7226; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7228 = 8'h6d == _T_442[7:0] ? 4'hf : _GEN_7227; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7229 = 8'h6e == _T_442[7:0] ? 4'hf : _GEN_7228; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7230 = 8'h6f == _T_442[7:0] ? 4'hf : _GEN_7229; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7231 = 8'h70 == _T_442[7:0] ? 4'h0 : _GEN_7230; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7232 = 8'h71 == _T_442[7:0] ? 4'h0 : _GEN_7231; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7233 = 8'h72 == _T_442[7:0] ? 4'h0 : _GEN_7232; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7234 = 8'h73 == _T_442[7:0] ? 4'h0 : _GEN_7233; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7235 = 8'h74 == _T_442[7:0] ? 4'h0 : _GEN_7234; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7236 = 8'h75 == _T_442[7:0] ? 4'h0 : _GEN_7235; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7237 = 8'h76 == _T_442[7:0] ? 4'h0 : _GEN_7236; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7238 = 8'h77 == _T_442[7:0] ? 4'h0 : _GEN_7237; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7239 = 8'h78 == _T_442[7:0] ? 4'hf : _GEN_7238; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7240 = 8'h79 == _T_442[7:0] ? 4'hf : _GEN_7239; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7241 = 8'h7a == _T_442[7:0] ? 4'hf : _GEN_7240; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7242 = 8'h7b == _T_442[7:0] ? 4'hf : _GEN_7241; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7243 = 8'h7c == _T_442[7:0] ? 4'hf : _GEN_7242; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7244 = 8'h7d == _T_442[7:0] ? 4'hf : _GEN_7243; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7245 = 8'h7e == _T_442[7:0] ? 4'hf : _GEN_7244; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7246 = 8'h7f == _T_442[7:0] ? 4'hf : _GEN_7245; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7247 = 8'h80 == _T_442[7:0] ? 4'h0 : _GEN_7246; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7248 = 8'h81 == _T_442[7:0] ? 4'h0 : _GEN_7247; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7249 = 8'h82 == _T_442[7:0] ? 4'h0 : _GEN_7248; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7250 = 8'h83 == _T_442[7:0] ? 4'h0 : _GEN_7249; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7251 = 8'h84 == _T_442[7:0] ? 4'h0 : _GEN_7250; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7252 = 8'h85 == _T_442[7:0] ? 4'h0 : _GEN_7251; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7253 = 8'h86 == _T_442[7:0] ? 4'h0 : _GEN_7252; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7254 = 8'h87 == _T_442[7:0] ? 4'h0 : _GEN_7253; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7255 = 8'h88 == _T_442[7:0] ? 4'hf : _GEN_7254; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7256 = 8'h89 == _T_442[7:0] ? 4'hf : _GEN_7255; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7257 = 8'h8a == _T_442[7:0] ? 4'hf : _GEN_7256; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7258 = 8'h8b == _T_442[7:0] ? 4'hf : _GEN_7257; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7259 = 8'h8c == _T_442[7:0] ? 4'hf : _GEN_7258; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7260 = 8'h8d == _T_442[7:0] ? 4'hf : _GEN_7259; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7261 = 8'h8e == _T_442[7:0] ? 4'hf : _GEN_7260; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7262 = 8'h8f == _T_442[7:0] ? 4'hf : _GEN_7261; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7263 = 8'h90 == _T_442[7:0] ? 4'h0 : _GEN_7262; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7264 = 8'h91 == _T_442[7:0] ? 4'h0 : _GEN_7263; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7265 = 8'h92 == _T_442[7:0] ? 4'h0 : _GEN_7264; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7266 = 8'h93 == _T_442[7:0] ? 4'h0 : _GEN_7265; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7267 = 8'h94 == _T_442[7:0] ? 4'h0 : _GEN_7266; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7268 = 8'h95 == _T_442[7:0] ? 4'h0 : _GEN_7267; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7269 = 8'h96 == _T_442[7:0] ? 4'h0 : _GEN_7268; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7270 = 8'h97 == _T_442[7:0] ? 4'h0 : _GEN_7269; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7271 = 8'h98 == _T_442[7:0] ? 4'hf : _GEN_7270; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7272 = 8'h99 == _T_442[7:0] ? 4'hf : _GEN_7271; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7273 = 8'h9a == _T_442[7:0] ? 4'hf : _GEN_7272; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7274 = 8'h9b == _T_442[7:0] ? 4'hf : _GEN_7273; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7275 = 8'h9c == _T_442[7:0] ? 4'hf : _GEN_7274; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7276 = 8'h9d == _T_442[7:0] ? 4'hf : _GEN_7275; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7277 = 8'h9e == _T_442[7:0] ? 4'hf : _GEN_7276; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7278 = 8'h9f == _T_442[7:0] ? 4'hf : _GEN_7277; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7279 = 8'ha0 == _T_442[7:0] ? 4'h0 : _GEN_7278; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7280 = 8'ha1 == _T_442[7:0] ? 4'h0 : _GEN_7279; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7281 = 8'ha2 == _T_442[7:0] ? 4'h0 : _GEN_7280; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7282 = 8'ha3 == _T_442[7:0] ? 4'h0 : _GEN_7281; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7283 = 8'ha4 == _T_442[7:0] ? 4'h0 : _GEN_7282; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7284 = 8'ha5 == _T_442[7:0] ? 4'h0 : _GEN_7283; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7285 = 8'ha6 == _T_442[7:0] ? 4'h0 : _GEN_7284; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7286 = 8'ha7 == _T_442[7:0] ? 4'h0 : _GEN_7285; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7287 = 8'ha8 == _T_442[7:0] ? 4'hf : _GEN_7286; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7288 = 8'ha9 == _T_442[7:0] ? 4'hf : _GEN_7287; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7289 = 8'haa == _T_442[7:0] ? 4'hf : _GEN_7288; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7290 = 8'hab == _T_442[7:0] ? 4'hf : _GEN_7289; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7291 = 8'hac == _T_442[7:0] ? 4'hf : _GEN_7290; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7292 = 8'had == _T_442[7:0] ? 4'hf : _GEN_7291; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7293 = 8'hae == _T_442[7:0] ? 4'hf : _GEN_7292; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7294 = 8'haf == _T_442[7:0] ? 4'hf : _GEN_7293; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7295 = 8'hb0 == _T_442[7:0] ? 4'h0 : _GEN_7294; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7296 = 8'hb1 == _T_442[7:0] ? 4'h0 : _GEN_7295; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7297 = 8'hb2 == _T_442[7:0] ? 4'h0 : _GEN_7296; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7298 = 8'hb3 == _T_442[7:0] ? 4'h0 : _GEN_7297; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7299 = 8'hb4 == _T_442[7:0] ? 4'h0 : _GEN_7298; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7300 = 8'hb5 == _T_442[7:0] ? 4'h0 : _GEN_7299; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7301 = 8'hb6 == _T_442[7:0] ? 4'h0 : _GEN_7300; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7302 = 8'hb7 == _T_442[7:0] ? 4'h0 : _GEN_7301; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7303 = 8'hb8 == _T_442[7:0] ? 4'hf : _GEN_7302; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7304 = 8'hb9 == _T_442[7:0] ? 4'hf : _GEN_7303; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7305 = 8'hba == _T_442[7:0] ? 4'hf : _GEN_7304; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7306 = 8'hbb == _T_442[7:0] ? 4'hf : _GEN_7305; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7307 = 8'hbc == _T_442[7:0] ? 4'hf : _GEN_7306; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7308 = 8'hbd == _T_442[7:0] ? 4'hf : _GEN_7307; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7309 = 8'hbe == _T_442[7:0] ? 4'hf : _GEN_7308; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7310 = 8'hbf == _T_442[7:0] ? 4'hf : _GEN_7309; // @[Filter.scala 160:62]
  wire [4:0] _GEN_9938 = {{1'd0}, _GEN_7310}; // @[Filter.scala 160:62]
  wire [8:0] _T_444 = _GEN_9938 * 5'h14; // @[Filter.scala 160:62]
  wire [3:0] _GEN_7407 = 8'h60 == _T_442[7:0] ? 4'hf : 4'h0; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7408 = 8'h61 == _T_442[7:0] ? 4'hf : _GEN_7407; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7409 = 8'h62 == _T_442[7:0] ? 4'hf : _GEN_7408; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7410 = 8'h63 == _T_442[7:0] ? 4'hf : _GEN_7409; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7411 = 8'h64 == _T_442[7:0] ? 4'hf : _GEN_7410; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7412 = 8'h65 == _T_442[7:0] ? 4'hf : _GEN_7411; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7413 = 8'h66 == _T_442[7:0] ? 4'hf : _GEN_7412; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7414 = 8'h67 == _T_442[7:0] ? 4'hf : _GEN_7413; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7415 = 8'h68 == _T_442[7:0] ? 4'hf : _GEN_7414; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7416 = 8'h69 == _T_442[7:0] ? 4'hf : _GEN_7415; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7417 = 8'h6a == _T_442[7:0] ? 4'hf : _GEN_7416; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7418 = 8'h6b == _T_442[7:0] ? 4'hf : _GEN_7417; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7419 = 8'h6c == _T_442[7:0] ? 4'hf : _GEN_7418; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7420 = 8'h6d == _T_442[7:0] ? 4'hf : _GEN_7419; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7421 = 8'h6e == _T_442[7:0] ? 4'hf : _GEN_7420; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7422 = 8'h6f == _T_442[7:0] ? 4'hf : _GEN_7421; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7423 = 8'h70 == _T_442[7:0] ? 4'hf : _GEN_7422; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7424 = 8'h71 == _T_442[7:0] ? 4'hf : _GEN_7423; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7425 = 8'h72 == _T_442[7:0] ? 4'hf : _GEN_7424; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7426 = 8'h73 == _T_442[7:0] ? 4'hf : _GEN_7425; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7427 = 8'h74 == _T_442[7:0] ? 4'hf : _GEN_7426; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7428 = 8'h75 == _T_442[7:0] ? 4'hf : _GEN_7427; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7429 = 8'h76 == _T_442[7:0] ? 4'hf : _GEN_7428; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7430 = 8'h77 == _T_442[7:0] ? 4'hf : _GEN_7429; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7431 = 8'h78 == _T_442[7:0] ? 4'hf : _GEN_7430; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7432 = 8'h79 == _T_442[7:0] ? 4'hf : _GEN_7431; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7433 = 8'h7a == _T_442[7:0] ? 4'hf : _GEN_7432; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7434 = 8'h7b == _T_442[7:0] ? 4'hf : _GEN_7433; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7435 = 8'h7c == _T_442[7:0] ? 4'hf : _GEN_7434; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7436 = 8'h7d == _T_442[7:0] ? 4'hf : _GEN_7435; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7437 = 8'h7e == _T_442[7:0] ? 4'hf : _GEN_7436; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7438 = 8'h7f == _T_442[7:0] ? 4'hf : _GEN_7437; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7439 = 8'h80 == _T_442[7:0] ? 4'hf : _GEN_7438; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7440 = 8'h81 == _T_442[7:0] ? 4'hf : _GEN_7439; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7441 = 8'h82 == _T_442[7:0] ? 4'hf : _GEN_7440; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7442 = 8'h83 == _T_442[7:0] ? 4'hf : _GEN_7441; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7443 = 8'h84 == _T_442[7:0] ? 4'hf : _GEN_7442; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7444 = 8'h85 == _T_442[7:0] ? 4'hf : _GEN_7443; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7445 = 8'h86 == _T_442[7:0] ? 4'hf : _GEN_7444; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7446 = 8'h87 == _T_442[7:0] ? 4'hf : _GEN_7445; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7447 = 8'h88 == _T_442[7:0] ? 4'hf : _GEN_7446; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7448 = 8'h89 == _T_442[7:0] ? 4'hf : _GEN_7447; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7449 = 8'h8a == _T_442[7:0] ? 4'hf : _GEN_7448; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7450 = 8'h8b == _T_442[7:0] ? 4'hf : _GEN_7449; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7451 = 8'h8c == _T_442[7:0] ? 4'hf : _GEN_7450; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7452 = 8'h8d == _T_442[7:0] ? 4'hf : _GEN_7451; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7453 = 8'h8e == _T_442[7:0] ? 4'hf : _GEN_7452; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7454 = 8'h8f == _T_442[7:0] ? 4'hf : _GEN_7453; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7455 = 8'h90 == _T_442[7:0] ? 4'hf : _GEN_7454; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7456 = 8'h91 == _T_442[7:0] ? 4'hf : _GEN_7455; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7457 = 8'h92 == _T_442[7:0] ? 4'hf : _GEN_7456; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7458 = 8'h93 == _T_442[7:0] ? 4'hf : _GEN_7457; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7459 = 8'h94 == _T_442[7:0] ? 4'hf : _GEN_7458; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7460 = 8'h95 == _T_442[7:0] ? 4'hf : _GEN_7459; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7461 = 8'h96 == _T_442[7:0] ? 4'hf : _GEN_7460; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7462 = 8'h97 == _T_442[7:0] ? 4'hf : _GEN_7461; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7463 = 8'h98 == _T_442[7:0] ? 4'hf : _GEN_7462; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7464 = 8'h99 == _T_442[7:0] ? 4'hf : _GEN_7463; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7465 = 8'h9a == _T_442[7:0] ? 4'hf : _GEN_7464; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7466 = 8'h9b == _T_442[7:0] ? 4'hf : _GEN_7465; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7467 = 8'h9c == _T_442[7:0] ? 4'hf : _GEN_7466; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7468 = 8'h9d == _T_442[7:0] ? 4'hf : _GEN_7467; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7469 = 8'h9e == _T_442[7:0] ? 4'hf : _GEN_7468; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7470 = 8'h9f == _T_442[7:0] ? 4'hf : _GEN_7469; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7471 = 8'ha0 == _T_442[7:0] ? 4'hf : _GEN_7470; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7472 = 8'ha1 == _T_442[7:0] ? 4'hf : _GEN_7471; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7473 = 8'ha2 == _T_442[7:0] ? 4'hf : _GEN_7472; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7474 = 8'ha3 == _T_442[7:0] ? 4'hf : _GEN_7473; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7475 = 8'ha4 == _T_442[7:0] ? 4'hf : _GEN_7474; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7476 = 8'ha5 == _T_442[7:0] ? 4'hf : _GEN_7475; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7477 = 8'ha6 == _T_442[7:0] ? 4'hf : _GEN_7476; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7478 = 8'ha7 == _T_442[7:0] ? 4'hf : _GEN_7477; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7479 = 8'ha8 == _T_442[7:0] ? 4'hf : _GEN_7478; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7480 = 8'ha9 == _T_442[7:0] ? 4'hf : _GEN_7479; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7481 = 8'haa == _T_442[7:0] ? 4'hf : _GEN_7480; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7482 = 8'hab == _T_442[7:0] ? 4'hf : _GEN_7481; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7483 = 8'hac == _T_442[7:0] ? 4'hf : _GEN_7482; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7484 = 8'had == _T_442[7:0] ? 4'hf : _GEN_7483; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7485 = 8'hae == _T_442[7:0] ? 4'hf : _GEN_7484; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7486 = 8'haf == _T_442[7:0] ? 4'hf : _GEN_7485; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7487 = 8'hb0 == _T_442[7:0] ? 4'hf : _GEN_7486; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7488 = 8'hb1 == _T_442[7:0] ? 4'hf : _GEN_7487; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7489 = 8'hb2 == _T_442[7:0] ? 4'hf : _GEN_7488; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7490 = 8'hb3 == _T_442[7:0] ? 4'hf : _GEN_7489; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7491 = 8'hb4 == _T_442[7:0] ? 4'hf : _GEN_7490; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7492 = 8'hb5 == _T_442[7:0] ? 4'hf : _GEN_7491; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7493 = 8'hb6 == _T_442[7:0] ? 4'hf : _GEN_7492; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7494 = 8'hb7 == _T_442[7:0] ? 4'hf : _GEN_7493; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7495 = 8'hb8 == _T_442[7:0] ? 4'hf : _GEN_7494; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7496 = 8'hb9 == _T_442[7:0] ? 4'hf : _GEN_7495; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7497 = 8'hba == _T_442[7:0] ? 4'hf : _GEN_7496; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7498 = 8'hbb == _T_442[7:0] ? 4'hf : _GEN_7497; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7499 = 8'hbc == _T_442[7:0] ? 4'hf : _GEN_7498; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7500 = 8'hbd == _T_442[7:0] ? 4'hf : _GEN_7499; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7501 = 8'hbe == _T_442[7:0] ? 4'hf : _GEN_7500; // @[Filter.scala 160:102]
  wire [3:0] _GEN_7502 = 8'hbf == _T_442[7:0] ? 4'hf : _GEN_7501; // @[Filter.scala 160:102]
  wire [6:0] _GEN_9940 = {{3'd0}, _GEN_7502}; // @[Filter.scala 160:102]
  wire [10:0] _T_449 = _GEN_9940 * 7'h46; // @[Filter.scala 160:102]
  wire [10:0] _GEN_9941 = {{2'd0}, _T_444}; // @[Filter.scala 160:69]
  wire [10:0] _T_451 = _GEN_9941 + _T_449; // @[Filter.scala 160:69]
  wire [3:0] _GEN_7511 = 8'h8 == _T_442[7:0] ? 4'hf : 4'h0; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7512 = 8'h9 == _T_442[7:0] ? 4'hf : _GEN_7511; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7513 = 8'ha == _T_442[7:0] ? 4'hf : _GEN_7512; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7514 = 8'hb == _T_442[7:0] ? 4'hf : _GEN_7513; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7515 = 8'hc == _T_442[7:0] ? 4'hf : _GEN_7514; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7516 = 8'hd == _T_442[7:0] ? 4'hf : _GEN_7515; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7517 = 8'he == _T_442[7:0] ? 4'hf : _GEN_7516; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7518 = 8'hf == _T_442[7:0] ? 4'hf : _GEN_7517; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7519 = 8'h10 == _T_442[7:0] ? 4'h0 : _GEN_7518; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7520 = 8'h11 == _T_442[7:0] ? 4'h0 : _GEN_7519; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7521 = 8'h12 == _T_442[7:0] ? 4'h0 : _GEN_7520; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7522 = 8'h13 == _T_442[7:0] ? 4'h0 : _GEN_7521; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7523 = 8'h14 == _T_442[7:0] ? 4'h0 : _GEN_7522; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7524 = 8'h15 == _T_442[7:0] ? 4'h0 : _GEN_7523; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7525 = 8'h16 == _T_442[7:0] ? 4'h0 : _GEN_7524; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7526 = 8'h17 == _T_442[7:0] ? 4'h0 : _GEN_7525; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7527 = 8'h18 == _T_442[7:0] ? 4'hf : _GEN_7526; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7528 = 8'h19 == _T_442[7:0] ? 4'hf : _GEN_7527; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7529 = 8'h1a == _T_442[7:0] ? 4'hf : _GEN_7528; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7530 = 8'h1b == _T_442[7:0] ? 4'hf : _GEN_7529; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7531 = 8'h1c == _T_442[7:0] ? 4'hf : _GEN_7530; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7532 = 8'h1d == _T_442[7:0] ? 4'hf : _GEN_7531; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7533 = 8'h1e == _T_442[7:0] ? 4'hf : _GEN_7532; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7534 = 8'h1f == _T_442[7:0] ? 4'hf : _GEN_7533; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7535 = 8'h20 == _T_442[7:0] ? 4'h0 : _GEN_7534; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7536 = 8'h21 == _T_442[7:0] ? 4'h0 : _GEN_7535; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7537 = 8'h22 == _T_442[7:0] ? 4'h0 : _GEN_7536; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7538 = 8'h23 == _T_442[7:0] ? 4'h0 : _GEN_7537; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7539 = 8'h24 == _T_442[7:0] ? 4'h0 : _GEN_7538; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7540 = 8'h25 == _T_442[7:0] ? 4'h0 : _GEN_7539; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7541 = 8'h26 == _T_442[7:0] ? 4'h0 : _GEN_7540; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7542 = 8'h27 == _T_442[7:0] ? 4'h0 : _GEN_7541; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7543 = 8'h28 == _T_442[7:0] ? 4'hf : _GEN_7542; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7544 = 8'h29 == _T_442[7:0] ? 4'hf : _GEN_7543; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7545 = 8'h2a == _T_442[7:0] ? 4'hf : _GEN_7544; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7546 = 8'h2b == _T_442[7:0] ? 4'hf : _GEN_7545; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7547 = 8'h2c == _T_442[7:0] ? 4'hf : _GEN_7546; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7548 = 8'h2d == _T_442[7:0] ? 4'hf : _GEN_7547; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7549 = 8'h2e == _T_442[7:0] ? 4'hf : _GEN_7548; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7550 = 8'h2f == _T_442[7:0] ? 4'hf : _GEN_7549; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7551 = 8'h30 == _T_442[7:0] ? 4'h0 : _GEN_7550; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7552 = 8'h31 == _T_442[7:0] ? 4'h0 : _GEN_7551; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7553 = 8'h32 == _T_442[7:0] ? 4'h0 : _GEN_7552; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7554 = 8'h33 == _T_442[7:0] ? 4'h0 : _GEN_7553; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7555 = 8'h34 == _T_442[7:0] ? 4'h0 : _GEN_7554; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7556 = 8'h35 == _T_442[7:0] ? 4'h0 : _GEN_7555; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7557 = 8'h36 == _T_442[7:0] ? 4'h0 : _GEN_7556; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7558 = 8'h37 == _T_442[7:0] ? 4'h0 : _GEN_7557; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7559 = 8'h38 == _T_442[7:0] ? 4'hf : _GEN_7558; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7560 = 8'h39 == _T_442[7:0] ? 4'hf : _GEN_7559; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7561 = 8'h3a == _T_442[7:0] ? 4'hf : _GEN_7560; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7562 = 8'h3b == _T_442[7:0] ? 4'hf : _GEN_7561; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7563 = 8'h3c == _T_442[7:0] ? 4'hf : _GEN_7562; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7564 = 8'h3d == _T_442[7:0] ? 4'hf : _GEN_7563; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7565 = 8'h3e == _T_442[7:0] ? 4'hf : _GEN_7564; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7566 = 8'h3f == _T_442[7:0] ? 4'hf : _GEN_7565; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7567 = 8'h40 == _T_442[7:0] ? 4'h0 : _GEN_7566; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7568 = 8'h41 == _T_442[7:0] ? 4'h0 : _GEN_7567; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7569 = 8'h42 == _T_442[7:0] ? 4'h0 : _GEN_7568; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7570 = 8'h43 == _T_442[7:0] ? 4'h0 : _GEN_7569; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7571 = 8'h44 == _T_442[7:0] ? 4'h0 : _GEN_7570; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7572 = 8'h45 == _T_442[7:0] ? 4'h0 : _GEN_7571; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7573 = 8'h46 == _T_442[7:0] ? 4'h0 : _GEN_7572; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7574 = 8'h47 == _T_442[7:0] ? 4'h0 : _GEN_7573; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7575 = 8'h48 == _T_442[7:0] ? 4'hf : _GEN_7574; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7576 = 8'h49 == _T_442[7:0] ? 4'hf : _GEN_7575; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7577 = 8'h4a == _T_442[7:0] ? 4'hf : _GEN_7576; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7578 = 8'h4b == _T_442[7:0] ? 4'hf : _GEN_7577; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7579 = 8'h4c == _T_442[7:0] ? 4'hf : _GEN_7578; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7580 = 8'h4d == _T_442[7:0] ? 4'hf : _GEN_7579; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7581 = 8'h4e == _T_442[7:0] ? 4'hf : _GEN_7580; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7582 = 8'h4f == _T_442[7:0] ? 4'hf : _GEN_7581; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7583 = 8'h50 == _T_442[7:0] ? 4'h0 : _GEN_7582; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7584 = 8'h51 == _T_442[7:0] ? 4'h0 : _GEN_7583; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7585 = 8'h52 == _T_442[7:0] ? 4'h0 : _GEN_7584; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7586 = 8'h53 == _T_442[7:0] ? 4'h0 : _GEN_7585; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7587 = 8'h54 == _T_442[7:0] ? 4'h0 : _GEN_7586; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7588 = 8'h55 == _T_442[7:0] ? 4'h0 : _GEN_7587; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7589 = 8'h56 == _T_442[7:0] ? 4'h0 : _GEN_7588; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7590 = 8'h57 == _T_442[7:0] ? 4'h0 : _GEN_7589; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7591 = 8'h58 == _T_442[7:0] ? 4'hf : _GEN_7590; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7592 = 8'h59 == _T_442[7:0] ? 4'hf : _GEN_7591; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7593 = 8'h5a == _T_442[7:0] ? 4'hf : _GEN_7592; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7594 = 8'h5b == _T_442[7:0] ? 4'hf : _GEN_7593; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7595 = 8'h5c == _T_442[7:0] ? 4'hf : _GEN_7594; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7596 = 8'h5d == _T_442[7:0] ? 4'hf : _GEN_7595; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7597 = 8'h5e == _T_442[7:0] ? 4'hf : _GEN_7596; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7598 = 8'h5f == _T_442[7:0] ? 4'hf : _GEN_7597; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7599 = 8'h60 == _T_442[7:0] ? 4'h0 : _GEN_7598; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7600 = 8'h61 == _T_442[7:0] ? 4'h0 : _GEN_7599; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7601 = 8'h62 == _T_442[7:0] ? 4'h0 : _GEN_7600; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7602 = 8'h63 == _T_442[7:0] ? 4'h0 : _GEN_7601; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7603 = 8'h64 == _T_442[7:0] ? 4'h0 : _GEN_7602; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7604 = 8'h65 == _T_442[7:0] ? 4'h0 : _GEN_7603; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7605 = 8'h66 == _T_442[7:0] ? 4'h0 : _GEN_7604; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7606 = 8'h67 == _T_442[7:0] ? 4'h0 : _GEN_7605; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7607 = 8'h68 == _T_442[7:0] ? 4'hf : _GEN_7606; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7608 = 8'h69 == _T_442[7:0] ? 4'hf : _GEN_7607; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7609 = 8'h6a == _T_442[7:0] ? 4'hf : _GEN_7608; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7610 = 8'h6b == _T_442[7:0] ? 4'hf : _GEN_7609; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7611 = 8'h6c == _T_442[7:0] ? 4'hf : _GEN_7610; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7612 = 8'h6d == _T_442[7:0] ? 4'hf : _GEN_7611; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7613 = 8'h6e == _T_442[7:0] ? 4'hf : _GEN_7612; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7614 = 8'h6f == _T_442[7:0] ? 4'hf : _GEN_7613; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7615 = 8'h70 == _T_442[7:0] ? 4'h0 : _GEN_7614; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7616 = 8'h71 == _T_442[7:0] ? 4'h0 : _GEN_7615; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7617 = 8'h72 == _T_442[7:0] ? 4'h0 : _GEN_7616; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7618 = 8'h73 == _T_442[7:0] ? 4'h0 : _GEN_7617; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7619 = 8'h74 == _T_442[7:0] ? 4'h0 : _GEN_7618; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7620 = 8'h75 == _T_442[7:0] ? 4'h0 : _GEN_7619; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7621 = 8'h76 == _T_442[7:0] ? 4'h0 : _GEN_7620; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7622 = 8'h77 == _T_442[7:0] ? 4'h0 : _GEN_7621; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7623 = 8'h78 == _T_442[7:0] ? 4'hf : _GEN_7622; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7624 = 8'h79 == _T_442[7:0] ? 4'hf : _GEN_7623; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7625 = 8'h7a == _T_442[7:0] ? 4'hf : _GEN_7624; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7626 = 8'h7b == _T_442[7:0] ? 4'hf : _GEN_7625; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7627 = 8'h7c == _T_442[7:0] ? 4'hf : _GEN_7626; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7628 = 8'h7d == _T_442[7:0] ? 4'hf : _GEN_7627; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7629 = 8'h7e == _T_442[7:0] ? 4'hf : _GEN_7628; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7630 = 8'h7f == _T_442[7:0] ? 4'hf : _GEN_7629; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7631 = 8'h80 == _T_442[7:0] ? 4'h0 : _GEN_7630; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7632 = 8'h81 == _T_442[7:0] ? 4'h0 : _GEN_7631; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7633 = 8'h82 == _T_442[7:0] ? 4'h0 : _GEN_7632; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7634 = 8'h83 == _T_442[7:0] ? 4'h0 : _GEN_7633; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7635 = 8'h84 == _T_442[7:0] ? 4'h0 : _GEN_7634; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7636 = 8'h85 == _T_442[7:0] ? 4'h0 : _GEN_7635; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7637 = 8'h86 == _T_442[7:0] ? 4'h0 : _GEN_7636; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7638 = 8'h87 == _T_442[7:0] ? 4'h0 : _GEN_7637; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7639 = 8'h88 == _T_442[7:0] ? 4'hf : _GEN_7638; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7640 = 8'h89 == _T_442[7:0] ? 4'hf : _GEN_7639; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7641 = 8'h8a == _T_442[7:0] ? 4'hf : _GEN_7640; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7642 = 8'h8b == _T_442[7:0] ? 4'hf : _GEN_7641; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7643 = 8'h8c == _T_442[7:0] ? 4'hf : _GEN_7642; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7644 = 8'h8d == _T_442[7:0] ? 4'hf : _GEN_7643; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7645 = 8'h8e == _T_442[7:0] ? 4'hf : _GEN_7644; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7646 = 8'h8f == _T_442[7:0] ? 4'hf : _GEN_7645; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7647 = 8'h90 == _T_442[7:0] ? 4'h0 : _GEN_7646; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7648 = 8'h91 == _T_442[7:0] ? 4'h0 : _GEN_7647; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7649 = 8'h92 == _T_442[7:0] ? 4'h0 : _GEN_7648; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7650 = 8'h93 == _T_442[7:0] ? 4'h0 : _GEN_7649; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7651 = 8'h94 == _T_442[7:0] ? 4'h0 : _GEN_7650; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7652 = 8'h95 == _T_442[7:0] ? 4'h0 : _GEN_7651; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7653 = 8'h96 == _T_442[7:0] ? 4'h0 : _GEN_7652; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7654 = 8'h97 == _T_442[7:0] ? 4'h0 : _GEN_7653; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7655 = 8'h98 == _T_442[7:0] ? 4'hf : _GEN_7654; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7656 = 8'h99 == _T_442[7:0] ? 4'hf : _GEN_7655; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7657 = 8'h9a == _T_442[7:0] ? 4'hf : _GEN_7656; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7658 = 8'h9b == _T_442[7:0] ? 4'hf : _GEN_7657; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7659 = 8'h9c == _T_442[7:0] ? 4'hf : _GEN_7658; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7660 = 8'h9d == _T_442[7:0] ? 4'hf : _GEN_7659; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7661 = 8'h9e == _T_442[7:0] ? 4'hf : _GEN_7660; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7662 = 8'h9f == _T_442[7:0] ? 4'hf : _GEN_7661; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7663 = 8'ha0 == _T_442[7:0] ? 4'h0 : _GEN_7662; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7664 = 8'ha1 == _T_442[7:0] ? 4'h0 : _GEN_7663; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7665 = 8'ha2 == _T_442[7:0] ? 4'h0 : _GEN_7664; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7666 = 8'ha3 == _T_442[7:0] ? 4'h0 : _GEN_7665; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7667 = 8'ha4 == _T_442[7:0] ? 4'h0 : _GEN_7666; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7668 = 8'ha5 == _T_442[7:0] ? 4'h0 : _GEN_7667; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7669 = 8'ha6 == _T_442[7:0] ? 4'h0 : _GEN_7668; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7670 = 8'ha7 == _T_442[7:0] ? 4'h0 : _GEN_7669; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7671 = 8'ha8 == _T_442[7:0] ? 4'hf : _GEN_7670; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7672 = 8'ha9 == _T_442[7:0] ? 4'hf : _GEN_7671; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7673 = 8'haa == _T_442[7:0] ? 4'hf : _GEN_7672; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7674 = 8'hab == _T_442[7:0] ? 4'hf : _GEN_7673; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7675 = 8'hac == _T_442[7:0] ? 4'hf : _GEN_7674; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7676 = 8'had == _T_442[7:0] ? 4'hf : _GEN_7675; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7677 = 8'hae == _T_442[7:0] ? 4'hf : _GEN_7676; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7678 = 8'haf == _T_442[7:0] ? 4'hf : _GEN_7677; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7679 = 8'hb0 == _T_442[7:0] ? 4'h0 : _GEN_7678; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7680 = 8'hb1 == _T_442[7:0] ? 4'h0 : _GEN_7679; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7681 = 8'hb2 == _T_442[7:0] ? 4'h0 : _GEN_7680; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7682 = 8'hb3 == _T_442[7:0] ? 4'h0 : _GEN_7681; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7683 = 8'hb4 == _T_442[7:0] ? 4'h0 : _GEN_7682; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7684 = 8'hb5 == _T_442[7:0] ? 4'h0 : _GEN_7683; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7685 = 8'hb6 == _T_442[7:0] ? 4'h0 : _GEN_7684; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7686 = 8'hb7 == _T_442[7:0] ? 4'h0 : _GEN_7685; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7687 = 8'hb8 == _T_442[7:0] ? 4'hf : _GEN_7686; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7688 = 8'hb9 == _T_442[7:0] ? 4'hf : _GEN_7687; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7689 = 8'hba == _T_442[7:0] ? 4'hf : _GEN_7688; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7690 = 8'hbb == _T_442[7:0] ? 4'hf : _GEN_7689; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7691 = 8'hbc == _T_442[7:0] ? 4'hf : _GEN_7690; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7692 = 8'hbd == _T_442[7:0] ? 4'hf : _GEN_7691; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7693 = 8'hbe == _T_442[7:0] ? 4'hf : _GEN_7692; // @[Filter.scala 160:142]
  wire [3:0] _GEN_7694 = 8'hbf == _T_442[7:0] ? 4'hf : _GEN_7693; // @[Filter.scala 160:142]
  wire [7:0] _T_456 = _GEN_7694 * 4'ha; // @[Filter.scala 160:142]
  wire [10:0] _GEN_9943 = {{3'd0}, _T_456}; // @[Filter.scala 160:109]
  wire [10:0] _T_458 = _T_451 + _GEN_9943; // @[Filter.scala 160:109]
  wire [10:0] _T_459 = _T_458 / 11'h64; // @[Filter.scala 160:150]
  wire  _T_461 = _T_432 >= 5'h10; // @[Filter.scala 163:31]
  wire  _T_465 = _T_439 >= 32'hc; // @[Filter.scala 163:63]
  wire  _T_466 = _T_461 | _T_465; // @[Filter.scala 163:58]
  wire [10:0] _GEN_7887 = io_SPI_distort ? _T_459 : {{7'd0}, _GEN_7310}; // @[Filter.scala 165:35]
  wire [10:0] _GEN_7888 = _T_466 ? 11'h0 : _GEN_7887; // @[Filter.scala 163:80]
  wire [10:0] _GEN_8081 = io_SPI_distort ? _T_459 : {{7'd0}, _GEN_7502}; // @[Filter.scala 165:35]
  wire [10:0] _GEN_8082 = _T_466 ? 11'h0 : _GEN_8081; // @[Filter.scala 163:80]
  wire [10:0] _GEN_8275 = io_SPI_distort ? _T_459 : {{7'd0}, _GEN_7694}; // @[Filter.scala 165:35]
  wire [10:0] _GEN_8276 = _T_466 ? 11'h0 : _GEN_8275; // @[Filter.scala 163:80]
  wire [31:0] _T_494 = pixelIndex + 32'h7; // @[Filter.scala 158:31]
  wire [31:0] _GEN_56 = _T_494 % 32'h10; // @[Filter.scala 158:38]
  wire [4:0] _T_495 = _GEN_56[4:0]; // @[Filter.scala 158:38]
  wire [4:0] _T_497 = _T_495 + _GEN_9863; // @[Filter.scala 158:53]
  wire [4:0] _T_499 = _T_497 - 5'h1; // @[Filter.scala 158:69]
  wire [31:0] _T_502 = _T_494 / 32'h10; // @[Filter.scala 159:38]
  wire [31:0] _T_504 = _T_502 + _GEN_9864; // @[Filter.scala 159:53]
  wire [31:0] _T_506 = _T_504 - 32'h1; // @[Filter.scala 159:69]
  wire [36:0] _T_507 = _T_506 * 32'h10; // @[Filter.scala 160:42]
  wire [36:0] _GEN_9949 = {{32'd0}, _T_499}; // @[Filter.scala 160:57]
  wire [36:0] _T_509 = _T_507 + _GEN_9949; // @[Filter.scala 160:57]
  wire [3:0] _GEN_8285 = 8'h8 == _T_509[7:0] ? 4'h0 : 4'hf; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8286 = 8'h9 == _T_509[7:0] ? 4'h0 : _GEN_8285; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8287 = 8'ha == _T_509[7:0] ? 4'h0 : _GEN_8286; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8288 = 8'hb == _T_509[7:0] ? 4'h0 : _GEN_8287; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8289 = 8'hc == _T_509[7:0] ? 4'h0 : _GEN_8288; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8290 = 8'hd == _T_509[7:0] ? 4'h0 : _GEN_8289; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8291 = 8'he == _T_509[7:0] ? 4'h0 : _GEN_8290; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8292 = 8'hf == _T_509[7:0] ? 4'h0 : _GEN_8291; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8293 = 8'h10 == _T_509[7:0] ? 4'hf : _GEN_8292; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8294 = 8'h11 == _T_509[7:0] ? 4'hf : _GEN_8293; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8295 = 8'h12 == _T_509[7:0] ? 4'hf : _GEN_8294; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8296 = 8'h13 == _T_509[7:0] ? 4'hf : _GEN_8295; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8297 = 8'h14 == _T_509[7:0] ? 4'hf : _GEN_8296; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8298 = 8'h15 == _T_509[7:0] ? 4'hf : _GEN_8297; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8299 = 8'h16 == _T_509[7:0] ? 4'hf : _GEN_8298; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8300 = 8'h17 == _T_509[7:0] ? 4'hf : _GEN_8299; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8301 = 8'h18 == _T_509[7:0] ? 4'h0 : _GEN_8300; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8302 = 8'h19 == _T_509[7:0] ? 4'h0 : _GEN_8301; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8303 = 8'h1a == _T_509[7:0] ? 4'h0 : _GEN_8302; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8304 = 8'h1b == _T_509[7:0] ? 4'h0 : _GEN_8303; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8305 = 8'h1c == _T_509[7:0] ? 4'h0 : _GEN_8304; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8306 = 8'h1d == _T_509[7:0] ? 4'h0 : _GEN_8305; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8307 = 8'h1e == _T_509[7:0] ? 4'h0 : _GEN_8306; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8308 = 8'h1f == _T_509[7:0] ? 4'h0 : _GEN_8307; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8309 = 8'h20 == _T_509[7:0] ? 4'hf : _GEN_8308; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8310 = 8'h21 == _T_509[7:0] ? 4'hf : _GEN_8309; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8311 = 8'h22 == _T_509[7:0] ? 4'hf : _GEN_8310; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8312 = 8'h23 == _T_509[7:0] ? 4'hf : _GEN_8311; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8313 = 8'h24 == _T_509[7:0] ? 4'hf : _GEN_8312; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8314 = 8'h25 == _T_509[7:0] ? 4'hf : _GEN_8313; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8315 = 8'h26 == _T_509[7:0] ? 4'hf : _GEN_8314; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8316 = 8'h27 == _T_509[7:0] ? 4'hf : _GEN_8315; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8317 = 8'h28 == _T_509[7:0] ? 4'h0 : _GEN_8316; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8318 = 8'h29 == _T_509[7:0] ? 4'h0 : _GEN_8317; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8319 = 8'h2a == _T_509[7:0] ? 4'h0 : _GEN_8318; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8320 = 8'h2b == _T_509[7:0] ? 4'h0 : _GEN_8319; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8321 = 8'h2c == _T_509[7:0] ? 4'h0 : _GEN_8320; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8322 = 8'h2d == _T_509[7:0] ? 4'h0 : _GEN_8321; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8323 = 8'h2e == _T_509[7:0] ? 4'h0 : _GEN_8322; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8324 = 8'h2f == _T_509[7:0] ? 4'h0 : _GEN_8323; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8325 = 8'h30 == _T_509[7:0] ? 4'hf : _GEN_8324; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8326 = 8'h31 == _T_509[7:0] ? 4'hf : _GEN_8325; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8327 = 8'h32 == _T_509[7:0] ? 4'hf : _GEN_8326; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8328 = 8'h33 == _T_509[7:0] ? 4'hf : _GEN_8327; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8329 = 8'h34 == _T_509[7:0] ? 4'hf : _GEN_8328; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8330 = 8'h35 == _T_509[7:0] ? 4'hf : _GEN_8329; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8331 = 8'h36 == _T_509[7:0] ? 4'hf : _GEN_8330; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8332 = 8'h37 == _T_509[7:0] ? 4'hf : _GEN_8331; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8333 = 8'h38 == _T_509[7:0] ? 4'h0 : _GEN_8332; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8334 = 8'h39 == _T_509[7:0] ? 4'h0 : _GEN_8333; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8335 = 8'h3a == _T_509[7:0] ? 4'h0 : _GEN_8334; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8336 = 8'h3b == _T_509[7:0] ? 4'h0 : _GEN_8335; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8337 = 8'h3c == _T_509[7:0] ? 4'h0 : _GEN_8336; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8338 = 8'h3d == _T_509[7:0] ? 4'h0 : _GEN_8337; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8339 = 8'h3e == _T_509[7:0] ? 4'h0 : _GEN_8338; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8340 = 8'h3f == _T_509[7:0] ? 4'h0 : _GEN_8339; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8341 = 8'h40 == _T_509[7:0] ? 4'hf : _GEN_8340; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8342 = 8'h41 == _T_509[7:0] ? 4'hf : _GEN_8341; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8343 = 8'h42 == _T_509[7:0] ? 4'hf : _GEN_8342; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8344 = 8'h43 == _T_509[7:0] ? 4'hf : _GEN_8343; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8345 = 8'h44 == _T_509[7:0] ? 4'hf : _GEN_8344; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8346 = 8'h45 == _T_509[7:0] ? 4'hf : _GEN_8345; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8347 = 8'h46 == _T_509[7:0] ? 4'hf : _GEN_8346; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8348 = 8'h47 == _T_509[7:0] ? 4'hf : _GEN_8347; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8349 = 8'h48 == _T_509[7:0] ? 4'h0 : _GEN_8348; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8350 = 8'h49 == _T_509[7:0] ? 4'h0 : _GEN_8349; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8351 = 8'h4a == _T_509[7:0] ? 4'h0 : _GEN_8350; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8352 = 8'h4b == _T_509[7:0] ? 4'h0 : _GEN_8351; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8353 = 8'h4c == _T_509[7:0] ? 4'h0 : _GEN_8352; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8354 = 8'h4d == _T_509[7:0] ? 4'h0 : _GEN_8353; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8355 = 8'h4e == _T_509[7:0] ? 4'h0 : _GEN_8354; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8356 = 8'h4f == _T_509[7:0] ? 4'h0 : _GEN_8355; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8357 = 8'h50 == _T_509[7:0] ? 4'hf : _GEN_8356; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8358 = 8'h51 == _T_509[7:0] ? 4'hf : _GEN_8357; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8359 = 8'h52 == _T_509[7:0] ? 4'hf : _GEN_8358; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8360 = 8'h53 == _T_509[7:0] ? 4'hf : _GEN_8359; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8361 = 8'h54 == _T_509[7:0] ? 4'hf : _GEN_8360; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8362 = 8'h55 == _T_509[7:0] ? 4'hf : _GEN_8361; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8363 = 8'h56 == _T_509[7:0] ? 4'hf : _GEN_8362; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8364 = 8'h57 == _T_509[7:0] ? 4'hf : _GEN_8363; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8365 = 8'h58 == _T_509[7:0] ? 4'h0 : _GEN_8364; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8366 = 8'h59 == _T_509[7:0] ? 4'h0 : _GEN_8365; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8367 = 8'h5a == _T_509[7:0] ? 4'h0 : _GEN_8366; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8368 = 8'h5b == _T_509[7:0] ? 4'h0 : _GEN_8367; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8369 = 8'h5c == _T_509[7:0] ? 4'h0 : _GEN_8368; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8370 = 8'h5d == _T_509[7:0] ? 4'h0 : _GEN_8369; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8371 = 8'h5e == _T_509[7:0] ? 4'h0 : _GEN_8370; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8372 = 8'h5f == _T_509[7:0] ? 4'h0 : _GEN_8371; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8373 = 8'h60 == _T_509[7:0] ? 4'h0 : _GEN_8372; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8374 = 8'h61 == _T_509[7:0] ? 4'h0 : _GEN_8373; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8375 = 8'h62 == _T_509[7:0] ? 4'h0 : _GEN_8374; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8376 = 8'h63 == _T_509[7:0] ? 4'h0 : _GEN_8375; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8377 = 8'h64 == _T_509[7:0] ? 4'h0 : _GEN_8376; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8378 = 8'h65 == _T_509[7:0] ? 4'h0 : _GEN_8377; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8379 = 8'h66 == _T_509[7:0] ? 4'h0 : _GEN_8378; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8380 = 8'h67 == _T_509[7:0] ? 4'h0 : _GEN_8379; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8381 = 8'h68 == _T_509[7:0] ? 4'hf : _GEN_8380; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8382 = 8'h69 == _T_509[7:0] ? 4'hf : _GEN_8381; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8383 = 8'h6a == _T_509[7:0] ? 4'hf : _GEN_8382; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8384 = 8'h6b == _T_509[7:0] ? 4'hf : _GEN_8383; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8385 = 8'h6c == _T_509[7:0] ? 4'hf : _GEN_8384; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8386 = 8'h6d == _T_509[7:0] ? 4'hf : _GEN_8385; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8387 = 8'h6e == _T_509[7:0] ? 4'hf : _GEN_8386; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8388 = 8'h6f == _T_509[7:0] ? 4'hf : _GEN_8387; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8389 = 8'h70 == _T_509[7:0] ? 4'h0 : _GEN_8388; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8390 = 8'h71 == _T_509[7:0] ? 4'h0 : _GEN_8389; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8391 = 8'h72 == _T_509[7:0] ? 4'h0 : _GEN_8390; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8392 = 8'h73 == _T_509[7:0] ? 4'h0 : _GEN_8391; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8393 = 8'h74 == _T_509[7:0] ? 4'h0 : _GEN_8392; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8394 = 8'h75 == _T_509[7:0] ? 4'h0 : _GEN_8393; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8395 = 8'h76 == _T_509[7:0] ? 4'h0 : _GEN_8394; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8396 = 8'h77 == _T_509[7:0] ? 4'h0 : _GEN_8395; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8397 = 8'h78 == _T_509[7:0] ? 4'hf : _GEN_8396; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8398 = 8'h79 == _T_509[7:0] ? 4'hf : _GEN_8397; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8399 = 8'h7a == _T_509[7:0] ? 4'hf : _GEN_8398; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8400 = 8'h7b == _T_509[7:0] ? 4'hf : _GEN_8399; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8401 = 8'h7c == _T_509[7:0] ? 4'hf : _GEN_8400; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8402 = 8'h7d == _T_509[7:0] ? 4'hf : _GEN_8401; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8403 = 8'h7e == _T_509[7:0] ? 4'hf : _GEN_8402; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8404 = 8'h7f == _T_509[7:0] ? 4'hf : _GEN_8403; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8405 = 8'h80 == _T_509[7:0] ? 4'h0 : _GEN_8404; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8406 = 8'h81 == _T_509[7:0] ? 4'h0 : _GEN_8405; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8407 = 8'h82 == _T_509[7:0] ? 4'h0 : _GEN_8406; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8408 = 8'h83 == _T_509[7:0] ? 4'h0 : _GEN_8407; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8409 = 8'h84 == _T_509[7:0] ? 4'h0 : _GEN_8408; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8410 = 8'h85 == _T_509[7:0] ? 4'h0 : _GEN_8409; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8411 = 8'h86 == _T_509[7:0] ? 4'h0 : _GEN_8410; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8412 = 8'h87 == _T_509[7:0] ? 4'h0 : _GEN_8411; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8413 = 8'h88 == _T_509[7:0] ? 4'hf : _GEN_8412; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8414 = 8'h89 == _T_509[7:0] ? 4'hf : _GEN_8413; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8415 = 8'h8a == _T_509[7:0] ? 4'hf : _GEN_8414; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8416 = 8'h8b == _T_509[7:0] ? 4'hf : _GEN_8415; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8417 = 8'h8c == _T_509[7:0] ? 4'hf : _GEN_8416; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8418 = 8'h8d == _T_509[7:0] ? 4'hf : _GEN_8417; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8419 = 8'h8e == _T_509[7:0] ? 4'hf : _GEN_8418; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8420 = 8'h8f == _T_509[7:0] ? 4'hf : _GEN_8419; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8421 = 8'h90 == _T_509[7:0] ? 4'h0 : _GEN_8420; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8422 = 8'h91 == _T_509[7:0] ? 4'h0 : _GEN_8421; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8423 = 8'h92 == _T_509[7:0] ? 4'h0 : _GEN_8422; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8424 = 8'h93 == _T_509[7:0] ? 4'h0 : _GEN_8423; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8425 = 8'h94 == _T_509[7:0] ? 4'h0 : _GEN_8424; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8426 = 8'h95 == _T_509[7:0] ? 4'h0 : _GEN_8425; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8427 = 8'h96 == _T_509[7:0] ? 4'h0 : _GEN_8426; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8428 = 8'h97 == _T_509[7:0] ? 4'h0 : _GEN_8427; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8429 = 8'h98 == _T_509[7:0] ? 4'hf : _GEN_8428; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8430 = 8'h99 == _T_509[7:0] ? 4'hf : _GEN_8429; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8431 = 8'h9a == _T_509[7:0] ? 4'hf : _GEN_8430; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8432 = 8'h9b == _T_509[7:0] ? 4'hf : _GEN_8431; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8433 = 8'h9c == _T_509[7:0] ? 4'hf : _GEN_8432; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8434 = 8'h9d == _T_509[7:0] ? 4'hf : _GEN_8433; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8435 = 8'h9e == _T_509[7:0] ? 4'hf : _GEN_8434; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8436 = 8'h9f == _T_509[7:0] ? 4'hf : _GEN_8435; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8437 = 8'ha0 == _T_509[7:0] ? 4'h0 : _GEN_8436; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8438 = 8'ha1 == _T_509[7:0] ? 4'h0 : _GEN_8437; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8439 = 8'ha2 == _T_509[7:0] ? 4'h0 : _GEN_8438; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8440 = 8'ha3 == _T_509[7:0] ? 4'h0 : _GEN_8439; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8441 = 8'ha4 == _T_509[7:0] ? 4'h0 : _GEN_8440; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8442 = 8'ha5 == _T_509[7:0] ? 4'h0 : _GEN_8441; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8443 = 8'ha6 == _T_509[7:0] ? 4'h0 : _GEN_8442; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8444 = 8'ha7 == _T_509[7:0] ? 4'h0 : _GEN_8443; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8445 = 8'ha8 == _T_509[7:0] ? 4'hf : _GEN_8444; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8446 = 8'ha9 == _T_509[7:0] ? 4'hf : _GEN_8445; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8447 = 8'haa == _T_509[7:0] ? 4'hf : _GEN_8446; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8448 = 8'hab == _T_509[7:0] ? 4'hf : _GEN_8447; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8449 = 8'hac == _T_509[7:0] ? 4'hf : _GEN_8448; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8450 = 8'had == _T_509[7:0] ? 4'hf : _GEN_8449; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8451 = 8'hae == _T_509[7:0] ? 4'hf : _GEN_8450; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8452 = 8'haf == _T_509[7:0] ? 4'hf : _GEN_8451; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8453 = 8'hb0 == _T_509[7:0] ? 4'h0 : _GEN_8452; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8454 = 8'hb1 == _T_509[7:0] ? 4'h0 : _GEN_8453; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8455 = 8'hb2 == _T_509[7:0] ? 4'h0 : _GEN_8454; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8456 = 8'hb3 == _T_509[7:0] ? 4'h0 : _GEN_8455; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8457 = 8'hb4 == _T_509[7:0] ? 4'h0 : _GEN_8456; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8458 = 8'hb5 == _T_509[7:0] ? 4'h0 : _GEN_8457; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8459 = 8'hb6 == _T_509[7:0] ? 4'h0 : _GEN_8458; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8460 = 8'hb7 == _T_509[7:0] ? 4'h0 : _GEN_8459; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8461 = 8'hb8 == _T_509[7:0] ? 4'hf : _GEN_8460; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8462 = 8'hb9 == _T_509[7:0] ? 4'hf : _GEN_8461; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8463 = 8'hba == _T_509[7:0] ? 4'hf : _GEN_8462; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8464 = 8'hbb == _T_509[7:0] ? 4'hf : _GEN_8463; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8465 = 8'hbc == _T_509[7:0] ? 4'hf : _GEN_8464; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8466 = 8'hbd == _T_509[7:0] ? 4'hf : _GEN_8465; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8467 = 8'hbe == _T_509[7:0] ? 4'hf : _GEN_8466; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8468 = 8'hbf == _T_509[7:0] ? 4'hf : _GEN_8467; // @[Filter.scala 160:62]
  wire [4:0] _GEN_9950 = {{1'd0}, _GEN_8468}; // @[Filter.scala 160:62]
  wire [8:0] _T_511 = _GEN_9950 * 5'h14; // @[Filter.scala 160:62]
  wire [3:0] _GEN_8565 = 8'h60 == _T_509[7:0] ? 4'hf : 4'h0; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8566 = 8'h61 == _T_509[7:0] ? 4'hf : _GEN_8565; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8567 = 8'h62 == _T_509[7:0] ? 4'hf : _GEN_8566; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8568 = 8'h63 == _T_509[7:0] ? 4'hf : _GEN_8567; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8569 = 8'h64 == _T_509[7:0] ? 4'hf : _GEN_8568; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8570 = 8'h65 == _T_509[7:0] ? 4'hf : _GEN_8569; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8571 = 8'h66 == _T_509[7:0] ? 4'hf : _GEN_8570; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8572 = 8'h67 == _T_509[7:0] ? 4'hf : _GEN_8571; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8573 = 8'h68 == _T_509[7:0] ? 4'hf : _GEN_8572; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8574 = 8'h69 == _T_509[7:0] ? 4'hf : _GEN_8573; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8575 = 8'h6a == _T_509[7:0] ? 4'hf : _GEN_8574; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8576 = 8'h6b == _T_509[7:0] ? 4'hf : _GEN_8575; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8577 = 8'h6c == _T_509[7:0] ? 4'hf : _GEN_8576; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8578 = 8'h6d == _T_509[7:0] ? 4'hf : _GEN_8577; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8579 = 8'h6e == _T_509[7:0] ? 4'hf : _GEN_8578; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8580 = 8'h6f == _T_509[7:0] ? 4'hf : _GEN_8579; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8581 = 8'h70 == _T_509[7:0] ? 4'hf : _GEN_8580; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8582 = 8'h71 == _T_509[7:0] ? 4'hf : _GEN_8581; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8583 = 8'h72 == _T_509[7:0] ? 4'hf : _GEN_8582; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8584 = 8'h73 == _T_509[7:0] ? 4'hf : _GEN_8583; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8585 = 8'h74 == _T_509[7:0] ? 4'hf : _GEN_8584; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8586 = 8'h75 == _T_509[7:0] ? 4'hf : _GEN_8585; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8587 = 8'h76 == _T_509[7:0] ? 4'hf : _GEN_8586; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8588 = 8'h77 == _T_509[7:0] ? 4'hf : _GEN_8587; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8589 = 8'h78 == _T_509[7:0] ? 4'hf : _GEN_8588; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8590 = 8'h79 == _T_509[7:0] ? 4'hf : _GEN_8589; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8591 = 8'h7a == _T_509[7:0] ? 4'hf : _GEN_8590; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8592 = 8'h7b == _T_509[7:0] ? 4'hf : _GEN_8591; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8593 = 8'h7c == _T_509[7:0] ? 4'hf : _GEN_8592; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8594 = 8'h7d == _T_509[7:0] ? 4'hf : _GEN_8593; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8595 = 8'h7e == _T_509[7:0] ? 4'hf : _GEN_8594; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8596 = 8'h7f == _T_509[7:0] ? 4'hf : _GEN_8595; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8597 = 8'h80 == _T_509[7:0] ? 4'hf : _GEN_8596; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8598 = 8'h81 == _T_509[7:0] ? 4'hf : _GEN_8597; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8599 = 8'h82 == _T_509[7:0] ? 4'hf : _GEN_8598; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8600 = 8'h83 == _T_509[7:0] ? 4'hf : _GEN_8599; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8601 = 8'h84 == _T_509[7:0] ? 4'hf : _GEN_8600; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8602 = 8'h85 == _T_509[7:0] ? 4'hf : _GEN_8601; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8603 = 8'h86 == _T_509[7:0] ? 4'hf : _GEN_8602; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8604 = 8'h87 == _T_509[7:0] ? 4'hf : _GEN_8603; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8605 = 8'h88 == _T_509[7:0] ? 4'hf : _GEN_8604; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8606 = 8'h89 == _T_509[7:0] ? 4'hf : _GEN_8605; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8607 = 8'h8a == _T_509[7:0] ? 4'hf : _GEN_8606; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8608 = 8'h8b == _T_509[7:0] ? 4'hf : _GEN_8607; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8609 = 8'h8c == _T_509[7:0] ? 4'hf : _GEN_8608; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8610 = 8'h8d == _T_509[7:0] ? 4'hf : _GEN_8609; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8611 = 8'h8e == _T_509[7:0] ? 4'hf : _GEN_8610; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8612 = 8'h8f == _T_509[7:0] ? 4'hf : _GEN_8611; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8613 = 8'h90 == _T_509[7:0] ? 4'hf : _GEN_8612; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8614 = 8'h91 == _T_509[7:0] ? 4'hf : _GEN_8613; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8615 = 8'h92 == _T_509[7:0] ? 4'hf : _GEN_8614; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8616 = 8'h93 == _T_509[7:0] ? 4'hf : _GEN_8615; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8617 = 8'h94 == _T_509[7:0] ? 4'hf : _GEN_8616; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8618 = 8'h95 == _T_509[7:0] ? 4'hf : _GEN_8617; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8619 = 8'h96 == _T_509[7:0] ? 4'hf : _GEN_8618; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8620 = 8'h97 == _T_509[7:0] ? 4'hf : _GEN_8619; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8621 = 8'h98 == _T_509[7:0] ? 4'hf : _GEN_8620; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8622 = 8'h99 == _T_509[7:0] ? 4'hf : _GEN_8621; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8623 = 8'h9a == _T_509[7:0] ? 4'hf : _GEN_8622; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8624 = 8'h9b == _T_509[7:0] ? 4'hf : _GEN_8623; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8625 = 8'h9c == _T_509[7:0] ? 4'hf : _GEN_8624; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8626 = 8'h9d == _T_509[7:0] ? 4'hf : _GEN_8625; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8627 = 8'h9e == _T_509[7:0] ? 4'hf : _GEN_8626; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8628 = 8'h9f == _T_509[7:0] ? 4'hf : _GEN_8627; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8629 = 8'ha0 == _T_509[7:0] ? 4'hf : _GEN_8628; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8630 = 8'ha1 == _T_509[7:0] ? 4'hf : _GEN_8629; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8631 = 8'ha2 == _T_509[7:0] ? 4'hf : _GEN_8630; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8632 = 8'ha3 == _T_509[7:0] ? 4'hf : _GEN_8631; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8633 = 8'ha4 == _T_509[7:0] ? 4'hf : _GEN_8632; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8634 = 8'ha5 == _T_509[7:0] ? 4'hf : _GEN_8633; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8635 = 8'ha6 == _T_509[7:0] ? 4'hf : _GEN_8634; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8636 = 8'ha7 == _T_509[7:0] ? 4'hf : _GEN_8635; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8637 = 8'ha8 == _T_509[7:0] ? 4'hf : _GEN_8636; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8638 = 8'ha9 == _T_509[7:0] ? 4'hf : _GEN_8637; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8639 = 8'haa == _T_509[7:0] ? 4'hf : _GEN_8638; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8640 = 8'hab == _T_509[7:0] ? 4'hf : _GEN_8639; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8641 = 8'hac == _T_509[7:0] ? 4'hf : _GEN_8640; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8642 = 8'had == _T_509[7:0] ? 4'hf : _GEN_8641; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8643 = 8'hae == _T_509[7:0] ? 4'hf : _GEN_8642; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8644 = 8'haf == _T_509[7:0] ? 4'hf : _GEN_8643; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8645 = 8'hb0 == _T_509[7:0] ? 4'hf : _GEN_8644; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8646 = 8'hb1 == _T_509[7:0] ? 4'hf : _GEN_8645; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8647 = 8'hb2 == _T_509[7:0] ? 4'hf : _GEN_8646; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8648 = 8'hb3 == _T_509[7:0] ? 4'hf : _GEN_8647; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8649 = 8'hb4 == _T_509[7:0] ? 4'hf : _GEN_8648; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8650 = 8'hb5 == _T_509[7:0] ? 4'hf : _GEN_8649; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8651 = 8'hb6 == _T_509[7:0] ? 4'hf : _GEN_8650; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8652 = 8'hb7 == _T_509[7:0] ? 4'hf : _GEN_8651; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8653 = 8'hb8 == _T_509[7:0] ? 4'hf : _GEN_8652; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8654 = 8'hb9 == _T_509[7:0] ? 4'hf : _GEN_8653; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8655 = 8'hba == _T_509[7:0] ? 4'hf : _GEN_8654; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8656 = 8'hbb == _T_509[7:0] ? 4'hf : _GEN_8655; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8657 = 8'hbc == _T_509[7:0] ? 4'hf : _GEN_8656; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8658 = 8'hbd == _T_509[7:0] ? 4'hf : _GEN_8657; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8659 = 8'hbe == _T_509[7:0] ? 4'hf : _GEN_8658; // @[Filter.scala 160:102]
  wire [3:0] _GEN_8660 = 8'hbf == _T_509[7:0] ? 4'hf : _GEN_8659; // @[Filter.scala 160:102]
  wire [6:0] _GEN_9952 = {{3'd0}, _GEN_8660}; // @[Filter.scala 160:102]
  wire [10:0] _T_516 = _GEN_9952 * 7'h46; // @[Filter.scala 160:102]
  wire [10:0] _GEN_9953 = {{2'd0}, _T_511}; // @[Filter.scala 160:69]
  wire [10:0] _T_518 = _GEN_9953 + _T_516; // @[Filter.scala 160:69]
  wire [3:0] _GEN_8669 = 8'h8 == _T_509[7:0] ? 4'hf : 4'h0; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8670 = 8'h9 == _T_509[7:0] ? 4'hf : _GEN_8669; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8671 = 8'ha == _T_509[7:0] ? 4'hf : _GEN_8670; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8672 = 8'hb == _T_509[7:0] ? 4'hf : _GEN_8671; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8673 = 8'hc == _T_509[7:0] ? 4'hf : _GEN_8672; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8674 = 8'hd == _T_509[7:0] ? 4'hf : _GEN_8673; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8675 = 8'he == _T_509[7:0] ? 4'hf : _GEN_8674; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8676 = 8'hf == _T_509[7:0] ? 4'hf : _GEN_8675; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8677 = 8'h10 == _T_509[7:0] ? 4'h0 : _GEN_8676; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8678 = 8'h11 == _T_509[7:0] ? 4'h0 : _GEN_8677; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8679 = 8'h12 == _T_509[7:0] ? 4'h0 : _GEN_8678; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8680 = 8'h13 == _T_509[7:0] ? 4'h0 : _GEN_8679; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8681 = 8'h14 == _T_509[7:0] ? 4'h0 : _GEN_8680; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8682 = 8'h15 == _T_509[7:0] ? 4'h0 : _GEN_8681; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8683 = 8'h16 == _T_509[7:0] ? 4'h0 : _GEN_8682; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8684 = 8'h17 == _T_509[7:0] ? 4'h0 : _GEN_8683; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8685 = 8'h18 == _T_509[7:0] ? 4'hf : _GEN_8684; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8686 = 8'h19 == _T_509[7:0] ? 4'hf : _GEN_8685; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8687 = 8'h1a == _T_509[7:0] ? 4'hf : _GEN_8686; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8688 = 8'h1b == _T_509[7:0] ? 4'hf : _GEN_8687; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8689 = 8'h1c == _T_509[7:0] ? 4'hf : _GEN_8688; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8690 = 8'h1d == _T_509[7:0] ? 4'hf : _GEN_8689; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8691 = 8'h1e == _T_509[7:0] ? 4'hf : _GEN_8690; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8692 = 8'h1f == _T_509[7:0] ? 4'hf : _GEN_8691; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8693 = 8'h20 == _T_509[7:0] ? 4'h0 : _GEN_8692; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8694 = 8'h21 == _T_509[7:0] ? 4'h0 : _GEN_8693; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8695 = 8'h22 == _T_509[7:0] ? 4'h0 : _GEN_8694; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8696 = 8'h23 == _T_509[7:0] ? 4'h0 : _GEN_8695; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8697 = 8'h24 == _T_509[7:0] ? 4'h0 : _GEN_8696; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8698 = 8'h25 == _T_509[7:0] ? 4'h0 : _GEN_8697; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8699 = 8'h26 == _T_509[7:0] ? 4'h0 : _GEN_8698; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8700 = 8'h27 == _T_509[7:0] ? 4'h0 : _GEN_8699; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8701 = 8'h28 == _T_509[7:0] ? 4'hf : _GEN_8700; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8702 = 8'h29 == _T_509[7:0] ? 4'hf : _GEN_8701; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8703 = 8'h2a == _T_509[7:0] ? 4'hf : _GEN_8702; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8704 = 8'h2b == _T_509[7:0] ? 4'hf : _GEN_8703; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8705 = 8'h2c == _T_509[7:0] ? 4'hf : _GEN_8704; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8706 = 8'h2d == _T_509[7:0] ? 4'hf : _GEN_8705; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8707 = 8'h2e == _T_509[7:0] ? 4'hf : _GEN_8706; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8708 = 8'h2f == _T_509[7:0] ? 4'hf : _GEN_8707; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8709 = 8'h30 == _T_509[7:0] ? 4'h0 : _GEN_8708; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8710 = 8'h31 == _T_509[7:0] ? 4'h0 : _GEN_8709; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8711 = 8'h32 == _T_509[7:0] ? 4'h0 : _GEN_8710; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8712 = 8'h33 == _T_509[7:0] ? 4'h0 : _GEN_8711; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8713 = 8'h34 == _T_509[7:0] ? 4'h0 : _GEN_8712; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8714 = 8'h35 == _T_509[7:0] ? 4'h0 : _GEN_8713; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8715 = 8'h36 == _T_509[7:0] ? 4'h0 : _GEN_8714; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8716 = 8'h37 == _T_509[7:0] ? 4'h0 : _GEN_8715; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8717 = 8'h38 == _T_509[7:0] ? 4'hf : _GEN_8716; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8718 = 8'h39 == _T_509[7:0] ? 4'hf : _GEN_8717; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8719 = 8'h3a == _T_509[7:0] ? 4'hf : _GEN_8718; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8720 = 8'h3b == _T_509[7:0] ? 4'hf : _GEN_8719; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8721 = 8'h3c == _T_509[7:0] ? 4'hf : _GEN_8720; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8722 = 8'h3d == _T_509[7:0] ? 4'hf : _GEN_8721; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8723 = 8'h3e == _T_509[7:0] ? 4'hf : _GEN_8722; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8724 = 8'h3f == _T_509[7:0] ? 4'hf : _GEN_8723; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8725 = 8'h40 == _T_509[7:0] ? 4'h0 : _GEN_8724; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8726 = 8'h41 == _T_509[7:0] ? 4'h0 : _GEN_8725; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8727 = 8'h42 == _T_509[7:0] ? 4'h0 : _GEN_8726; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8728 = 8'h43 == _T_509[7:0] ? 4'h0 : _GEN_8727; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8729 = 8'h44 == _T_509[7:0] ? 4'h0 : _GEN_8728; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8730 = 8'h45 == _T_509[7:0] ? 4'h0 : _GEN_8729; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8731 = 8'h46 == _T_509[7:0] ? 4'h0 : _GEN_8730; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8732 = 8'h47 == _T_509[7:0] ? 4'h0 : _GEN_8731; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8733 = 8'h48 == _T_509[7:0] ? 4'hf : _GEN_8732; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8734 = 8'h49 == _T_509[7:0] ? 4'hf : _GEN_8733; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8735 = 8'h4a == _T_509[7:0] ? 4'hf : _GEN_8734; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8736 = 8'h4b == _T_509[7:0] ? 4'hf : _GEN_8735; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8737 = 8'h4c == _T_509[7:0] ? 4'hf : _GEN_8736; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8738 = 8'h4d == _T_509[7:0] ? 4'hf : _GEN_8737; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8739 = 8'h4e == _T_509[7:0] ? 4'hf : _GEN_8738; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8740 = 8'h4f == _T_509[7:0] ? 4'hf : _GEN_8739; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8741 = 8'h50 == _T_509[7:0] ? 4'h0 : _GEN_8740; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8742 = 8'h51 == _T_509[7:0] ? 4'h0 : _GEN_8741; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8743 = 8'h52 == _T_509[7:0] ? 4'h0 : _GEN_8742; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8744 = 8'h53 == _T_509[7:0] ? 4'h0 : _GEN_8743; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8745 = 8'h54 == _T_509[7:0] ? 4'h0 : _GEN_8744; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8746 = 8'h55 == _T_509[7:0] ? 4'h0 : _GEN_8745; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8747 = 8'h56 == _T_509[7:0] ? 4'h0 : _GEN_8746; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8748 = 8'h57 == _T_509[7:0] ? 4'h0 : _GEN_8747; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8749 = 8'h58 == _T_509[7:0] ? 4'hf : _GEN_8748; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8750 = 8'h59 == _T_509[7:0] ? 4'hf : _GEN_8749; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8751 = 8'h5a == _T_509[7:0] ? 4'hf : _GEN_8750; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8752 = 8'h5b == _T_509[7:0] ? 4'hf : _GEN_8751; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8753 = 8'h5c == _T_509[7:0] ? 4'hf : _GEN_8752; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8754 = 8'h5d == _T_509[7:0] ? 4'hf : _GEN_8753; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8755 = 8'h5e == _T_509[7:0] ? 4'hf : _GEN_8754; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8756 = 8'h5f == _T_509[7:0] ? 4'hf : _GEN_8755; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8757 = 8'h60 == _T_509[7:0] ? 4'h0 : _GEN_8756; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8758 = 8'h61 == _T_509[7:0] ? 4'h0 : _GEN_8757; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8759 = 8'h62 == _T_509[7:0] ? 4'h0 : _GEN_8758; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8760 = 8'h63 == _T_509[7:0] ? 4'h0 : _GEN_8759; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8761 = 8'h64 == _T_509[7:0] ? 4'h0 : _GEN_8760; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8762 = 8'h65 == _T_509[7:0] ? 4'h0 : _GEN_8761; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8763 = 8'h66 == _T_509[7:0] ? 4'h0 : _GEN_8762; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8764 = 8'h67 == _T_509[7:0] ? 4'h0 : _GEN_8763; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8765 = 8'h68 == _T_509[7:0] ? 4'hf : _GEN_8764; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8766 = 8'h69 == _T_509[7:0] ? 4'hf : _GEN_8765; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8767 = 8'h6a == _T_509[7:0] ? 4'hf : _GEN_8766; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8768 = 8'h6b == _T_509[7:0] ? 4'hf : _GEN_8767; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8769 = 8'h6c == _T_509[7:0] ? 4'hf : _GEN_8768; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8770 = 8'h6d == _T_509[7:0] ? 4'hf : _GEN_8769; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8771 = 8'h6e == _T_509[7:0] ? 4'hf : _GEN_8770; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8772 = 8'h6f == _T_509[7:0] ? 4'hf : _GEN_8771; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8773 = 8'h70 == _T_509[7:0] ? 4'h0 : _GEN_8772; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8774 = 8'h71 == _T_509[7:0] ? 4'h0 : _GEN_8773; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8775 = 8'h72 == _T_509[7:0] ? 4'h0 : _GEN_8774; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8776 = 8'h73 == _T_509[7:0] ? 4'h0 : _GEN_8775; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8777 = 8'h74 == _T_509[7:0] ? 4'h0 : _GEN_8776; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8778 = 8'h75 == _T_509[7:0] ? 4'h0 : _GEN_8777; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8779 = 8'h76 == _T_509[7:0] ? 4'h0 : _GEN_8778; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8780 = 8'h77 == _T_509[7:0] ? 4'h0 : _GEN_8779; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8781 = 8'h78 == _T_509[7:0] ? 4'hf : _GEN_8780; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8782 = 8'h79 == _T_509[7:0] ? 4'hf : _GEN_8781; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8783 = 8'h7a == _T_509[7:0] ? 4'hf : _GEN_8782; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8784 = 8'h7b == _T_509[7:0] ? 4'hf : _GEN_8783; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8785 = 8'h7c == _T_509[7:0] ? 4'hf : _GEN_8784; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8786 = 8'h7d == _T_509[7:0] ? 4'hf : _GEN_8785; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8787 = 8'h7e == _T_509[7:0] ? 4'hf : _GEN_8786; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8788 = 8'h7f == _T_509[7:0] ? 4'hf : _GEN_8787; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8789 = 8'h80 == _T_509[7:0] ? 4'h0 : _GEN_8788; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8790 = 8'h81 == _T_509[7:0] ? 4'h0 : _GEN_8789; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8791 = 8'h82 == _T_509[7:0] ? 4'h0 : _GEN_8790; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8792 = 8'h83 == _T_509[7:0] ? 4'h0 : _GEN_8791; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8793 = 8'h84 == _T_509[7:0] ? 4'h0 : _GEN_8792; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8794 = 8'h85 == _T_509[7:0] ? 4'h0 : _GEN_8793; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8795 = 8'h86 == _T_509[7:0] ? 4'h0 : _GEN_8794; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8796 = 8'h87 == _T_509[7:0] ? 4'h0 : _GEN_8795; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8797 = 8'h88 == _T_509[7:0] ? 4'hf : _GEN_8796; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8798 = 8'h89 == _T_509[7:0] ? 4'hf : _GEN_8797; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8799 = 8'h8a == _T_509[7:0] ? 4'hf : _GEN_8798; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8800 = 8'h8b == _T_509[7:0] ? 4'hf : _GEN_8799; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8801 = 8'h8c == _T_509[7:0] ? 4'hf : _GEN_8800; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8802 = 8'h8d == _T_509[7:0] ? 4'hf : _GEN_8801; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8803 = 8'h8e == _T_509[7:0] ? 4'hf : _GEN_8802; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8804 = 8'h8f == _T_509[7:0] ? 4'hf : _GEN_8803; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8805 = 8'h90 == _T_509[7:0] ? 4'h0 : _GEN_8804; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8806 = 8'h91 == _T_509[7:0] ? 4'h0 : _GEN_8805; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8807 = 8'h92 == _T_509[7:0] ? 4'h0 : _GEN_8806; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8808 = 8'h93 == _T_509[7:0] ? 4'h0 : _GEN_8807; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8809 = 8'h94 == _T_509[7:0] ? 4'h0 : _GEN_8808; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8810 = 8'h95 == _T_509[7:0] ? 4'h0 : _GEN_8809; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8811 = 8'h96 == _T_509[7:0] ? 4'h0 : _GEN_8810; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8812 = 8'h97 == _T_509[7:0] ? 4'h0 : _GEN_8811; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8813 = 8'h98 == _T_509[7:0] ? 4'hf : _GEN_8812; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8814 = 8'h99 == _T_509[7:0] ? 4'hf : _GEN_8813; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8815 = 8'h9a == _T_509[7:0] ? 4'hf : _GEN_8814; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8816 = 8'h9b == _T_509[7:0] ? 4'hf : _GEN_8815; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8817 = 8'h9c == _T_509[7:0] ? 4'hf : _GEN_8816; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8818 = 8'h9d == _T_509[7:0] ? 4'hf : _GEN_8817; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8819 = 8'h9e == _T_509[7:0] ? 4'hf : _GEN_8818; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8820 = 8'h9f == _T_509[7:0] ? 4'hf : _GEN_8819; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8821 = 8'ha0 == _T_509[7:0] ? 4'h0 : _GEN_8820; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8822 = 8'ha1 == _T_509[7:0] ? 4'h0 : _GEN_8821; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8823 = 8'ha2 == _T_509[7:0] ? 4'h0 : _GEN_8822; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8824 = 8'ha3 == _T_509[7:0] ? 4'h0 : _GEN_8823; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8825 = 8'ha4 == _T_509[7:0] ? 4'h0 : _GEN_8824; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8826 = 8'ha5 == _T_509[7:0] ? 4'h0 : _GEN_8825; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8827 = 8'ha6 == _T_509[7:0] ? 4'h0 : _GEN_8826; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8828 = 8'ha7 == _T_509[7:0] ? 4'h0 : _GEN_8827; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8829 = 8'ha8 == _T_509[7:0] ? 4'hf : _GEN_8828; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8830 = 8'ha9 == _T_509[7:0] ? 4'hf : _GEN_8829; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8831 = 8'haa == _T_509[7:0] ? 4'hf : _GEN_8830; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8832 = 8'hab == _T_509[7:0] ? 4'hf : _GEN_8831; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8833 = 8'hac == _T_509[7:0] ? 4'hf : _GEN_8832; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8834 = 8'had == _T_509[7:0] ? 4'hf : _GEN_8833; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8835 = 8'hae == _T_509[7:0] ? 4'hf : _GEN_8834; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8836 = 8'haf == _T_509[7:0] ? 4'hf : _GEN_8835; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8837 = 8'hb0 == _T_509[7:0] ? 4'h0 : _GEN_8836; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8838 = 8'hb1 == _T_509[7:0] ? 4'h0 : _GEN_8837; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8839 = 8'hb2 == _T_509[7:0] ? 4'h0 : _GEN_8838; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8840 = 8'hb3 == _T_509[7:0] ? 4'h0 : _GEN_8839; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8841 = 8'hb4 == _T_509[7:0] ? 4'h0 : _GEN_8840; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8842 = 8'hb5 == _T_509[7:0] ? 4'h0 : _GEN_8841; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8843 = 8'hb6 == _T_509[7:0] ? 4'h0 : _GEN_8842; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8844 = 8'hb7 == _T_509[7:0] ? 4'h0 : _GEN_8843; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8845 = 8'hb8 == _T_509[7:0] ? 4'hf : _GEN_8844; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8846 = 8'hb9 == _T_509[7:0] ? 4'hf : _GEN_8845; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8847 = 8'hba == _T_509[7:0] ? 4'hf : _GEN_8846; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8848 = 8'hbb == _T_509[7:0] ? 4'hf : _GEN_8847; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8849 = 8'hbc == _T_509[7:0] ? 4'hf : _GEN_8848; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8850 = 8'hbd == _T_509[7:0] ? 4'hf : _GEN_8849; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8851 = 8'hbe == _T_509[7:0] ? 4'hf : _GEN_8850; // @[Filter.scala 160:142]
  wire [3:0] _GEN_8852 = 8'hbf == _T_509[7:0] ? 4'hf : _GEN_8851; // @[Filter.scala 160:142]
  wire [7:0] _T_523 = _GEN_8852 * 4'ha; // @[Filter.scala 160:142]
  wire [10:0] _GEN_9955 = {{3'd0}, _T_523}; // @[Filter.scala 160:109]
  wire [10:0] _T_525 = _T_518 + _GEN_9955; // @[Filter.scala 160:109]
  wire [10:0] _T_526 = _T_525 / 11'h64; // @[Filter.scala 160:150]
  wire  _T_528 = _T_499 >= 5'h10; // @[Filter.scala 163:31]
  wire  _T_532 = _T_506 >= 32'hc; // @[Filter.scala 163:63]
  wire  _T_533 = _T_528 | _T_532; // @[Filter.scala 163:58]
  wire [10:0] _GEN_9045 = io_SPI_distort ? _T_526 : {{7'd0}, _GEN_8468}; // @[Filter.scala 165:35]
  wire [10:0] _GEN_9046 = _T_533 ? 11'h0 : _GEN_9045; // @[Filter.scala 163:80]
  wire [10:0] _GEN_9239 = io_SPI_distort ? _T_526 : {{7'd0}, _GEN_8660}; // @[Filter.scala 165:35]
  wire [10:0] _GEN_9240 = _T_533 ? 11'h0 : _GEN_9239; // @[Filter.scala 163:80]
  wire [10:0] _GEN_9433 = io_SPI_distort ? _T_526 : {{7'd0}, _GEN_8852}; // @[Filter.scala 165:35]
  wire [10:0] _GEN_9434 = _T_533 ? 11'h0 : _GEN_9433; // @[Filter.scala 163:80]
  wire [7:0] _GEN_9436 = 3'h1 == io_SPI_filterIndex[2:0] ? $signed(8'sh9) : $signed(8'sh1); // @[Filter.scala 177:61]
  wire [7:0] _GEN_9437 = 3'h2 == io_SPI_filterIndex[2:0] ? $signed(8'sh10) : $signed(_GEN_9436); // @[Filter.scala 177:61]
  wire [7:0] _GEN_9438 = 3'h3 == io_SPI_filterIndex[2:0] ? $signed(8'sh1) : $signed(_GEN_9437); // @[Filter.scala 177:61]
  wire [7:0] _GEN_9439 = 3'h4 == io_SPI_filterIndex[2:0] ? $signed(8'sh1) : $signed(_GEN_9438); // @[Filter.scala 177:61]
  wire [7:0] _GEN_9440 = 3'h5 == io_SPI_filterIndex[2:0] ? $signed(8'sh1) : $signed(_GEN_9439); // @[Filter.scala 177:61]
  wire [8:0] _GEN_9959 = {{1{_GEN_9440[7]}},_GEN_9440}; // @[Filter.scala 177:61]
  wire [9:0] _T_561 = $signed(KernelConvolution_io_pixelVal_out_0) / $signed(_GEN_9959); // @[Filter.scala 177:61]
  wire  _T_562 = $signed(_T_561) < 10'sh0; // @[Filter.scala 179:24]
  wire  _T_565 = $signed(_T_561) > 10'shf; // @[Filter.scala 184:30]
  wire [9:0] _T_568 = $signed(KernelConvolution_io_pixelVal_out_0) / $signed(_GEN_9959); // @[Filter.scala 189:52]
  wire [9:0] _GEN_9442 = _T_565 ? 10'hf : _T_568; // @[Filter.scala 186:38]
  wire [9:0] _GEN_9444 = _T_562 ? 10'h0 : _GEN_9442; // @[Filter.scala 181:37]
  wire [9:0] _T_572 = $signed(KernelConvolution_io_pixelVal_out_1) / $signed(_GEN_9959); // @[Filter.scala 177:61]
  wire  _T_573 = $signed(_T_572) < 10'sh0; // @[Filter.scala 179:24]
  wire  _T_576 = $signed(_T_572) > 10'shf; // @[Filter.scala 184:30]
  wire [9:0] _T_579 = $signed(KernelConvolution_io_pixelVal_out_1) / $signed(_GEN_9959); // @[Filter.scala 189:52]
  wire [9:0] _GEN_9447 = _T_576 ? 10'hf : _T_579; // @[Filter.scala 186:38]
  wire [9:0] _GEN_9449 = _T_573 ? 10'h0 : _GEN_9447; // @[Filter.scala 181:37]
  wire [9:0] _T_583 = $signed(KernelConvolution_io_pixelVal_out_2) / $signed(_GEN_9959); // @[Filter.scala 177:61]
  wire  _T_584 = $signed(_T_583) < 10'sh0; // @[Filter.scala 179:24]
  wire  _T_587 = $signed(_T_583) > 10'shf; // @[Filter.scala 184:30]
  wire [9:0] _T_590 = $signed(KernelConvolution_io_pixelVal_out_2) / $signed(_GEN_9959); // @[Filter.scala 189:52]
  wire [9:0] _GEN_9452 = _T_587 ? 10'hf : _T_590; // @[Filter.scala 186:38]
  wire [9:0] _GEN_9454 = _T_584 ? 10'h0 : _GEN_9452; // @[Filter.scala 181:37]
  wire [9:0] _T_594 = $signed(KernelConvolution_io_pixelVal_out_3) / $signed(_GEN_9959); // @[Filter.scala 177:61]
  wire  _T_595 = $signed(_T_594) < 10'sh0; // @[Filter.scala 179:24]
  wire  _T_598 = $signed(_T_594) > 10'shf; // @[Filter.scala 184:30]
  wire [9:0] _T_601 = $signed(KernelConvolution_io_pixelVal_out_3) / $signed(_GEN_9959); // @[Filter.scala 189:52]
  wire [9:0] _GEN_9457 = _T_598 ? 10'hf : _T_601; // @[Filter.scala 186:38]
  wire [9:0] _GEN_9459 = _T_595 ? 10'h0 : _GEN_9457; // @[Filter.scala 181:37]
  wire [9:0] _T_605 = $signed(KernelConvolution_io_pixelVal_out_4) / $signed(_GEN_9959); // @[Filter.scala 177:61]
  wire  _T_606 = $signed(_T_605) < 10'sh0; // @[Filter.scala 179:24]
  wire  _T_609 = $signed(_T_605) > 10'shf; // @[Filter.scala 184:30]
  wire [9:0] _T_612 = $signed(KernelConvolution_io_pixelVal_out_4) / $signed(_GEN_9959); // @[Filter.scala 189:52]
  wire [9:0] _GEN_9462 = _T_609 ? 10'hf : _T_612; // @[Filter.scala 186:38]
  wire [9:0] _GEN_9464 = _T_606 ? 10'h0 : _GEN_9462; // @[Filter.scala 181:37]
  wire [9:0] _T_616 = $signed(KernelConvolution_io_pixelVal_out_5) / $signed(_GEN_9959); // @[Filter.scala 177:61]
  wire  _T_617 = $signed(_T_616) < 10'sh0; // @[Filter.scala 179:24]
  wire  _T_620 = $signed(_T_616) > 10'shf; // @[Filter.scala 184:30]
  wire [9:0] _T_623 = $signed(KernelConvolution_io_pixelVal_out_5) / $signed(_GEN_9959); // @[Filter.scala 189:52]
  wire [9:0] _GEN_9467 = _T_620 ? 10'hf : _T_623; // @[Filter.scala 186:38]
  wire [9:0] _GEN_9469 = _T_617 ? 10'h0 : _GEN_9467; // @[Filter.scala 181:37]
  wire [9:0] _T_627 = $signed(KernelConvolution_io_pixelVal_out_6) / $signed(_GEN_9959); // @[Filter.scala 177:61]
  wire  _T_628 = $signed(_T_627) < 10'sh0; // @[Filter.scala 179:24]
  wire  _T_631 = $signed(_T_627) > 10'shf; // @[Filter.scala 184:30]
  wire [9:0] _T_634 = $signed(KernelConvolution_io_pixelVal_out_6) / $signed(_GEN_9959); // @[Filter.scala 189:52]
  wire [9:0] _GEN_9472 = _T_631 ? 10'hf : _T_634; // @[Filter.scala 186:38]
  wire [9:0] _GEN_9474 = _T_628 ? 10'h0 : _GEN_9472; // @[Filter.scala 181:37]
  wire [9:0] _T_638 = $signed(KernelConvolution_io_pixelVal_out_7) / $signed(_GEN_9959); // @[Filter.scala 177:61]
  wire  _T_639 = $signed(_T_638) < 10'sh0; // @[Filter.scala 179:24]
  wire  _T_642 = $signed(_T_638) > 10'shf; // @[Filter.scala 184:30]
  wire [9:0] _T_645 = $signed(KernelConvolution_io_pixelVal_out_7) / $signed(_GEN_9959); // @[Filter.scala 189:52]
  wire [9:0] _GEN_9477 = _T_642 ? 10'hf : _T_645; // @[Filter.scala 186:38]
  wire [9:0] _GEN_9479 = _T_639 ? 10'h0 : _GEN_9477; // @[Filter.scala 181:37]
  wire [9:0] _T_649 = $signed(KernelConvolution_1_io_pixelVal_out_0) / $signed(_GEN_9959); // @[Filter.scala 177:61]
  wire  _T_650 = $signed(_T_649) < 10'sh0; // @[Filter.scala 179:24]
  wire  _T_653 = $signed(_T_649) > 10'shf; // @[Filter.scala 184:30]
  wire [9:0] _T_656 = $signed(KernelConvolution_1_io_pixelVal_out_0) / $signed(_GEN_9959); // @[Filter.scala 189:52]
  wire [9:0] _GEN_9482 = _T_653 ? 10'hf : _T_656; // @[Filter.scala 186:38]
  wire [9:0] _GEN_9484 = _T_650 ? 10'h0 : _GEN_9482; // @[Filter.scala 181:37]
  wire [9:0] _T_660 = $signed(KernelConvolution_1_io_pixelVal_out_1) / $signed(_GEN_9959); // @[Filter.scala 177:61]
  wire  _T_661 = $signed(_T_660) < 10'sh0; // @[Filter.scala 179:24]
  wire  _T_664 = $signed(_T_660) > 10'shf; // @[Filter.scala 184:30]
  wire [9:0] _T_667 = $signed(KernelConvolution_1_io_pixelVal_out_1) / $signed(_GEN_9959); // @[Filter.scala 189:52]
  wire [9:0] _GEN_9487 = _T_664 ? 10'hf : _T_667; // @[Filter.scala 186:38]
  wire [9:0] _GEN_9489 = _T_661 ? 10'h0 : _GEN_9487; // @[Filter.scala 181:37]
  wire [9:0] _T_671 = $signed(KernelConvolution_1_io_pixelVal_out_2) / $signed(_GEN_9959); // @[Filter.scala 177:61]
  wire  _T_672 = $signed(_T_671) < 10'sh0; // @[Filter.scala 179:24]
  wire  _T_675 = $signed(_T_671) > 10'shf; // @[Filter.scala 184:30]
  wire [9:0] _T_678 = $signed(KernelConvolution_1_io_pixelVal_out_2) / $signed(_GEN_9959); // @[Filter.scala 189:52]
  wire [9:0] _GEN_9492 = _T_675 ? 10'hf : _T_678; // @[Filter.scala 186:38]
  wire [9:0] _GEN_9494 = _T_672 ? 10'h0 : _GEN_9492; // @[Filter.scala 181:37]
  wire [9:0] _T_682 = $signed(KernelConvolution_1_io_pixelVal_out_3) / $signed(_GEN_9959); // @[Filter.scala 177:61]
  wire  _T_683 = $signed(_T_682) < 10'sh0; // @[Filter.scala 179:24]
  wire  _T_686 = $signed(_T_682) > 10'shf; // @[Filter.scala 184:30]
  wire [9:0] _T_689 = $signed(KernelConvolution_1_io_pixelVal_out_3) / $signed(_GEN_9959); // @[Filter.scala 189:52]
  wire [9:0] _GEN_9497 = _T_686 ? 10'hf : _T_689; // @[Filter.scala 186:38]
  wire [9:0] _GEN_9499 = _T_683 ? 10'h0 : _GEN_9497; // @[Filter.scala 181:37]
  wire [9:0] _T_693 = $signed(KernelConvolution_1_io_pixelVal_out_4) / $signed(_GEN_9959); // @[Filter.scala 177:61]
  wire  _T_694 = $signed(_T_693) < 10'sh0; // @[Filter.scala 179:24]
  wire  _T_697 = $signed(_T_693) > 10'shf; // @[Filter.scala 184:30]
  wire [9:0] _T_700 = $signed(KernelConvolution_1_io_pixelVal_out_4) / $signed(_GEN_9959); // @[Filter.scala 189:52]
  wire [9:0] _GEN_9502 = _T_697 ? 10'hf : _T_700; // @[Filter.scala 186:38]
  wire [9:0] _GEN_9504 = _T_694 ? 10'h0 : _GEN_9502; // @[Filter.scala 181:37]
  wire [9:0] _T_704 = $signed(KernelConvolution_1_io_pixelVal_out_5) / $signed(_GEN_9959); // @[Filter.scala 177:61]
  wire  _T_705 = $signed(_T_704) < 10'sh0; // @[Filter.scala 179:24]
  wire  _T_708 = $signed(_T_704) > 10'shf; // @[Filter.scala 184:30]
  wire [9:0] _T_711 = $signed(KernelConvolution_1_io_pixelVal_out_5) / $signed(_GEN_9959); // @[Filter.scala 189:52]
  wire [9:0] _GEN_9507 = _T_708 ? 10'hf : _T_711; // @[Filter.scala 186:38]
  wire [9:0] _GEN_9509 = _T_705 ? 10'h0 : _GEN_9507; // @[Filter.scala 181:37]
  wire [9:0] _T_715 = $signed(KernelConvolution_1_io_pixelVal_out_6) / $signed(_GEN_9959); // @[Filter.scala 177:61]
  wire  _T_716 = $signed(_T_715) < 10'sh0; // @[Filter.scala 179:24]
  wire  _T_719 = $signed(_T_715) > 10'shf; // @[Filter.scala 184:30]
  wire [9:0] _T_722 = $signed(KernelConvolution_1_io_pixelVal_out_6) / $signed(_GEN_9959); // @[Filter.scala 189:52]
  wire [9:0] _GEN_9512 = _T_719 ? 10'hf : _T_722; // @[Filter.scala 186:38]
  wire [9:0] _GEN_9514 = _T_716 ? 10'h0 : _GEN_9512; // @[Filter.scala 181:37]
  wire [9:0] _T_726 = $signed(KernelConvolution_1_io_pixelVal_out_7) / $signed(_GEN_9959); // @[Filter.scala 177:61]
  wire  _T_727 = $signed(_T_726) < 10'sh0; // @[Filter.scala 179:24]
  wire  _T_730 = $signed(_T_726) > 10'shf; // @[Filter.scala 184:30]
  wire [9:0] _T_733 = $signed(KernelConvolution_1_io_pixelVal_out_7) / $signed(_GEN_9959); // @[Filter.scala 189:52]
  wire [9:0] _GEN_9517 = _T_730 ? 10'hf : _T_733; // @[Filter.scala 186:38]
  wire [9:0] _GEN_9519 = _T_727 ? 10'h0 : _GEN_9517; // @[Filter.scala 181:37]
  wire [9:0] _T_737 = $signed(KernelConvolution_2_io_pixelVal_out_0) / $signed(_GEN_9959); // @[Filter.scala 177:61]
  wire  _T_738 = $signed(_T_737) < 10'sh0; // @[Filter.scala 179:24]
  wire  _T_741 = $signed(_T_737) > 10'shf; // @[Filter.scala 184:30]
  wire [9:0] _T_744 = $signed(KernelConvolution_2_io_pixelVal_out_0) / $signed(_GEN_9959); // @[Filter.scala 189:52]
  wire [9:0] _GEN_9522 = _T_741 ? 10'hf : _T_744; // @[Filter.scala 186:38]
  wire [9:0] _GEN_9524 = _T_738 ? 10'h0 : _GEN_9522; // @[Filter.scala 181:37]
  wire [9:0] _T_748 = $signed(KernelConvolution_2_io_pixelVal_out_1) / $signed(_GEN_9959); // @[Filter.scala 177:61]
  wire  _T_749 = $signed(_T_748) < 10'sh0; // @[Filter.scala 179:24]
  wire  _T_752 = $signed(_T_748) > 10'shf; // @[Filter.scala 184:30]
  wire [9:0] _T_755 = $signed(KernelConvolution_2_io_pixelVal_out_1) / $signed(_GEN_9959); // @[Filter.scala 189:52]
  wire [9:0] _GEN_9527 = _T_752 ? 10'hf : _T_755; // @[Filter.scala 186:38]
  wire [9:0] _GEN_9529 = _T_749 ? 10'h0 : _GEN_9527; // @[Filter.scala 181:37]
  wire [9:0] _T_759 = $signed(KernelConvolution_2_io_pixelVal_out_2) / $signed(_GEN_9959); // @[Filter.scala 177:61]
  wire  _T_760 = $signed(_T_759) < 10'sh0; // @[Filter.scala 179:24]
  wire  _T_763 = $signed(_T_759) > 10'shf; // @[Filter.scala 184:30]
  wire [9:0] _T_766 = $signed(KernelConvolution_2_io_pixelVal_out_2) / $signed(_GEN_9959); // @[Filter.scala 189:52]
  wire [9:0] _GEN_9532 = _T_763 ? 10'hf : _T_766; // @[Filter.scala 186:38]
  wire [9:0] _GEN_9534 = _T_760 ? 10'h0 : _GEN_9532; // @[Filter.scala 181:37]
  wire [9:0] _T_770 = $signed(KernelConvolution_2_io_pixelVal_out_3) / $signed(_GEN_9959); // @[Filter.scala 177:61]
  wire  _T_771 = $signed(_T_770) < 10'sh0; // @[Filter.scala 179:24]
  wire  _T_774 = $signed(_T_770) > 10'shf; // @[Filter.scala 184:30]
  wire [9:0] _T_777 = $signed(KernelConvolution_2_io_pixelVal_out_3) / $signed(_GEN_9959); // @[Filter.scala 189:52]
  wire [9:0] _GEN_9537 = _T_774 ? 10'hf : _T_777; // @[Filter.scala 186:38]
  wire [9:0] _GEN_9539 = _T_771 ? 10'h0 : _GEN_9537; // @[Filter.scala 181:37]
  wire [9:0] _T_781 = $signed(KernelConvolution_2_io_pixelVal_out_4) / $signed(_GEN_9959); // @[Filter.scala 177:61]
  wire  _T_782 = $signed(_T_781) < 10'sh0; // @[Filter.scala 179:24]
  wire  _T_785 = $signed(_T_781) > 10'shf; // @[Filter.scala 184:30]
  wire [9:0] _T_788 = $signed(KernelConvolution_2_io_pixelVal_out_4) / $signed(_GEN_9959); // @[Filter.scala 189:52]
  wire [9:0] _GEN_9542 = _T_785 ? 10'hf : _T_788; // @[Filter.scala 186:38]
  wire [9:0] _GEN_9544 = _T_782 ? 10'h0 : _GEN_9542; // @[Filter.scala 181:37]
  wire [9:0] _T_792 = $signed(KernelConvolution_2_io_pixelVal_out_5) / $signed(_GEN_9959); // @[Filter.scala 177:61]
  wire  _T_793 = $signed(_T_792) < 10'sh0; // @[Filter.scala 179:24]
  wire  _T_796 = $signed(_T_792) > 10'shf; // @[Filter.scala 184:30]
  wire [9:0] _T_799 = $signed(KernelConvolution_2_io_pixelVal_out_5) / $signed(_GEN_9959); // @[Filter.scala 189:52]
  wire [9:0] _GEN_9547 = _T_796 ? 10'hf : _T_799; // @[Filter.scala 186:38]
  wire [9:0] _GEN_9549 = _T_793 ? 10'h0 : _GEN_9547; // @[Filter.scala 181:37]
  wire [9:0] _T_803 = $signed(KernelConvolution_2_io_pixelVal_out_6) / $signed(_GEN_9959); // @[Filter.scala 177:61]
  wire  _T_804 = $signed(_T_803) < 10'sh0; // @[Filter.scala 179:24]
  wire  _T_807 = $signed(_T_803) > 10'shf; // @[Filter.scala 184:30]
  wire [9:0] _T_810 = $signed(KernelConvolution_2_io_pixelVal_out_6) / $signed(_GEN_9959); // @[Filter.scala 189:52]
  wire [9:0] _GEN_9552 = _T_807 ? 10'hf : _T_810; // @[Filter.scala 186:38]
  wire [9:0] _GEN_9554 = _T_804 ? 10'h0 : _GEN_9552; // @[Filter.scala 181:37]
  wire [9:0] _T_814 = $signed(KernelConvolution_2_io_pixelVal_out_7) / $signed(_GEN_9959); // @[Filter.scala 177:61]
  wire  _T_815 = $signed(_T_814) < 10'sh0; // @[Filter.scala 179:24]
  wire  _T_818 = $signed(_T_814) > 10'shf; // @[Filter.scala 184:30]
  wire [9:0] _T_821 = $signed(KernelConvolution_2_io_pixelVal_out_7) / $signed(_GEN_9959); // @[Filter.scala 189:52]
  wire [9:0] _GEN_9557 = _T_818 ? 10'hf : _T_821; // @[Filter.scala 186:38]
  wire [9:0] _GEN_9559 = _T_815 ? 10'h0 : _GEN_9557; // @[Filter.scala 181:37]
  wire [31:0] _T_826 = pixelIndex + 32'h8; // @[Filter.scala 199:34]
  wire [8:0] _T_827 = 5'h10 * 5'hc; // @[Filter.scala 200:42]
  wire [31:0] _GEN_9983 = {{23'd0}, _T_827}; // @[Filter.scala 200:25]
  wire  _T_828 = pixelIndex == _GEN_9983; // @[Filter.scala 200:25]
  KernelConvolution KernelConvolution ( // @[Filter.scala 142:36]
    .clock(KernelConvolution_clock),
    .reset(KernelConvolution_reset),
    .io_kernelVal_in(KernelConvolution_io_kernelVal_in),
    .io_pixelVal_in_0(KernelConvolution_io_pixelVal_in_0),
    .io_pixelVal_in_1(KernelConvolution_io_pixelVal_in_1),
    .io_pixelVal_in_2(KernelConvolution_io_pixelVal_in_2),
    .io_pixelVal_in_3(KernelConvolution_io_pixelVal_in_3),
    .io_pixelVal_in_4(KernelConvolution_io_pixelVal_in_4),
    .io_pixelVal_in_5(KernelConvolution_io_pixelVal_in_5),
    .io_pixelVal_in_6(KernelConvolution_io_pixelVal_in_6),
    .io_pixelVal_in_7(KernelConvolution_io_pixelVal_in_7),
    .io_pixelVal_out_0(KernelConvolution_io_pixelVal_out_0),
    .io_pixelVal_out_1(KernelConvolution_io_pixelVal_out_1),
    .io_pixelVal_out_2(KernelConvolution_io_pixelVal_out_2),
    .io_pixelVal_out_3(KernelConvolution_io_pixelVal_out_3),
    .io_pixelVal_out_4(KernelConvolution_io_pixelVal_out_4),
    .io_pixelVal_out_5(KernelConvolution_io_pixelVal_out_5),
    .io_pixelVal_out_6(KernelConvolution_io_pixelVal_out_6),
    .io_pixelVal_out_7(KernelConvolution_io_pixelVal_out_7),
    .io_valid_out(KernelConvolution_io_valid_out)
  );
  KernelConvolution KernelConvolution_1 ( // @[Filter.scala 143:36]
    .clock(KernelConvolution_1_clock),
    .reset(KernelConvolution_1_reset),
    .io_kernelVal_in(KernelConvolution_1_io_kernelVal_in),
    .io_pixelVal_in_0(KernelConvolution_1_io_pixelVal_in_0),
    .io_pixelVal_in_1(KernelConvolution_1_io_pixelVal_in_1),
    .io_pixelVal_in_2(KernelConvolution_1_io_pixelVal_in_2),
    .io_pixelVal_in_3(KernelConvolution_1_io_pixelVal_in_3),
    .io_pixelVal_in_4(KernelConvolution_1_io_pixelVal_in_4),
    .io_pixelVal_in_5(KernelConvolution_1_io_pixelVal_in_5),
    .io_pixelVal_in_6(KernelConvolution_1_io_pixelVal_in_6),
    .io_pixelVal_in_7(KernelConvolution_1_io_pixelVal_in_7),
    .io_pixelVal_out_0(KernelConvolution_1_io_pixelVal_out_0),
    .io_pixelVal_out_1(KernelConvolution_1_io_pixelVal_out_1),
    .io_pixelVal_out_2(KernelConvolution_1_io_pixelVal_out_2),
    .io_pixelVal_out_3(KernelConvolution_1_io_pixelVal_out_3),
    .io_pixelVal_out_4(KernelConvolution_1_io_pixelVal_out_4),
    .io_pixelVal_out_5(KernelConvolution_1_io_pixelVal_out_5),
    .io_pixelVal_out_6(KernelConvolution_1_io_pixelVal_out_6),
    .io_pixelVal_out_7(KernelConvolution_1_io_pixelVal_out_7),
    .io_valid_out(KernelConvolution_1_io_valid_out)
  );
  KernelConvolution KernelConvolution_2 ( // @[Filter.scala 144:36]
    .clock(KernelConvolution_2_clock),
    .reset(KernelConvolution_2_reset),
    .io_kernelVal_in(KernelConvolution_2_io_kernelVal_in),
    .io_pixelVal_in_0(KernelConvolution_2_io_pixelVal_in_0),
    .io_pixelVal_in_1(KernelConvolution_2_io_pixelVal_in_1),
    .io_pixelVal_in_2(KernelConvolution_2_io_pixelVal_in_2),
    .io_pixelVal_in_3(KernelConvolution_2_io_pixelVal_in_3),
    .io_pixelVal_in_4(KernelConvolution_2_io_pixelVal_in_4),
    .io_pixelVal_in_5(KernelConvolution_2_io_pixelVal_in_5),
    .io_pixelVal_in_6(KernelConvolution_2_io_pixelVal_in_6),
    .io_pixelVal_in_7(KernelConvolution_2_io_pixelVal_in_7),
    .io_pixelVal_out_0(KernelConvolution_2_io_pixelVal_out_0),
    .io_pixelVal_out_1(KernelConvolution_2_io_pixelVal_out_1),
    .io_pixelVal_out_2(KernelConvolution_2_io_pixelVal_out_2),
    .io_pixelVal_out_3(KernelConvolution_2_io_pixelVal_out_3),
    .io_pixelVal_out_4(KernelConvolution_2_io_pixelVal_out_4),
    .io_pixelVal_out_5(KernelConvolution_2_io_pixelVal_out_5),
    .io_pixelVal_out_6(KernelConvolution_2_io_pixelVal_out_6),
    .io_pixelVal_out_7(KernelConvolution_2_io_pixelVal_out_7),
    .io_valid_out(KernelConvolution_2_io_valid_out)
  );
  assign io_pixelVal_out_0_0 = _GEN_9444[3:0]; // @[Filter.scala 180:35 Filter.scala 182:37 Filter.scala 185:35 Filter.scala 187:35 Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_0_1 = _GEN_9449[3:0]; // @[Filter.scala 180:35 Filter.scala 182:37 Filter.scala 185:35 Filter.scala 187:35 Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_0_2 = _GEN_9454[3:0]; // @[Filter.scala 180:35 Filter.scala 182:37 Filter.scala 185:35 Filter.scala 187:35 Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_0_3 = _GEN_9459[3:0]; // @[Filter.scala 180:35 Filter.scala 182:37 Filter.scala 185:35 Filter.scala 187:35 Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_0_4 = _GEN_9464[3:0]; // @[Filter.scala 180:35 Filter.scala 182:37 Filter.scala 185:35 Filter.scala 187:35 Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_0_5 = _GEN_9469[3:0]; // @[Filter.scala 180:35 Filter.scala 182:37 Filter.scala 185:35 Filter.scala 187:35 Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_0_6 = _GEN_9474[3:0]; // @[Filter.scala 180:35 Filter.scala 182:37 Filter.scala 185:35 Filter.scala 187:35 Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_0_7 = _GEN_9479[3:0]; // @[Filter.scala 180:35 Filter.scala 182:37 Filter.scala 185:35 Filter.scala 187:35 Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_1_0 = _GEN_9484[3:0]; // @[Filter.scala 180:35 Filter.scala 182:37 Filter.scala 185:35 Filter.scala 187:35 Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_1_1 = _GEN_9489[3:0]; // @[Filter.scala 180:35 Filter.scala 182:37 Filter.scala 185:35 Filter.scala 187:35 Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_1_2 = _GEN_9494[3:0]; // @[Filter.scala 180:35 Filter.scala 182:37 Filter.scala 185:35 Filter.scala 187:35 Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_1_3 = _GEN_9499[3:0]; // @[Filter.scala 180:35 Filter.scala 182:37 Filter.scala 185:35 Filter.scala 187:35 Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_1_4 = _GEN_9504[3:0]; // @[Filter.scala 180:35 Filter.scala 182:37 Filter.scala 185:35 Filter.scala 187:35 Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_1_5 = _GEN_9509[3:0]; // @[Filter.scala 180:35 Filter.scala 182:37 Filter.scala 185:35 Filter.scala 187:35 Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_1_6 = _GEN_9514[3:0]; // @[Filter.scala 180:35 Filter.scala 182:37 Filter.scala 185:35 Filter.scala 187:35 Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_1_7 = _GEN_9519[3:0]; // @[Filter.scala 180:35 Filter.scala 182:37 Filter.scala 185:35 Filter.scala 187:35 Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_2_0 = _GEN_9524[3:0]; // @[Filter.scala 180:35 Filter.scala 182:37 Filter.scala 185:35 Filter.scala 187:35 Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_2_1 = _GEN_9529[3:0]; // @[Filter.scala 180:35 Filter.scala 182:37 Filter.scala 185:35 Filter.scala 187:35 Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_2_2 = _GEN_9534[3:0]; // @[Filter.scala 180:35 Filter.scala 182:37 Filter.scala 185:35 Filter.scala 187:35 Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_2_3 = _GEN_9539[3:0]; // @[Filter.scala 180:35 Filter.scala 182:37 Filter.scala 185:35 Filter.scala 187:35 Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_2_4 = _GEN_9544[3:0]; // @[Filter.scala 180:35 Filter.scala 182:37 Filter.scala 185:35 Filter.scala 187:35 Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_2_5 = _GEN_9549[3:0]; // @[Filter.scala 180:35 Filter.scala 182:37 Filter.scala 185:35 Filter.scala 187:35 Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_2_6 = _GEN_9554[3:0]; // @[Filter.scala 180:35 Filter.scala 182:37 Filter.scala 185:35 Filter.scala 187:35 Filter.scala 189:35 Filter.scala 191:35]
  assign io_pixelVal_out_2_7 = _GEN_9559[3:0]; // @[Filter.scala 180:35 Filter.scala 182:37 Filter.scala 185:35 Filter.scala 187:35 Filter.scala 189:35 Filter.scala 191:35]
  assign io_valid_out = KernelConvolution_io_valid_out; // @[Filter.scala 196:18]
  assign KernelConvolution_clock = clock;
  assign KernelConvolution_reset = reset;
  assign KernelConvolution_io_kernelVal_in = _GEN_9645 & _GEN_9572 ? $signed(5'sh0) : $signed(_GEN_55); // @[Filter.scala 150:41]
  assign KernelConvolution_io_pixelVal_in_0 = _GEN_940[3:0]; // @[Filter.scala 164:53 Filter.scala 166:51 Filter.scala 168:51]
  assign KernelConvolution_io_pixelVal_in_1 = _GEN_2098[3:0]; // @[Filter.scala 164:53 Filter.scala 166:51 Filter.scala 168:51]
  assign KernelConvolution_io_pixelVal_in_2 = _GEN_3256[3:0]; // @[Filter.scala 164:53 Filter.scala 166:51 Filter.scala 168:51]
  assign KernelConvolution_io_pixelVal_in_3 = _GEN_4414[3:0]; // @[Filter.scala 164:53 Filter.scala 166:51 Filter.scala 168:51]
  assign KernelConvolution_io_pixelVal_in_4 = _GEN_5572[3:0]; // @[Filter.scala 164:53 Filter.scala 166:51 Filter.scala 168:51]
  assign KernelConvolution_io_pixelVal_in_5 = _GEN_6730[3:0]; // @[Filter.scala 164:53 Filter.scala 166:51 Filter.scala 168:51]
  assign KernelConvolution_io_pixelVal_in_6 = _GEN_7888[3:0]; // @[Filter.scala 164:53 Filter.scala 166:51 Filter.scala 168:51]
  assign KernelConvolution_io_pixelVal_in_7 = _GEN_9046[3:0]; // @[Filter.scala 164:53 Filter.scala 166:51 Filter.scala 168:51]
  assign KernelConvolution_1_clock = clock;
  assign KernelConvolution_1_reset = reset;
  assign KernelConvolution_1_io_kernelVal_in = _GEN_9645 & _GEN_9572 ? $signed(5'sh0) : $signed(_GEN_55); // @[Filter.scala 150:41]
  assign KernelConvolution_1_io_pixelVal_in_0 = _GEN_1134[3:0]; // @[Filter.scala 164:53 Filter.scala 166:51 Filter.scala 168:51]
  assign KernelConvolution_1_io_pixelVal_in_1 = _GEN_2292[3:0]; // @[Filter.scala 164:53 Filter.scala 166:51 Filter.scala 168:51]
  assign KernelConvolution_1_io_pixelVal_in_2 = _GEN_3450[3:0]; // @[Filter.scala 164:53 Filter.scala 166:51 Filter.scala 168:51]
  assign KernelConvolution_1_io_pixelVal_in_3 = _GEN_4608[3:0]; // @[Filter.scala 164:53 Filter.scala 166:51 Filter.scala 168:51]
  assign KernelConvolution_1_io_pixelVal_in_4 = _GEN_5766[3:0]; // @[Filter.scala 164:53 Filter.scala 166:51 Filter.scala 168:51]
  assign KernelConvolution_1_io_pixelVal_in_5 = _GEN_6924[3:0]; // @[Filter.scala 164:53 Filter.scala 166:51 Filter.scala 168:51]
  assign KernelConvolution_1_io_pixelVal_in_6 = _GEN_8082[3:0]; // @[Filter.scala 164:53 Filter.scala 166:51 Filter.scala 168:51]
  assign KernelConvolution_1_io_pixelVal_in_7 = _GEN_9240[3:0]; // @[Filter.scala 164:53 Filter.scala 166:51 Filter.scala 168:51]
  assign KernelConvolution_2_clock = clock;
  assign KernelConvolution_2_reset = reset;
  assign KernelConvolution_2_io_kernelVal_in = _GEN_9645 & _GEN_9572 ? $signed(5'sh0) : $signed(_GEN_55); // @[Filter.scala 150:41]
  assign KernelConvolution_2_io_pixelVal_in_0 = _GEN_1328[3:0]; // @[Filter.scala 164:53 Filter.scala 166:51 Filter.scala 168:51]
  assign KernelConvolution_2_io_pixelVal_in_1 = _GEN_2486[3:0]; // @[Filter.scala 164:53 Filter.scala 166:51 Filter.scala 168:51]
  assign KernelConvolution_2_io_pixelVal_in_2 = _GEN_3644[3:0]; // @[Filter.scala 164:53 Filter.scala 166:51 Filter.scala 168:51]
  assign KernelConvolution_2_io_pixelVal_in_3 = _GEN_4802[3:0]; // @[Filter.scala 164:53 Filter.scala 166:51 Filter.scala 168:51]
  assign KernelConvolution_2_io_pixelVal_in_4 = _GEN_5960[3:0]; // @[Filter.scala 164:53 Filter.scala 166:51 Filter.scala 168:51]
  assign KernelConvolution_2_io_pixelVal_in_5 = _GEN_7118[3:0]; // @[Filter.scala 164:53 Filter.scala 166:51 Filter.scala 168:51]
  assign KernelConvolution_2_io_pixelVal_in_6 = _GEN_8276[3:0]; // @[Filter.scala 164:53 Filter.scala 166:51 Filter.scala 168:51]
  assign KernelConvolution_2_io_pixelVal_in_7 = _GEN_9434[3:0]; // @[Filter.scala 164:53 Filter.scala 166:51 Filter.scala 168:51]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  kernelCounter = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  imageCounterX = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  imageCounterY = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  pixelIndex = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      kernelCounter <= 4'h0;
    end else if (kernelCountReset) begin
      kernelCounter <= 4'h0;
    end else begin
      kernelCounter <= _T_14;
    end
    if (reset) begin
      imageCounterX <= 2'h0;
    end else if (imageCounterXReset) begin
      imageCounterX <= 2'h0;
    end else begin
      imageCounterX <= _T_20;
    end
    if (reset) begin
      imageCounterY <= 2'h0;
    end else if (imageCounterXReset) begin
      if (_T_21) begin
        imageCounterY <= 2'h0;
      end else begin
        imageCounterY <= _T_23;
      end
    end
    if (reset) begin
      pixelIndex <= 32'h0;
    end else if (kernelCountReset) begin
      if (_T_828) begin
        pixelIndex <= 32'h0;
      end else begin
        pixelIndex <= _T_826;
      end
    end
  end
endmodule
module VideoBuffer(
  input         clock,
  input         reset,
  input  [3:0]  io_pixelVal_in_0_0,
  input  [3:0]  io_pixelVal_in_0_1,
  input  [3:0]  io_pixelVal_in_0_2,
  input  [3:0]  io_pixelVal_in_0_3,
  input  [3:0]  io_pixelVal_in_0_4,
  input  [3:0]  io_pixelVal_in_0_5,
  input  [3:0]  io_pixelVal_in_0_6,
  input  [3:0]  io_pixelVal_in_0_7,
  input  [3:0]  io_pixelVal_in_1_0,
  input  [3:0]  io_pixelVal_in_1_1,
  input  [3:0]  io_pixelVal_in_1_2,
  input  [3:0]  io_pixelVal_in_1_3,
  input  [3:0]  io_pixelVal_in_1_4,
  input  [3:0]  io_pixelVal_in_1_5,
  input  [3:0]  io_pixelVal_in_1_6,
  input  [3:0]  io_pixelVal_in_1_7,
  input  [3:0]  io_pixelVal_in_2_0,
  input  [3:0]  io_pixelVal_in_2_1,
  input  [3:0]  io_pixelVal_in_2_2,
  input  [3:0]  io_pixelVal_in_2_3,
  input  [3:0]  io_pixelVal_in_2_4,
  input  [3:0]  io_pixelVal_in_2_5,
  input  [3:0]  io_pixelVal_in_2_6,
  input  [3:0]  io_pixelVal_in_2_7,
  input         io_valid_in,
  input  [10:0] io_rowIndex,
  input  [10:0] io_colIndex,
  output [3:0]  io_pixelVal_out_0,
  output [3:0]  io_pixelVal_out_1,
  output [3:0]  io_pixelVal_out_2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] image_0_0; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_1; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_2; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_3; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_4; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_5; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_6; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_7; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_8; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_9; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_10; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_11; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_12; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_13; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_14; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_15; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_16; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_17; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_18; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_19; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_20; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_21; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_22; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_23; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_24; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_25; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_26; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_27; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_28; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_29; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_30; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_31; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_32; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_33; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_34; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_35; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_36; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_37; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_38; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_39; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_40; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_41; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_42; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_43; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_44; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_45; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_46; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_47; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_48; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_49; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_50; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_51; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_52; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_53; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_54; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_55; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_56; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_57; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_58; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_59; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_60; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_61; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_62; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_63; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_64; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_65; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_66; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_67; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_68; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_69; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_70; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_71; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_72; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_73; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_74; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_75; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_76; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_77; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_78; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_79; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_80; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_81; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_82; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_83; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_84; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_85; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_86; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_87; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_88; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_89; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_90; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_91; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_92; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_93; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_94; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_95; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_96; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_97; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_98; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_99; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_100; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_101; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_102; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_103; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_104; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_105; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_106; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_107; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_108; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_109; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_110; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_111; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_112; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_113; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_114; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_115; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_116; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_117; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_118; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_119; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_120; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_121; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_122; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_123; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_124; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_125; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_126; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_127; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_128; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_129; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_130; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_131; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_132; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_133; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_134; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_135; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_136; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_137; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_138; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_139; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_140; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_141; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_142; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_143; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_144; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_145; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_146; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_147; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_148; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_149; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_150; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_151; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_152; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_153; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_154; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_155; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_156; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_157; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_158; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_159; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_160; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_161; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_162; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_163; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_164; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_165; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_166; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_167; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_168; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_169; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_170; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_171; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_172; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_173; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_174; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_175; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_176; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_177; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_178; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_179; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_180; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_181; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_182; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_183; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_184; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_185; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_186; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_187; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_188; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_189; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_190; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_191; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_1_0; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_1; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_2; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_3; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_4; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_5; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_6; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_7; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_8; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_9; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_10; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_11; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_12; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_13; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_14; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_15; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_16; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_17; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_18; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_19; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_20; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_21; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_22; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_23; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_24; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_25; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_26; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_27; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_28; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_29; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_30; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_31; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_32; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_33; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_34; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_35; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_36; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_37; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_38; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_39; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_40; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_41; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_42; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_43; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_44; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_45; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_46; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_47; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_48; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_49; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_50; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_51; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_52; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_53; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_54; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_55; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_56; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_57; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_58; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_59; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_60; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_61; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_62; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_63; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_64; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_65; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_66; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_67; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_68; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_69; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_70; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_71; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_72; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_73; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_74; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_75; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_76; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_77; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_78; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_79; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_80; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_81; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_82; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_83; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_84; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_85; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_86; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_87; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_88; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_89; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_90; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_91; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_92; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_93; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_94; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_95; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_96; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_97; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_98; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_99; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_100; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_101; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_102; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_103; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_104; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_105; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_106; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_107; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_108; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_109; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_110; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_111; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_112; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_113; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_114; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_115; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_116; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_117; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_118; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_119; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_120; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_121; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_122; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_123; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_124; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_125; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_126; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_127; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_128; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_129; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_130; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_131; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_132; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_133; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_134; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_135; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_136; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_137; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_138; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_139; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_140; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_141; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_142; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_143; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_144; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_145; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_146; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_147; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_148; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_149; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_150; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_151; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_152; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_153; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_154; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_155; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_156; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_157; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_158; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_159; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_160; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_161; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_162; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_163; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_164; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_165; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_166; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_167; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_168; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_169; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_170; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_171; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_172; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_173; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_174; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_175; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_176; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_177; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_178; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_179; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_180; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_181; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_182; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_183; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_184; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_185; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_186; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_187; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_188; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_189; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_190; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_191; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_2_0; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_1; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_2; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_3; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_4; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_5; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_6; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_7; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_8; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_9; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_10; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_11; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_12; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_13; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_14; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_15; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_16; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_17; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_18; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_19; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_20; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_21; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_22; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_23; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_24; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_25; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_26; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_27; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_28; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_29; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_30; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_31; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_32; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_33; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_34; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_35; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_36; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_37; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_38; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_39; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_40; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_41; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_42; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_43; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_44; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_45; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_46; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_47; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_48; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_49; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_50; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_51; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_52; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_53; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_54; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_55; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_56; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_57; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_58; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_59; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_60; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_61; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_62; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_63; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_64; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_65; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_66; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_67; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_68; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_69; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_70; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_71; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_72; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_73; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_74; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_75; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_76; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_77; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_78; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_79; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_80; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_81; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_82; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_83; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_84; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_85; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_86; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_87; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_88; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_89; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_90; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_91; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_92; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_93; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_94; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_95; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_96; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_97; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_98; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_99; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_100; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_101; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_102; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_103; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_104; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_105; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_106; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_107; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_108; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_109; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_110; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_111; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_112; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_113; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_114; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_115; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_116; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_117; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_118; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_119; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_120; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_121; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_122; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_123; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_124; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_125; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_126; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_127; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_128; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_129; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_130; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_131; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_132; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_133; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_134; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_135; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_136; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_137; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_138; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_139; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_140; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_141; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_142; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_143; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_144; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_145; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_146; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_147; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_148; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_149; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_150; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_151; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_152; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_153; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_154; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_155; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_156; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_157; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_158; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_159; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_160; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_161; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_162; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_163; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_164; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_165; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_166; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_167; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_168; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_169; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_170; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_171; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_172; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_173; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_174; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_175; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_176; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_177; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_178; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_179; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_180; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_181; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_182; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_183; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_184; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_185; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_186; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_187; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_188; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_189; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_190; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_191; // @[VideoBuffer.scala 21:25]
  reg [31:0] pixelIndex; // @[VideoBuffer.scala 24:33]
  wire [15:0] _T_3 = io_rowIndex * 11'h10; // @[VideoBuffer.scala 27:54]
  wire [15:0] _GEN_5762 = {{5'd0}, io_colIndex}; // @[VideoBuffer.scala 27:69]
  wire [15:0] _T_5 = _T_3 + _GEN_5762; // @[VideoBuffer.scala 27:69]
  wire [3:0] _GEN_1 = 8'h1 == _T_5[7:0] ? image_0_1 : image_0_0; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2 = 8'h2 == _T_5[7:0] ? image_0_2 : _GEN_1; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3 = 8'h3 == _T_5[7:0] ? image_0_3 : _GEN_2; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4 = 8'h4 == _T_5[7:0] ? image_0_4 : _GEN_3; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_5 = 8'h5 == _T_5[7:0] ? image_0_5 : _GEN_4; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_6 = 8'h6 == _T_5[7:0] ? image_0_6 : _GEN_5; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_7 = 8'h7 == _T_5[7:0] ? image_0_7 : _GEN_6; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_8 = 8'h8 == _T_5[7:0] ? image_0_8 : _GEN_7; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_9 = 8'h9 == _T_5[7:0] ? image_0_9 : _GEN_8; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_10 = 8'ha == _T_5[7:0] ? image_0_10 : _GEN_9; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_11 = 8'hb == _T_5[7:0] ? image_0_11 : _GEN_10; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_12 = 8'hc == _T_5[7:0] ? image_0_12 : _GEN_11; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_13 = 8'hd == _T_5[7:0] ? image_0_13 : _GEN_12; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_14 = 8'he == _T_5[7:0] ? image_0_14 : _GEN_13; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_15 = 8'hf == _T_5[7:0] ? image_0_15 : _GEN_14; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_16 = 8'h10 == _T_5[7:0] ? image_0_16 : _GEN_15; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_17 = 8'h11 == _T_5[7:0] ? image_0_17 : _GEN_16; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_18 = 8'h12 == _T_5[7:0] ? image_0_18 : _GEN_17; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_19 = 8'h13 == _T_5[7:0] ? image_0_19 : _GEN_18; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_20 = 8'h14 == _T_5[7:0] ? image_0_20 : _GEN_19; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_21 = 8'h15 == _T_5[7:0] ? image_0_21 : _GEN_20; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_22 = 8'h16 == _T_5[7:0] ? image_0_22 : _GEN_21; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_23 = 8'h17 == _T_5[7:0] ? image_0_23 : _GEN_22; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_24 = 8'h18 == _T_5[7:0] ? image_0_24 : _GEN_23; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_25 = 8'h19 == _T_5[7:0] ? image_0_25 : _GEN_24; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_26 = 8'h1a == _T_5[7:0] ? image_0_26 : _GEN_25; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_27 = 8'h1b == _T_5[7:0] ? image_0_27 : _GEN_26; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_28 = 8'h1c == _T_5[7:0] ? image_0_28 : _GEN_27; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_29 = 8'h1d == _T_5[7:0] ? image_0_29 : _GEN_28; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_30 = 8'h1e == _T_5[7:0] ? image_0_30 : _GEN_29; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_31 = 8'h1f == _T_5[7:0] ? image_0_31 : _GEN_30; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_32 = 8'h20 == _T_5[7:0] ? image_0_32 : _GEN_31; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_33 = 8'h21 == _T_5[7:0] ? image_0_33 : _GEN_32; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_34 = 8'h22 == _T_5[7:0] ? image_0_34 : _GEN_33; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_35 = 8'h23 == _T_5[7:0] ? image_0_35 : _GEN_34; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_36 = 8'h24 == _T_5[7:0] ? image_0_36 : _GEN_35; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_37 = 8'h25 == _T_5[7:0] ? image_0_37 : _GEN_36; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_38 = 8'h26 == _T_5[7:0] ? image_0_38 : _GEN_37; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_39 = 8'h27 == _T_5[7:0] ? image_0_39 : _GEN_38; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_40 = 8'h28 == _T_5[7:0] ? image_0_40 : _GEN_39; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_41 = 8'h29 == _T_5[7:0] ? image_0_41 : _GEN_40; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_42 = 8'h2a == _T_5[7:0] ? image_0_42 : _GEN_41; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_43 = 8'h2b == _T_5[7:0] ? image_0_43 : _GEN_42; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_44 = 8'h2c == _T_5[7:0] ? image_0_44 : _GEN_43; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_45 = 8'h2d == _T_5[7:0] ? image_0_45 : _GEN_44; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_46 = 8'h2e == _T_5[7:0] ? image_0_46 : _GEN_45; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_47 = 8'h2f == _T_5[7:0] ? image_0_47 : _GEN_46; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_48 = 8'h30 == _T_5[7:0] ? image_0_48 : _GEN_47; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_49 = 8'h31 == _T_5[7:0] ? image_0_49 : _GEN_48; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_50 = 8'h32 == _T_5[7:0] ? image_0_50 : _GEN_49; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_51 = 8'h33 == _T_5[7:0] ? image_0_51 : _GEN_50; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_52 = 8'h34 == _T_5[7:0] ? image_0_52 : _GEN_51; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_53 = 8'h35 == _T_5[7:0] ? image_0_53 : _GEN_52; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_54 = 8'h36 == _T_5[7:0] ? image_0_54 : _GEN_53; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_55 = 8'h37 == _T_5[7:0] ? image_0_55 : _GEN_54; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_56 = 8'h38 == _T_5[7:0] ? image_0_56 : _GEN_55; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_57 = 8'h39 == _T_5[7:0] ? image_0_57 : _GEN_56; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_58 = 8'h3a == _T_5[7:0] ? image_0_58 : _GEN_57; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_59 = 8'h3b == _T_5[7:0] ? image_0_59 : _GEN_58; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_60 = 8'h3c == _T_5[7:0] ? image_0_60 : _GEN_59; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_61 = 8'h3d == _T_5[7:0] ? image_0_61 : _GEN_60; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_62 = 8'h3e == _T_5[7:0] ? image_0_62 : _GEN_61; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_63 = 8'h3f == _T_5[7:0] ? image_0_63 : _GEN_62; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_64 = 8'h40 == _T_5[7:0] ? image_0_64 : _GEN_63; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_65 = 8'h41 == _T_5[7:0] ? image_0_65 : _GEN_64; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_66 = 8'h42 == _T_5[7:0] ? image_0_66 : _GEN_65; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_67 = 8'h43 == _T_5[7:0] ? image_0_67 : _GEN_66; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_68 = 8'h44 == _T_5[7:0] ? image_0_68 : _GEN_67; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_69 = 8'h45 == _T_5[7:0] ? image_0_69 : _GEN_68; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_70 = 8'h46 == _T_5[7:0] ? image_0_70 : _GEN_69; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_71 = 8'h47 == _T_5[7:0] ? image_0_71 : _GEN_70; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_72 = 8'h48 == _T_5[7:0] ? image_0_72 : _GEN_71; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_73 = 8'h49 == _T_5[7:0] ? image_0_73 : _GEN_72; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_74 = 8'h4a == _T_5[7:0] ? image_0_74 : _GEN_73; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_75 = 8'h4b == _T_5[7:0] ? image_0_75 : _GEN_74; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_76 = 8'h4c == _T_5[7:0] ? image_0_76 : _GEN_75; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_77 = 8'h4d == _T_5[7:0] ? image_0_77 : _GEN_76; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_78 = 8'h4e == _T_5[7:0] ? image_0_78 : _GEN_77; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_79 = 8'h4f == _T_5[7:0] ? image_0_79 : _GEN_78; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_80 = 8'h50 == _T_5[7:0] ? image_0_80 : _GEN_79; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_81 = 8'h51 == _T_5[7:0] ? image_0_81 : _GEN_80; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_82 = 8'h52 == _T_5[7:0] ? image_0_82 : _GEN_81; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_83 = 8'h53 == _T_5[7:0] ? image_0_83 : _GEN_82; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_84 = 8'h54 == _T_5[7:0] ? image_0_84 : _GEN_83; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_85 = 8'h55 == _T_5[7:0] ? image_0_85 : _GEN_84; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_86 = 8'h56 == _T_5[7:0] ? image_0_86 : _GEN_85; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_87 = 8'h57 == _T_5[7:0] ? image_0_87 : _GEN_86; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_88 = 8'h58 == _T_5[7:0] ? image_0_88 : _GEN_87; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_89 = 8'h59 == _T_5[7:0] ? image_0_89 : _GEN_88; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_90 = 8'h5a == _T_5[7:0] ? image_0_90 : _GEN_89; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_91 = 8'h5b == _T_5[7:0] ? image_0_91 : _GEN_90; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_92 = 8'h5c == _T_5[7:0] ? image_0_92 : _GEN_91; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_93 = 8'h5d == _T_5[7:0] ? image_0_93 : _GEN_92; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_94 = 8'h5e == _T_5[7:0] ? image_0_94 : _GEN_93; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_95 = 8'h5f == _T_5[7:0] ? image_0_95 : _GEN_94; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_96 = 8'h60 == _T_5[7:0] ? image_0_96 : _GEN_95; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_97 = 8'h61 == _T_5[7:0] ? image_0_97 : _GEN_96; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_98 = 8'h62 == _T_5[7:0] ? image_0_98 : _GEN_97; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_99 = 8'h63 == _T_5[7:0] ? image_0_99 : _GEN_98; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_100 = 8'h64 == _T_5[7:0] ? image_0_100 : _GEN_99; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_101 = 8'h65 == _T_5[7:0] ? image_0_101 : _GEN_100; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_102 = 8'h66 == _T_5[7:0] ? image_0_102 : _GEN_101; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_103 = 8'h67 == _T_5[7:0] ? image_0_103 : _GEN_102; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_104 = 8'h68 == _T_5[7:0] ? image_0_104 : _GEN_103; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_105 = 8'h69 == _T_5[7:0] ? image_0_105 : _GEN_104; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_106 = 8'h6a == _T_5[7:0] ? image_0_106 : _GEN_105; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_107 = 8'h6b == _T_5[7:0] ? image_0_107 : _GEN_106; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_108 = 8'h6c == _T_5[7:0] ? image_0_108 : _GEN_107; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_109 = 8'h6d == _T_5[7:0] ? image_0_109 : _GEN_108; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_110 = 8'h6e == _T_5[7:0] ? image_0_110 : _GEN_109; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_111 = 8'h6f == _T_5[7:0] ? image_0_111 : _GEN_110; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_112 = 8'h70 == _T_5[7:0] ? image_0_112 : _GEN_111; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_113 = 8'h71 == _T_5[7:0] ? image_0_113 : _GEN_112; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_114 = 8'h72 == _T_5[7:0] ? image_0_114 : _GEN_113; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_115 = 8'h73 == _T_5[7:0] ? image_0_115 : _GEN_114; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_116 = 8'h74 == _T_5[7:0] ? image_0_116 : _GEN_115; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_117 = 8'h75 == _T_5[7:0] ? image_0_117 : _GEN_116; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_118 = 8'h76 == _T_5[7:0] ? image_0_118 : _GEN_117; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_119 = 8'h77 == _T_5[7:0] ? image_0_119 : _GEN_118; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_120 = 8'h78 == _T_5[7:0] ? image_0_120 : _GEN_119; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_121 = 8'h79 == _T_5[7:0] ? image_0_121 : _GEN_120; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_122 = 8'h7a == _T_5[7:0] ? image_0_122 : _GEN_121; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_123 = 8'h7b == _T_5[7:0] ? image_0_123 : _GEN_122; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_124 = 8'h7c == _T_5[7:0] ? image_0_124 : _GEN_123; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_125 = 8'h7d == _T_5[7:0] ? image_0_125 : _GEN_124; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_126 = 8'h7e == _T_5[7:0] ? image_0_126 : _GEN_125; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_127 = 8'h7f == _T_5[7:0] ? image_0_127 : _GEN_126; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_128 = 8'h80 == _T_5[7:0] ? image_0_128 : _GEN_127; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_129 = 8'h81 == _T_5[7:0] ? image_0_129 : _GEN_128; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_130 = 8'h82 == _T_5[7:0] ? image_0_130 : _GEN_129; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_131 = 8'h83 == _T_5[7:0] ? image_0_131 : _GEN_130; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_132 = 8'h84 == _T_5[7:0] ? image_0_132 : _GEN_131; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_133 = 8'h85 == _T_5[7:0] ? image_0_133 : _GEN_132; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_134 = 8'h86 == _T_5[7:0] ? image_0_134 : _GEN_133; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_135 = 8'h87 == _T_5[7:0] ? image_0_135 : _GEN_134; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_136 = 8'h88 == _T_5[7:0] ? image_0_136 : _GEN_135; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_137 = 8'h89 == _T_5[7:0] ? image_0_137 : _GEN_136; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_138 = 8'h8a == _T_5[7:0] ? image_0_138 : _GEN_137; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_139 = 8'h8b == _T_5[7:0] ? image_0_139 : _GEN_138; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_140 = 8'h8c == _T_5[7:0] ? image_0_140 : _GEN_139; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_141 = 8'h8d == _T_5[7:0] ? image_0_141 : _GEN_140; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_142 = 8'h8e == _T_5[7:0] ? image_0_142 : _GEN_141; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_143 = 8'h8f == _T_5[7:0] ? image_0_143 : _GEN_142; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_144 = 8'h90 == _T_5[7:0] ? image_0_144 : _GEN_143; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_145 = 8'h91 == _T_5[7:0] ? image_0_145 : _GEN_144; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_146 = 8'h92 == _T_5[7:0] ? image_0_146 : _GEN_145; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_147 = 8'h93 == _T_5[7:0] ? image_0_147 : _GEN_146; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_148 = 8'h94 == _T_5[7:0] ? image_0_148 : _GEN_147; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_149 = 8'h95 == _T_5[7:0] ? image_0_149 : _GEN_148; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_150 = 8'h96 == _T_5[7:0] ? image_0_150 : _GEN_149; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_151 = 8'h97 == _T_5[7:0] ? image_0_151 : _GEN_150; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_152 = 8'h98 == _T_5[7:0] ? image_0_152 : _GEN_151; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_153 = 8'h99 == _T_5[7:0] ? image_0_153 : _GEN_152; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_154 = 8'h9a == _T_5[7:0] ? image_0_154 : _GEN_153; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_155 = 8'h9b == _T_5[7:0] ? image_0_155 : _GEN_154; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_156 = 8'h9c == _T_5[7:0] ? image_0_156 : _GEN_155; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_157 = 8'h9d == _T_5[7:0] ? image_0_157 : _GEN_156; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_158 = 8'h9e == _T_5[7:0] ? image_0_158 : _GEN_157; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_159 = 8'h9f == _T_5[7:0] ? image_0_159 : _GEN_158; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_160 = 8'ha0 == _T_5[7:0] ? image_0_160 : _GEN_159; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_161 = 8'ha1 == _T_5[7:0] ? image_0_161 : _GEN_160; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_162 = 8'ha2 == _T_5[7:0] ? image_0_162 : _GEN_161; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_163 = 8'ha3 == _T_5[7:0] ? image_0_163 : _GEN_162; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_164 = 8'ha4 == _T_5[7:0] ? image_0_164 : _GEN_163; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_165 = 8'ha5 == _T_5[7:0] ? image_0_165 : _GEN_164; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_166 = 8'ha6 == _T_5[7:0] ? image_0_166 : _GEN_165; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_167 = 8'ha7 == _T_5[7:0] ? image_0_167 : _GEN_166; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_168 = 8'ha8 == _T_5[7:0] ? image_0_168 : _GEN_167; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_169 = 8'ha9 == _T_5[7:0] ? image_0_169 : _GEN_168; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_170 = 8'haa == _T_5[7:0] ? image_0_170 : _GEN_169; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_171 = 8'hab == _T_5[7:0] ? image_0_171 : _GEN_170; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_172 = 8'hac == _T_5[7:0] ? image_0_172 : _GEN_171; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_173 = 8'had == _T_5[7:0] ? image_0_173 : _GEN_172; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_174 = 8'hae == _T_5[7:0] ? image_0_174 : _GEN_173; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_175 = 8'haf == _T_5[7:0] ? image_0_175 : _GEN_174; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_176 = 8'hb0 == _T_5[7:0] ? image_0_176 : _GEN_175; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_177 = 8'hb1 == _T_5[7:0] ? image_0_177 : _GEN_176; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_178 = 8'hb2 == _T_5[7:0] ? image_0_178 : _GEN_177; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_179 = 8'hb3 == _T_5[7:0] ? image_0_179 : _GEN_178; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_180 = 8'hb4 == _T_5[7:0] ? image_0_180 : _GEN_179; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_181 = 8'hb5 == _T_5[7:0] ? image_0_181 : _GEN_180; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_182 = 8'hb6 == _T_5[7:0] ? image_0_182 : _GEN_181; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_183 = 8'hb7 == _T_5[7:0] ? image_0_183 : _GEN_182; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_184 = 8'hb8 == _T_5[7:0] ? image_0_184 : _GEN_183; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_185 = 8'hb9 == _T_5[7:0] ? image_0_185 : _GEN_184; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_186 = 8'hba == _T_5[7:0] ? image_0_186 : _GEN_185; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_187 = 8'hbb == _T_5[7:0] ? image_0_187 : _GEN_186; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_188 = 8'hbc == _T_5[7:0] ? image_0_188 : _GEN_187; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_189 = 8'hbd == _T_5[7:0] ? image_0_189 : _GEN_188; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_190 = 8'hbe == _T_5[7:0] ? image_0_190 : _GEN_189; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_193 = 8'h1 == _T_5[7:0] ? image_1_1 : image_1_0; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_194 = 8'h2 == _T_5[7:0] ? image_1_2 : _GEN_193; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_195 = 8'h3 == _T_5[7:0] ? image_1_3 : _GEN_194; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_196 = 8'h4 == _T_5[7:0] ? image_1_4 : _GEN_195; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_197 = 8'h5 == _T_5[7:0] ? image_1_5 : _GEN_196; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_198 = 8'h6 == _T_5[7:0] ? image_1_6 : _GEN_197; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_199 = 8'h7 == _T_5[7:0] ? image_1_7 : _GEN_198; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_200 = 8'h8 == _T_5[7:0] ? image_1_8 : _GEN_199; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_201 = 8'h9 == _T_5[7:0] ? image_1_9 : _GEN_200; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_202 = 8'ha == _T_5[7:0] ? image_1_10 : _GEN_201; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_203 = 8'hb == _T_5[7:0] ? image_1_11 : _GEN_202; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_204 = 8'hc == _T_5[7:0] ? image_1_12 : _GEN_203; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_205 = 8'hd == _T_5[7:0] ? image_1_13 : _GEN_204; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_206 = 8'he == _T_5[7:0] ? image_1_14 : _GEN_205; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_207 = 8'hf == _T_5[7:0] ? image_1_15 : _GEN_206; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_208 = 8'h10 == _T_5[7:0] ? image_1_16 : _GEN_207; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_209 = 8'h11 == _T_5[7:0] ? image_1_17 : _GEN_208; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_210 = 8'h12 == _T_5[7:0] ? image_1_18 : _GEN_209; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_211 = 8'h13 == _T_5[7:0] ? image_1_19 : _GEN_210; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_212 = 8'h14 == _T_5[7:0] ? image_1_20 : _GEN_211; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_213 = 8'h15 == _T_5[7:0] ? image_1_21 : _GEN_212; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_214 = 8'h16 == _T_5[7:0] ? image_1_22 : _GEN_213; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_215 = 8'h17 == _T_5[7:0] ? image_1_23 : _GEN_214; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_216 = 8'h18 == _T_5[7:0] ? image_1_24 : _GEN_215; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_217 = 8'h19 == _T_5[7:0] ? image_1_25 : _GEN_216; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_218 = 8'h1a == _T_5[7:0] ? image_1_26 : _GEN_217; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_219 = 8'h1b == _T_5[7:0] ? image_1_27 : _GEN_218; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_220 = 8'h1c == _T_5[7:0] ? image_1_28 : _GEN_219; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_221 = 8'h1d == _T_5[7:0] ? image_1_29 : _GEN_220; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_222 = 8'h1e == _T_5[7:0] ? image_1_30 : _GEN_221; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_223 = 8'h1f == _T_5[7:0] ? image_1_31 : _GEN_222; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_224 = 8'h20 == _T_5[7:0] ? image_1_32 : _GEN_223; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_225 = 8'h21 == _T_5[7:0] ? image_1_33 : _GEN_224; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_226 = 8'h22 == _T_5[7:0] ? image_1_34 : _GEN_225; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_227 = 8'h23 == _T_5[7:0] ? image_1_35 : _GEN_226; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_228 = 8'h24 == _T_5[7:0] ? image_1_36 : _GEN_227; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_229 = 8'h25 == _T_5[7:0] ? image_1_37 : _GEN_228; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_230 = 8'h26 == _T_5[7:0] ? image_1_38 : _GEN_229; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_231 = 8'h27 == _T_5[7:0] ? image_1_39 : _GEN_230; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_232 = 8'h28 == _T_5[7:0] ? image_1_40 : _GEN_231; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_233 = 8'h29 == _T_5[7:0] ? image_1_41 : _GEN_232; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_234 = 8'h2a == _T_5[7:0] ? image_1_42 : _GEN_233; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_235 = 8'h2b == _T_5[7:0] ? image_1_43 : _GEN_234; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_236 = 8'h2c == _T_5[7:0] ? image_1_44 : _GEN_235; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_237 = 8'h2d == _T_5[7:0] ? image_1_45 : _GEN_236; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_238 = 8'h2e == _T_5[7:0] ? image_1_46 : _GEN_237; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_239 = 8'h2f == _T_5[7:0] ? image_1_47 : _GEN_238; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_240 = 8'h30 == _T_5[7:0] ? image_1_48 : _GEN_239; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_241 = 8'h31 == _T_5[7:0] ? image_1_49 : _GEN_240; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_242 = 8'h32 == _T_5[7:0] ? image_1_50 : _GEN_241; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_243 = 8'h33 == _T_5[7:0] ? image_1_51 : _GEN_242; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_244 = 8'h34 == _T_5[7:0] ? image_1_52 : _GEN_243; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_245 = 8'h35 == _T_5[7:0] ? image_1_53 : _GEN_244; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_246 = 8'h36 == _T_5[7:0] ? image_1_54 : _GEN_245; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_247 = 8'h37 == _T_5[7:0] ? image_1_55 : _GEN_246; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_248 = 8'h38 == _T_5[7:0] ? image_1_56 : _GEN_247; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_249 = 8'h39 == _T_5[7:0] ? image_1_57 : _GEN_248; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_250 = 8'h3a == _T_5[7:0] ? image_1_58 : _GEN_249; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_251 = 8'h3b == _T_5[7:0] ? image_1_59 : _GEN_250; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_252 = 8'h3c == _T_5[7:0] ? image_1_60 : _GEN_251; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_253 = 8'h3d == _T_5[7:0] ? image_1_61 : _GEN_252; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_254 = 8'h3e == _T_5[7:0] ? image_1_62 : _GEN_253; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_255 = 8'h3f == _T_5[7:0] ? image_1_63 : _GEN_254; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_256 = 8'h40 == _T_5[7:0] ? image_1_64 : _GEN_255; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_257 = 8'h41 == _T_5[7:0] ? image_1_65 : _GEN_256; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_258 = 8'h42 == _T_5[7:0] ? image_1_66 : _GEN_257; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_259 = 8'h43 == _T_5[7:0] ? image_1_67 : _GEN_258; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_260 = 8'h44 == _T_5[7:0] ? image_1_68 : _GEN_259; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_261 = 8'h45 == _T_5[7:0] ? image_1_69 : _GEN_260; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_262 = 8'h46 == _T_5[7:0] ? image_1_70 : _GEN_261; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_263 = 8'h47 == _T_5[7:0] ? image_1_71 : _GEN_262; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_264 = 8'h48 == _T_5[7:0] ? image_1_72 : _GEN_263; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_265 = 8'h49 == _T_5[7:0] ? image_1_73 : _GEN_264; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_266 = 8'h4a == _T_5[7:0] ? image_1_74 : _GEN_265; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_267 = 8'h4b == _T_5[7:0] ? image_1_75 : _GEN_266; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_268 = 8'h4c == _T_5[7:0] ? image_1_76 : _GEN_267; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_269 = 8'h4d == _T_5[7:0] ? image_1_77 : _GEN_268; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_270 = 8'h4e == _T_5[7:0] ? image_1_78 : _GEN_269; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_271 = 8'h4f == _T_5[7:0] ? image_1_79 : _GEN_270; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_272 = 8'h50 == _T_5[7:0] ? image_1_80 : _GEN_271; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_273 = 8'h51 == _T_5[7:0] ? image_1_81 : _GEN_272; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_274 = 8'h52 == _T_5[7:0] ? image_1_82 : _GEN_273; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_275 = 8'h53 == _T_5[7:0] ? image_1_83 : _GEN_274; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_276 = 8'h54 == _T_5[7:0] ? image_1_84 : _GEN_275; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_277 = 8'h55 == _T_5[7:0] ? image_1_85 : _GEN_276; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_278 = 8'h56 == _T_5[7:0] ? image_1_86 : _GEN_277; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_279 = 8'h57 == _T_5[7:0] ? image_1_87 : _GEN_278; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_280 = 8'h58 == _T_5[7:0] ? image_1_88 : _GEN_279; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_281 = 8'h59 == _T_5[7:0] ? image_1_89 : _GEN_280; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_282 = 8'h5a == _T_5[7:0] ? image_1_90 : _GEN_281; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_283 = 8'h5b == _T_5[7:0] ? image_1_91 : _GEN_282; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_284 = 8'h5c == _T_5[7:0] ? image_1_92 : _GEN_283; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_285 = 8'h5d == _T_5[7:0] ? image_1_93 : _GEN_284; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_286 = 8'h5e == _T_5[7:0] ? image_1_94 : _GEN_285; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_287 = 8'h5f == _T_5[7:0] ? image_1_95 : _GEN_286; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_288 = 8'h60 == _T_5[7:0] ? image_1_96 : _GEN_287; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_289 = 8'h61 == _T_5[7:0] ? image_1_97 : _GEN_288; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_290 = 8'h62 == _T_5[7:0] ? image_1_98 : _GEN_289; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_291 = 8'h63 == _T_5[7:0] ? image_1_99 : _GEN_290; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_292 = 8'h64 == _T_5[7:0] ? image_1_100 : _GEN_291; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_293 = 8'h65 == _T_5[7:0] ? image_1_101 : _GEN_292; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_294 = 8'h66 == _T_5[7:0] ? image_1_102 : _GEN_293; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_295 = 8'h67 == _T_5[7:0] ? image_1_103 : _GEN_294; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_296 = 8'h68 == _T_5[7:0] ? image_1_104 : _GEN_295; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_297 = 8'h69 == _T_5[7:0] ? image_1_105 : _GEN_296; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_298 = 8'h6a == _T_5[7:0] ? image_1_106 : _GEN_297; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_299 = 8'h6b == _T_5[7:0] ? image_1_107 : _GEN_298; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_300 = 8'h6c == _T_5[7:0] ? image_1_108 : _GEN_299; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_301 = 8'h6d == _T_5[7:0] ? image_1_109 : _GEN_300; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_302 = 8'h6e == _T_5[7:0] ? image_1_110 : _GEN_301; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_303 = 8'h6f == _T_5[7:0] ? image_1_111 : _GEN_302; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_304 = 8'h70 == _T_5[7:0] ? image_1_112 : _GEN_303; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_305 = 8'h71 == _T_5[7:0] ? image_1_113 : _GEN_304; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_306 = 8'h72 == _T_5[7:0] ? image_1_114 : _GEN_305; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_307 = 8'h73 == _T_5[7:0] ? image_1_115 : _GEN_306; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_308 = 8'h74 == _T_5[7:0] ? image_1_116 : _GEN_307; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_309 = 8'h75 == _T_5[7:0] ? image_1_117 : _GEN_308; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_310 = 8'h76 == _T_5[7:0] ? image_1_118 : _GEN_309; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_311 = 8'h77 == _T_5[7:0] ? image_1_119 : _GEN_310; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_312 = 8'h78 == _T_5[7:0] ? image_1_120 : _GEN_311; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_313 = 8'h79 == _T_5[7:0] ? image_1_121 : _GEN_312; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_314 = 8'h7a == _T_5[7:0] ? image_1_122 : _GEN_313; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_315 = 8'h7b == _T_5[7:0] ? image_1_123 : _GEN_314; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_316 = 8'h7c == _T_5[7:0] ? image_1_124 : _GEN_315; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_317 = 8'h7d == _T_5[7:0] ? image_1_125 : _GEN_316; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_318 = 8'h7e == _T_5[7:0] ? image_1_126 : _GEN_317; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_319 = 8'h7f == _T_5[7:0] ? image_1_127 : _GEN_318; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_320 = 8'h80 == _T_5[7:0] ? image_1_128 : _GEN_319; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_321 = 8'h81 == _T_5[7:0] ? image_1_129 : _GEN_320; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_322 = 8'h82 == _T_5[7:0] ? image_1_130 : _GEN_321; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_323 = 8'h83 == _T_5[7:0] ? image_1_131 : _GEN_322; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_324 = 8'h84 == _T_5[7:0] ? image_1_132 : _GEN_323; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_325 = 8'h85 == _T_5[7:0] ? image_1_133 : _GEN_324; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_326 = 8'h86 == _T_5[7:0] ? image_1_134 : _GEN_325; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_327 = 8'h87 == _T_5[7:0] ? image_1_135 : _GEN_326; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_328 = 8'h88 == _T_5[7:0] ? image_1_136 : _GEN_327; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_329 = 8'h89 == _T_5[7:0] ? image_1_137 : _GEN_328; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_330 = 8'h8a == _T_5[7:0] ? image_1_138 : _GEN_329; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_331 = 8'h8b == _T_5[7:0] ? image_1_139 : _GEN_330; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_332 = 8'h8c == _T_5[7:0] ? image_1_140 : _GEN_331; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_333 = 8'h8d == _T_5[7:0] ? image_1_141 : _GEN_332; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_334 = 8'h8e == _T_5[7:0] ? image_1_142 : _GEN_333; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_335 = 8'h8f == _T_5[7:0] ? image_1_143 : _GEN_334; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_336 = 8'h90 == _T_5[7:0] ? image_1_144 : _GEN_335; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_337 = 8'h91 == _T_5[7:0] ? image_1_145 : _GEN_336; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_338 = 8'h92 == _T_5[7:0] ? image_1_146 : _GEN_337; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_339 = 8'h93 == _T_5[7:0] ? image_1_147 : _GEN_338; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_340 = 8'h94 == _T_5[7:0] ? image_1_148 : _GEN_339; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_341 = 8'h95 == _T_5[7:0] ? image_1_149 : _GEN_340; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_342 = 8'h96 == _T_5[7:0] ? image_1_150 : _GEN_341; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_343 = 8'h97 == _T_5[7:0] ? image_1_151 : _GEN_342; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_344 = 8'h98 == _T_5[7:0] ? image_1_152 : _GEN_343; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_345 = 8'h99 == _T_5[7:0] ? image_1_153 : _GEN_344; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_346 = 8'h9a == _T_5[7:0] ? image_1_154 : _GEN_345; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_347 = 8'h9b == _T_5[7:0] ? image_1_155 : _GEN_346; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_348 = 8'h9c == _T_5[7:0] ? image_1_156 : _GEN_347; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_349 = 8'h9d == _T_5[7:0] ? image_1_157 : _GEN_348; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_350 = 8'h9e == _T_5[7:0] ? image_1_158 : _GEN_349; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_351 = 8'h9f == _T_5[7:0] ? image_1_159 : _GEN_350; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_352 = 8'ha0 == _T_5[7:0] ? image_1_160 : _GEN_351; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_353 = 8'ha1 == _T_5[7:0] ? image_1_161 : _GEN_352; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_354 = 8'ha2 == _T_5[7:0] ? image_1_162 : _GEN_353; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_355 = 8'ha3 == _T_5[7:0] ? image_1_163 : _GEN_354; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_356 = 8'ha4 == _T_5[7:0] ? image_1_164 : _GEN_355; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_357 = 8'ha5 == _T_5[7:0] ? image_1_165 : _GEN_356; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_358 = 8'ha6 == _T_5[7:0] ? image_1_166 : _GEN_357; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_359 = 8'ha7 == _T_5[7:0] ? image_1_167 : _GEN_358; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_360 = 8'ha8 == _T_5[7:0] ? image_1_168 : _GEN_359; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_361 = 8'ha9 == _T_5[7:0] ? image_1_169 : _GEN_360; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_362 = 8'haa == _T_5[7:0] ? image_1_170 : _GEN_361; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_363 = 8'hab == _T_5[7:0] ? image_1_171 : _GEN_362; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_364 = 8'hac == _T_5[7:0] ? image_1_172 : _GEN_363; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_365 = 8'had == _T_5[7:0] ? image_1_173 : _GEN_364; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_366 = 8'hae == _T_5[7:0] ? image_1_174 : _GEN_365; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_367 = 8'haf == _T_5[7:0] ? image_1_175 : _GEN_366; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_368 = 8'hb0 == _T_5[7:0] ? image_1_176 : _GEN_367; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_369 = 8'hb1 == _T_5[7:0] ? image_1_177 : _GEN_368; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_370 = 8'hb2 == _T_5[7:0] ? image_1_178 : _GEN_369; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_371 = 8'hb3 == _T_5[7:0] ? image_1_179 : _GEN_370; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_372 = 8'hb4 == _T_5[7:0] ? image_1_180 : _GEN_371; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_373 = 8'hb5 == _T_5[7:0] ? image_1_181 : _GEN_372; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_374 = 8'hb6 == _T_5[7:0] ? image_1_182 : _GEN_373; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_375 = 8'hb7 == _T_5[7:0] ? image_1_183 : _GEN_374; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_376 = 8'hb8 == _T_5[7:0] ? image_1_184 : _GEN_375; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_377 = 8'hb9 == _T_5[7:0] ? image_1_185 : _GEN_376; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_378 = 8'hba == _T_5[7:0] ? image_1_186 : _GEN_377; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_379 = 8'hbb == _T_5[7:0] ? image_1_187 : _GEN_378; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_380 = 8'hbc == _T_5[7:0] ? image_1_188 : _GEN_379; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_381 = 8'hbd == _T_5[7:0] ? image_1_189 : _GEN_380; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_382 = 8'hbe == _T_5[7:0] ? image_1_190 : _GEN_381; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_385 = 8'h1 == _T_5[7:0] ? image_2_1 : image_2_0; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_386 = 8'h2 == _T_5[7:0] ? image_2_2 : _GEN_385; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_387 = 8'h3 == _T_5[7:0] ? image_2_3 : _GEN_386; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_388 = 8'h4 == _T_5[7:0] ? image_2_4 : _GEN_387; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_389 = 8'h5 == _T_5[7:0] ? image_2_5 : _GEN_388; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_390 = 8'h6 == _T_5[7:0] ? image_2_6 : _GEN_389; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_391 = 8'h7 == _T_5[7:0] ? image_2_7 : _GEN_390; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_392 = 8'h8 == _T_5[7:0] ? image_2_8 : _GEN_391; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_393 = 8'h9 == _T_5[7:0] ? image_2_9 : _GEN_392; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_394 = 8'ha == _T_5[7:0] ? image_2_10 : _GEN_393; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_395 = 8'hb == _T_5[7:0] ? image_2_11 : _GEN_394; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_396 = 8'hc == _T_5[7:0] ? image_2_12 : _GEN_395; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_397 = 8'hd == _T_5[7:0] ? image_2_13 : _GEN_396; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_398 = 8'he == _T_5[7:0] ? image_2_14 : _GEN_397; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_399 = 8'hf == _T_5[7:0] ? image_2_15 : _GEN_398; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_400 = 8'h10 == _T_5[7:0] ? image_2_16 : _GEN_399; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_401 = 8'h11 == _T_5[7:0] ? image_2_17 : _GEN_400; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_402 = 8'h12 == _T_5[7:0] ? image_2_18 : _GEN_401; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_403 = 8'h13 == _T_5[7:0] ? image_2_19 : _GEN_402; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_404 = 8'h14 == _T_5[7:0] ? image_2_20 : _GEN_403; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_405 = 8'h15 == _T_5[7:0] ? image_2_21 : _GEN_404; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_406 = 8'h16 == _T_5[7:0] ? image_2_22 : _GEN_405; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_407 = 8'h17 == _T_5[7:0] ? image_2_23 : _GEN_406; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_408 = 8'h18 == _T_5[7:0] ? image_2_24 : _GEN_407; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_409 = 8'h19 == _T_5[7:0] ? image_2_25 : _GEN_408; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_410 = 8'h1a == _T_5[7:0] ? image_2_26 : _GEN_409; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_411 = 8'h1b == _T_5[7:0] ? image_2_27 : _GEN_410; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_412 = 8'h1c == _T_5[7:0] ? image_2_28 : _GEN_411; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_413 = 8'h1d == _T_5[7:0] ? image_2_29 : _GEN_412; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_414 = 8'h1e == _T_5[7:0] ? image_2_30 : _GEN_413; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_415 = 8'h1f == _T_5[7:0] ? image_2_31 : _GEN_414; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_416 = 8'h20 == _T_5[7:0] ? image_2_32 : _GEN_415; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_417 = 8'h21 == _T_5[7:0] ? image_2_33 : _GEN_416; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_418 = 8'h22 == _T_5[7:0] ? image_2_34 : _GEN_417; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_419 = 8'h23 == _T_5[7:0] ? image_2_35 : _GEN_418; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_420 = 8'h24 == _T_5[7:0] ? image_2_36 : _GEN_419; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_421 = 8'h25 == _T_5[7:0] ? image_2_37 : _GEN_420; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_422 = 8'h26 == _T_5[7:0] ? image_2_38 : _GEN_421; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_423 = 8'h27 == _T_5[7:0] ? image_2_39 : _GEN_422; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_424 = 8'h28 == _T_5[7:0] ? image_2_40 : _GEN_423; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_425 = 8'h29 == _T_5[7:0] ? image_2_41 : _GEN_424; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_426 = 8'h2a == _T_5[7:0] ? image_2_42 : _GEN_425; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_427 = 8'h2b == _T_5[7:0] ? image_2_43 : _GEN_426; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_428 = 8'h2c == _T_5[7:0] ? image_2_44 : _GEN_427; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_429 = 8'h2d == _T_5[7:0] ? image_2_45 : _GEN_428; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_430 = 8'h2e == _T_5[7:0] ? image_2_46 : _GEN_429; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_431 = 8'h2f == _T_5[7:0] ? image_2_47 : _GEN_430; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_432 = 8'h30 == _T_5[7:0] ? image_2_48 : _GEN_431; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_433 = 8'h31 == _T_5[7:0] ? image_2_49 : _GEN_432; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_434 = 8'h32 == _T_5[7:0] ? image_2_50 : _GEN_433; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_435 = 8'h33 == _T_5[7:0] ? image_2_51 : _GEN_434; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_436 = 8'h34 == _T_5[7:0] ? image_2_52 : _GEN_435; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_437 = 8'h35 == _T_5[7:0] ? image_2_53 : _GEN_436; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_438 = 8'h36 == _T_5[7:0] ? image_2_54 : _GEN_437; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_439 = 8'h37 == _T_5[7:0] ? image_2_55 : _GEN_438; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_440 = 8'h38 == _T_5[7:0] ? image_2_56 : _GEN_439; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_441 = 8'h39 == _T_5[7:0] ? image_2_57 : _GEN_440; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_442 = 8'h3a == _T_5[7:0] ? image_2_58 : _GEN_441; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_443 = 8'h3b == _T_5[7:0] ? image_2_59 : _GEN_442; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_444 = 8'h3c == _T_5[7:0] ? image_2_60 : _GEN_443; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_445 = 8'h3d == _T_5[7:0] ? image_2_61 : _GEN_444; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_446 = 8'h3e == _T_5[7:0] ? image_2_62 : _GEN_445; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_447 = 8'h3f == _T_5[7:0] ? image_2_63 : _GEN_446; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_448 = 8'h40 == _T_5[7:0] ? image_2_64 : _GEN_447; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_449 = 8'h41 == _T_5[7:0] ? image_2_65 : _GEN_448; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_450 = 8'h42 == _T_5[7:0] ? image_2_66 : _GEN_449; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_451 = 8'h43 == _T_5[7:0] ? image_2_67 : _GEN_450; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_452 = 8'h44 == _T_5[7:0] ? image_2_68 : _GEN_451; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_453 = 8'h45 == _T_5[7:0] ? image_2_69 : _GEN_452; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_454 = 8'h46 == _T_5[7:0] ? image_2_70 : _GEN_453; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_455 = 8'h47 == _T_5[7:0] ? image_2_71 : _GEN_454; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_456 = 8'h48 == _T_5[7:0] ? image_2_72 : _GEN_455; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_457 = 8'h49 == _T_5[7:0] ? image_2_73 : _GEN_456; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_458 = 8'h4a == _T_5[7:0] ? image_2_74 : _GEN_457; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_459 = 8'h4b == _T_5[7:0] ? image_2_75 : _GEN_458; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_460 = 8'h4c == _T_5[7:0] ? image_2_76 : _GEN_459; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_461 = 8'h4d == _T_5[7:0] ? image_2_77 : _GEN_460; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_462 = 8'h4e == _T_5[7:0] ? image_2_78 : _GEN_461; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_463 = 8'h4f == _T_5[7:0] ? image_2_79 : _GEN_462; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_464 = 8'h50 == _T_5[7:0] ? image_2_80 : _GEN_463; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_465 = 8'h51 == _T_5[7:0] ? image_2_81 : _GEN_464; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_466 = 8'h52 == _T_5[7:0] ? image_2_82 : _GEN_465; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_467 = 8'h53 == _T_5[7:0] ? image_2_83 : _GEN_466; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_468 = 8'h54 == _T_5[7:0] ? image_2_84 : _GEN_467; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_469 = 8'h55 == _T_5[7:0] ? image_2_85 : _GEN_468; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_470 = 8'h56 == _T_5[7:0] ? image_2_86 : _GEN_469; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_471 = 8'h57 == _T_5[7:0] ? image_2_87 : _GEN_470; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_472 = 8'h58 == _T_5[7:0] ? image_2_88 : _GEN_471; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_473 = 8'h59 == _T_5[7:0] ? image_2_89 : _GEN_472; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_474 = 8'h5a == _T_5[7:0] ? image_2_90 : _GEN_473; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_475 = 8'h5b == _T_5[7:0] ? image_2_91 : _GEN_474; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_476 = 8'h5c == _T_5[7:0] ? image_2_92 : _GEN_475; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_477 = 8'h5d == _T_5[7:0] ? image_2_93 : _GEN_476; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_478 = 8'h5e == _T_5[7:0] ? image_2_94 : _GEN_477; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_479 = 8'h5f == _T_5[7:0] ? image_2_95 : _GEN_478; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_480 = 8'h60 == _T_5[7:0] ? image_2_96 : _GEN_479; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_481 = 8'h61 == _T_5[7:0] ? image_2_97 : _GEN_480; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_482 = 8'h62 == _T_5[7:0] ? image_2_98 : _GEN_481; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_483 = 8'h63 == _T_5[7:0] ? image_2_99 : _GEN_482; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_484 = 8'h64 == _T_5[7:0] ? image_2_100 : _GEN_483; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_485 = 8'h65 == _T_5[7:0] ? image_2_101 : _GEN_484; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_486 = 8'h66 == _T_5[7:0] ? image_2_102 : _GEN_485; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_487 = 8'h67 == _T_5[7:0] ? image_2_103 : _GEN_486; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_488 = 8'h68 == _T_5[7:0] ? image_2_104 : _GEN_487; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_489 = 8'h69 == _T_5[7:0] ? image_2_105 : _GEN_488; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_490 = 8'h6a == _T_5[7:0] ? image_2_106 : _GEN_489; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_491 = 8'h6b == _T_5[7:0] ? image_2_107 : _GEN_490; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_492 = 8'h6c == _T_5[7:0] ? image_2_108 : _GEN_491; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_493 = 8'h6d == _T_5[7:0] ? image_2_109 : _GEN_492; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_494 = 8'h6e == _T_5[7:0] ? image_2_110 : _GEN_493; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_495 = 8'h6f == _T_5[7:0] ? image_2_111 : _GEN_494; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_496 = 8'h70 == _T_5[7:0] ? image_2_112 : _GEN_495; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_497 = 8'h71 == _T_5[7:0] ? image_2_113 : _GEN_496; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_498 = 8'h72 == _T_5[7:0] ? image_2_114 : _GEN_497; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_499 = 8'h73 == _T_5[7:0] ? image_2_115 : _GEN_498; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_500 = 8'h74 == _T_5[7:0] ? image_2_116 : _GEN_499; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_501 = 8'h75 == _T_5[7:0] ? image_2_117 : _GEN_500; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_502 = 8'h76 == _T_5[7:0] ? image_2_118 : _GEN_501; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_503 = 8'h77 == _T_5[7:0] ? image_2_119 : _GEN_502; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_504 = 8'h78 == _T_5[7:0] ? image_2_120 : _GEN_503; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_505 = 8'h79 == _T_5[7:0] ? image_2_121 : _GEN_504; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_506 = 8'h7a == _T_5[7:0] ? image_2_122 : _GEN_505; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_507 = 8'h7b == _T_5[7:0] ? image_2_123 : _GEN_506; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_508 = 8'h7c == _T_5[7:0] ? image_2_124 : _GEN_507; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_509 = 8'h7d == _T_5[7:0] ? image_2_125 : _GEN_508; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_510 = 8'h7e == _T_5[7:0] ? image_2_126 : _GEN_509; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_511 = 8'h7f == _T_5[7:0] ? image_2_127 : _GEN_510; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_512 = 8'h80 == _T_5[7:0] ? image_2_128 : _GEN_511; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_513 = 8'h81 == _T_5[7:0] ? image_2_129 : _GEN_512; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_514 = 8'h82 == _T_5[7:0] ? image_2_130 : _GEN_513; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_515 = 8'h83 == _T_5[7:0] ? image_2_131 : _GEN_514; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_516 = 8'h84 == _T_5[7:0] ? image_2_132 : _GEN_515; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_517 = 8'h85 == _T_5[7:0] ? image_2_133 : _GEN_516; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_518 = 8'h86 == _T_5[7:0] ? image_2_134 : _GEN_517; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_519 = 8'h87 == _T_5[7:0] ? image_2_135 : _GEN_518; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_520 = 8'h88 == _T_5[7:0] ? image_2_136 : _GEN_519; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_521 = 8'h89 == _T_5[7:0] ? image_2_137 : _GEN_520; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_522 = 8'h8a == _T_5[7:0] ? image_2_138 : _GEN_521; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_523 = 8'h8b == _T_5[7:0] ? image_2_139 : _GEN_522; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_524 = 8'h8c == _T_5[7:0] ? image_2_140 : _GEN_523; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_525 = 8'h8d == _T_5[7:0] ? image_2_141 : _GEN_524; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_526 = 8'h8e == _T_5[7:0] ? image_2_142 : _GEN_525; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_527 = 8'h8f == _T_5[7:0] ? image_2_143 : _GEN_526; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_528 = 8'h90 == _T_5[7:0] ? image_2_144 : _GEN_527; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_529 = 8'h91 == _T_5[7:0] ? image_2_145 : _GEN_528; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_530 = 8'h92 == _T_5[7:0] ? image_2_146 : _GEN_529; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_531 = 8'h93 == _T_5[7:0] ? image_2_147 : _GEN_530; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_532 = 8'h94 == _T_5[7:0] ? image_2_148 : _GEN_531; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_533 = 8'h95 == _T_5[7:0] ? image_2_149 : _GEN_532; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_534 = 8'h96 == _T_5[7:0] ? image_2_150 : _GEN_533; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_535 = 8'h97 == _T_5[7:0] ? image_2_151 : _GEN_534; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_536 = 8'h98 == _T_5[7:0] ? image_2_152 : _GEN_535; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_537 = 8'h99 == _T_5[7:0] ? image_2_153 : _GEN_536; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_538 = 8'h9a == _T_5[7:0] ? image_2_154 : _GEN_537; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_539 = 8'h9b == _T_5[7:0] ? image_2_155 : _GEN_538; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_540 = 8'h9c == _T_5[7:0] ? image_2_156 : _GEN_539; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_541 = 8'h9d == _T_5[7:0] ? image_2_157 : _GEN_540; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_542 = 8'h9e == _T_5[7:0] ? image_2_158 : _GEN_541; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_543 = 8'h9f == _T_5[7:0] ? image_2_159 : _GEN_542; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_544 = 8'ha0 == _T_5[7:0] ? image_2_160 : _GEN_543; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_545 = 8'ha1 == _T_5[7:0] ? image_2_161 : _GEN_544; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_546 = 8'ha2 == _T_5[7:0] ? image_2_162 : _GEN_545; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_547 = 8'ha3 == _T_5[7:0] ? image_2_163 : _GEN_546; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_548 = 8'ha4 == _T_5[7:0] ? image_2_164 : _GEN_547; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_549 = 8'ha5 == _T_5[7:0] ? image_2_165 : _GEN_548; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_550 = 8'ha6 == _T_5[7:0] ? image_2_166 : _GEN_549; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_551 = 8'ha7 == _T_5[7:0] ? image_2_167 : _GEN_550; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_552 = 8'ha8 == _T_5[7:0] ? image_2_168 : _GEN_551; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_553 = 8'ha9 == _T_5[7:0] ? image_2_169 : _GEN_552; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_554 = 8'haa == _T_5[7:0] ? image_2_170 : _GEN_553; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_555 = 8'hab == _T_5[7:0] ? image_2_171 : _GEN_554; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_556 = 8'hac == _T_5[7:0] ? image_2_172 : _GEN_555; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_557 = 8'had == _T_5[7:0] ? image_2_173 : _GEN_556; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_558 = 8'hae == _T_5[7:0] ? image_2_174 : _GEN_557; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_559 = 8'haf == _T_5[7:0] ? image_2_175 : _GEN_558; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_560 = 8'hb0 == _T_5[7:0] ? image_2_176 : _GEN_559; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_561 = 8'hb1 == _T_5[7:0] ? image_2_177 : _GEN_560; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_562 = 8'hb2 == _T_5[7:0] ? image_2_178 : _GEN_561; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_563 = 8'hb3 == _T_5[7:0] ? image_2_179 : _GEN_562; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_564 = 8'hb4 == _T_5[7:0] ? image_2_180 : _GEN_563; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_565 = 8'hb5 == _T_5[7:0] ? image_2_181 : _GEN_564; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_566 = 8'hb6 == _T_5[7:0] ? image_2_182 : _GEN_565; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_567 = 8'hb7 == _T_5[7:0] ? image_2_183 : _GEN_566; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_568 = 8'hb8 == _T_5[7:0] ? image_2_184 : _GEN_567; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_569 = 8'hb9 == _T_5[7:0] ? image_2_185 : _GEN_568; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_570 = 8'hba == _T_5[7:0] ? image_2_186 : _GEN_569; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_571 = 8'hbb == _T_5[7:0] ? image_2_187 : _GEN_570; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_572 = 8'hbc == _T_5[7:0] ? image_2_188 : _GEN_571; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_573 = 8'hbd == _T_5[7:0] ? image_2_189 : _GEN_572; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_574 = 8'hbe == _T_5[7:0] ? image_2_190 : _GEN_573; // @[VideoBuffer.scala 27:30]
  wire [32:0] _T_15 = {{1'd0}, pixelIndex}; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_19 = pixelIndex + 32'h1; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_22 = pixelIndex + 32'h2; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_25 = pixelIndex + 32'h3; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_28 = pixelIndex + 32'h4; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_31 = pixelIndex + 32'h5; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_34 = pixelIndex + 32'h6; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_37 = pixelIndex + 32'h7; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_88 = pixelIndex + 32'h8; // @[VideoBuffer.scala 36:34]
  wire [8:0] _T_89 = 5'h10 * 5'hc; // @[VideoBuffer.scala 37:42]
  wire [31:0] _GEN_5765 = {{23'd0}, _T_89}; // @[VideoBuffer.scala 37:25]
  wire  _T_90 = pixelIndex == _GEN_5765; // @[VideoBuffer.scala 37:25]
  assign io_pixelVal_out_0 = 8'hbf == _T_5[7:0] ? image_0_191 : _GEN_190; // @[VideoBuffer.scala 27:30]
  assign io_pixelVal_out_1 = 8'hbf == _T_5[7:0] ? image_1_191 : _GEN_382; // @[VideoBuffer.scala 27:30]
  assign io_pixelVal_out_2 = 8'hbf == _T_5[7:0] ? image_2_191 : _GEN_574; // @[VideoBuffer.scala 27:30]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  image_0_0 = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  image_0_1 = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  image_0_2 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  image_0_3 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  image_0_4 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  image_0_5 = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  image_0_6 = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  image_0_7 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  image_0_8 = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  image_0_9 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  image_0_10 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  image_0_11 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  image_0_12 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  image_0_13 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  image_0_14 = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  image_0_15 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  image_0_16 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  image_0_17 = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  image_0_18 = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  image_0_19 = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  image_0_20 = _RAND_20[3:0];
  _RAND_21 = {1{`RANDOM}};
  image_0_21 = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  image_0_22 = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  image_0_23 = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  image_0_24 = _RAND_24[3:0];
  _RAND_25 = {1{`RANDOM}};
  image_0_25 = _RAND_25[3:0];
  _RAND_26 = {1{`RANDOM}};
  image_0_26 = _RAND_26[3:0];
  _RAND_27 = {1{`RANDOM}};
  image_0_27 = _RAND_27[3:0];
  _RAND_28 = {1{`RANDOM}};
  image_0_28 = _RAND_28[3:0];
  _RAND_29 = {1{`RANDOM}};
  image_0_29 = _RAND_29[3:0];
  _RAND_30 = {1{`RANDOM}};
  image_0_30 = _RAND_30[3:0];
  _RAND_31 = {1{`RANDOM}};
  image_0_31 = _RAND_31[3:0];
  _RAND_32 = {1{`RANDOM}};
  image_0_32 = _RAND_32[3:0];
  _RAND_33 = {1{`RANDOM}};
  image_0_33 = _RAND_33[3:0];
  _RAND_34 = {1{`RANDOM}};
  image_0_34 = _RAND_34[3:0];
  _RAND_35 = {1{`RANDOM}};
  image_0_35 = _RAND_35[3:0];
  _RAND_36 = {1{`RANDOM}};
  image_0_36 = _RAND_36[3:0];
  _RAND_37 = {1{`RANDOM}};
  image_0_37 = _RAND_37[3:0];
  _RAND_38 = {1{`RANDOM}};
  image_0_38 = _RAND_38[3:0];
  _RAND_39 = {1{`RANDOM}};
  image_0_39 = _RAND_39[3:0];
  _RAND_40 = {1{`RANDOM}};
  image_0_40 = _RAND_40[3:0];
  _RAND_41 = {1{`RANDOM}};
  image_0_41 = _RAND_41[3:0];
  _RAND_42 = {1{`RANDOM}};
  image_0_42 = _RAND_42[3:0];
  _RAND_43 = {1{`RANDOM}};
  image_0_43 = _RAND_43[3:0];
  _RAND_44 = {1{`RANDOM}};
  image_0_44 = _RAND_44[3:0];
  _RAND_45 = {1{`RANDOM}};
  image_0_45 = _RAND_45[3:0];
  _RAND_46 = {1{`RANDOM}};
  image_0_46 = _RAND_46[3:0];
  _RAND_47 = {1{`RANDOM}};
  image_0_47 = _RAND_47[3:0];
  _RAND_48 = {1{`RANDOM}};
  image_0_48 = _RAND_48[3:0];
  _RAND_49 = {1{`RANDOM}};
  image_0_49 = _RAND_49[3:0];
  _RAND_50 = {1{`RANDOM}};
  image_0_50 = _RAND_50[3:0];
  _RAND_51 = {1{`RANDOM}};
  image_0_51 = _RAND_51[3:0];
  _RAND_52 = {1{`RANDOM}};
  image_0_52 = _RAND_52[3:0];
  _RAND_53 = {1{`RANDOM}};
  image_0_53 = _RAND_53[3:0];
  _RAND_54 = {1{`RANDOM}};
  image_0_54 = _RAND_54[3:0];
  _RAND_55 = {1{`RANDOM}};
  image_0_55 = _RAND_55[3:0];
  _RAND_56 = {1{`RANDOM}};
  image_0_56 = _RAND_56[3:0];
  _RAND_57 = {1{`RANDOM}};
  image_0_57 = _RAND_57[3:0];
  _RAND_58 = {1{`RANDOM}};
  image_0_58 = _RAND_58[3:0];
  _RAND_59 = {1{`RANDOM}};
  image_0_59 = _RAND_59[3:0];
  _RAND_60 = {1{`RANDOM}};
  image_0_60 = _RAND_60[3:0];
  _RAND_61 = {1{`RANDOM}};
  image_0_61 = _RAND_61[3:0];
  _RAND_62 = {1{`RANDOM}};
  image_0_62 = _RAND_62[3:0];
  _RAND_63 = {1{`RANDOM}};
  image_0_63 = _RAND_63[3:0];
  _RAND_64 = {1{`RANDOM}};
  image_0_64 = _RAND_64[3:0];
  _RAND_65 = {1{`RANDOM}};
  image_0_65 = _RAND_65[3:0];
  _RAND_66 = {1{`RANDOM}};
  image_0_66 = _RAND_66[3:0];
  _RAND_67 = {1{`RANDOM}};
  image_0_67 = _RAND_67[3:0];
  _RAND_68 = {1{`RANDOM}};
  image_0_68 = _RAND_68[3:0];
  _RAND_69 = {1{`RANDOM}};
  image_0_69 = _RAND_69[3:0];
  _RAND_70 = {1{`RANDOM}};
  image_0_70 = _RAND_70[3:0];
  _RAND_71 = {1{`RANDOM}};
  image_0_71 = _RAND_71[3:0];
  _RAND_72 = {1{`RANDOM}};
  image_0_72 = _RAND_72[3:0];
  _RAND_73 = {1{`RANDOM}};
  image_0_73 = _RAND_73[3:0];
  _RAND_74 = {1{`RANDOM}};
  image_0_74 = _RAND_74[3:0];
  _RAND_75 = {1{`RANDOM}};
  image_0_75 = _RAND_75[3:0];
  _RAND_76 = {1{`RANDOM}};
  image_0_76 = _RAND_76[3:0];
  _RAND_77 = {1{`RANDOM}};
  image_0_77 = _RAND_77[3:0];
  _RAND_78 = {1{`RANDOM}};
  image_0_78 = _RAND_78[3:0];
  _RAND_79 = {1{`RANDOM}};
  image_0_79 = _RAND_79[3:0];
  _RAND_80 = {1{`RANDOM}};
  image_0_80 = _RAND_80[3:0];
  _RAND_81 = {1{`RANDOM}};
  image_0_81 = _RAND_81[3:0];
  _RAND_82 = {1{`RANDOM}};
  image_0_82 = _RAND_82[3:0];
  _RAND_83 = {1{`RANDOM}};
  image_0_83 = _RAND_83[3:0];
  _RAND_84 = {1{`RANDOM}};
  image_0_84 = _RAND_84[3:0];
  _RAND_85 = {1{`RANDOM}};
  image_0_85 = _RAND_85[3:0];
  _RAND_86 = {1{`RANDOM}};
  image_0_86 = _RAND_86[3:0];
  _RAND_87 = {1{`RANDOM}};
  image_0_87 = _RAND_87[3:0];
  _RAND_88 = {1{`RANDOM}};
  image_0_88 = _RAND_88[3:0];
  _RAND_89 = {1{`RANDOM}};
  image_0_89 = _RAND_89[3:0];
  _RAND_90 = {1{`RANDOM}};
  image_0_90 = _RAND_90[3:0];
  _RAND_91 = {1{`RANDOM}};
  image_0_91 = _RAND_91[3:0];
  _RAND_92 = {1{`RANDOM}};
  image_0_92 = _RAND_92[3:0];
  _RAND_93 = {1{`RANDOM}};
  image_0_93 = _RAND_93[3:0];
  _RAND_94 = {1{`RANDOM}};
  image_0_94 = _RAND_94[3:0];
  _RAND_95 = {1{`RANDOM}};
  image_0_95 = _RAND_95[3:0];
  _RAND_96 = {1{`RANDOM}};
  image_0_96 = _RAND_96[3:0];
  _RAND_97 = {1{`RANDOM}};
  image_0_97 = _RAND_97[3:0];
  _RAND_98 = {1{`RANDOM}};
  image_0_98 = _RAND_98[3:0];
  _RAND_99 = {1{`RANDOM}};
  image_0_99 = _RAND_99[3:0];
  _RAND_100 = {1{`RANDOM}};
  image_0_100 = _RAND_100[3:0];
  _RAND_101 = {1{`RANDOM}};
  image_0_101 = _RAND_101[3:0];
  _RAND_102 = {1{`RANDOM}};
  image_0_102 = _RAND_102[3:0];
  _RAND_103 = {1{`RANDOM}};
  image_0_103 = _RAND_103[3:0];
  _RAND_104 = {1{`RANDOM}};
  image_0_104 = _RAND_104[3:0];
  _RAND_105 = {1{`RANDOM}};
  image_0_105 = _RAND_105[3:0];
  _RAND_106 = {1{`RANDOM}};
  image_0_106 = _RAND_106[3:0];
  _RAND_107 = {1{`RANDOM}};
  image_0_107 = _RAND_107[3:0];
  _RAND_108 = {1{`RANDOM}};
  image_0_108 = _RAND_108[3:0];
  _RAND_109 = {1{`RANDOM}};
  image_0_109 = _RAND_109[3:0];
  _RAND_110 = {1{`RANDOM}};
  image_0_110 = _RAND_110[3:0];
  _RAND_111 = {1{`RANDOM}};
  image_0_111 = _RAND_111[3:0];
  _RAND_112 = {1{`RANDOM}};
  image_0_112 = _RAND_112[3:0];
  _RAND_113 = {1{`RANDOM}};
  image_0_113 = _RAND_113[3:0];
  _RAND_114 = {1{`RANDOM}};
  image_0_114 = _RAND_114[3:0];
  _RAND_115 = {1{`RANDOM}};
  image_0_115 = _RAND_115[3:0];
  _RAND_116 = {1{`RANDOM}};
  image_0_116 = _RAND_116[3:0];
  _RAND_117 = {1{`RANDOM}};
  image_0_117 = _RAND_117[3:0];
  _RAND_118 = {1{`RANDOM}};
  image_0_118 = _RAND_118[3:0];
  _RAND_119 = {1{`RANDOM}};
  image_0_119 = _RAND_119[3:0];
  _RAND_120 = {1{`RANDOM}};
  image_0_120 = _RAND_120[3:0];
  _RAND_121 = {1{`RANDOM}};
  image_0_121 = _RAND_121[3:0];
  _RAND_122 = {1{`RANDOM}};
  image_0_122 = _RAND_122[3:0];
  _RAND_123 = {1{`RANDOM}};
  image_0_123 = _RAND_123[3:0];
  _RAND_124 = {1{`RANDOM}};
  image_0_124 = _RAND_124[3:0];
  _RAND_125 = {1{`RANDOM}};
  image_0_125 = _RAND_125[3:0];
  _RAND_126 = {1{`RANDOM}};
  image_0_126 = _RAND_126[3:0];
  _RAND_127 = {1{`RANDOM}};
  image_0_127 = _RAND_127[3:0];
  _RAND_128 = {1{`RANDOM}};
  image_0_128 = _RAND_128[3:0];
  _RAND_129 = {1{`RANDOM}};
  image_0_129 = _RAND_129[3:0];
  _RAND_130 = {1{`RANDOM}};
  image_0_130 = _RAND_130[3:0];
  _RAND_131 = {1{`RANDOM}};
  image_0_131 = _RAND_131[3:0];
  _RAND_132 = {1{`RANDOM}};
  image_0_132 = _RAND_132[3:0];
  _RAND_133 = {1{`RANDOM}};
  image_0_133 = _RAND_133[3:0];
  _RAND_134 = {1{`RANDOM}};
  image_0_134 = _RAND_134[3:0];
  _RAND_135 = {1{`RANDOM}};
  image_0_135 = _RAND_135[3:0];
  _RAND_136 = {1{`RANDOM}};
  image_0_136 = _RAND_136[3:0];
  _RAND_137 = {1{`RANDOM}};
  image_0_137 = _RAND_137[3:0];
  _RAND_138 = {1{`RANDOM}};
  image_0_138 = _RAND_138[3:0];
  _RAND_139 = {1{`RANDOM}};
  image_0_139 = _RAND_139[3:0];
  _RAND_140 = {1{`RANDOM}};
  image_0_140 = _RAND_140[3:0];
  _RAND_141 = {1{`RANDOM}};
  image_0_141 = _RAND_141[3:0];
  _RAND_142 = {1{`RANDOM}};
  image_0_142 = _RAND_142[3:0];
  _RAND_143 = {1{`RANDOM}};
  image_0_143 = _RAND_143[3:0];
  _RAND_144 = {1{`RANDOM}};
  image_0_144 = _RAND_144[3:0];
  _RAND_145 = {1{`RANDOM}};
  image_0_145 = _RAND_145[3:0];
  _RAND_146 = {1{`RANDOM}};
  image_0_146 = _RAND_146[3:0];
  _RAND_147 = {1{`RANDOM}};
  image_0_147 = _RAND_147[3:0];
  _RAND_148 = {1{`RANDOM}};
  image_0_148 = _RAND_148[3:0];
  _RAND_149 = {1{`RANDOM}};
  image_0_149 = _RAND_149[3:0];
  _RAND_150 = {1{`RANDOM}};
  image_0_150 = _RAND_150[3:0];
  _RAND_151 = {1{`RANDOM}};
  image_0_151 = _RAND_151[3:0];
  _RAND_152 = {1{`RANDOM}};
  image_0_152 = _RAND_152[3:0];
  _RAND_153 = {1{`RANDOM}};
  image_0_153 = _RAND_153[3:0];
  _RAND_154 = {1{`RANDOM}};
  image_0_154 = _RAND_154[3:0];
  _RAND_155 = {1{`RANDOM}};
  image_0_155 = _RAND_155[3:0];
  _RAND_156 = {1{`RANDOM}};
  image_0_156 = _RAND_156[3:0];
  _RAND_157 = {1{`RANDOM}};
  image_0_157 = _RAND_157[3:0];
  _RAND_158 = {1{`RANDOM}};
  image_0_158 = _RAND_158[3:0];
  _RAND_159 = {1{`RANDOM}};
  image_0_159 = _RAND_159[3:0];
  _RAND_160 = {1{`RANDOM}};
  image_0_160 = _RAND_160[3:0];
  _RAND_161 = {1{`RANDOM}};
  image_0_161 = _RAND_161[3:0];
  _RAND_162 = {1{`RANDOM}};
  image_0_162 = _RAND_162[3:0];
  _RAND_163 = {1{`RANDOM}};
  image_0_163 = _RAND_163[3:0];
  _RAND_164 = {1{`RANDOM}};
  image_0_164 = _RAND_164[3:0];
  _RAND_165 = {1{`RANDOM}};
  image_0_165 = _RAND_165[3:0];
  _RAND_166 = {1{`RANDOM}};
  image_0_166 = _RAND_166[3:0];
  _RAND_167 = {1{`RANDOM}};
  image_0_167 = _RAND_167[3:0];
  _RAND_168 = {1{`RANDOM}};
  image_0_168 = _RAND_168[3:0];
  _RAND_169 = {1{`RANDOM}};
  image_0_169 = _RAND_169[3:0];
  _RAND_170 = {1{`RANDOM}};
  image_0_170 = _RAND_170[3:0];
  _RAND_171 = {1{`RANDOM}};
  image_0_171 = _RAND_171[3:0];
  _RAND_172 = {1{`RANDOM}};
  image_0_172 = _RAND_172[3:0];
  _RAND_173 = {1{`RANDOM}};
  image_0_173 = _RAND_173[3:0];
  _RAND_174 = {1{`RANDOM}};
  image_0_174 = _RAND_174[3:0];
  _RAND_175 = {1{`RANDOM}};
  image_0_175 = _RAND_175[3:0];
  _RAND_176 = {1{`RANDOM}};
  image_0_176 = _RAND_176[3:0];
  _RAND_177 = {1{`RANDOM}};
  image_0_177 = _RAND_177[3:0];
  _RAND_178 = {1{`RANDOM}};
  image_0_178 = _RAND_178[3:0];
  _RAND_179 = {1{`RANDOM}};
  image_0_179 = _RAND_179[3:0];
  _RAND_180 = {1{`RANDOM}};
  image_0_180 = _RAND_180[3:0];
  _RAND_181 = {1{`RANDOM}};
  image_0_181 = _RAND_181[3:0];
  _RAND_182 = {1{`RANDOM}};
  image_0_182 = _RAND_182[3:0];
  _RAND_183 = {1{`RANDOM}};
  image_0_183 = _RAND_183[3:0];
  _RAND_184 = {1{`RANDOM}};
  image_0_184 = _RAND_184[3:0];
  _RAND_185 = {1{`RANDOM}};
  image_0_185 = _RAND_185[3:0];
  _RAND_186 = {1{`RANDOM}};
  image_0_186 = _RAND_186[3:0];
  _RAND_187 = {1{`RANDOM}};
  image_0_187 = _RAND_187[3:0];
  _RAND_188 = {1{`RANDOM}};
  image_0_188 = _RAND_188[3:0];
  _RAND_189 = {1{`RANDOM}};
  image_0_189 = _RAND_189[3:0];
  _RAND_190 = {1{`RANDOM}};
  image_0_190 = _RAND_190[3:0];
  _RAND_191 = {1{`RANDOM}};
  image_0_191 = _RAND_191[3:0];
  _RAND_192 = {1{`RANDOM}};
  image_1_0 = _RAND_192[3:0];
  _RAND_193 = {1{`RANDOM}};
  image_1_1 = _RAND_193[3:0];
  _RAND_194 = {1{`RANDOM}};
  image_1_2 = _RAND_194[3:0];
  _RAND_195 = {1{`RANDOM}};
  image_1_3 = _RAND_195[3:0];
  _RAND_196 = {1{`RANDOM}};
  image_1_4 = _RAND_196[3:0];
  _RAND_197 = {1{`RANDOM}};
  image_1_5 = _RAND_197[3:0];
  _RAND_198 = {1{`RANDOM}};
  image_1_6 = _RAND_198[3:0];
  _RAND_199 = {1{`RANDOM}};
  image_1_7 = _RAND_199[3:0];
  _RAND_200 = {1{`RANDOM}};
  image_1_8 = _RAND_200[3:0];
  _RAND_201 = {1{`RANDOM}};
  image_1_9 = _RAND_201[3:0];
  _RAND_202 = {1{`RANDOM}};
  image_1_10 = _RAND_202[3:0];
  _RAND_203 = {1{`RANDOM}};
  image_1_11 = _RAND_203[3:0];
  _RAND_204 = {1{`RANDOM}};
  image_1_12 = _RAND_204[3:0];
  _RAND_205 = {1{`RANDOM}};
  image_1_13 = _RAND_205[3:0];
  _RAND_206 = {1{`RANDOM}};
  image_1_14 = _RAND_206[3:0];
  _RAND_207 = {1{`RANDOM}};
  image_1_15 = _RAND_207[3:0];
  _RAND_208 = {1{`RANDOM}};
  image_1_16 = _RAND_208[3:0];
  _RAND_209 = {1{`RANDOM}};
  image_1_17 = _RAND_209[3:0];
  _RAND_210 = {1{`RANDOM}};
  image_1_18 = _RAND_210[3:0];
  _RAND_211 = {1{`RANDOM}};
  image_1_19 = _RAND_211[3:0];
  _RAND_212 = {1{`RANDOM}};
  image_1_20 = _RAND_212[3:0];
  _RAND_213 = {1{`RANDOM}};
  image_1_21 = _RAND_213[3:0];
  _RAND_214 = {1{`RANDOM}};
  image_1_22 = _RAND_214[3:0];
  _RAND_215 = {1{`RANDOM}};
  image_1_23 = _RAND_215[3:0];
  _RAND_216 = {1{`RANDOM}};
  image_1_24 = _RAND_216[3:0];
  _RAND_217 = {1{`RANDOM}};
  image_1_25 = _RAND_217[3:0];
  _RAND_218 = {1{`RANDOM}};
  image_1_26 = _RAND_218[3:0];
  _RAND_219 = {1{`RANDOM}};
  image_1_27 = _RAND_219[3:0];
  _RAND_220 = {1{`RANDOM}};
  image_1_28 = _RAND_220[3:0];
  _RAND_221 = {1{`RANDOM}};
  image_1_29 = _RAND_221[3:0];
  _RAND_222 = {1{`RANDOM}};
  image_1_30 = _RAND_222[3:0];
  _RAND_223 = {1{`RANDOM}};
  image_1_31 = _RAND_223[3:0];
  _RAND_224 = {1{`RANDOM}};
  image_1_32 = _RAND_224[3:0];
  _RAND_225 = {1{`RANDOM}};
  image_1_33 = _RAND_225[3:0];
  _RAND_226 = {1{`RANDOM}};
  image_1_34 = _RAND_226[3:0];
  _RAND_227 = {1{`RANDOM}};
  image_1_35 = _RAND_227[3:0];
  _RAND_228 = {1{`RANDOM}};
  image_1_36 = _RAND_228[3:0];
  _RAND_229 = {1{`RANDOM}};
  image_1_37 = _RAND_229[3:0];
  _RAND_230 = {1{`RANDOM}};
  image_1_38 = _RAND_230[3:0];
  _RAND_231 = {1{`RANDOM}};
  image_1_39 = _RAND_231[3:0];
  _RAND_232 = {1{`RANDOM}};
  image_1_40 = _RAND_232[3:0];
  _RAND_233 = {1{`RANDOM}};
  image_1_41 = _RAND_233[3:0];
  _RAND_234 = {1{`RANDOM}};
  image_1_42 = _RAND_234[3:0];
  _RAND_235 = {1{`RANDOM}};
  image_1_43 = _RAND_235[3:0];
  _RAND_236 = {1{`RANDOM}};
  image_1_44 = _RAND_236[3:0];
  _RAND_237 = {1{`RANDOM}};
  image_1_45 = _RAND_237[3:0];
  _RAND_238 = {1{`RANDOM}};
  image_1_46 = _RAND_238[3:0];
  _RAND_239 = {1{`RANDOM}};
  image_1_47 = _RAND_239[3:0];
  _RAND_240 = {1{`RANDOM}};
  image_1_48 = _RAND_240[3:0];
  _RAND_241 = {1{`RANDOM}};
  image_1_49 = _RAND_241[3:0];
  _RAND_242 = {1{`RANDOM}};
  image_1_50 = _RAND_242[3:0];
  _RAND_243 = {1{`RANDOM}};
  image_1_51 = _RAND_243[3:0];
  _RAND_244 = {1{`RANDOM}};
  image_1_52 = _RAND_244[3:0];
  _RAND_245 = {1{`RANDOM}};
  image_1_53 = _RAND_245[3:0];
  _RAND_246 = {1{`RANDOM}};
  image_1_54 = _RAND_246[3:0];
  _RAND_247 = {1{`RANDOM}};
  image_1_55 = _RAND_247[3:0];
  _RAND_248 = {1{`RANDOM}};
  image_1_56 = _RAND_248[3:0];
  _RAND_249 = {1{`RANDOM}};
  image_1_57 = _RAND_249[3:0];
  _RAND_250 = {1{`RANDOM}};
  image_1_58 = _RAND_250[3:0];
  _RAND_251 = {1{`RANDOM}};
  image_1_59 = _RAND_251[3:0];
  _RAND_252 = {1{`RANDOM}};
  image_1_60 = _RAND_252[3:0];
  _RAND_253 = {1{`RANDOM}};
  image_1_61 = _RAND_253[3:0];
  _RAND_254 = {1{`RANDOM}};
  image_1_62 = _RAND_254[3:0];
  _RAND_255 = {1{`RANDOM}};
  image_1_63 = _RAND_255[3:0];
  _RAND_256 = {1{`RANDOM}};
  image_1_64 = _RAND_256[3:0];
  _RAND_257 = {1{`RANDOM}};
  image_1_65 = _RAND_257[3:0];
  _RAND_258 = {1{`RANDOM}};
  image_1_66 = _RAND_258[3:0];
  _RAND_259 = {1{`RANDOM}};
  image_1_67 = _RAND_259[3:0];
  _RAND_260 = {1{`RANDOM}};
  image_1_68 = _RAND_260[3:0];
  _RAND_261 = {1{`RANDOM}};
  image_1_69 = _RAND_261[3:0];
  _RAND_262 = {1{`RANDOM}};
  image_1_70 = _RAND_262[3:0];
  _RAND_263 = {1{`RANDOM}};
  image_1_71 = _RAND_263[3:0];
  _RAND_264 = {1{`RANDOM}};
  image_1_72 = _RAND_264[3:0];
  _RAND_265 = {1{`RANDOM}};
  image_1_73 = _RAND_265[3:0];
  _RAND_266 = {1{`RANDOM}};
  image_1_74 = _RAND_266[3:0];
  _RAND_267 = {1{`RANDOM}};
  image_1_75 = _RAND_267[3:0];
  _RAND_268 = {1{`RANDOM}};
  image_1_76 = _RAND_268[3:0];
  _RAND_269 = {1{`RANDOM}};
  image_1_77 = _RAND_269[3:0];
  _RAND_270 = {1{`RANDOM}};
  image_1_78 = _RAND_270[3:0];
  _RAND_271 = {1{`RANDOM}};
  image_1_79 = _RAND_271[3:0];
  _RAND_272 = {1{`RANDOM}};
  image_1_80 = _RAND_272[3:0];
  _RAND_273 = {1{`RANDOM}};
  image_1_81 = _RAND_273[3:0];
  _RAND_274 = {1{`RANDOM}};
  image_1_82 = _RAND_274[3:0];
  _RAND_275 = {1{`RANDOM}};
  image_1_83 = _RAND_275[3:0];
  _RAND_276 = {1{`RANDOM}};
  image_1_84 = _RAND_276[3:0];
  _RAND_277 = {1{`RANDOM}};
  image_1_85 = _RAND_277[3:0];
  _RAND_278 = {1{`RANDOM}};
  image_1_86 = _RAND_278[3:0];
  _RAND_279 = {1{`RANDOM}};
  image_1_87 = _RAND_279[3:0];
  _RAND_280 = {1{`RANDOM}};
  image_1_88 = _RAND_280[3:0];
  _RAND_281 = {1{`RANDOM}};
  image_1_89 = _RAND_281[3:0];
  _RAND_282 = {1{`RANDOM}};
  image_1_90 = _RAND_282[3:0];
  _RAND_283 = {1{`RANDOM}};
  image_1_91 = _RAND_283[3:0];
  _RAND_284 = {1{`RANDOM}};
  image_1_92 = _RAND_284[3:0];
  _RAND_285 = {1{`RANDOM}};
  image_1_93 = _RAND_285[3:0];
  _RAND_286 = {1{`RANDOM}};
  image_1_94 = _RAND_286[3:0];
  _RAND_287 = {1{`RANDOM}};
  image_1_95 = _RAND_287[3:0];
  _RAND_288 = {1{`RANDOM}};
  image_1_96 = _RAND_288[3:0];
  _RAND_289 = {1{`RANDOM}};
  image_1_97 = _RAND_289[3:0];
  _RAND_290 = {1{`RANDOM}};
  image_1_98 = _RAND_290[3:0];
  _RAND_291 = {1{`RANDOM}};
  image_1_99 = _RAND_291[3:0];
  _RAND_292 = {1{`RANDOM}};
  image_1_100 = _RAND_292[3:0];
  _RAND_293 = {1{`RANDOM}};
  image_1_101 = _RAND_293[3:0];
  _RAND_294 = {1{`RANDOM}};
  image_1_102 = _RAND_294[3:0];
  _RAND_295 = {1{`RANDOM}};
  image_1_103 = _RAND_295[3:0];
  _RAND_296 = {1{`RANDOM}};
  image_1_104 = _RAND_296[3:0];
  _RAND_297 = {1{`RANDOM}};
  image_1_105 = _RAND_297[3:0];
  _RAND_298 = {1{`RANDOM}};
  image_1_106 = _RAND_298[3:0];
  _RAND_299 = {1{`RANDOM}};
  image_1_107 = _RAND_299[3:0];
  _RAND_300 = {1{`RANDOM}};
  image_1_108 = _RAND_300[3:0];
  _RAND_301 = {1{`RANDOM}};
  image_1_109 = _RAND_301[3:0];
  _RAND_302 = {1{`RANDOM}};
  image_1_110 = _RAND_302[3:0];
  _RAND_303 = {1{`RANDOM}};
  image_1_111 = _RAND_303[3:0];
  _RAND_304 = {1{`RANDOM}};
  image_1_112 = _RAND_304[3:0];
  _RAND_305 = {1{`RANDOM}};
  image_1_113 = _RAND_305[3:0];
  _RAND_306 = {1{`RANDOM}};
  image_1_114 = _RAND_306[3:0];
  _RAND_307 = {1{`RANDOM}};
  image_1_115 = _RAND_307[3:0];
  _RAND_308 = {1{`RANDOM}};
  image_1_116 = _RAND_308[3:0];
  _RAND_309 = {1{`RANDOM}};
  image_1_117 = _RAND_309[3:0];
  _RAND_310 = {1{`RANDOM}};
  image_1_118 = _RAND_310[3:0];
  _RAND_311 = {1{`RANDOM}};
  image_1_119 = _RAND_311[3:0];
  _RAND_312 = {1{`RANDOM}};
  image_1_120 = _RAND_312[3:0];
  _RAND_313 = {1{`RANDOM}};
  image_1_121 = _RAND_313[3:0];
  _RAND_314 = {1{`RANDOM}};
  image_1_122 = _RAND_314[3:0];
  _RAND_315 = {1{`RANDOM}};
  image_1_123 = _RAND_315[3:0];
  _RAND_316 = {1{`RANDOM}};
  image_1_124 = _RAND_316[3:0];
  _RAND_317 = {1{`RANDOM}};
  image_1_125 = _RAND_317[3:0];
  _RAND_318 = {1{`RANDOM}};
  image_1_126 = _RAND_318[3:0];
  _RAND_319 = {1{`RANDOM}};
  image_1_127 = _RAND_319[3:0];
  _RAND_320 = {1{`RANDOM}};
  image_1_128 = _RAND_320[3:0];
  _RAND_321 = {1{`RANDOM}};
  image_1_129 = _RAND_321[3:0];
  _RAND_322 = {1{`RANDOM}};
  image_1_130 = _RAND_322[3:0];
  _RAND_323 = {1{`RANDOM}};
  image_1_131 = _RAND_323[3:0];
  _RAND_324 = {1{`RANDOM}};
  image_1_132 = _RAND_324[3:0];
  _RAND_325 = {1{`RANDOM}};
  image_1_133 = _RAND_325[3:0];
  _RAND_326 = {1{`RANDOM}};
  image_1_134 = _RAND_326[3:0];
  _RAND_327 = {1{`RANDOM}};
  image_1_135 = _RAND_327[3:0];
  _RAND_328 = {1{`RANDOM}};
  image_1_136 = _RAND_328[3:0];
  _RAND_329 = {1{`RANDOM}};
  image_1_137 = _RAND_329[3:0];
  _RAND_330 = {1{`RANDOM}};
  image_1_138 = _RAND_330[3:0];
  _RAND_331 = {1{`RANDOM}};
  image_1_139 = _RAND_331[3:0];
  _RAND_332 = {1{`RANDOM}};
  image_1_140 = _RAND_332[3:0];
  _RAND_333 = {1{`RANDOM}};
  image_1_141 = _RAND_333[3:0];
  _RAND_334 = {1{`RANDOM}};
  image_1_142 = _RAND_334[3:0];
  _RAND_335 = {1{`RANDOM}};
  image_1_143 = _RAND_335[3:0];
  _RAND_336 = {1{`RANDOM}};
  image_1_144 = _RAND_336[3:0];
  _RAND_337 = {1{`RANDOM}};
  image_1_145 = _RAND_337[3:0];
  _RAND_338 = {1{`RANDOM}};
  image_1_146 = _RAND_338[3:0];
  _RAND_339 = {1{`RANDOM}};
  image_1_147 = _RAND_339[3:0];
  _RAND_340 = {1{`RANDOM}};
  image_1_148 = _RAND_340[3:0];
  _RAND_341 = {1{`RANDOM}};
  image_1_149 = _RAND_341[3:0];
  _RAND_342 = {1{`RANDOM}};
  image_1_150 = _RAND_342[3:0];
  _RAND_343 = {1{`RANDOM}};
  image_1_151 = _RAND_343[3:0];
  _RAND_344 = {1{`RANDOM}};
  image_1_152 = _RAND_344[3:0];
  _RAND_345 = {1{`RANDOM}};
  image_1_153 = _RAND_345[3:0];
  _RAND_346 = {1{`RANDOM}};
  image_1_154 = _RAND_346[3:0];
  _RAND_347 = {1{`RANDOM}};
  image_1_155 = _RAND_347[3:0];
  _RAND_348 = {1{`RANDOM}};
  image_1_156 = _RAND_348[3:0];
  _RAND_349 = {1{`RANDOM}};
  image_1_157 = _RAND_349[3:0];
  _RAND_350 = {1{`RANDOM}};
  image_1_158 = _RAND_350[3:0];
  _RAND_351 = {1{`RANDOM}};
  image_1_159 = _RAND_351[3:0];
  _RAND_352 = {1{`RANDOM}};
  image_1_160 = _RAND_352[3:0];
  _RAND_353 = {1{`RANDOM}};
  image_1_161 = _RAND_353[3:0];
  _RAND_354 = {1{`RANDOM}};
  image_1_162 = _RAND_354[3:0];
  _RAND_355 = {1{`RANDOM}};
  image_1_163 = _RAND_355[3:0];
  _RAND_356 = {1{`RANDOM}};
  image_1_164 = _RAND_356[3:0];
  _RAND_357 = {1{`RANDOM}};
  image_1_165 = _RAND_357[3:0];
  _RAND_358 = {1{`RANDOM}};
  image_1_166 = _RAND_358[3:0];
  _RAND_359 = {1{`RANDOM}};
  image_1_167 = _RAND_359[3:0];
  _RAND_360 = {1{`RANDOM}};
  image_1_168 = _RAND_360[3:0];
  _RAND_361 = {1{`RANDOM}};
  image_1_169 = _RAND_361[3:0];
  _RAND_362 = {1{`RANDOM}};
  image_1_170 = _RAND_362[3:0];
  _RAND_363 = {1{`RANDOM}};
  image_1_171 = _RAND_363[3:0];
  _RAND_364 = {1{`RANDOM}};
  image_1_172 = _RAND_364[3:0];
  _RAND_365 = {1{`RANDOM}};
  image_1_173 = _RAND_365[3:0];
  _RAND_366 = {1{`RANDOM}};
  image_1_174 = _RAND_366[3:0];
  _RAND_367 = {1{`RANDOM}};
  image_1_175 = _RAND_367[3:0];
  _RAND_368 = {1{`RANDOM}};
  image_1_176 = _RAND_368[3:0];
  _RAND_369 = {1{`RANDOM}};
  image_1_177 = _RAND_369[3:0];
  _RAND_370 = {1{`RANDOM}};
  image_1_178 = _RAND_370[3:0];
  _RAND_371 = {1{`RANDOM}};
  image_1_179 = _RAND_371[3:0];
  _RAND_372 = {1{`RANDOM}};
  image_1_180 = _RAND_372[3:0];
  _RAND_373 = {1{`RANDOM}};
  image_1_181 = _RAND_373[3:0];
  _RAND_374 = {1{`RANDOM}};
  image_1_182 = _RAND_374[3:0];
  _RAND_375 = {1{`RANDOM}};
  image_1_183 = _RAND_375[3:0];
  _RAND_376 = {1{`RANDOM}};
  image_1_184 = _RAND_376[3:0];
  _RAND_377 = {1{`RANDOM}};
  image_1_185 = _RAND_377[3:0];
  _RAND_378 = {1{`RANDOM}};
  image_1_186 = _RAND_378[3:0];
  _RAND_379 = {1{`RANDOM}};
  image_1_187 = _RAND_379[3:0];
  _RAND_380 = {1{`RANDOM}};
  image_1_188 = _RAND_380[3:0];
  _RAND_381 = {1{`RANDOM}};
  image_1_189 = _RAND_381[3:0];
  _RAND_382 = {1{`RANDOM}};
  image_1_190 = _RAND_382[3:0];
  _RAND_383 = {1{`RANDOM}};
  image_1_191 = _RAND_383[3:0];
  _RAND_384 = {1{`RANDOM}};
  image_2_0 = _RAND_384[3:0];
  _RAND_385 = {1{`RANDOM}};
  image_2_1 = _RAND_385[3:0];
  _RAND_386 = {1{`RANDOM}};
  image_2_2 = _RAND_386[3:0];
  _RAND_387 = {1{`RANDOM}};
  image_2_3 = _RAND_387[3:0];
  _RAND_388 = {1{`RANDOM}};
  image_2_4 = _RAND_388[3:0];
  _RAND_389 = {1{`RANDOM}};
  image_2_5 = _RAND_389[3:0];
  _RAND_390 = {1{`RANDOM}};
  image_2_6 = _RAND_390[3:0];
  _RAND_391 = {1{`RANDOM}};
  image_2_7 = _RAND_391[3:0];
  _RAND_392 = {1{`RANDOM}};
  image_2_8 = _RAND_392[3:0];
  _RAND_393 = {1{`RANDOM}};
  image_2_9 = _RAND_393[3:0];
  _RAND_394 = {1{`RANDOM}};
  image_2_10 = _RAND_394[3:0];
  _RAND_395 = {1{`RANDOM}};
  image_2_11 = _RAND_395[3:0];
  _RAND_396 = {1{`RANDOM}};
  image_2_12 = _RAND_396[3:0];
  _RAND_397 = {1{`RANDOM}};
  image_2_13 = _RAND_397[3:0];
  _RAND_398 = {1{`RANDOM}};
  image_2_14 = _RAND_398[3:0];
  _RAND_399 = {1{`RANDOM}};
  image_2_15 = _RAND_399[3:0];
  _RAND_400 = {1{`RANDOM}};
  image_2_16 = _RAND_400[3:0];
  _RAND_401 = {1{`RANDOM}};
  image_2_17 = _RAND_401[3:0];
  _RAND_402 = {1{`RANDOM}};
  image_2_18 = _RAND_402[3:0];
  _RAND_403 = {1{`RANDOM}};
  image_2_19 = _RAND_403[3:0];
  _RAND_404 = {1{`RANDOM}};
  image_2_20 = _RAND_404[3:0];
  _RAND_405 = {1{`RANDOM}};
  image_2_21 = _RAND_405[3:0];
  _RAND_406 = {1{`RANDOM}};
  image_2_22 = _RAND_406[3:0];
  _RAND_407 = {1{`RANDOM}};
  image_2_23 = _RAND_407[3:0];
  _RAND_408 = {1{`RANDOM}};
  image_2_24 = _RAND_408[3:0];
  _RAND_409 = {1{`RANDOM}};
  image_2_25 = _RAND_409[3:0];
  _RAND_410 = {1{`RANDOM}};
  image_2_26 = _RAND_410[3:0];
  _RAND_411 = {1{`RANDOM}};
  image_2_27 = _RAND_411[3:0];
  _RAND_412 = {1{`RANDOM}};
  image_2_28 = _RAND_412[3:0];
  _RAND_413 = {1{`RANDOM}};
  image_2_29 = _RAND_413[3:0];
  _RAND_414 = {1{`RANDOM}};
  image_2_30 = _RAND_414[3:0];
  _RAND_415 = {1{`RANDOM}};
  image_2_31 = _RAND_415[3:0];
  _RAND_416 = {1{`RANDOM}};
  image_2_32 = _RAND_416[3:0];
  _RAND_417 = {1{`RANDOM}};
  image_2_33 = _RAND_417[3:0];
  _RAND_418 = {1{`RANDOM}};
  image_2_34 = _RAND_418[3:0];
  _RAND_419 = {1{`RANDOM}};
  image_2_35 = _RAND_419[3:0];
  _RAND_420 = {1{`RANDOM}};
  image_2_36 = _RAND_420[3:0];
  _RAND_421 = {1{`RANDOM}};
  image_2_37 = _RAND_421[3:0];
  _RAND_422 = {1{`RANDOM}};
  image_2_38 = _RAND_422[3:0];
  _RAND_423 = {1{`RANDOM}};
  image_2_39 = _RAND_423[3:0];
  _RAND_424 = {1{`RANDOM}};
  image_2_40 = _RAND_424[3:0];
  _RAND_425 = {1{`RANDOM}};
  image_2_41 = _RAND_425[3:0];
  _RAND_426 = {1{`RANDOM}};
  image_2_42 = _RAND_426[3:0];
  _RAND_427 = {1{`RANDOM}};
  image_2_43 = _RAND_427[3:0];
  _RAND_428 = {1{`RANDOM}};
  image_2_44 = _RAND_428[3:0];
  _RAND_429 = {1{`RANDOM}};
  image_2_45 = _RAND_429[3:0];
  _RAND_430 = {1{`RANDOM}};
  image_2_46 = _RAND_430[3:0];
  _RAND_431 = {1{`RANDOM}};
  image_2_47 = _RAND_431[3:0];
  _RAND_432 = {1{`RANDOM}};
  image_2_48 = _RAND_432[3:0];
  _RAND_433 = {1{`RANDOM}};
  image_2_49 = _RAND_433[3:0];
  _RAND_434 = {1{`RANDOM}};
  image_2_50 = _RAND_434[3:0];
  _RAND_435 = {1{`RANDOM}};
  image_2_51 = _RAND_435[3:0];
  _RAND_436 = {1{`RANDOM}};
  image_2_52 = _RAND_436[3:0];
  _RAND_437 = {1{`RANDOM}};
  image_2_53 = _RAND_437[3:0];
  _RAND_438 = {1{`RANDOM}};
  image_2_54 = _RAND_438[3:0];
  _RAND_439 = {1{`RANDOM}};
  image_2_55 = _RAND_439[3:0];
  _RAND_440 = {1{`RANDOM}};
  image_2_56 = _RAND_440[3:0];
  _RAND_441 = {1{`RANDOM}};
  image_2_57 = _RAND_441[3:0];
  _RAND_442 = {1{`RANDOM}};
  image_2_58 = _RAND_442[3:0];
  _RAND_443 = {1{`RANDOM}};
  image_2_59 = _RAND_443[3:0];
  _RAND_444 = {1{`RANDOM}};
  image_2_60 = _RAND_444[3:0];
  _RAND_445 = {1{`RANDOM}};
  image_2_61 = _RAND_445[3:0];
  _RAND_446 = {1{`RANDOM}};
  image_2_62 = _RAND_446[3:0];
  _RAND_447 = {1{`RANDOM}};
  image_2_63 = _RAND_447[3:0];
  _RAND_448 = {1{`RANDOM}};
  image_2_64 = _RAND_448[3:0];
  _RAND_449 = {1{`RANDOM}};
  image_2_65 = _RAND_449[3:0];
  _RAND_450 = {1{`RANDOM}};
  image_2_66 = _RAND_450[3:0];
  _RAND_451 = {1{`RANDOM}};
  image_2_67 = _RAND_451[3:0];
  _RAND_452 = {1{`RANDOM}};
  image_2_68 = _RAND_452[3:0];
  _RAND_453 = {1{`RANDOM}};
  image_2_69 = _RAND_453[3:0];
  _RAND_454 = {1{`RANDOM}};
  image_2_70 = _RAND_454[3:0];
  _RAND_455 = {1{`RANDOM}};
  image_2_71 = _RAND_455[3:0];
  _RAND_456 = {1{`RANDOM}};
  image_2_72 = _RAND_456[3:0];
  _RAND_457 = {1{`RANDOM}};
  image_2_73 = _RAND_457[3:0];
  _RAND_458 = {1{`RANDOM}};
  image_2_74 = _RAND_458[3:0];
  _RAND_459 = {1{`RANDOM}};
  image_2_75 = _RAND_459[3:0];
  _RAND_460 = {1{`RANDOM}};
  image_2_76 = _RAND_460[3:0];
  _RAND_461 = {1{`RANDOM}};
  image_2_77 = _RAND_461[3:0];
  _RAND_462 = {1{`RANDOM}};
  image_2_78 = _RAND_462[3:0];
  _RAND_463 = {1{`RANDOM}};
  image_2_79 = _RAND_463[3:0];
  _RAND_464 = {1{`RANDOM}};
  image_2_80 = _RAND_464[3:0];
  _RAND_465 = {1{`RANDOM}};
  image_2_81 = _RAND_465[3:0];
  _RAND_466 = {1{`RANDOM}};
  image_2_82 = _RAND_466[3:0];
  _RAND_467 = {1{`RANDOM}};
  image_2_83 = _RAND_467[3:0];
  _RAND_468 = {1{`RANDOM}};
  image_2_84 = _RAND_468[3:0];
  _RAND_469 = {1{`RANDOM}};
  image_2_85 = _RAND_469[3:0];
  _RAND_470 = {1{`RANDOM}};
  image_2_86 = _RAND_470[3:0];
  _RAND_471 = {1{`RANDOM}};
  image_2_87 = _RAND_471[3:0];
  _RAND_472 = {1{`RANDOM}};
  image_2_88 = _RAND_472[3:0];
  _RAND_473 = {1{`RANDOM}};
  image_2_89 = _RAND_473[3:0];
  _RAND_474 = {1{`RANDOM}};
  image_2_90 = _RAND_474[3:0];
  _RAND_475 = {1{`RANDOM}};
  image_2_91 = _RAND_475[3:0];
  _RAND_476 = {1{`RANDOM}};
  image_2_92 = _RAND_476[3:0];
  _RAND_477 = {1{`RANDOM}};
  image_2_93 = _RAND_477[3:0];
  _RAND_478 = {1{`RANDOM}};
  image_2_94 = _RAND_478[3:0];
  _RAND_479 = {1{`RANDOM}};
  image_2_95 = _RAND_479[3:0];
  _RAND_480 = {1{`RANDOM}};
  image_2_96 = _RAND_480[3:0];
  _RAND_481 = {1{`RANDOM}};
  image_2_97 = _RAND_481[3:0];
  _RAND_482 = {1{`RANDOM}};
  image_2_98 = _RAND_482[3:0];
  _RAND_483 = {1{`RANDOM}};
  image_2_99 = _RAND_483[3:0];
  _RAND_484 = {1{`RANDOM}};
  image_2_100 = _RAND_484[3:0];
  _RAND_485 = {1{`RANDOM}};
  image_2_101 = _RAND_485[3:0];
  _RAND_486 = {1{`RANDOM}};
  image_2_102 = _RAND_486[3:0];
  _RAND_487 = {1{`RANDOM}};
  image_2_103 = _RAND_487[3:0];
  _RAND_488 = {1{`RANDOM}};
  image_2_104 = _RAND_488[3:0];
  _RAND_489 = {1{`RANDOM}};
  image_2_105 = _RAND_489[3:0];
  _RAND_490 = {1{`RANDOM}};
  image_2_106 = _RAND_490[3:0];
  _RAND_491 = {1{`RANDOM}};
  image_2_107 = _RAND_491[3:0];
  _RAND_492 = {1{`RANDOM}};
  image_2_108 = _RAND_492[3:0];
  _RAND_493 = {1{`RANDOM}};
  image_2_109 = _RAND_493[3:0];
  _RAND_494 = {1{`RANDOM}};
  image_2_110 = _RAND_494[3:0];
  _RAND_495 = {1{`RANDOM}};
  image_2_111 = _RAND_495[3:0];
  _RAND_496 = {1{`RANDOM}};
  image_2_112 = _RAND_496[3:0];
  _RAND_497 = {1{`RANDOM}};
  image_2_113 = _RAND_497[3:0];
  _RAND_498 = {1{`RANDOM}};
  image_2_114 = _RAND_498[3:0];
  _RAND_499 = {1{`RANDOM}};
  image_2_115 = _RAND_499[3:0];
  _RAND_500 = {1{`RANDOM}};
  image_2_116 = _RAND_500[3:0];
  _RAND_501 = {1{`RANDOM}};
  image_2_117 = _RAND_501[3:0];
  _RAND_502 = {1{`RANDOM}};
  image_2_118 = _RAND_502[3:0];
  _RAND_503 = {1{`RANDOM}};
  image_2_119 = _RAND_503[3:0];
  _RAND_504 = {1{`RANDOM}};
  image_2_120 = _RAND_504[3:0];
  _RAND_505 = {1{`RANDOM}};
  image_2_121 = _RAND_505[3:0];
  _RAND_506 = {1{`RANDOM}};
  image_2_122 = _RAND_506[3:0];
  _RAND_507 = {1{`RANDOM}};
  image_2_123 = _RAND_507[3:0];
  _RAND_508 = {1{`RANDOM}};
  image_2_124 = _RAND_508[3:0];
  _RAND_509 = {1{`RANDOM}};
  image_2_125 = _RAND_509[3:0];
  _RAND_510 = {1{`RANDOM}};
  image_2_126 = _RAND_510[3:0];
  _RAND_511 = {1{`RANDOM}};
  image_2_127 = _RAND_511[3:0];
  _RAND_512 = {1{`RANDOM}};
  image_2_128 = _RAND_512[3:0];
  _RAND_513 = {1{`RANDOM}};
  image_2_129 = _RAND_513[3:0];
  _RAND_514 = {1{`RANDOM}};
  image_2_130 = _RAND_514[3:0];
  _RAND_515 = {1{`RANDOM}};
  image_2_131 = _RAND_515[3:0];
  _RAND_516 = {1{`RANDOM}};
  image_2_132 = _RAND_516[3:0];
  _RAND_517 = {1{`RANDOM}};
  image_2_133 = _RAND_517[3:0];
  _RAND_518 = {1{`RANDOM}};
  image_2_134 = _RAND_518[3:0];
  _RAND_519 = {1{`RANDOM}};
  image_2_135 = _RAND_519[3:0];
  _RAND_520 = {1{`RANDOM}};
  image_2_136 = _RAND_520[3:0];
  _RAND_521 = {1{`RANDOM}};
  image_2_137 = _RAND_521[3:0];
  _RAND_522 = {1{`RANDOM}};
  image_2_138 = _RAND_522[3:0];
  _RAND_523 = {1{`RANDOM}};
  image_2_139 = _RAND_523[3:0];
  _RAND_524 = {1{`RANDOM}};
  image_2_140 = _RAND_524[3:0];
  _RAND_525 = {1{`RANDOM}};
  image_2_141 = _RAND_525[3:0];
  _RAND_526 = {1{`RANDOM}};
  image_2_142 = _RAND_526[3:0];
  _RAND_527 = {1{`RANDOM}};
  image_2_143 = _RAND_527[3:0];
  _RAND_528 = {1{`RANDOM}};
  image_2_144 = _RAND_528[3:0];
  _RAND_529 = {1{`RANDOM}};
  image_2_145 = _RAND_529[3:0];
  _RAND_530 = {1{`RANDOM}};
  image_2_146 = _RAND_530[3:0];
  _RAND_531 = {1{`RANDOM}};
  image_2_147 = _RAND_531[3:0];
  _RAND_532 = {1{`RANDOM}};
  image_2_148 = _RAND_532[3:0];
  _RAND_533 = {1{`RANDOM}};
  image_2_149 = _RAND_533[3:0];
  _RAND_534 = {1{`RANDOM}};
  image_2_150 = _RAND_534[3:0];
  _RAND_535 = {1{`RANDOM}};
  image_2_151 = _RAND_535[3:0];
  _RAND_536 = {1{`RANDOM}};
  image_2_152 = _RAND_536[3:0];
  _RAND_537 = {1{`RANDOM}};
  image_2_153 = _RAND_537[3:0];
  _RAND_538 = {1{`RANDOM}};
  image_2_154 = _RAND_538[3:0];
  _RAND_539 = {1{`RANDOM}};
  image_2_155 = _RAND_539[3:0];
  _RAND_540 = {1{`RANDOM}};
  image_2_156 = _RAND_540[3:0];
  _RAND_541 = {1{`RANDOM}};
  image_2_157 = _RAND_541[3:0];
  _RAND_542 = {1{`RANDOM}};
  image_2_158 = _RAND_542[3:0];
  _RAND_543 = {1{`RANDOM}};
  image_2_159 = _RAND_543[3:0];
  _RAND_544 = {1{`RANDOM}};
  image_2_160 = _RAND_544[3:0];
  _RAND_545 = {1{`RANDOM}};
  image_2_161 = _RAND_545[3:0];
  _RAND_546 = {1{`RANDOM}};
  image_2_162 = _RAND_546[3:0];
  _RAND_547 = {1{`RANDOM}};
  image_2_163 = _RAND_547[3:0];
  _RAND_548 = {1{`RANDOM}};
  image_2_164 = _RAND_548[3:0];
  _RAND_549 = {1{`RANDOM}};
  image_2_165 = _RAND_549[3:0];
  _RAND_550 = {1{`RANDOM}};
  image_2_166 = _RAND_550[3:0];
  _RAND_551 = {1{`RANDOM}};
  image_2_167 = _RAND_551[3:0];
  _RAND_552 = {1{`RANDOM}};
  image_2_168 = _RAND_552[3:0];
  _RAND_553 = {1{`RANDOM}};
  image_2_169 = _RAND_553[3:0];
  _RAND_554 = {1{`RANDOM}};
  image_2_170 = _RAND_554[3:0];
  _RAND_555 = {1{`RANDOM}};
  image_2_171 = _RAND_555[3:0];
  _RAND_556 = {1{`RANDOM}};
  image_2_172 = _RAND_556[3:0];
  _RAND_557 = {1{`RANDOM}};
  image_2_173 = _RAND_557[3:0];
  _RAND_558 = {1{`RANDOM}};
  image_2_174 = _RAND_558[3:0];
  _RAND_559 = {1{`RANDOM}};
  image_2_175 = _RAND_559[3:0];
  _RAND_560 = {1{`RANDOM}};
  image_2_176 = _RAND_560[3:0];
  _RAND_561 = {1{`RANDOM}};
  image_2_177 = _RAND_561[3:0];
  _RAND_562 = {1{`RANDOM}};
  image_2_178 = _RAND_562[3:0];
  _RAND_563 = {1{`RANDOM}};
  image_2_179 = _RAND_563[3:0];
  _RAND_564 = {1{`RANDOM}};
  image_2_180 = _RAND_564[3:0];
  _RAND_565 = {1{`RANDOM}};
  image_2_181 = _RAND_565[3:0];
  _RAND_566 = {1{`RANDOM}};
  image_2_182 = _RAND_566[3:0];
  _RAND_567 = {1{`RANDOM}};
  image_2_183 = _RAND_567[3:0];
  _RAND_568 = {1{`RANDOM}};
  image_2_184 = _RAND_568[3:0];
  _RAND_569 = {1{`RANDOM}};
  image_2_185 = _RAND_569[3:0];
  _RAND_570 = {1{`RANDOM}};
  image_2_186 = _RAND_570[3:0];
  _RAND_571 = {1{`RANDOM}};
  image_2_187 = _RAND_571[3:0];
  _RAND_572 = {1{`RANDOM}};
  image_2_188 = _RAND_572[3:0];
  _RAND_573 = {1{`RANDOM}};
  image_2_189 = _RAND_573[3:0];
  _RAND_574 = {1{`RANDOM}};
  image_2_190 = _RAND_574[3:0];
  _RAND_575 = {1{`RANDOM}};
  image_2_191 = _RAND_575[3:0];
  _RAND_576 = {1{`RANDOM}};
  pixelIndex = _RAND_576[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      image_0_0 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h0 == _T_37[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_7;
      end else if (8'h0 == _T_34[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_6;
      end else if (8'h0 == _T_31[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_5;
      end else if (8'h0 == _T_28[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_4;
      end else if (8'h0 == _T_25[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_3;
      end else if (8'h0 == _T_22[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_2;
      end else if (8'h0 == _T_19[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_1;
      end else if (8'h0 == _T_15[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_1 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1 == _T_37[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_7;
      end else if (8'h1 == _T_34[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_6;
      end else if (8'h1 == _T_31[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_5;
      end else if (8'h1 == _T_28[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_4;
      end else if (8'h1 == _T_25[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_3;
      end else if (8'h1 == _T_22[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_2;
      end else if (8'h1 == _T_19[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_1;
      end else if (8'h1 == _T_15[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_2 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2 == _T_37[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_7;
      end else if (8'h2 == _T_34[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_6;
      end else if (8'h2 == _T_31[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_5;
      end else if (8'h2 == _T_28[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_4;
      end else if (8'h2 == _T_25[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_3;
      end else if (8'h2 == _T_22[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_2;
      end else if (8'h2 == _T_19[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_1;
      end else if (8'h2 == _T_15[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_3 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3 == _T_37[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_7;
      end else if (8'h3 == _T_34[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_6;
      end else if (8'h3 == _T_31[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_5;
      end else if (8'h3 == _T_28[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_4;
      end else if (8'h3 == _T_25[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_3;
      end else if (8'h3 == _T_22[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_2;
      end else if (8'h3 == _T_19[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_1;
      end else if (8'h3 == _T_15[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_4 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4 == _T_37[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_7;
      end else if (8'h4 == _T_34[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_6;
      end else if (8'h4 == _T_31[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_5;
      end else if (8'h4 == _T_28[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_4;
      end else if (8'h4 == _T_25[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_3;
      end else if (8'h4 == _T_22[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_2;
      end else if (8'h4 == _T_19[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_1;
      end else if (8'h4 == _T_15[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_5 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5 == _T_37[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_7;
      end else if (8'h5 == _T_34[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_6;
      end else if (8'h5 == _T_31[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_5;
      end else if (8'h5 == _T_28[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_4;
      end else if (8'h5 == _T_25[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_3;
      end else if (8'h5 == _T_22[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_2;
      end else if (8'h5 == _T_19[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_1;
      end else if (8'h5 == _T_15[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_6 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6 == _T_37[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_7;
      end else if (8'h6 == _T_34[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_6;
      end else if (8'h6 == _T_31[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_5;
      end else if (8'h6 == _T_28[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_4;
      end else if (8'h6 == _T_25[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_3;
      end else if (8'h6 == _T_22[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_2;
      end else if (8'h6 == _T_19[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_1;
      end else if (8'h6 == _T_15[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_7 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7 == _T_37[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_7;
      end else if (8'h7 == _T_34[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_6;
      end else if (8'h7 == _T_31[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_5;
      end else if (8'h7 == _T_28[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_4;
      end else if (8'h7 == _T_25[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_3;
      end else if (8'h7 == _T_22[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_2;
      end else if (8'h7 == _T_19[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_1;
      end else if (8'h7 == _T_15[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_8 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8 == _T_37[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_7;
      end else if (8'h8 == _T_34[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_6;
      end else if (8'h8 == _T_31[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_5;
      end else if (8'h8 == _T_28[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_4;
      end else if (8'h8 == _T_25[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_3;
      end else if (8'h8 == _T_22[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_2;
      end else if (8'h8 == _T_19[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_1;
      end else if (8'h8 == _T_15[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_9 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h9 == _T_37[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_7;
      end else if (8'h9 == _T_34[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_6;
      end else if (8'h9 == _T_31[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_5;
      end else if (8'h9 == _T_28[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_4;
      end else if (8'h9 == _T_25[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_3;
      end else if (8'h9 == _T_22[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_2;
      end else if (8'h9 == _T_19[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_1;
      end else if (8'h9 == _T_15[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_10 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha == _T_37[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_7;
      end else if (8'ha == _T_34[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_6;
      end else if (8'ha == _T_31[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_5;
      end else if (8'ha == _T_28[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_4;
      end else if (8'ha == _T_25[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_3;
      end else if (8'ha == _T_22[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_2;
      end else if (8'ha == _T_19[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_1;
      end else if (8'ha == _T_15[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_11 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb == _T_37[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_7;
      end else if (8'hb == _T_34[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_6;
      end else if (8'hb == _T_31[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_5;
      end else if (8'hb == _T_28[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_4;
      end else if (8'hb == _T_25[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_3;
      end else if (8'hb == _T_22[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_2;
      end else if (8'hb == _T_19[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_1;
      end else if (8'hb == _T_15[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_12 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hc == _T_37[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_7;
      end else if (8'hc == _T_34[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_6;
      end else if (8'hc == _T_31[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_5;
      end else if (8'hc == _T_28[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_4;
      end else if (8'hc == _T_25[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_3;
      end else if (8'hc == _T_22[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_2;
      end else if (8'hc == _T_19[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_1;
      end else if (8'hc == _T_15[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_13 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hd == _T_37[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_7;
      end else if (8'hd == _T_34[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_6;
      end else if (8'hd == _T_31[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_5;
      end else if (8'hd == _T_28[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_4;
      end else if (8'hd == _T_25[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_3;
      end else if (8'hd == _T_22[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_2;
      end else if (8'hd == _T_19[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_1;
      end else if (8'hd == _T_15[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_14 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'he == _T_37[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_7;
      end else if (8'he == _T_34[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_6;
      end else if (8'he == _T_31[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_5;
      end else if (8'he == _T_28[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_4;
      end else if (8'he == _T_25[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_3;
      end else if (8'he == _T_22[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_2;
      end else if (8'he == _T_19[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_1;
      end else if (8'he == _T_15[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_15 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hf == _T_37[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_7;
      end else if (8'hf == _T_34[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_6;
      end else if (8'hf == _T_31[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_5;
      end else if (8'hf == _T_28[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_4;
      end else if (8'hf == _T_25[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_3;
      end else if (8'hf == _T_22[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_2;
      end else if (8'hf == _T_19[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_1;
      end else if (8'hf == _T_15[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_16 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h10 == _T_37[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_7;
      end else if (8'h10 == _T_34[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_6;
      end else if (8'h10 == _T_31[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_5;
      end else if (8'h10 == _T_28[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_4;
      end else if (8'h10 == _T_25[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_3;
      end else if (8'h10 == _T_22[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_2;
      end else if (8'h10 == _T_19[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_1;
      end else if (8'h10 == _T_15[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_17 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h11 == _T_37[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_7;
      end else if (8'h11 == _T_34[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_6;
      end else if (8'h11 == _T_31[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_5;
      end else if (8'h11 == _T_28[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_4;
      end else if (8'h11 == _T_25[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_3;
      end else if (8'h11 == _T_22[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_2;
      end else if (8'h11 == _T_19[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_1;
      end else if (8'h11 == _T_15[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_18 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h12 == _T_37[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_7;
      end else if (8'h12 == _T_34[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_6;
      end else if (8'h12 == _T_31[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_5;
      end else if (8'h12 == _T_28[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_4;
      end else if (8'h12 == _T_25[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_3;
      end else if (8'h12 == _T_22[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_2;
      end else if (8'h12 == _T_19[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_1;
      end else if (8'h12 == _T_15[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_19 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h13 == _T_37[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_7;
      end else if (8'h13 == _T_34[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_6;
      end else if (8'h13 == _T_31[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_5;
      end else if (8'h13 == _T_28[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_4;
      end else if (8'h13 == _T_25[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_3;
      end else if (8'h13 == _T_22[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_2;
      end else if (8'h13 == _T_19[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_1;
      end else if (8'h13 == _T_15[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_20 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h14 == _T_37[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_7;
      end else if (8'h14 == _T_34[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_6;
      end else if (8'h14 == _T_31[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_5;
      end else if (8'h14 == _T_28[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_4;
      end else if (8'h14 == _T_25[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_3;
      end else if (8'h14 == _T_22[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_2;
      end else if (8'h14 == _T_19[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_1;
      end else if (8'h14 == _T_15[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_21 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h15 == _T_37[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_7;
      end else if (8'h15 == _T_34[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_6;
      end else if (8'h15 == _T_31[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_5;
      end else if (8'h15 == _T_28[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_4;
      end else if (8'h15 == _T_25[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_3;
      end else if (8'h15 == _T_22[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_2;
      end else if (8'h15 == _T_19[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_1;
      end else if (8'h15 == _T_15[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_22 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h16 == _T_37[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_7;
      end else if (8'h16 == _T_34[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_6;
      end else if (8'h16 == _T_31[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_5;
      end else if (8'h16 == _T_28[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_4;
      end else if (8'h16 == _T_25[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_3;
      end else if (8'h16 == _T_22[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_2;
      end else if (8'h16 == _T_19[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_1;
      end else if (8'h16 == _T_15[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_23 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h17 == _T_37[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_7;
      end else if (8'h17 == _T_34[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_6;
      end else if (8'h17 == _T_31[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_5;
      end else if (8'h17 == _T_28[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_4;
      end else if (8'h17 == _T_25[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_3;
      end else if (8'h17 == _T_22[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_2;
      end else if (8'h17 == _T_19[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_1;
      end else if (8'h17 == _T_15[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_24 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h18 == _T_37[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_7;
      end else if (8'h18 == _T_34[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_6;
      end else if (8'h18 == _T_31[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_5;
      end else if (8'h18 == _T_28[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_4;
      end else if (8'h18 == _T_25[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_3;
      end else if (8'h18 == _T_22[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_2;
      end else if (8'h18 == _T_19[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_1;
      end else if (8'h18 == _T_15[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_25 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h19 == _T_37[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_7;
      end else if (8'h19 == _T_34[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_6;
      end else if (8'h19 == _T_31[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_5;
      end else if (8'h19 == _T_28[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_4;
      end else if (8'h19 == _T_25[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_3;
      end else if (8'h19 == _T_22[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_2;
      end else if (8'h19 == _T_19[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_1;
      end else if (8'h19 == _T_15[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_26 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1a == _T_37[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_7;
      end else if (8'h1a == _T_34[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_6;
      end else if (8'h1a == _T_31[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_5;
      end else if (8'h1a == _T_28[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_4;
      end else if (8'h1a == _T_25[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_3;
      end else if (8'h1a == _T_22[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_2;
      end else if (8'h1a == _T_19[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_1;
      end else if (8'h1a == _T_15[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_27 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1b == _T_37[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_7;
      end else if (8'h1b == _T_34[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_6;
      end else if (8'h1b == _T_31[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_5;
      end else if (8'h1b == _T_28[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_4;
      end else if (8'h1b == _T_25[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_3;
      end else if (8'h1b == _T_22[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_2;
      end else if (8'h1b == _T_19[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_1;
      end else if (8'h1b == _T_15[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_28 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1c == _T_37[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_7;
      end else if (8'h1c == _T_34[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_6;
      end else if (8'h1c == _T_31[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_5;
      end else if (8'h1c == _T_28[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_4;
      end else if (8'h1c == _T_25[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_3;
      end else if (8'h1c == _T_22[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_2;
      end else if (8'h1c == _T_19[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_1;
      end else if (8'h1c == _T_15[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_29 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1d == _T_37[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_7;
      end else if (8'h1d == _T_34[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_6;
      end else if (8'h1d == _T_31[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_5;
      end else if (8'h1d == _T_28[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_4;
      end else if (8'h1d == _T_25[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_3;
      end else if (8'h1d == _T_22[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_2;
      end else if (8'h1d == _T_19[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_1;
      end else if (8'h1d == _T_15[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_30 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1e == _T_37[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_7;
      end else if (8'h1e == _T_34[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_6;
      end else if (8'h1e == _T_31[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_5;
      end else if (8'h1e == _T_28[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_4;
      end else if (8'h1e == _T_25[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_3;
      end else if (8'h1e == _T_22[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_2;
      end else if (8'h1e == _T_19[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_1;
      end else if (8'h1e == _T_15[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_31 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1f == _T_37[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_7;
      end else if (8'h1f == _T_34[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_6;
      end else if (8'h1f == _T_31[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_5;
      end else if (8'h1f == _T_28[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_4;
      end else if (8'h1f == _T_25[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_3;
      end else if (8'h1f == _T_22[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_2;
      end else if (8'h1f == _T_19[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_1;
      end else if (8'h1f == _T_15[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_32 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h20 == _T_37[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_7;
      end else if (8'h20 == _T_34[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_6;
      end else if (8'h20 == _T_31[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_5;
      end else if (8'h20 == _T_28[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_4;
      end else if (8'h20 == _T_25[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_3;
      end else if (8'h20 == _T_22[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_2;
      end else if (8'h20 == _T_19[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_1;
      end else if (8'h20 == _T_15[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_33 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h21 == _T_37[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_7;
      end else if (8'h21 == _T_34[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_6;
      end else if (8'h21 == _T_31[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_5;
      end else if (8'h21 == _T_28[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_4;
      end else if (8'h21 == _T_25[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_3;
      end else if (8'h21 == _T_22[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_2;
      end else if (8'h21 == _T_19[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_1;
      end else if (8'h21 == _T_15[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_34 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h22 == _T_37[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_7;
      end else if (8'h22 == _T_34[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_6;
      end else if (8'h22 == _T_31[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_5;
      end else if (8'h22 == _T_28[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_4;
      end else if (8'h22 == _T_25[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_3;
      end else if (8'h22 == _T_22[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_2;
      end else if (8'h22 == _T_19[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_1;
      end else if (8'h22 == _T_15[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_35 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h23 == _T_37[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_7;
      end else if (8'h23 == _T_34[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_6;
      end else if (8'h23 == _T_31[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_5;
      end else if (8'h23 == _T_28[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_4;
      end else if (8'h23 == _T_25[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_3;
      end else if (8'h23 == _T_22[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_2;
      end else if (8'h23 == _T_19[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_1;
      end else if (8'h23 == _T_15[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_36 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h24 == _T_37[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_7;
      end else if (8'h24 == _T_34[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_6;
      end else if (8'h24 == _T_31[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_5;
      end else if (8'h24 == _T_28[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_4;
      end else if (8'h24 == _T_25[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_3;
      end else if (8'h24 == _T_22[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_2;
      end else if (8'h24 == _T_19[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_1;
      end else if (8'h24 == _T_15[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_37 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h25 == _T_37[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_7;
      end else if (8'h25 == _T_34[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_6;
      end else if (8'h25 == _T_31[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_5;
      end else if (8'h25 == _T_28[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_4;
      end else if (8'h25 == _T_25[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_3;
      end else if (8'h25 == _T_22[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_2;
      end else if (8'h25 == _T_19[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_1;
      end else if (8'h25 == _T_15[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_38 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h26 == _T_37[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_7;
      end else if (8'h26 == _T_34[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_6;
      end else if (8'h26 == _T_31[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_5;
      end else if (8'h26 == _T_28[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_4;
      end else if (8'h26 == _T_25[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_3;
      end else if (8'h26 == _T_22[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_2;
      end else if (8'h26 == _T_19[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_1;
      end else if (8'h26 == _T_15[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_39 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h27 == _T_37[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_7;
      end else if (8'h27 == _T_34[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_6;
      end else if (8'h27 == _T_31[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_5;
      end else if (8'h27 == _T_28[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_4;
      end else if (8'h27 == _T_25[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_3;
      end else if (8'h27 == _T_22[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_2;
      end else if (8'h27 == _T_19[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_1;
      end else if (8'h27 == _T_15[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_40 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h28 == _T_37[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_7;
      end else if (8'h28 == _T_34[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_6;
      end else if (8'h28 == _T_31[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_5;
      end else if (8'h28 == _T_28[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_4;
      end else if (8'h28 == _T_25[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_3;
      end else if (8'h28 == _T_22[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_2;
      end else if (8'h28 == _T_19[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_1;
      end else if (8'h28 == _T_15[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_41 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h29 == _T_37[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_7;
      end else if (8'h29 == _T_34[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_6;
      end else if (8'h29 == _T_31[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_5;
      end else if (8'h29 == _T_28[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_4;
      end else if (8'h29 == _T_25[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_3;
      end else if (8'h29 == _T_22[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_2;
      end else if (8'h29 == _T_19[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_1;
      end else if (8'h29 == _T_15[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_42 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2a == _T_37[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_7;
      end else if (8'h2a == _T_34[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_6;
      end else if (8'h2a == _T_31[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_5;
      end else if (8'h2a == _T_28[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_4;
      end else if (8'h2a == _T_25[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_3;
      end else if (8'h2a == _T_22[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_2;
      end else if (8'h2a == _T_19[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_1;
      end else if (8'h2a == _T_15[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_43 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2b == _T_37[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_7;
      end else if (8'h2b == _T_34[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_6;
      end else if (8'h2b == _T_31[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_5;
      end else if (8'h2b == _T_28[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_4;
      end else if (8'h2b == _T_25[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_3;
      end else if (8'h2b == _T_22[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_2;
      end else if (8'h2b == _T_19[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_1;
      end else if (8'h2b == _T_15[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_44 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2c == _T_37[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_7;
      end else if (8'h2c == _T_34[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_6;
      end else if (8'h2c == _T_31[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_5;
      end else if (8'h2c == _T_28[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_4;
      end else if (8'h2c == _T_25[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_3;
      end else if (8'h2c == _T_22[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_2;
      end else if (8'h2c == _T_19[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_1;
      end else if (8'h2c == _T_15[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_45 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2d == _T_37[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_7;
      end else if (8'h2d == _T_34[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_6;
      end else if (8'h2d == _T_31[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_5;
      end else if (8'h2d == _T_28[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_4;
      end else if (8'h2d == _T_25[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_3;
      end else if (8'h2d == _T_22[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_2;
      end else if (8'h2d == _T_19[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_1;
      end else if (8'h2d == _T_15[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_46 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2e == _T_37[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_7;
      end else if (8'h2e == _T_34[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_6;
      end else if (8'h2e == _T_31[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_5;
      end else if (8'h2e == _T_28[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_4;
      end else if (8'h2e == _T_25[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_3;
      end else if (8'h2e == _T_22[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_2;
      end else if (8'h2e == _T_19[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_1;
      end else if (8'h2e == _T_15[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_47 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2f == _T_37[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_7;
      end else if (8'h2f == _T_34[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_6;
      end else if (8'h2f == _T_31[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_5;
      end else if (8'h2f == _T_28[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_4;
      end else if (8'h2f == _T_25[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_3;
      end else if (8'h2f == _T_22[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_2;
      end else if (8'h2f == _T_19[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_1;
      end else if (8'h2f == _T_15[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_48 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h30 == _T_37[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_7;
      end else if (8'h30 == _T_34[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_6;
      end else if (8'h30 == _T_31[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_5;
      end else if (8'h30 == _T_28[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_4;
      end else if (8'h30 == _T_25[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_3;
      end else if (8'h30 == _T_22[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_2;
      end else if (8'h30 == _T_19[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_1;
      end else if (8'h30 == _T_15[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_49 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h31 == _T_37[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_7;
      end else if (8'h31 == _T_34[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_6;
      end else if (8'h31 == _T_31[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_5;
      end else if (8'h31 == _T_28[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_4;
      end else if (8'h31 == _T_25[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_3;
      end else if (8'h31 == _T_22[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_2;
      end else if (8'h31 == _T_19[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_1;
      end else if (8'h31 == _T_15[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_50 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h32 == _T_37[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_7;
      end else if (8'h32 == _T_34[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_6;
      end else if (8'h32 == _T_31[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_5;
      end else if (8'h32 == _T_28[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_4;
      end else if (8'h32 == _T_25[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_3;
      end else if (8'h32 == _T_22[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_2;
      end else if (8'h32 == _T_19[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_1;
      end else if (8'h32 == _T_15[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_51 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h33 == _T_37[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_7;
      end else if (8'h33 == _T_34[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_6;
      end else if (8'h33 == _T_31[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_5;
      end else if (8'h33 == _T_28[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_4;
      end else if (8'h33 == _T_25[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_3;
      end else if (8'h33 == _T_22[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_2;
      end else if (8'h33 == _T_19[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_1;
      end else if (8'h33 == _T_15[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_52 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h34 == _T_37[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_7;
      end else if (8'h34 == _T_34[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_6;
      end else if (8'h34 == _T_31[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_5;
      end else if (8'h34 == _T_28[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_4;
      end else if (8'h34 == _T_25[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_3;
      end else if (8'h34 == _T_22[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_2;
      end else if (8'h34 == _T_19[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_1;
      end else if (8'h34 == _T_15[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_53 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h35 == _T_37[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_7;
      end else if (8'h35 == _T_34[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_6;
      end else if (8'h35 == _T_31[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_5;
      end else if (8'h35 == _T_28[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_4;
      end else if (8'h35 == _T_25[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_3;
      end else if (8'h35 == _T_22[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_2;
      end else if (8'h35 == _T_19[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_1;
      end else if (8'h35 == _T_15[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_54 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h36 == _T_37[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_7;
      end else if (8'h36 == _T_34[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_6;
      end else if (8'h36 == _T_31[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_5;
      end else if (8'h36 == _T_28[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_4;
      end else if (8'h36 == _T_25[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_3;
      end else if (8'h36 == _T_22[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_2;
      end else if (8'h36 == _T_19[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_1;
      end else if (8'h36 == _T_15[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_55 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h37 == _T_37[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_7;
      end else if (8'h37 == _T_34[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_6;
      end else if (8'h37 == _T_31[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_5;
      end else if (8'h37 == _T_28[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_4;
      end else if (8'h37 == _T_25[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_3;
      end else if (8'h37 == _T_22[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_2;
      end else if (8'h37 == _T_19[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_1;
      end else if (8'h37 == _T_15[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_56 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h38 == _T_37[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_7;
      end else if (8'h38 == _T_34[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_6;
      end else if (8'h38 == _T_31[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_5;
      end else if (8'h38 == _T_28[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_4;
      end else if (8'h38 == _T_25[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_3;
      end else if (8'h38 == _T_22[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_2;
      end else if (8'h38 == _T_19[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_1;
      end else if (8'h38 == _T_15[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_57 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h39 == _T_37[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_7;
      end else if (8'h39 == _T_34[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_6;
      end else if (8'h39 == _T_31[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_5;
      end else if (8'h39 == _T_28[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_4;
      end else if (8'h39 == _T_25[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_3;
      end else if (8'h39 == _T_22[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_2;
      end else if (8'h39 == _T_19[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_1;
      end else if (8'h39 == _T_15[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_58 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3a == _T_37[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_7;
      end else if (8'h3a == _T_34[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_6;
      end else if (8'h3a == _T_31[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_5;
      end else if (8'h3a == _T_28[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_4;
      end else if (8'h3a == _T_25[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_3;
      end else if (8'h3a == _T_22[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_2;
      end else if (8'h3a == _T_19[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_1;
      end else if (8'h3a == _T_15[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_59 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3b == _T_37[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_7;
      end else if (8'h3b == _T_34[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_6;
      end else if (8'h3b == _T_31[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_5;
      end else if (8'h3b == _T_28[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_4;
      end else if (8'h3b == _T_25[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_3;
      end else if (8'h3b == _T_22[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_2;
      end else if (8'h3b == _T_19[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_1;
      end else if (8'h3b == _T_15[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_60 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3c == _T_37[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_7;
      end else if (8'h3c == _T_34[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_6;
      end else if (8'h3c == _T_31[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_5;
      end else if (8'h3c == _T_28[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_4;
      end else if (8'h3c == _T_25[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_3;
      end else if (8'h3c == _T_22[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_2;
      end else if (8'h3c == _T_19[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_1;
      end else if (8'h3c == _T_15[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_61 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3d == _T_37[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_7;
      end else if (8'h3d == _T_34[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_6;
      end else if (8'h3d == _T_31[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_5;
      end else if (8'h3d == _T_28[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_4;
      end else if (8'h3d == _T_25[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_3;
      end else if (8'h3d == _T_22[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_2;
      end else if (8'h3d == _T_19[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_1;
      end else if (8'h3d == _T_15[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_62 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3e == _T_37[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_7;
      end else if (8'h3e == _T_34[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_6;
      end else if (8'h3e == _T_31[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_5;
      end else if (8'h3e == _T_28[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_4;
      end else if (8'h3e == _T_25[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_3;
      end else if (8'h3e == _T_22[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_2;
      end else if (8'h3e == _T_19[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_1;
      end else if (8'h3e == _T_15[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_63 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3f == _T_37[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_7;
      end else if (8'h3f == _T_34[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_6;
      end else if (8'h3f == _T_31[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_5;
      end else if (8'h3f == _T_28[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_4;
      end else if (8'h3f == _T_25[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_3;
      end else if (8'h3f == _T_22[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_2;
      end else if (8'h3f == _T_19[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_1;
      end else if (8'h3f == _T_15[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_64 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h40 == _T_37[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_7;
      end else if (8'h40 == _T_34[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_6;
      end else if (8'h40 == _T_31[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_5;
      end else if (8'h40 == _T_28[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_4;
      end else if (8'h40 == _T_25[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_3;
      end else if (8'h40 == _T_22[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_2;
      end else if (8'h40 == _T_19[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_1;
      end else if (8'h40 == _T_15[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_65 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h41 == _T_37[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_7;
      end else if (8'h41 == _T_34[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_6;
      end else if (8'h41 == _T_31[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_5;
      end else if (8'h41 == _T_28[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_4;
      end else if (8'h41 == _T_25[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_3;
      end else if (8'h41 == _T_22[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_2;
      end else if (8'h41 == _T_19[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_1;
      end else if (8'h41 == _T_15[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_66 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h42 == _T_37[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_7;
      end else if (8'h42 == _T_34[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_6;
      end else if (8'h42 == _T_31[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_5;
      end else if (8'h42 == _T_28[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_4;
      end else if (8'h42 == _T_25[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_3;
      end else if (8'h42 == _T_22[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_2;
      end else if (8'h42 == _T_19[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_1;
      end else if (8'h42 == _T_15[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_67 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h43 == _T_37[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_7;
      end else if (8'h43 == _T_34[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_6;
      end else if (8'h43 == _T_31[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_5;
      end else if (8'h43 == _T_28[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_4;
      end else if (8'h43 == _T_25[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_3;
      end else if (8'h43 == _T_22[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_2;
      end else if (8'h43 == _T_19[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_1;
      end else if (8'h43 == _T_15[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_68 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h44 == _T_37[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_7;
      end else if (8'h44 == _T_34[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_6;
      end else if (8'h44 == _T_31[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_5;
      end else if (8'h44 == _T_28[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_4;
      end else if (8'h44 == _T_25[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_3;
      end else if (8'h44 == _T_22[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_2;
      end else if (8'h44 == _T_19[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_1;
      end else if (8'h44 == _T_15[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_69 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h45 == _T_37[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_7;
      end else if (8'h45 == _T_34[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_6;
      end else if (8'h45 == _T_31[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_5;
      end else if (8'h45 == _T_28[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_4;
      end else if (8'h45 == _T_25[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_3;
      end else if (8'h45 == _T_22[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_2;
      end else if (8'h45 == _T_19[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_1;
      end else if (8'h45 == _T_15[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_70 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h46 == _T_37[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_7;
      end else if (8'h46 == _T_34[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_6;
      end else if (8'h46 == _T_31[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_5;
      end else if (8'h46 == _T_28[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_4;
      end else if (8'h46 == _T_25[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_3;
      end else if (8'h46 == _T_22[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_2;
      end else if (8'h46 == _T_19[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_1;
      end else if (8'h46 == _T_15[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_71 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h47 == _T_37[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_7;
      end else if (8'h47 == _T_34[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_6;
      end else if (8'h47 == _T_31[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_5;
      end else if (8'h47 == _T_28[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_4;
      end else if (8'h47 == _T_25[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_3;
      end else if (8'h47 == _T_22[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_2;
      end else if (8'h47 == _T_19[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_1;
      end else if (8'h47 == _T_15[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_72 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h48 == _T_37[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_7;
      end else if (8'h48 == _T_34[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_6;
      end else if (8'h48 == _T_31[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_5;
      end else if (8'h48 == _T_28[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_4;
      end else if (8'h48 == _T_25[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_3;
      end else if (8'h48 == _T_22[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_2;
      end else if (8'h48 == _T_19[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_1;
      end else if (8'h48 == _T_15[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_73 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h49 == _T_37[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_7;
      end else if (8'h49 == _T_34[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_6;
      end else if (8'h49 == _T_31[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_5;
      end else if (8'h49 == _T_28[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_4;
      end else if (8'h49 == _T_25[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_3;
      end else if (8'h49 == _T_22[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_2;
      end else if (8'h49 == _T_19[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_1;
      end else if (8'h49 == _T_15[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_74 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4a == _T_37[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_7;
      end else if (8'h4a == _T_34[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_6;
      end else if (8'h4a == _T_31[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_5;
      end else if (8'h4a == _T_28[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_4;
      end else if (8'h4a == _T_25[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_3;
      end else if (8'h4a == _T_22[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_2;
      end else if (8'h4a == _T_19[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_1;
      end else if (8'h4a == _T_15[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_75 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4b == _T_37[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_7;
      end else if (8'h4b == _T_34[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_6;
      end else if (8'h4b == _T_31[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_5;
      end else if (8'h4b == _T_28[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_4;
      end else if (8'h4b == _T_25[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_3;
      end else if (8'h4b == _T_22[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_2;
      end else if (8'h4b == _T_19[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_1;
      end else if (8'h4b == _T_15[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_76 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4c == _T_37[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_7;
      end else if (8'h4c == _T_34[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_6;
      end else if (8'h4c == _T_31[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_5;
      end else if (8'h4c == _T_28[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_4;
      end else if (8'h4c == _T_25[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_3;
      end else if (8'h4c == _T_22[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_2;
      end else if (8'h4c == _T_19[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_1;
      end else if (8'h4c == _T_15[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_77 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4d == _T_37[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_7;
      end else if (8'h4d == _T_34[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_6;
      end else if (8'h4d == _T_31[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_5;
      end else if (8'h4d == _T_28[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_4;
      end else if (8'h4d == _T_25[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_3;
      end else if (8'h4d == _T_22[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_2;
      end else if (8'h4d == _T_19[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_1;
      end else if (8'h4d == _T_15[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_78 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4e == _T_37[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_7;
      end else if (8'h4e == _T_34[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_6;
      end else if (8'h4e == _T_31[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_5;
      end else if (8'h4e == _T_28[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_4;
      end else if (8'h4e == _T_25[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_3;
      end else if (8'h4e == _T_22[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_2;
      end else if (8'h4e == _T_19[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_1;
      end else if (8'h4e == _T_15[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_79 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4f == _T_37[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_7;
      end else if (8'h4f == _T_34[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_6;
      end else if (8'h4f == _T_31[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_5;
      end else if (8'h4f == _T_28[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_4;
      end else if (8'h4f == _T_25[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_3;
      end else if (8'h4f == _T_22[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_2;
      end else if (8'h4f == _T_19[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_1;
      end else if (8'h4f == _T_15[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_80 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h50 == _T_37[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_7;
      end else if (8'h50 == _T_34[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_6;
      end else if (8'h50 == _T_31[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_5;
      end else if (8'h50 == _T_28[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_4;
      end else if (8'h50 == _T_25[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_3;
      end else if (8'h50 == _T_22[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_2;
      end else if (8'h50 == _T_19[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_1;
      end else if (8'h50 == _T_15[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_81 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h51 == _T_37[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_7;
      end else if (8'h51 == _T_34[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_6;
      end else if (8'h51 == _T_31[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_5;
      end else if (8'h51 == _T_28[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_4;
      end else if (8'h51 == _T_25[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_3;
      end else if (8'h51 == _T_22[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_2;
      end else if (8'h51 == _T_19[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_1;
      end else if (8'h51 == _T_15[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_82 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h52 == _T_37[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_7;
      end else if (8'h52 == _T_34[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_6;
      end else if (8'h52 == _T_31[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_5;
      end else if (8'h52 == _T_28[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_4;
      end else if (8'h52 == _T_25[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_3;
      end else if (8'h52 == _T_22[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_2;
      end else if (8'h52 == _T_19[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_1;
      end else if (8'h52 == _T_15[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_83 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h53 == _T_37[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_7;
      end else if (8'h53 == _T_34[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_6;
      end else if (8'h53 == _T_31[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_5;
      end else if (8'h53 == _T_28[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_4;
      end else if (8'h53 == _T_25[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_3;
      end else if (8'h53 == _T_22[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_2;
      end else if (8'h53 == _T_19[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_1;
      end else if (8'h53 == _T_15[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_84 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h54 == _T_37[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_7;
      end else if (8'h54 == _T_34[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_6;
      end else if (8'h54 == _T_31[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_5;
      end else if (8'h54 == _T_28[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_4;
      end else if (8'h54 == _T_25[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_3;
      end else if (8'h54 == _T_22[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_2;
      end else if (8'h54 == _T_19[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_1;
      end else if (8'h54 == _T_15[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_85 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h55 == _T_37[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_7;
      end else if (8'h55 == _T_34[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_6;
      end else if (8'h55 == _T_31[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_5;
      end else if (8'h55 == _T_28[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_4;
      end else if (8'h55 == _T_25[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_3;
      end else if (8'h55 == _T_22[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_2;
      end else if (8'h55 == _T_19[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_1;
      end else if (8'h55 == _T_15[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_86 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h56 == _T_37[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_7;
      end else if (8'h56 == _T_34[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_6;
      end else if (8'h56 == _T_31[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_5;
      end else if (8'h56 == _T_28[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_4;
      end else if (8'h56 == _T_25[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_3;
      end else if (8'h56 == _T_22[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_2;
      end else if (8'h56 == _T_19[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_1;
      end else if (8'h56 == _T_15[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_87 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h57 == _T_37[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_7;
      end else if (8'h57 == _T_34[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_6;
      end else if (8'h57 == _T_31[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_5;
      end else if (8'h57 == _T_28[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_4;
      end else if (8'h57 == _T_25[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_3;
      end else if (8'h57 == _T_22[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_2;
      end else if (8'h57 == _T_19[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_1;
      end else if (8'h57 == _T_15[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_88 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h58 == _T_37[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_7;
      end else if (8'h58 == _T_34[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_6;
      end else if (8'h58 == _T_31[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_5;
      end else if (8'h58 == _T_28[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_4;
      end else if (8'h58 == _T_25[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_3;
      end else if (8'h58 == _T_22[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_2;
      end else if (8'h58 == _T_19[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_1;
      end else if (8'h58 == _T_15[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_89 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h59 == _T_37[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_7;
      end else if (8'h59 == _T_34[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_6;
      end else if (8'h59 == _T_31[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_5;
      end else if (8'h59 == _T_28[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_4;
      end else if (8'h59 == _T_25[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_3;
      end else if (8'h59 == _T_22[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_2;
      end else if (8'h59 == _T_19[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_1;
      end else if (8'h59 == _T_15[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_90 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5a == _T_37[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_7;
      end else if (8'h5a == _T_34[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_6;
      end else if (8'h5a == _T_31[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_5;
      end else if (8'h5a == _T_28[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_4;
      end else if (8'h5a == _T_25[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_3;
      end else if (8'h5a == _T_22[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_2;
      end else if (8'h5a == _T_19[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_1;
      end else if (8'h5a == _T_15[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_91 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5b == _T_37[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_7;
      end else if (8'h5b == _T_34[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_6;
      end else if (8'h5b == _T_31[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_5;
      end else if (8'h5b == _T_28[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_4;
      end else if (8'h5b == _T_25[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_3;
      end else if (8'h5b == _T_22[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_2;
      end else if (8'h5b == _T_19[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_1;
      end else if (8'h5b == _T_15[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_92 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5c == _T_37[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_7;
      end else if (8'h5c == _T_34[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_6;
      end else if (8'h5c == _T_31[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_5;
      end else if (8'h5c == _T_28[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_4;
      end else if (8'h5c == _T_25[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_3;
      end else if (8'h5c == _T_22[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_2;
      end else if (8'h5c == _T_19[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_1;
      end else if (8'h5c == _T_15[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_93 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5d == _T_37[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_7;
      end else if (8'h5d == _T_34[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_6;
      end else if (8'h5d == _T_31[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_5;
      end else if (8'h5d == _T_28[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_4;
      end else if (8'h5d == _T_25[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_3;
      end else if (8'h5d == _T_22[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_2;
      end else if (8'h5d == _T_19[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_1;
      end else if (8'h5d == _T_15[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_94 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5e == _T_37[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_7;
      end else if (8'h5e == _T_34[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_6;
      end else if (8'h5e == _T_31[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_5;
      end else if (8'h5e == _T_28[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_4;
      end else if (8'h5e == _T_25[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_3;
      end else if (8'h5e == _T_22[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_2;
      end else if (8'h5e == _T_19[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_1;
      end else if (8'h5e == _T_15[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_95 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5f == _T_37[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_7;
      end else if (8'h5f == _T_34[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_6;
      end else if (8'h5f == _T_31[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_5;
      end else if (8'h5f == _T_28[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_4;
      end else if (8'h5f == _T_25[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_3;
      end else if (8'h5f == _T_22[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_2;
      end else if (8'h5f == _T_19[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_1;
      end else if (8'h5f == _T_15[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_96 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h60 == _T_37[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_7;
      end else if (8'h60 == _T_34[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_6;
      end else if (8'h60 == _T_31[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_5;
      end else if (8'h60 == _T_28[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_4;
      end else if (8'h60 == _T_25[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_3;
      end else if (8'h60 == _T_22[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_2;
      end else if (8'h60 == _T_19[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_1;
      end else if (8'h60 == _T_15[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_97 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h61 == _T_37[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_7;
      end else if (8'h61 == _T_34[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_6;
      end else if (8'h61 == _T_31[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_5;
      end else if (8'h61 == _T_28[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_4;
      end else if (8'h61 == _T_25[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_3;
      end else if (8'h61 == _T_22[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_2;
      end else if (8'h61 == _T_19[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_1;
      end else if (8'h61 == _T_15[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_98 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h62 == _T_37[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_7;
      end else if (8'h62 == _T_34[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_6;
      end else if (8'h62 == _T_31[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_5;
      end else if (8'h62 == _T_28[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_4;
      end else if (8'h62 == _T_25[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_3;
      end else if (8'h62 == _T_22[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_2;
      end else if (8'h62 == _T_19[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_1;
      end else if (8'h62 == _T_15[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_99 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h63 == _T_37[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_7;
      end else if (8'h63 == _T_34[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_6;
      end else if (8'h63 == _T_31[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_5;
      end else if (8'h63 == _T_28[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_4;
      end else if (8'h63 == _T_25[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_3;
      end else if (8'h63 == _T_22[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_2;
      end else if (8'h63 == _T_19[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_1;
      end else if (8'h63 == _T_15[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_100 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h64 == _T_37[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_7;
      end else if (8'h64 == _T_34[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_6;
      end else if (8'h64 == _T_31[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_5;
      end else if (8'h64 == _T_28[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_4;
      end else if (8'h64 == _T_25[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_3;
      end else if (8'h64 == _T_22[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_2;
      end else if (8'h64 == _T_19[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_1;
      end else if (8'h64 == _T_15[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_101 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h65 == _T_37[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_7;
      end else if (8'h65 == _T_34[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_6;
      end else if (8'h65 == _T_31[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_5;
      end else if (8'h65 == _T_28[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_4;
      end else if (8'h65 == _T_25[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_3;
      end else if (8'h65 == _T_22[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_2;
      end else if (8'h65 == _T_19[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_1;
      end else if (8'h65 == _T_15[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_102 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h66 == _T_37[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_7;
      end else if (8'h66 == _T_34[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_6;
      end else if (8'h66 == _T_31[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_5;
      end else if (8'h66 == _T_28[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_4;
      end else if (8'h66 == _T_25[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_3;
      end else if (8'h66 == _T_22[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_2;
      end else if (8'h66 == _T_19[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_1;
      end else if (8'h66 == _T_15[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_103 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h67 == _T_37[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_7;
      end else if (8'h67 == _T_34[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_6;
      end else if (8'h67 == _T_31[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_5;
      end else if (8'h67 == _T_28[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_4;
      end else if (8'h67 == _T_25[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_3;
      end else if (8'h67 == _T_22[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_2;
      end else if (8'h67 == _T_19[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_1;
      end else if (8'h67 == _T_15[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_104 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h68 == _T_37[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_7;
      end else if (8'h68 == _T_34[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_6;
      end else if (8'h68 == _T_31[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_5;
      end else if (8'h68 == _T_28[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_4;
      end else if (8'h68 == _T_25[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_3;
      end else if (8'h68 == _T_22[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_2;
      end else if (8'h68 == _T_19[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_1;
      end else if (8'h68 == _T_15[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_105 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h69 == _T_37[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_7;
      end else if (8'h69 == _T_34[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_6;
      end else if (8'h69 == _T_31[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_5;
      end else if (8'h69 == _T_28[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_4;
      end else if (8'h69 == _T_25[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_3;
      end else if (8'h69 == _T_22[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_2;
      end else if (8'h69 == _T_19[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_1;
      end else if (8'h69 == _T_15[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_106 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6a == _T_37[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_7;
      end else if (8'h6a == _T_34[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_6;
      end else if (8'h6a == _T_31[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_5;
      end else if (8'h6a == _T_28[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_4;
      end else if (8'h6a == _T_25[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_3;
      end else if (8'h6a == _T_22[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_2;
      end else if (8'h6a == _T_19[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_1;
      end else if (8'h6a == _T_15[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_107 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6b == _T_37[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_7;
      end else if (8'h6b == _T_34[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_6;
      end else if (8'h6b == _T_31[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_5;
      end else if (8'h6b == _T_28[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_4;
      end else if (8'h6b == _T_25[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_3;
      end else if (8'h6b == _T_22[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_2;
      end else if (8'h6b == _T_19[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_1;
      end else if (8'h6b == _T_15[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_108 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6c == _T_37[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_7;
      end else if (8'h6c == _T_34[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_6;
      end else if (8'h6c == _T_31[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_5;
      end else if (8'h6c == _T_28[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_4;
      end else if (8'h6c == _T_25[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_3;
      end else if (8'h6c == _T_22[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_2;
      end else if (8'h6c == _T_19[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_1;
      end else if (8'h6c == _T_15[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_109 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6d == _T_37[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_7;
      end else if (8'h6d == _T_34[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_6;
      end else if (8'h6d == _T_31[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_5;
      end else if (8'h6d == _T_28[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_4;
      end else if (8'h6d == _T_25[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_3;
      end else if (8'h6d == _T_22[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_2;
      end else if (8'h6d == _T_19[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_1;
      end else if (8'h6d == _T_15[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_110 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6e == _T_37[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_7;
      end else if (8'h6e == _T_34[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_6;
      end else if (8'h6e == _T_31[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_5;
      end else if (8'h6e == _T_28[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_4;
      end else if (8'h6e == _T_25[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_3;
      end else if (8'h6e == _T_22[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_2;
      end else if (8'h6e == _T_19[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_1;
      end else if (8'h6e == _T_15[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_111 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6f == _T_37[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_7;
      end else if (8'h6f == _T_34[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_6;
      end else if (8'h6f == _T_31[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_5;
      end else if (8'h6f == _T_28[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_4;
      end else if (8'h6f == _T_25[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_3;
      end else if (8'h6f == _T_22[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_2;
      end else if (8'h6f == _T_19[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_1;
      end else if (8'h6f == _T_15[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_112 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h70 == _T_37[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_7;
      end else if (8'h70 == _T_34[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_6;
      end else if (8'h70 == _T_31[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_5;
      end else if (8'h70 == _T_28[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_4;
      end else if (8'h70 == _T_25[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_3;
      end else if (8'h70 == _T_22[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_2;
      end else if (8'h70 == _T_19[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_1;
      end else if (8'h70 == _T_15[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_113 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h71 == _T_37[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_7;
      end else if (8'h71 == _T_34[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_6;
      end else if (8'h71 == _T_31[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_5;
      end else if (8'h71 == _T_28[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_4;
      end else if (8'h71 == _T_25[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_3;
      end else if (8'h71 == _T_22[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_2;
      end else if (8'h71 == _T_19[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_1;
      end else if (8'h71 == _T_15[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_114 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h72 == _T_37[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_7;
      end else if (8'h72 == _T_34[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_6;
      end else if (8'h72 == _T_31[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_5;
      end else if (8'h72 == _T_28[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_4;
      end else if (8'h72 == _T_25[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_3;
      end else if (8'h72 == _T_22[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_2;
      end else if (8'h72 == _T_19[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_1;
      end else if (8'h72 == _T_15[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_115 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h73 == _T_37[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_7;
      end else if (8'h73 == _T_34[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_6;
      end else if (8'h73 == _T_31[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_5;
      end else if (8'h73 == _T_28[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_4;
      end else if (8'h73 == _T_25[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_3;
      end else if (8'h73 == _T_22[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_2;
      end else if (8'h73 == _T_19[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_1;
      end else if (8'h73 == _T_15[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_116 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h74 == _T_37[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_7;
      end else if (8'h74 == _T_34[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_6;
      end else if (8'h74 == _T_31[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_5;
      end else if (8'h74 == _T_28[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_4;
      end else if (8'h74 == _T_25[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_3;
      end else if (8'h74 == _T_22[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_2;
      end else if (8'h74 == _T_19[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_1;
      end else if (8'h74 == _T_15[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_117 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h75 == _T_37[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_7;
      end else if (8'h75 == _T_34[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_6;
      end else if (8'h75 == _T_31[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_5;
      end else if (8'h75 == _T_28[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_4;
      end else if (8'h75 == _T_25[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_3;
      end else if (8'h75 == _T_22[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_2;
      end else if (8'h75 == _T_19[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_1;
      end else if (8'h75 == _T_15[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_118 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h76 == _T_37[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_7;
      end else if (8'h76 == _T_34[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_6;
      end else if (8'h76 == _T_31[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_5;
      end else if (8'h76 == _T_28[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_4;
      end else if (8'h76 == _T_25[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_3;
      end else if (8'h76 == _T_22[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_2;
      end else if (8'h76 == _T_19[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_1;
      end else if (8'h76 == _T_15[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_119 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h77 == _T_37[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_7;
      end else if (8'h77 == _T_34[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_6;
      end else if (8'h77 == _T_31[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_5;
      end else if (8'h77 == _T_28[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_4;
      end else if (8'h77 == _T_25[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_3;
      end else if (8'h77 == _T_22[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_2;
      end else if (8'h77 == _T_19[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_1;
      end else if (8'h77 == _T_15[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_120 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h78 == _T_37[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_7;
      end else if (8'h78 == _T_34[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_6;
      end else if (8'h78 == _T_31[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_5;
      end else if (8'h78 == _T_28[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_4;
      end else if (8'h78 == _T_25[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_3;
      end else if (8'h78 == _T_22[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_2;
      end else if (8'h78 == _T_19[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_1;
      end else if (8'h78 == _T_15[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_121 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h79 == _T_37[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_7;
      end else if (8'h79 == _T_34[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_6;
      end else if (8'h79 == _T_31[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_5;
      end else if (8'h79 == _T_28[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_4;
      end else if (8'h79 == _T_25[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_3;
      end else if (8'h79 == _T_22[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_2;
      end else if (8'h79 == _T_19[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_1;
      end else if (8'h79 == _T_15[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_122 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7a == _T_37[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_7;
      end else if (8'h7a == _T_34[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_6;
      end else if (8'h7a == _T_31[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_5;
      end else if (8'h7a == _T_28[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_4;
      end else if (8'h7a == _T_25[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_3;
      end else if (8'h7a == _T_22[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_2;
      end else if (8'h7a == _T_19[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_1;
      end else if (8'h7a == _T_15[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_123 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7b == _T_37[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_7;
      end else if (8'h7b == _T_34[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_6;
      end else if (8'h7b == _T_31[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_5;
      end else if (8'h7b == _T_28[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_4;
      end else if (8'h7b == _T_25[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_3;
      end else if (8'h7b == _T_22[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_2;
      end else if (8'h7b == _T_19[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_1;
      end else if (8'h7b == _T_15[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_124 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7c == _T_37[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_7;
      end else if (8'h7c == _T_34[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_6;
      end else if (8'h7c == _T_31[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_5;
      end else if (8'h7c == _T_28[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_4;
      end else if (8'h7c == _T_25[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_3;
      end else if (8'h7c == _T_22[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_2;
      end else if (8'h7c == _T_19[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_1;
      end else if (8'h7c == _T_15[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_125 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7d == _T_37[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_7;
      end else if (8'h7d == _T_34[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_6;
      end else if (8'h7d == _T_31[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_5;
      end else if (8'h7d == _T_28[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_4;
      end else if (8'h7d == _T_25[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_3;
      end else if (8'h7d == _T_22[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_2;
      end else if (8'h7d == _T_19[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_1;
      end else if (8'h7d == _T_15[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_126 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7e == _T_37[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_7;
      end else if (8'h7e == _T_34[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_6;
      end else if (8'h7e == _T_31[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_5;
      end else if (8'h7e == _T_28[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_4;
      end else if (8'h7e == _T_25[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_3;
      end else if (8'h7e == _T_22[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_2;
      end else if (8'h7e == _T_19[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_1;
      end else if (8'h7e == _T_15[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_127 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7f == _T_37[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_7;
      end else if (8'h7f == _T_34[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_6;
      end else if (8'h7f == _T_31[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_5;
      end else if (8'h7f == _T_28[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_4;
      end else if (8'h7f == _T_25[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_3;
      end else if (8'h7f == _T_22[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_2;
      end else if (8'h7f == _T_19[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_1;
      end else if (8'h7f == _T_15[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_128 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h80 == _T_37[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_7;
      end else if (8'h80 == _T_34[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_6;
      end else if (8'h80 == _T_31[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_5;
      end else if (8'h80 == _T_28[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_4;
      end else if (8'h80 == _T_25[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_3;
      end else if (8'h80 == _T_22[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_2;
      end else if (8'h80 == _T_19[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_1;
      end else if (8'h80 == _T_15[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_129 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h81 == _T_37[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_7;
      end else if (8'h81 == _T_34[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_6;
      end else if (8'h81 == _T_31[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_5;
      end else if (8'h81 == _T_28[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_4;
      end else if (8'h81 == _T_25[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_3;
      end else if (8'h81 == _T_22[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_2;
      end else if (8'h81 == _T_19[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_1;
      end else if (8'h81 == _T_15[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_130 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h82 == _T_37[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_7;
      end else if (8'h82 == _T_34[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_6;
      end else if (8'h82 == _T_31[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_5;
      end else if (8'h82 == _T_28[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_4;
      end else if (8'h82 == _T_25[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_3;
      end else if (8'h82 == _T_22[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_2;
      end else if (8'h82 == _T_19[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_1;
      end else if (8'h82 == _T_15[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_131 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h83 == _T_37[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_7;
      end else if (8'h83 == _T_34[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_6;
      end else if (8'h83 == _T_31[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_5;
      end else if (8'h83 == _T_28[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_4;
      end else if (8'h83 == _T_25[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_3;
      end else if (8'h83 == _T_22[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_2;
      end else if (8'h83 == _T_19[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_1;
      end else if (8'h83 == _T_15[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_132 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h84 == _T_37[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_7;
      end else if (8'h84 == _T_34[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_6;
      end else if (8'h84 == _T_31[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_5;
      end else if (8'h84 == _T_28[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_4;
      end else if (8'h84 == _T_25[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_3;
      end else if (8'h84 == _T_22[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_2;
      end else if (8'h84 == _T_19[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_1;
      end else if (8'h84 == _T_15[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_133 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h85 == _T_37[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_7;
      end else if (8'h85 == _T_34[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_6;
      end else if (8'h85 == _T_31[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_5;
      end else if (8'h85 == _T_28[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_4;
      end else if (8'h85 == _T_25[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_3;
      end else if (8'h85 == _T_22[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_2;
      end else if (8'h85 == _T_19[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_1;
      end else if (8'h85 == _T_15[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_134 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h86 == _T_37[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_7;
      end else if (8'h86 == _T_34[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_6;
      end else if (8'h86 == _T_31[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_5;
      end else if (8'h86 == _T_28[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_4;
      end else if (8'h86 == _T_25[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_3;
      end else if (8'h86 == _T_22[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_2;
      end else if (8'h86 == _T_19[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_1;
      end else if (8'h86 == _T_15[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_135 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h87 == _T_37[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_7;
      end else if (8'h87 == _T_34[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_6;
      end else if (8'h87 == _T_31[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_5;
      end else if (8'h87 == _T_28[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_4;
      end else if (8'h87 == _T_25[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_3;
      end else if (8'h87 == _T_22[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_2;
      end else if (8'h87 == _T_19[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_1;
      end else if (8'h87 == _T_15[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_136 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h88 == _T_37[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_7;
      end else if (8'h88 == _T_34[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_6;
      end else if (8'h88 == _T_31[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_5;
      end else if (8'h88 == _T_28[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_4;
      end else if (8'h88 == _T_25[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_3;
      end else if (8'h88 == _T_22[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_2;
      end else if (8'h88 == _T_19[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_1;
      end else if (8'h88 == _T_15[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_137 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h89 == _T_37[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_7;
      end else if (8'h89 == _T_34[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_6;
      end else if (8'h89 == _T_31[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_5;
      end else if (8'h89 == _T_28[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_4;
      end else if (8'h89 == _T_25[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_3;
      end else if (8'h89 == _T_22[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_2;
      end else if (8'h89 == _T_19[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_1;
      end else if (8'h89 == _T_15[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_138 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8a == _T_37[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_7;
      end else if (8'h8a == _T_34[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_6;
      end else if (8'h8a == _T_31[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_5;
      end else if (8'h8a == _T_28[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_4;
      end else if (8'h8a == _T_25[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_3;
      end else if (8'h8a == _T_22[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_2;
      end else if (8'h8a == _T_19[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_1;
      end else if (8'h8a == _T_15[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_139 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8b == _T_37[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_7;
      end else if (8'h8b == _T_34[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_6;
      end else if (8'h8b == _T_31[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_5;
      end else if (8'h8b == _T_28[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_4;
      end else if (8'h8b == _T_25[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_3;
      end else if (8'h8b == _T_22[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_2;
      end else if (8'h8b == _T_19[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_1;
      end else if (8'h8b == _T_15[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_140 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8c == _T_37[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_7;
      end else if (8'h8c == _T_34[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_6;
      end else if (8'h8c == _T_31[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_5;
      end else if (8'h8c == _T_28[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_4;
      end else if (8'h8c == _T_25[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_3;
      end else if (8'h8c == _T_22[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_2;
      end else if (8'h8c == _T_19[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_1;
      end else if (8'h8c == _T_15[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_141 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8d == _T_37[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_7;
      end else if (8'h8d == _T_34[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_6;
      end else if (8'h8d == _T_31[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_5;
      end else if (8'h8d == _T_28[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_4;
      end else if (8'h8d == _T_25[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_3;
      end else if (8'h8d == _T_22[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_2;
      end else if (8'h8d == _T_19[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_1;
      end else if (8'h8d == _T_15[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_142 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8e == _T_37[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_7;
      end else if (8'h8e == _T_34[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_6;
      end else if (8'h8e == _T_31[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_5;
      end else if (8'h8e == _T_28[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_4;
      end else if (8'h8e == _T_25[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_3;
      end else if (8'h8e == _T_22[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_2;
      end else if (8'h8e == _T_19[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_1;
      end else if (8'h8e == _T_15[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_143 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8f == _T_37[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_7;
      end else if (8'h8f == _T_34[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_6;
      end else if (8'h8f == _T_31[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_5;
      end else if (8'h8f == _T_28[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_4;
      end else if (8'h8f == _T_25[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_3;
      end else if (8'h8f == _T_22[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_2;
      end else if (8'h8f == _T_19[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_1;
      end else if (8'h8f == _T_15[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_144 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h90 == _T_37[7:0]) begin
        image_0_144 <= io_pixelVal_in_0_7;
      end else if (8'h90 == _T_34[7:0]) begin
        image_0_144 <= io_pixelVal_in_0_6;
      end else if (8'h90 == _T_31[7:0]) begin
        image_0_144 <= io_pixelVal_in_0_5;
      end else if (8'h90 == _T_28[7:0]) begin
        image_0_144 <= io_pixelVal_in_0_4;
      end else if (8'h90 == _T_25[7:0]) begin
        image_0_144 <= io_pixelVal_in_0_3;
      end else if (8'h90 == _T_22[7:0]) begin
        image_0_144 <= io_pixelVal_in_0_2;
      end else if (8'h90 == _T_19[7:0]) begin
        image_0_144 <= io_pixelVal_in_0_1;
      end else if (8'h90 == _T_15[7:0]) begin
        image_0_144 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_145 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h91 == _T_37[7:0]) begin
        image_0_145 <= io_pixelVal_in_0_7;
      end else if (8'h91 == _T_34[7:0]) begin
        image_0_145 <= io_pixelVal_in_0_6;
      end else if (8'h91 == _T_31[7:0]) begin
        image_0_145 <= io_pixelVal_in_0_5;
      end else if (8'h91 == _T_28[7:0]) begin
        image_0_145 <= io_pixelVal_in_0_4;
      end else if (8'h91 == _T_25[7:0]) begin
        image_0_145 <= io_pixelVal_in_0_3;
      end else if (8'h91 == _T_22[7:0]) begin
        image_0_145 <= io_pixelVal_in_0_2;
      end else if (8'h91 == _T_19[7:0]) begin
        image_0_145 <= io_pixelVal_in_0_1;
      end else if (8'h91 == _T_15[7:0]) begin
        image_0_145 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_146 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h92 == _T_37[7:0]) begin
        image_0_146 <= io_pixelVal_in_0_7;
      end else if (8'h92 == _T_34[7:0]) begin
        image_0_146 <= io_pixelVal_in_0_6;
      end else if (8'h92 == _T_31[7:0]) begin
        image_0_146 <= io_pixelVal_in_0_5;
      end else if (8'h92 == _T_28[7:0]) begin
        image_0_146 <= io_pixelVal_in_0_4;
      end else if (8'h92 == _T_25[7:0]) begin
        image_0_146 <= io_pixelVal_in_0_3;
      end else if (8'h92 == _T_22[7:0]) begin
        image_0_146 <= io_pixelVal_in_0_2;
      end else if (8'h92 == _T_19[7:0]) begin
        image_0_146 <= io_pixelVal_in_0_1;
      end else if (8'h92 == _T_15[7:0]) begin
        image_0_146 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_147 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h93 == _T_37[7:0]) begin
        image_0_147 <= io_pixelVal_in_0_7;
      end else if (8'h93 == _T_34[7:0]) begin
        image_0_147 <= io_pixelVal_in_0_6;
      end else if (8'h93 == _T_31[7:0]) begin
        image_0_147 <= io_pixelVal_in_0_5;
      end else if (8'h93 == _T_28[7:0]) begin
        image_0_147 <= io_pixelVal_in_0_4;
      end else if (8'h93 == _T_25[7:0]) begin
        image_0_147 <= io_pixelVal_in_0_3;
      end else if (8'h93 == _T_22[7:0]) begin
        image_0_147 <= io_pixelVal_in_0_2;
      end else if (8'h93 == _T_19[7:0]) begin
        image_0_147 <= io_pixelVal_in_0_1;
      end else if (8'h93 == _T_15[7:0]) begin
        image_0_147 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_148 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h94 == _T_37[7:0]) begin
        image_0_148 <= io_pixelVal_in_0_7;
      end else if (8'h94 == _T_34[7:0]) begin
        image_0_148 <= io_pixelVal_in_0_6;
      end else if (8'h94 == _T_31[7:0]) begin
        image_0_148 <= io_pixelVal_in_0_5;
      end else if (8'h94 == _T_28[7:0]) begin
        image_0_148 <= io_pixelVal_in_0_4;
      end else if (8'h94 == _T_25[7:0]) begin
        image_0_148 <= io_pixelVal_in_0_3;
      end else if (8'h94 == _T_22[7:0]) begin
        image_0_148 <= io_pixelVal_in_0_2;
      end else if (8'h94 == _T_19[7:0]) begin
        image_0_148 <= io_pixelVal_in_0_1;
      end else if (8'h94 == _T_15[7:0]) begin
        image_0_148 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_149 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h95 == _T_37[7:0]) begin
        image_0_149 <= io_pixelVal_in_0_7;
      end else if (8'h95 == _T_34[7:0]) begin
        image_0_149 <= io_pixelVal_in_0_6;
      end else if (8'h95 == _T_31[7:0]) begin
        image_0_149 <= io_pixelVal_in_0_5;
      end else if (8'h95 == _T_28[7:0]) begin
        image_0_149 <= io_pixelVal_in_0_4;
      end else if (8'h95 == _T_25[7:0]) begin
        image_0_149 <= io_pixelVal_in_0_3;
      end else if (8'h95 == _T_22[7:0]) begin
        image_0_149 <= io_pixelVal_in_0_2;
      end else if (8'h95 == _T_19[7:0]) begin
        image_0_149 <= io_pixelVal_in_0_1;
      end else if (8'h95 == _T_15[7:0]) begin
        image_0_149 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_150 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h96 == _T_37[7:0]) begin
        image_0_150 <= io_pixelVal_in_0_7;
      end else if (8'h96 == _T_34[7:0]) begin
        image_0_150 <= io_pixelVal_in_0_6;
      end else if (8'h96 == _T_31[7:0]) begin
        image_0_150 <= io_pixelVal_in_0_5;
      end else if (8'h96 == _T_28[7:0]) begin
        image_0_150 <= io_pixelVal_in_0_4;
      end else if (8'h96 == _T_25[7:0]) begin
        image_0_150 <= io_pixelVal_in_0_3;
      end else if (8'h96 == _T_22[7:0]) begin
        image_0_150 <= io_pixelVal_in_0_2;
      end else if (8'h96 == _T_19[7:0]) begin
        image_0_150 <= io_pixelVal_in_0_1;
      end else if (8'h96 == _T_15[7:0]) begin
        image_0_150 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_151 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h97 == _T_37[7:0]) begin
        image_0_151 <= io_pixelVal_in_0_7;
      end else if (8'h97 == _T_34[7:0]) begin
        image_0_151 <= io_pixelVal_in_0_6;
      end else if (8'h97 == _T_31[7:0]) begin
        image_0_151 <= io_pixelVal_in_0_5;
      end else if (8'h97 == _T_28[7:0]) begin
        image_0_151 <= io_pixelVal_in_0_4;
      end else if (8'h97 == _T_25[7:0]) begin
        image_0_151 <= io_pixelVal_in_0_3;
      end else if (8'h97 == _T_22[7:0]) begin
        image_0_151 <= io_pixelVal_in_0_2;
      end else if (8'h97 == _T_19[7:0]) begin
        image_0_151 <= io_pixelVal_in_0_1;
      end else if (8'h97 == _T_15[7:0]) begin
        image_0_151 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_152 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h98 == _T_37[7:0]) begin
        image_0_152 <= io_pixelVal_in_0_7;
      end else if (8'h98 == _T_34[7:0]) begin
        image_0_152 <= io_pixelVal_in_0_6;
      end else if (8'h98 == _T_31[7:0]) begin
        image_0_152 <= io_pixelVal_in_0_5;
      end else if (8'h98 == _T_28[7:0]) begin
        image_0_152 <= io_pixelVal_in_0_4;
      end else if (8'h98 == _T_25[7:0]) begin
        image_0_152 <= io_pixelVal_in_0_3;
      end else if (8'h98 == _T_22[7:0]) begin
        image_0_152 <= io_pixelVal_in_0_2;
      end else if (8'h98 == _T_19[7:0]) begin
        image_0_152 <= io_pixelVal_in_0_1;
      end else if (8'h98 == _T_15[7:0]) begin
        image_0_152 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_153 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h99 == _T_37[7:0]) begin
        image_0_153 <= io_pixelVal_in_0_7;
      end else if (8'h99 == _T_34[7:0]) begin
        image_0_153 <= io_pixelVal_in_0_6;
      end else if (8'h99 == _T_31[7:0]) begin
        image_0_153 <= io_pixelVal_in_0_5;
      end else if (8'h99 == _T_28[7:0]) begin
        image_0_153 <= io_pixelVal_in_0_4;
      end else if (8'h99 == _T_25[7:0]) begin
        image_0_153 <= io_pixelVal_in_0_3;
      end else if (8'h99 == _T_22[7:0]) begin
        image_0_153 <= io_pixelVal_in_0_2;
      end else if (8'h99 == _T_19[7:0]) begin
        image_0_153 <= io_pixelVal_in_0_1;
      end else if (8'h99 == _T_15[7:0]) begin
        image_0_153 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_154 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h9a == _T_37[7:0]) begin
        image_0_154 <= io_pixelVal_in_0_7;
      end else if (8'h9a == _T_34[7:0]) begin
        image_0_154 <= io_pixelVal_in_0_6;
      end else if (8'h9a == _T_31[7:0]) begin
        image_0_154 <= io_pixelVal_in_0_5;
      end else if (8'h9a == _T_28[7:0]) begin
        image_0_154 <= io_pixelVal_in_0_4;
      end else if (8'h9a == _T_25[7:0]) begin
        image_0_154 <= io_pixelVal_in_0_3;
      end else if (8'h9a == _T_22[7:0]) begin
        image_0_154 <= io_pixelVal_in_0_2;
      end else if (8'h9a == _T_19[7:0]) begin
        image_0_154 <= io_pixelVal_in_0_1;
      end else if (8'h9a == _T_15[7:0]) begin
        image_0_154 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_155 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h9b == _T_37[7:0]) begin
        image_0_155 <= io_pixelVal_in_0_7;
      end else if (8'h9b == _T_34[7:0]) begin
        image_0_155 <= io_pixelVal_in_0_6;
      end else if (8'h9b == _T_31[7:0]) begin
        image_0_155 <= io_pixelVal_in_0_5;
      end else if (8'h9b == _T_28[7:0]) begin
        image_0_155 <= io_pixelVal_in_0_4;
      end else if (8'h9b == _T_25[7:0]) begin
        image_0_155 <= io_pixelVal_in_0_3;
      end else if (8'h9b == _T_22[7:0]) begin
        image_0_155 <= io_pixelVal_in_0_2;
      end else if (8'h9b == _T_19[7:0]) begin
        image_0_155 <= io_pixelVal_in_0_1;
      end else if (8'h9b == _T_15[7:0]) begin
        image_0_155 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_156 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h9c == _T_37[7:0]) begin
        image_0_156 <= io_pixelVal_in_0_7;
      end else if (8'h9c == _T_34[7:0]) begin
        image_0_156 <= io_pixelVal_in_0_6;
      end else if (8'h9c == _T_31[7:0]) begin
        image_0_156 <= io_pixelVal_in_0_5;
      end else if (8'h9c == _T_28[7:0]) begin
        image_0_156 <= io_pixelVal_in_0_4;
      end else if (8'h9c == _T_25[7:0]) begin
        image_0_156 <= io_pixelVal_in_0_3;
      end else if (8'h9c == _T_22[7:0]) begin
        image_0_156 <= io_pixelVal_in_0_2;
      end else if (8'h9c == _T_19[7:0]) begin
        image_0_156 <= io_pixelVal_in_0_1;
      end else if (8'h9c == _T_15[7:0]) begin
        image_0_156 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_157 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h9d == _T_37[7:0]) begin
        image_0_157 <= io_pixelVal_in_0_7;
      end else if (8'h9d == _T_34[7:0]) begin
        image_0_157 <= io_pixelVal_in_0_6;
      end else if (8'h9d == _T_31[7:0]) begin
        image_0_157 <= io_pixelVal_in_0_5;
      end else if (8'h9d == _T_28[7:0]) begin
        image_0_157 <= io_pixelVal_in_0_4;
      end else if (8'h9d == _T_25[7:0]) begin
        image_0_157 <= io_pixelVal_in_0_3;
      end else if (8'h9d == _T_22[7:0]) begin
        image_0_157 <= io_pixelVal_in_0_2;
      end else if (8'h9d == _T_19[7:0]) begin
        image_0_157 <= io_pixelVal_in_0_1;
      end else if (8'h9d == _T_15[7:0]) begin
        image_0_157 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_158 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h9e == _T_37[7:0]) begin
        image_0_158 <= io_pixelVal_in_0_7;
      end else if (8'h9e == _T_34[7:0]) begin
        image_0_158 <= io_pixelVal_in_0_6;
      end else if (8'h9e == _T_31[7:0]) begin
        image_0_158 <= io_pixelVal_in_0_5;
      end else if (8'h9e == _T_28[7:0]) begin
        image_0_158 <= io_pixelVal_in_0_4;
      end else if (8'h9e == _T_25[7:0]) begin
        image_0_158 <= io_pixelVal_in_0_3;
      end else if (8'h9e == _T_22[7:0]) begin
        image_0_158 <= io_pixelVal_in_0_2;
      end else if (8'h9e == _T_19[7:0]) begin
        image_0_158 <= io_pixelVal_in_0_1;
      end else if (8'h9e == _T_15[7:0]) begin
        image_0_158 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_159 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h9f == _T_37[7:0]) begin
        image_0_159 <= io_pixelVal_in_0_7;
      end else if (8'h9f == _T_34[7:0]) begin
        image_0_159 <= io_pixelVal_in_0_6;
      end else if (8'h9f == _T_31[7:0]) begin
        image_0_159 <= io_pixelVal_in_0_5;
      end else if (8'h9f == _T_28[7:0]) begin
        image_0_159 <= io_pixelVal_in_0_4;
      end else if (8'h9f == _T_25[7:0]) begin
        image_0_159 <= io_pixelVal_in_0_3;
      end else if (8'h9f == _T_22[7:0]) begin
        image_0_159 <= io_pixelVal_in_0_2;
      end else if (8'h9f == _T_19[7:0]) begin
        image_0_159 <= io_pixelVal_in_0_1;
      end else if (8'h9f == _T_15[7:0]) begin
        image_0_159 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_160 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha0 == _T_37[7:0]) begin
        image_0_160 <= io_pixelVal_in_0_7;
      end else if (8'ha0 == _T_34[7:0]) begin
        image_0_160 <= io_pixelVal_in_0_6;
      end else if (8'ha0 == _T_31[7:0]) begin
        image_0_160 <= io_pixelVal_in_0_5;
      end else if (8'ha0 == _T_28[7:0]) begin
        image_0_160 <= io_pixelVal_in_0_4;
      end else if (8'ha0 == _T_25[7:0]) begin
        image_0_160 <= io_pixelVal_in_0_3;
      end else if (8'ha0 == _T_22[7:0]) begin
        image_0_160 <= io_pixelVal_in_0_2;
      end else if (8'ha0 == _T_19[7:0]) begin
        image_0_160 <= io_pixelVal_in_0_1;
      end else if (8'ha0 == _T_15[7:0]) begin
        image_0_160 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_161 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha1 == _T_37[7:0]) begin
        image_0_161 <= io_pixelVal_in_0_7;
      end else if (8'ha1 == _T_34[7:0]) begin
        image_0_161 <= io_pixelVal_in_0_6;
      end else if (8'ha1 == _T_31[7:0]) begin
        image_0_161 <= io_pixelVal_in_0_5;
      end else if (8'ha1 == _T_28[7:0]) begin
        image_0_161 <= io_pixelVal_in_0_4;
      end else if (8'ha1 == _T_25[7:0]) begin
        image_0_161 <= io_pixelVal_in_0_3;
      end else if (8'ha1 == _T_22[7:0]) begin
        image_0_161 <= io_pixelVal_in_0_2;
      end else if (8'ha1 == _T_19[7:0]) begin
        image_0_161 <= io_pixelVal_in_0_1;
      end else if (8'ha1 == _T_15[7:0]) begin
        image_0_161 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_162 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha2 == _T_37[7:0]) begin
        image_0_162 <= io_pixelVal_in_0_7;
      end else if (8'ha2 == _T_34[7:0]) begin
        image_0_162 <= io_pixelVal_in_0_6;
      end else if (8'ha2 == _T_31[7:0]) begin
        image_0_162 <= io_pixelVal_in_0_5;
      end else if (8'ha2 == _T_28[7:0]) begin
        image_0_162 <= io_pixelVal_in_0_4;
      end else if (8'ha2 == _T_25[7:0]) begin
        image_0_162 <= io_pixelVal_in_0_3;
      end else if (8'ha2 == _T_22[7:0]) begin
        image_0_162 <= io_pixelVal_in_0_2;
      end else if (8'ha2 == _T_19[7:0]) begin
        image_0_162 <= io_pixelVal_in_0_1;
      end else if (8'ha2 == _T_15[7:0]) begin
        image_0_162 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_163 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha3 == _T_37[7:0]) begin
        image_0_163 <= io_pixelVal_in_0_7;
      end else if (8'ha3 == _T_34[7:0]) begin
        image_0_163 <= io_pixelVal_in_0_6;
      end else if (8'ha3 == _T_31[7:0]) begin
        image_0_163 <= io_pixelVal_in_0_5;
      end else if (8'ha3 == _T_28[7:0]) begin
        image_0_163 <= io_pixelVal_in_0_4;
      end else if (8'ha3 == _T_25[7:0]) begin
        image_0_163 <= io_pixelVal_in_0_3;
      end else if (8'ha3 == _T_22[7:0]) begin
        image_0_163 <= io_pixelVal_in_0_2;
      end else if (8'ha3 == _T_19[7:0]) begin
        image_0_163 <= io_pixelVal_in_0_1;
      end else if (8'ha3 == _T_15[7:0]) begin
        image_0_163 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_164 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha4 == _T_37[7:0]) begin
        image_0_164 <= io_pixelVal_in_0_7;
      end else if (8'ha4 == _T_34[7:0]) begin
        image_0_164 <= io_pixelVal_in_0_6;
      end else if (8'ha4 == _T_31[7:0]) begin
        image_0_164 <= io_pixelVal_in_0_5;
      end else if (8'ha4 == _T_28[7:0]) begin
        image_0_164 <= io_pixelVal_in_0_4;
      end else if (8'ha4 == _T_25[7:0]) begin
        image_0_164 <= io_pixelVal_in_0_3;
      end else if (8'ha4 == _T_22[7:0]) begin
        image_0_164 <= io_pixelVal_in_0_2;
      end else if (8'ha4 == _T_19[7:0]) begin
        image_0_164 <= io_pixelVal_in_0_1;
      end else if (8'ha4 == _T_15[7:0]) begin
        image_0_164 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_165 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha5 == _T_37[7:0]) begin
        image_0_165 <= io_pixelVal_in_0_7;
      end else if (8'ha5 == _T_34[7:0]) begin
        image_0_165 <= io_pixelVal_in_0_6;
      end else if (8'ha5 == _T_31[7:0]) begin
        image_0_165 <= io_pixelVal_in_0_5;
      end else if (8'ha5 == _T_28[7:0]) begin
        image_0_165 <= io_pixelVal_in_0_4;
      end else if (8'ha5 == _T_25[7:0]) begin
        image_0_165 <= io_pixelVal_in_0_3;
      end else if (8'ha5 == _T_22[7:0]) begin
        image_0_165 <= io_pixelVal_in_0_2;
      end else if (8'ha5 == _T_19[7:0]) begin
        image_0_165 <= io_pixelVal_in_0_1;
      end else if (8'ha5 == _T_15[7:0]) begin
        image_0_165 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_166 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha6 == _T_37[7:0]) begin
        image_0_166 <= io_pixelVal_in_0_7;
      end else if (8'ha6 == _T_34[7:0]) begin
        image_0_166 <= io_pixelVal_in_0_6;
      end else if (8'ha6 == _T_31[7:0]) begin
        image_0_166 <= io_pixelVal_in_0_5;
      end else if (8'ha6 == _T_28[7:0]) begin
        image_0_166 <= io_pixelVal_in_0_4;
      end else if (8'ha6 == _T_25[7:0]) begin
        image_0_166 <= io_pixelVal_in_0_3;
      end else if (8'ha6 == _T_22[7:0]) begin
        image_0_166 <= io_pixelVal_in_0_2;
      end else if (8'ha6 == _T_19[7:0]) begin
        image_0_166 <= io_pixelVal_in_0_1;
      end else if (8'ha6 == _T_15[7:0]) begin
        image_0_166 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_167 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha7 == _T_37[7:0]) begin
        image_0_167 <= io_pixelVal_in_0_7;
      end else if (8'ha7 == _T_34[7:0]) begin
        image_0_167 <= io_pixelVal_in_0_6;
      end else if (8'ha7 == _T_31[7:0]) begin
        image_0_167 <= io_pixelVal_in_0_5;
      end else if (8'ha7 == _T_28[7:0]) begin
        image_0_167 <= io_pixelVal_in_0_4;
      end else if (8'ha7 == _T_25[7:0]) begin
        image_0_167 <= io_pixelVal_in_0_3;
      end else if (8'ha7 == _T_22[7:0]) begin
        image_0_167 <= io_pixelVal_in_0_2;
      end else if (8'ha7 == _T_19[7:0]) begin
        image_0_167 <= io_pixelVal_in_0_1;
      end else if (8'ha7 == _T_15[7:0]) begin
        image_0_167 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_168 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha8 == _T_37[7:0]) begin
        image_0_168 <= io_pixelVal_in_0_7;
      end else if (8'ha8 == _T_34[7:0]) begin
        image_0_168 <= io_pixelVal_in_0_6;
      end else if (8'ha8 == _T_31[7:0]) begin
        image_0_168 <= io_pixelVal_in_0_5;
      end else if (8'ha8 == _T_28[7:0]) begin
        image_0_168 <= io_pixelVal_in_0_4;
      end else if (8'ha8 == _T_25[7:0]) begin
        image_0_168 <= io_pixelVal_in_0_3;
      end else if (8'ha8 == _T_22[7:0]) begin
        image_0_168 <= io_pixelVal_in_0_2;
      end else if (8'ha8 == _T_19[7:0]) begin
        image_0_168 <= io_pixelVal_in_0_1;
      end else if (8'ha8 == _T_15[7:0]) begin
        image_0_168 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_169 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha9 == _T_37[7:0]) begin
        image_0_169 <= io_pixelVal_in_0_7;
      end else if (8'ha9 == _T_34[7:0]) begin
        image_0_169 <= io_pixelVal_in_0_6;
      end else if (8'ha9 == _T_31[7:0]) begin
        image_0_169 <= io_pixelVal_in_0_5;
      end else if (8'ha9 == _T_28[7:0]) begin
        image_0_169 <= io_pixelVal_in_0_4;
      end else if (8'ha9 == _T_25[7:0]) begin
        image_0_169 <= io_pixelVal_in_0_3;
      end else if (8'ha9 == _T_22[7:0]) begin
        image_0_169 <= io_pixelVal_in_0_2;
      end else if (8'ha9 == _T_19[7:0]) begin
        image_0_169 <= io_pixelVal_in_0_1;
      end else if (8'ha9 == _T_15[7:0]) begin
        image_0_169 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_170 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'haa == _T_37[7:0]) begin
        image_0_170 <= io_pixelVal_in_0_7;
      end else if (8'haa == _T_34[7:0]) begin
        image_0_170 <= io_pixelVal_in_0_6;
      end else if (8'haa == _T_31[7:0]) begin
        image_0_170 <= io_pixelVal_in_0_5;
      end else if (8'haa == _T_28[7:0]) begin
        image_0_170 <= io_pixelVal_in_0_4;
      end else if (8'haa == _T_25[7:0]) begin
        image_0_170 <= io_pixelVal_in_0_3;
      end else if (8'haa == _T_22[7:0]) begin
        image_0_170 <= io_pixelVal_in_0_2;
      end else if (8'haa == _T_19[7:0]) begin
        image_0_170 <= io_pixelVal_in_0_1;
      end else if (8'haa == _T_15[7:0]) begin
        image_0_170 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_171 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hab == _T_37[7:0]) begin
        image_0_171 <= io_pixelVal_in_0_7;
      end else if (8'hab == _T_34[7:0]) begin
        image_0_171 <= io_pixelVal_in_0_6;
      end else if (8'hab == _T_31[7:0]) begin
        image_0_171 <= io_pixelVal_in_0_5;
      end else if (8'hab == _T_28[7:0]) begin
        image_0_171 <= io_pixelVal_in_0_4;
      end else if (8'hab == _T_25[7:0]) begin
        image_0_171 <= io_pixelVal_in_0_3;
      end else if (8'hab == _T_22[7:0]) begin
        image_0_171 <= io_pixelVal_in_0_2;
      end else if (8'hab == _T_19[7:0]) begin
        image_0_171 <= io_pixelVal_in_0_1;
      end else if (8'hab == _T_15[7:0]) begin
        image_0_171 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_172 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hac == _T_37[7:0]) begin
        image_0_172 <= io_pixelVal_in_0_7;
      end else if (8'hac == _T_34[7:0]) begin
        image_0_172 <= io_pixelVal_in_0_6;
      end else if (8'hac == _T_31[7:0]) begin
        image_0_172 <= io_pixelVal_in_0_5;
      end else if (8'hac == _T_28[7:0]) begin
        image_0_172 <= io_pixelVal_in_0_4;
      end else if (8'hac == _T_25[7:0]) begin
        image_0_172 <= io_pixelVal_in_0_3;
      end else if (8'hac == _T_22[7:0]) begin
        image_0_172 <= io_pixelVal_in_0_2;
      end else if (8'hac == _T_19[7:0]) begin
        image_0_172 <= io_pixelVal_in_0_1;
      end else if (8'hac == _T_15[7:0]) begin
        image_0_172 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_173 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'had == _T_37[7:0]) begin
        image_0_173 <= io_pixelVal_in_0_7;
      end else if (8'had == _T_34[7:0]) begin
        image_0_173 <= io_pixelVal_in_0_6;
      end else if (8'had == _T_31[7:0]) begin
        image_0_173 <= io_pixelVal_in_0_5;
      end else if (8'had == _T_28[7:0]) begin
        image_0_173 <= io_pixelVal_in_0_4;
      end else if (8'had == _T_25[7:0]) begin
        image_0_173 <= io_pixelVal_in_0_3;
      end else if (8'had == _T_22[7:0]) begin
        image_0_173 <= io_pixelVal_in_0_2;
      end else if (8'had == _T_19[7:0]) begin
        image_0_173 <= io_pixelVal_in_0_1;
      end else if (8'had == _T_15[7:0]) begin
        image_0_173 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_174 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hae == _T_37[7:0]) begin
        image_0_174 <= io_pixelVal_in_0_7;
      end else if (8'hae == _T_34[7:0]) begin
        image_0_174 <= io_pixelVal_in_0_6;
      end else if (8'hae == _T_31[7:0]) begin
        image_0_174 <= io_pixelVal_in_0_5;
      end else if (8'hae == _T_28[7:0]) begin
        image_0_174 <= io_pixelVal_in_0_4;
      end else if (8'hae == _T_25[7:0]) begin
        image_0_174 <= io_pixelVal_in_0_3;
      end else if (8'hae == _T_22[7:0]) begin
        image_0_174 <= io_pixelVal_in_0_2;
      end else if (8'hae == _T_19[7:0]) begin
        image_0_174 <= io_pixelVal_in_0_1;
      end else if (8'hae == _T_15[7:0]) begin
        image_0_174 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_175 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'haf == _T_37[7:0]) begin
        image_0_175 <= io_pixelVal_in_0_7;
      end else if (8'haf == _T_34[7:0]) begin
        image_0_175 <= io_pixelVal_in_0_6;
      end else if (8'haf == _T_31[7:0]) begin
        image_0_175 <= io_pixelVal_in_0_5;
      end else if (8'haf == _T_28[7:0]) begin
        image_0_175 <= io_pixelVal_in_0_4;
      end else if (8'haf == _T_25[7:0]) begin
        image_0_175 <= io_pixelVal_in_0_3;
      end else if (8'haf == _T_22[7:0]) begin
        image_0_175 <= io_pixelVal_in_0_2;
      end else if (8'haf == _T_19[7:0]) begin
        image_0_175 <= io_pixelVal_in_0_1;
      end else if (8'haf == _T_15[7:0]) begin
        image_0_175 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_176 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb0 == _T_37[7:0]) begin
        image_0_176 <= io_pixelVal_in_0_7;
      end else if (8'hb0 == _T_34[7:0]) begin
        image_0_176 <= io_pixelVal_in_0_6;
      end else if (8'hb0 == _T_31[7:0]) begin
        image_0_176 <= io_pixelVal_in_0_5;
      end else if (8'hb0 == _T_28[7:0]) begin
        image_0_176 <= io_pixelVal_in_0_4;
      end else if (8'hb0 == _T_25[7:0]) begin
        image_0_176 <= io_pixelVal_in_0_3;
      end else if (8'hb0 == _T_22[7:0]) begin
        image_0_176 <= io_pixelVal_in_0_2;
      end else if (8'hb0 == _T_19[7:0]) begin
        image_0_176 <= io_pixelVal_in_0_1;
      end else if (8'hb0 == _T_15[7:0]) begin
        image_0_176 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_177 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb1 == _T_37[7:0]) begin
        image_0_177 <= io_pixelVal_in_0_7;
      end else if (8'hb1 == _T_34[7:0]) begin
        image_0_177 <= io_pixelVal_in_0_6;
      end else if (8'hb1 == _T_31[7:0]) begin
        image_0_177 <= io_pixelVal_in_0_5;
      end else if (8'hb1 == _T_28[7:0]) begin
        image_0_177 <= io_pixelVal_in_0_4;
      end else if (8'hb1 == _T_25[7:0]) begin
        image_0_177 <= io_pixelVal_in_0_3;
      end else if (8'hb1 == _T_22[7:0]) begin
        image_0_177 <= io_pixelVal_in_0_2;
      end else if (8'hb1 == _T_19[7:0]) begin
        image_0_177 <= io_pixelVal_in_0_1;
      end else if (8'hb1 == _T_15[7:0]) begin
        image_0_177 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_178 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb2 == _T_37[7:0]) begin
        image_0_178 <= io_pixelVal_in_0_7;
      end else if (8'hb2 == _T_34[7:0]) begin
        image_0_178 <= io_pixelVal_in_0_6;
      end else if (8'hb2 == _T_31[7:0]) begin
        image_0_178 <= io_pixelVal_in_0_5;
      end else if (8'hb2 == _T_28[7:0]) begin
        image_0_178 <= io_pixelVal_in_0_4;
      end else if (8'hb2 == _T_25[7:0]) begin
        image_0_178 <= io_pixelVal_in_0_3;
      end else if (8'hb2 == _T_22[7:0]) begin
        image_0_178 <= io_pixelVal_in_0_2;
      end else if (8'hb2 == _T_19[7:0]) begin
        image_0_178 <= io_pixelVal_in_0_1;
      end else if (8'hb2 == _T_15[7:0]) begin
        image_0_178 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_179 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb3 == _T_37[7:0]) begin
        image_0_179 <= io_pixelVal_in_0_7;
      end else if (8'hb3 == _T_34[7:0]) begin
        image_0_179 <= io_pixelVal_in_0_6;
      end else if (8'hb3 == _T_31[7:0]) begin
        image_0_179 <= io_pixelVal_in_0_5;
      end else if (8'hb3 == _T_28[7:0]) begin
        image_0_179 <= io_pixelVal_in_0_4;
      end else if (8'hb3 == _T_25[7:0]) begin
        image_0_179 <= io_pixelVal_in_0_3;
      end else if (8'hb3 == _T_22[7:0]) begin
        image_0_179 <= io_pixelVal_in_0_2;
      end else if (8'hb3 == _T_19[7:0]) begin
        image_0_179 <= io_pixelVal_in_0_1;
      end else if (8'hb3 == _T_15[7:0]) begin
        image_0_179 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_180 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb4 == _T_37[7:0]) begin
        image_0_180 <= io_pixelVal_in_0_7;
      end else if (8'hb4 == _T_34[7:0]) begin
        image_0_180 <= io_pixelVal_in_0_6;
      end else if (8'hb4 == _T_31[7:0]) begin
        image_0_180 <= io_pixelVal_in_0_5;
      end else if (8'hb4 == _T_28[7:0]) begin
        image_0_180 <= io_pixelVal_in_0_4;
      end else if (8'hb4 == _T_25[7:0]) begin
        image_0_180 <= io_pixelVal_in_0_3;
      end else if (8'hb4 == _T_22[7:0]) begin
        image_0_180 <= io_pixelVal_in_0_2;
      end else if (8'hb4 == _T_19[7:0]) begin
        image_0_180 <= io_pixelVal_in_0_1;
      end else if (8'hb4 == _T_15[7:0]) begin
        image_0_180 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_181 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb5 == _T_37[7:0]) begin
        image_0_181 <= io_pixelVal_in_0_7;
      end else if (8'hb5 == _T_34[7:0]) begin
        image_0_181 <= io_pixelVal_in_0_6;
      end else if (8'hb5 == _T_31[7:0]) begin
        image_0_181 <= io_pixelVal_in_0_5;
      end else if (8'hb5 == _T_28[7:0]) begin
        image_0_181 <= io_pixelVal_in_0_4;
      end else if (8'hb5 == _T_25[7:0]) begin
        image_0_181 <= io_pixelVal_in_0_3;
      end else if (8'hb5 == _T_22[7:0]) begin
        image_0_181 <= io_pixelVal_in_0_2;
      end else if (8'hb5 == _T_19[7:0]) begin
        image_0_181 <= io_pixelVal_in_0_1;
      end else if (8'hb5 == _T_15[7:0]) begin
        image_0_181 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_182 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb6 == _T_37[7:0]) begin
        image_0_182 <= io_pixelVal_in_0_7;
      end else if (8'hb6 == _T_34[7:0]) begin
        image_0_182 <= io_pixelVal_in_0_6;
      end else if (8'hb6 == _T_31[7:0]) begin
        image_0_182 <= io_pixelVal_in_0_5;
      end else if (8'hb6 == _T_28[7:0]) begin
        image_0_182 <= io_pixelVal_in_0_4;
      end else if (8'hb6 == _T_25[7:0]) begin
        image_0_182 <= io_pixelVal_in_0_3;
      end else if (8'hb6 == _T_22[7:0]) begin
        image_0_182 <= io_pixelVal_in_0_2;
      end else if (8'hb6 == _T_19[7:0]) begin
        image_0_182 <= io_pixelVal_in_0_1;
      end else if (8'hb6 == _T_15[7:0]) begin
        image_0_182 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_183 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb7 == _T_37[7:0]) begin
        image_0_183 <= io_pixelVal_in_0_7;
      end else if (8'hb7 == _T_34[7:0]) begin
        image_0_183 <= io_pixelVal_in_0_6;
      end else if (8'hb7 == _T_31[7:0]) begin
        image_0_183 <= io_pixelVal_in_0_5;
      end else if (8'hb7 == _T_28[7:0]) begin
        image_0_183 <= io_pixelVal_in_0_4;
      end else if (8'hb7 == _T_25[7:0]) begin
        image_0_183 <= io_pixelVal_in_0_3;
      end else if (8'hb7 == _T_22[7:0]) begin
        image_0_183 <= io_pixelVal_in_0_2;
      end else if (8'hb7 == _T_19[7:0]) begin
        image_0_183 <= io_pixelVal_in_0_1;
      end else if (8'hb7 == _T_15[7:0]) begin
        image_0_183 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_184 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb8 == _T_37[7:0]) begin
        image_0_184 <= io_pixelVal_in_0_7;
      end else if (8'hb8 == _T_34[7:0]) begin
        image_0_184 <= io_pixelVal_in_0_6;
      end else if (8'hb8 == _T_31[7:0]) begin
        image_0_184 <= io_pixelVal_in_0_5;
      end else if (8'hb8 == _T_28[7:0]) begin
        image_0_184 <= io_pixelVal_in_0_4;
      end else if (8'hb8 == _T_25[7:0]) begin
        image_0_184 <= io_pixelVal_in_0_3;
      end else if (8'hb8 == _T_22[7:0]) begin
        image_0_184 <= io_pixelVal_in_0_2;
      end else if (8'hb8 == _T_19[7:0]) begin
        image_0_184 <= io_pixelVal_in_0_1;
      end else if (8'hb8 == _T_15[7:0]) begin
        image_0_184 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_185 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb9 == _T_37[7:0]) begin
        image_0_185 <= io_pixelVal_in_0_7;
      end else if (8'hb9 == _T_34[7:0]) begin
        image_0_185 <= io_pixelVal_in_0_6;
      end else if (8'hb9 == _T_31[7:0]) begin
        image_0_185 <= io_pixelVal_in_0_5;
      end else if (8'hb9 == _T_28[7:0]) begin
        image_0_185 <= io_pixelVal_in_0_4;
      end else if (8'hb9 == _T_25[7:0]) begin
        image_0_185 <= io_pixelVal_in_0_3;
      end else if (8'hb9 == _T_22[7:0]) begin
        image_0_185 <= io_pixelVal_in_0_2;
      end else if (8'hb9 == _T_19[7:0]) begin
        image_0_185 <= io_pixelVal_in_0_1;
      end else if (8'hb9 == _T_15[7:0]) begin
        image_0_185 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_186 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hba == _T_37[7:0]) begin
        image_0_186 <= io_pixelVal_in_0_7;
      end else if (8'hba == _T_34[7:0]) begin
        image_0_186 <= io_pixelVal_in_0_6;
      end else if (8'hba == _T_31[7:0]) begin
        image_0_186 <= io_pixelVal_in_0_5;
      end else if (8'hba == _T_28[7:0]) begin
        image_0_186 <= io_pixelVal_in_0_4;
      end else if (8'hba == _T_25[7:0]) begin
        image_0_186 <= io_pixelVal_in_0_3;
      end else if (8'hba == _T_22[7:0]) begin
        image_0_186 <= io_pixelVal_in_0_2;
      end else if (8'hba == _T_19[7:0]) begin
        image_0_186 <= io_pixelVal_in_0_1;
      end else if (8'hba == _T_15[7:0]) begin
        image_0_186 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_187 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hbb == _T_37[7:0]) begin
        image_0_187 <= io_pixelVal_in_0_7;
      end else if (8'hbb == _T_34[7:0]) begin
        image_0_187 <= io_pixelVal_in_0_6;
      end else if (8'hbb == _T_31[7:0]) begin
        image_0_187 <= io_pixelVal_in_0_5;
      end else if (8'hbb == _T_28[7:0]) begin
        image_0_187 <= io_pixelVal_in_0_4;
      end else if (8'hbb == _T_25[7:0]) begin
        image_0_187 <= io_pixelVal_in_0_3;
      end else if (8'hbb == _T_22[7:0]) begin
        image_0_187 <= io_pixelVal_in_0_2;
      end else if (8'hbb == _T_19[7:0]) begin
        image_0_187 <= io_pixelVal_in_0_1;
      end else if (8'hbb == _T_15[7:0]) begin
        image_0_187 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_188 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hbc == _T_37[7:0]) begin
        image_0_188 <= io_pixelVal_in_0_7;
      end else if (8'hbc == _T_34[7:0]) begin
        image_0_188 <= io_pixelVal_in_0_6;
      end else if (8'hbc == _T_31[7:0]) begin
        image_0_188 <= io_pixelVal_in_0_5;
      end else if (8'hbc == _T_28[7:0]) begin
        image_0_188 <= io_pixelVal_in_0_4;
      end else if (8'hbc == _T_25[7:0]) begin
        image_0_188 <= io_pixelVal_in_0_3;
      end else if (8'hbc == _T_22[7:0]) begin
        image_0_188 <= io_pixelVal_in_0_2;
      end else if (8'hbc == _T_19[7:0]) begin
        image_0_188 <= io_pixelVal_in_0_1;
      end else if (8'hbc == _T_15[7:0]) begin
        image_0_188 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_189 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hbd == _T_37[7:0]) begin
        image_0_189 <= io_pixelVal_in_0_7;
      end else if (8'hbd == _T_34[7:0]) begin
        image_0_189 <= io_pixelVal_in_0_6;
      end else if (8'hbd == _T_31[7:0]) begin
        image_0_189 <= io_pixelVal_in_0_5;
      end else if (8'hbd == _T_28[7:0]) begin
        image_0_189 <= io_pixelVal_in_0_4;
      end else if (8'hbd == _T_25[7:0]) begin
        image_0_189 <= io_pixelVal_in_0_3;
      end else if (8'hbd == _T_22[7:0]) begin
        image_0_189 <= io_pixelVal_in_0_2;
      end else if (8'hbd == _T_19[7:0]) begin
        image_0_189 <= io_pixelVal_in_0_1;
      end else if (8'hbd == _T_15[7:0]) begin
        image_0_189 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_190 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hbe == _T_37[7:0]) begin
        image_0_190 <= io_pixelVal_in_0_7;
      end else if (8'hbe == _T_34[7:0]) begin
        image_0_190 <= io_pixelVal_in_0_6;
      end else if (8'hbe == _T_31[7:0]) begin
        image_0_190 <= io_pixelVal_in_0_5;
      end else if (8'hbe == _T_28[7:0]) begin
        image_0_190 <= io_pixelVal_in_0_4;
      end else if (8'hbe == _T_25[7:0]) begin
        image_0_190 <= io_pixelVal_in_0_3;
      end else if (8'hbe == _T_22[7:0]) begin
        image_0_190 <= io_pixelVal_in_0_2;
      end else if (8'hbe == _T_19[7:0]) begin
        image_0_190 <= io_pixelVal_in_0_1;
      end else if (8'hbe == _T_15[7:0]) begin
        image_0_190 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_191 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hbf == _T_37[7:0]) begin
        image_0_191 <= io_pixelVal_in_0_7;
      end else if (8'hbf == _T_34[7:0]) begin
        image_0_191 <= io_pixelVal_in_0_6;
      end else if (8'hbf == _T_31[7:0]) begin
        image_0_191 <= io_pixelVal_in_0_5;
      end else if (8'hbf == _T_28[7:0]) begin
        image_0_191 <= io_pixelVal_in_0_4;
      end else if (8'hbf == _T_25[7:0]) begin
        image_0_191 <= io_pixelVal_in_0_3;
      end else if (8'hbf == _T_22[7:0]) begin
        image_0_191 <= io_pixelVal_in_0_2;
      end else if (8'hbf == _T_19[7:0]) begin
        image_0_191 <= io_pixelVal_in_0_1;
      end else if (8'hbf == _T_15[7:0]) begin
        image_0_191 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_1_0 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h0 == _T_37[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_7;
      end else if (8'h0 == _T_34[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_6;
      end else if (8'h0 == _T_31[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_5;
      end else if (8'h0 == _T_28[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_4;
      end else if (8'h0 == _T_25[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_3;
      end else if (8'h0 == _T_22[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_2;
      end else if (8'h0 == _T_19[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_1;
      end else if (8'h0 == _T_15[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_1 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1 == _T_37[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_7;
      end else if (8'h1 == _T_34[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_6;
      end else if (8'h1 == _T_31[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_5;
      end else if (8'h1 == _T_28[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_4;
      end else if (8'h1 == _T_25[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_3;
      end else if (8'h1 == _T_22[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_2;
      end else if (8'h1 == _T_19[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_1;
      end else if (8'h1 == _T_15[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_2 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2 == _T_37[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_7;
      end else if (8'h2 == _T_34[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_6;
      end else if (8'h2 == _T_31[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_5;
      end else if (8'h2 == _T_28[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_4;
      end else if (8'h2 == _T_25[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_3;
      end else if (8'h2 == _T_22[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_2;
      end else if (8'h2 == _T_19[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_1;
      end else if (8'h2 == _T_15[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_3 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3 == _T_37[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_7;
      end else if (8'h3 == _T_34[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_6;
      end else if (8'h3 == _T_31[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_5;
      end else if (8'h3 == _T_28[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_4;
      end else if (8'h3 == _T_25[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_3;
      end else if (8'h3 == _T_22[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_2;
      end else if (8'h3 == _T_19[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_1;
      end else if (8'h3 == _T_15[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_4 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4 == _T_37[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_7;
      end else if (8'h4 == _T_34[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_6;
      end else if (8'h4 == _T_31[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_5;
      end else if (8'h4 == _T_28[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_4;
      end else if (8'h4 == _T_25[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_3;
      end else if (8'h4 == _T_22[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_2;
      end else if (8'h4 == _T_19[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_1;
      end else if (8'h4 == _T_15[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_5 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5 == _T_37[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_7;
      end else if (8'h5 == _T_34[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_6;
      end else if (8'h5 == _T_31[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_5;
      end else if (8'h5 == _T_28[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_4;
      end else if (8'h5 == _T_25[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_3;
      end else if (8'h5 == _T_22[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_2;
      end else if (8'h5 == _T_19[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_1;
      end else if (8'h5 == _T_15[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_6 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6 == _T_37[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_7;
      end else if (8'h6 == _T_34[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_6;
      end else if (8'h6 == _T_31[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_5;
      end else if (8'h6 == _T_28[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_4;
      end else if (8'h6 == _T_25[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_3;
      end else if (8'h6 == _T_22[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_2;
      end else if (8'h6 == _T_19[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_1;
      end else if (8'h6 == _T_15[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_7 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7 == _T_37[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_7;
      end else if (8'h7 == _T_34[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_6;
      end else if (8'h7 == _T_31[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_5;
      end else if (8'h7 == _T_28[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_4;
      end else if (8'h7 == _T_25[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_3;
      end else if (8'h7 == _T_22[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_2;
      end else if (8'h7 == _T_19[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_1;
      end else if (8'h7 == _T_15[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_8 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8 == _T_37[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_7;
      end else if (8'h8 == _T_34[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_6;
      end else if (8'h8 == _T_31[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_5;
      end else if (8'h8 == _T_28[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_4;
      end else if (8'h8 == _T_25[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_3;
      end else if (8'h8 == _T_22[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_2;
      end else if (8'h8 == _T_19[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_1;
      end else if (8'h8 == _T_15[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_9 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9 == _T_37[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_7;
      end else if (8'h9 == _T_34[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_6;
      end else if (8'h9 == _T_31[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_5;
      end else if (8'h9 == _T_28[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_4;
      end else if (8'h9 == _T_25[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_3;
      end else if (8'h9 == _T_22[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_2;
      end else if (8'h9 == _T_19[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_1;
      end else if (8'h9 == _T_15[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_10 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha == _T_37[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_7;
      end else if (8'ha == _T_34[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_6;
      end else if (8'ha == _T_31[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_5;
      end else if (8'ha == _T_28[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_4;
      end else if (8'ha == _T_25[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_3;
      end else if (8'ha == _T_22[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_2;
      end else if (8'ha == _T_19[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_1;
      end else if (8'ha == _T_15[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_11 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb == _T_37[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_7;
      end else if (8'hb == _T_34[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_6;
      end else if (8'hb == _T_31[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_5;
      end else if (8'hb == _T_28[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_4;
      end else if (8'hb == _T_25[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_3;
      end else if (8'hb == _T_22[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_2;
      end else if (8'hb == _T_19[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_1;
      end else if (8'hb == _T_15[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_12 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc == _T_37[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_7;
      end else if (8'hc == _T_34[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_6;
      end else if (8'hc == _T_31[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_5;
      end else if (8'hc == _T_28[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_4;
      end else if (8'hc == _T_25[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_3;
      end else if (8'hc == _T_22[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_2;
      end else if (8'hc == _T_19[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_1;
      end else if (8'hc == _T_15[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_13 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd == _T_37[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_7;
      end else if (8'hd == _T_34[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_6;
      end else if (8'hd == _T_31[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_5;
      end else if (8'hd == _T_28[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_4;
      end else if (8'hd == _T_25[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_3;
      end else if (8'hd == _T_22[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_2;
      end else if (8'hd == _T_19[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_1;
      end else if (8'hd == _T_15[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_14 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he == _T_37[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_7;
      end else if (8'he == _T_34[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_6;
      end else if (8'he == _T_31[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_5;
      end else if (8'he == _T_28[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_4;
      end else if (8'he == _T_25[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_3;
      end else if (8'he == _T_22[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_2;
      end else if (8'he == _T_19[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_1;
      end else if (8'he == _T_15[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_15 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf == _T_37[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_7;
      end else if (8'hf == _T_34[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_6;
      end else if (8'hf == _T_31[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_5;
      end else if (8'hf == _T_28[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_4;
      end else if (8'hf == _T_25[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_3;
      end else if (8'hf == _T_22[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_2;
      end else if (8'hf == _T_19[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_1;
      end else if (8'hf == _T_15[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_16 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h10 == _T_37[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_7;
      end else if (8'h10 == _T_34[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_6;
      end else if (8'h10 == _T_31[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_5;
      end else if (8'h10 == _T_28[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_4;
      end else if (8'h10 == _T_25[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_3;
      end else if (8'h10 == _T_22[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_2;
      end else if (8'h10 == _T_19[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_1;
      end else if (8'h10 == _T_15[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_17 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h11 == _T_37[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_7;
      end else if (8'h11 == _T_34[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_6;
      end else if (8'h11 == _T_31[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_5;
      end else if (8'h11 == _T_28[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_4;
      end else if (8'h11 == _T_25[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_3;
      end else if (8'h11 == _T_22[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_2;
      end else if (8'h11 == _T_19[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_1;
      end else if (8'h11 == _T_15[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_18 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h12 == _T_37[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_7;
      end else if (8'h12 == _T_34[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_6;
      end else if (8'h12 == _T_31[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_5;
      end else if (8'h12 == _T_28[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_4;
      end else if (8'h12 == _T_25[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_3;
      end else if (8'h12 == _T_22[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_2;
      end else if (8'h12 == _T_19[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_1;
      end else if (8'h12 == _T_15[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_19 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h13 == _T_37[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_7;
      end else if (8'h13 == _T_34[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_6;
      end else if (8'h13 == _T_31[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_5;
      end else if (8'h13 == _T_28[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_4;
      end else if (8'h13 == _T_25[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_3;
      end else if (8'h13 == _T_22[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_2;
      end else if (8'h13 == _T_19[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_1;
      end else if (8'h13 == _T_15[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_20 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h14 == _T_37[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_7;
      end else if (8'h14 == _T_34[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_6;
      end else if (8'h14 == _T_31[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_5;
      end else if (8'h14 == _T_28[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_4;
      end else if (8'h14 == _T_25[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_3;
      end else if (8'h14 == _T_22[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_2;
      end else if (8'h14 == _T_19[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_1;
      end else if (8'h14 == _T_15[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_21 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h15 == _T_37[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_7;
      end else if (8'h15 == _T_34[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_6;
      end else if (8'h15 == _T_31[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_5;
      end else if (8'h15 == _T_28[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_4;
      end else if (8'h15 == _T_25[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_3;
      end else if (8'h15 == _T_22[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_2;
      end else if (8'h15 == _T_19[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_1;
      end else if (8'h15 == _T_15[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_22 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h16 == _T_37[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_7;
      end else if (8'h16 == _T_34[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_6;
      end else if (8'h16 == _T_31[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_5;
      end else if (8'h16 == _T_28[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_4;
      end else if (8'h16 == _T_25[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_3;
      end else if (8'h16 == _T_22[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_2;
      end else if (8'h16 == _T_19[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_1;
      end else if (8'h16 == _T_15[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_23 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h17 == _T_37[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_7;
      end else if (8'h17 == _T_34[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_6;
      end else if (8'h17 == _T_31[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_5;
      end else if (8'h17 == _T_28[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_4;
      end else if (8'h17 == _T_25[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_3;
      end else if (8'h17 == _T_22[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_2;
      end else if (8'h17 == _T_19[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_1;
      end else if (8'h17 == _T_15[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_24 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h18 == _T_37[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_7;
      end else if (8'h18 == _T_34[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_6;
      end else if (8'h18 == _T_31[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_5;
      end else if (8'h18 == _T_28[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_4;
      end else if (8'h18 == _T_25[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_3;
      end else if (8'h18 == _T_22[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_2;
      end else if (8'h18 == _T_19[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_1;
      end else if (8'h18 == _T_15[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_25 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h19 == _T_37[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_7;
      end else if (8'h19 == _T_34[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_6;
      end else if (8'h19 == _T_31[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_5;
      end else if (8'h19 == _T_28[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_4;
      end else if (8'h19 == _T_25[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_3;
      end else if (8'h19 == _T_22[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_2;
      end else if (8'h19 == _T_19[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_1;
      end else if (8'h19 == _T_15[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_26 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1a == _T_37[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_7;
      end else if (8'h1a == _T_34[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_6;
      end else if (8'h1a == _T_31[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_5;
      end else if (8'h1a == _T_28[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_4;
      end else if (8'h1a == _T_25[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_3;
      end else if (8'h1a == _T_22[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_2;
      end else if (8'h1a == _T_19[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_1;
      end else if (8'h1a == _T_15[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_27 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1b == _T_37[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_7;
      end else if (8'h1b == _T_34[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_6;
      end else if (8'h1b == _T_31[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_5;
      end else if (8'h1b == _T_28[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_4;
      end else if (8'h1b == _T_25[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_3;
      end else if (8'h1b == _T_22[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_2;
      end else if (8'h1b == _T_19[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_1;
      end else if (8'h1b == _T_15[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_28 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1c == _T_37[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_7;
      end else if (8'h1c == _T_34[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_6;
      end else if (8'h1c == _T_31[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_5;
      end else if (8'h1c == _T_28[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_4;
      end else if (8'h1c == _T_25[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_3;
      end else if (8'h1c == _T_22[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_2;
      end else if (8'h1c == _T_19[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_1;
      end else if (8'h1c == _T_15[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_29 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1d == _T_37[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_7;
      end else if (8'h1d == _T_34[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_6;
      end else if (8'h1d == _T_31[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_5;
      end else if (8'h1d == _T_28[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_4;
      end else if (8'h1d == _T_25[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_3;
      end else if (8'h1d == _T_22[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_2;
      end else if (8'h1d == _T_19[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_1;
      end else if (8'h1d == _T_15[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_30 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1e == _T_37[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_7;
      end else if (8'h1e == _T_34[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_6;
      end else if (8'h1e == _T_31[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_5;
      end else if (8'h1e == _T_28[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_4;
      end else if (8'h1e == _T_25[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_3;
      end else if (8'h1e == _T_22[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_2;
      end else if (8'h1e == _T_19[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_1;
      end else if (8'h1e == _T_15[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_31 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1f == _T_37[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_7;
      end else if (8'h1f == _T_34[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_6;
      end else if (8'h1f == _T_31[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_5;
      end else if (8'h1f == _T_28[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_4;
      end else if (8'h1f == _T_25[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_3;
      end else if (8'h1f == _T_22[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_2;
      end else if (8'h1f == _T_19[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_1;
      end else if (8'h1f == _T_15[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_32 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h20 == _T_37[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_7;
      end else if (8'h20 == _T_34[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_6;
      end else if (8'h20 == _T_31[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_5;
      end else if (8'h20 == _T_28[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_4;
      end else if (8'h20 == _T_25[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_3;
      end else if (8'h20 == _T_22[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_2;
      end else if (8'h20 == _T_19[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_1;
      end else if (8'h20 == _T_15[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_33 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h21 == _T_37[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_7;
      end else if (8'h21 == _T_34[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_6;
      end else if (8'h21 == _T_31[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_5;
      end else if (8'h21 == _T_28[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_4;
      end else if (8'h21 == _T_25[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_3;
      end else if (8'h21 == _T_22[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_2;
      end else if (8'h21 == _T_19[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_1;
      end else if (8'h21 == _T_15[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_34 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h22 == _T_37[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_7;
      end else if (8'h22 == _T_34[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_6;
      end else if (8'h22 == _T_31[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_5;
      end else if (8'h22 == _T_28[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_4;
      end else if (8'h22 == _T_25[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_3;
      end else if (8'h22 == _T_22[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_2;
      end else if (8'h22 == _T_19[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_1;
      end else if (8'h22 == _T_15[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_35 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h23 == _T_37[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_7;
      end else if (8'h23 == _T_34[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_6;
      end else if (8'h23 == _T_31[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_5;
      end else if (8'h23 == _T_28[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_4;
      end else if (8'h23 == _T_25[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_3;
      end else if (8'h23 == _T_22[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_2;
      end else if (8'h23 == _T_19[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_1;
      end else if (8'h23 == _T_15[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_36 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h24 == _T_37[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_7;
      end else if (8'h24 == _T_34[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_6;
      end else if (8'h24 == _T_31[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_5;
      end else if (8'h24 == _T_28[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_4;
      end else if (8'h24 == _T_25[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_3;
      end else if (8'h24 == _T_22[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_2;
      end else if (8'h24 == _T_19[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_1;
      end else if (8'h24 == _T_15[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_37 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h25 == _T_37[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_7;
      end else if (8'h25 == _T_34[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_6;
      end else if (8'h25 == _T_31[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_5;
      end else if (8'h25 == _T_28[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_4;
      end else if (8'h25 == _T_25[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_3;
      end else if (8'h25 == _T_22[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_2;
      end else if (8'h25 == _T_19[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_1;
      end else if (8'h25 == _T_15[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_38 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h26 == _T_37[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_7;
      end else if (8'h26 == _T_34[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_6;
      end else if (8'h26 == _T_31[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_5;
      end else if (8'h26 == _T_28[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_4;
      end else if (8'h26 == _T_25[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_3;
      end else if (8'h26 == _T_22[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_2;
      end else if (8'h26 == _T_19[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_1;
      end else if (8'h26 == _T_15[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_39 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h27 == _T_37[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_7;
      end else if (8'h27 == _T_34[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_6;
      end else if (8'h27 == _T_31[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_5;
      end else if (8'h27 == _T_28[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_4;
      end else if (8'h27 == _T_25[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_3;
      end else if (8'h27 == _T_22[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_2;
      end else if (8'h27 == _T_19[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_1;
      end else if (8'h27 == _T_15[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_40 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h28 == _T_37[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_7;
      end else if (8'h28 == _T_34[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_6;
      end else if (8'h28 == _T_31[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_5;
      end else if (8'h28 == _T_28[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_4;
      end else if (8'h28 == _T_25[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_3;
      end else if (8'h28 == _T_22[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_2;
      end else if (8'h28 == _T_19[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_1;
      end else if (8'h28 == _T_15[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_41 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h29 == _T_37[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_7;
      end else if (8'h29 == _T_34[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_6;
      end else if (8'h29 == _T_31[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_5;
      end else if (8'h29 == _T_28[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_4;
      end else if (8'h29 == _T_25[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_3;
      end else if (8'h29 == _T_22[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_2;
      end else if (8'h29 == _T_19[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_1;
      end else if (8'h29 == _T_15[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_42 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2a == _T_37[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_7;
      end else if (8'h2a == _T_34[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_6;
      end else if (8'h2a == _T_31[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_5;
      end else if (8'h2a == _T_28[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_4;
      end else if (8'h2a == _T_25[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_3;
      end else if (8'h2a == _T_22[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_2;
      end else if (8'h2a == _T_19[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_1;
      end else if (8'h2a == _T_15[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_43 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2b == _T_37[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_7;
      end else if (8'h2b == _T_34[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_6;
      end else if (8'h2b == _T_31[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_5;
      end else if (8'h2b == _T_28[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_4;
      end else if (8'h2b == _T_25[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_3;
      end else if (8'h2b == _T_22[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_2;
      end else if (8'h2b == _T_19[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_1;
      end else if (8'h2b == _T_15[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_44 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2c == _T_37[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_7;
      end else if (8'h2c == _T_34[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_6;
      end else if (8'h2c == _T_31[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_5;
      end else if (8'h2c == _T_28[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_4;
      end else if (8'h2c == _T_25[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_3;
      end else if (8'h2c == _T_22[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_2;
      end else if (8'h2c == _T_19[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_1;
      end else if (8'h2c == _T_15[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_45 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2d == _T_37[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_7;
      end else if (8'h2d == _T_34[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_6;
      end else if (8'h2d == _T_31[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_5;
      end else if (8'h2d == _T_28[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_4;
      end else if (8'h2d == _T_25[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_3;
      end else if (8'h2d == _T_22[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_2;
      end else if (8'h2d == _T_19[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_1;
      end else if (8'h2d == _T_15[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_46 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2e == _T_37[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_7;
      end else if (8'h2e == _T_34[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_6;
      end else if (8'h2e == _T_31[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_5;
      end else if (8'h2e == _T_28[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_4;
      end else if (8'h2e == _T_25[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_3;
      end else if (8'h2e == _T_22[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_2;
      end else if (8'h2e == _T_19[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_1;
      end else if (8'h2e == _T_15[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_47 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2f == _T_37[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_7;
      end else if (8'h2f == _T_34[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_6;
      end else if (8'h2f == _T_31[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_5;
      end else if (8'h2f == _T_28[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_4;
      end else if (8'h2f == _T_25[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_3;
      end else if (8'h2f == _T_22[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_2;
      end else if (8'h2f == _T_19[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_1;
      end else if (8'h2f == _T_15[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_48 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h30 == _T_37[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_7;
      end else if (8'h30 == _T_34[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_6;
      end else if (8'h30 == _T_31[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_5;
      end else if (8'h30 == _T_28[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_4;
      end else if (8'h30 == _T_25[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_3;
      end else if (8'h30 == _T_22[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_2;
      end else if (8'h30 == _T_19[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_1;
      end else if (8'h30 == _T_15[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_49 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h31 == _T_37[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_7;
      end else if (8'h31 == _T_34[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_6;
      end else if (8'h31 == _T_31[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_5;
      end else if (8'h31 == _T_28[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_4;
      end else if (8'h31 == _T_25[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_3;
      end else if (8'h31 == _T_22[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_2;
      end else if (8'h31 == _T_19[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_1;
      end else if (8'h31 == _T_15[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_50 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h32 == _T_37[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_7;
      end else if (8'h32 == _T_34[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_6;
      end else if (8'h32 == _T_31[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_5;
      end else if (8'h32 == _T_28[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_4;
      end else if (8'h32 == _T_25[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_3;
      end else if (8'h32 == _T_22[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_2;
      end else if (8'h32 == _T_19[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_1;
      end else if (8'h32 == _T_15[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_51 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h33 == _T_37[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_7;
      end else if (8'h33 == _T_34[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_6;
      end else if (8'h33 == _T_31[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_5;
      end else if (8'h33 == _T_28[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_4;
      end else if (8'h33 == _T_25[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_3;
      end else if (8'h33 == _T_22[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_2;
      end else if (8'h33 == _T_19[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_1;
      end else if (8'h33 == _T_15[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_52 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h34 == _T_37[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_7;
      end else if (8'h34 == _T_34[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_6;
      end else if (8'h34 == _T_31[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_5;
      end else if (8'h34 == _T_28[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_4;
      end else if (8'h34 == _T_25[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_3;
      end else if (8'h34 == _T_22[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_2;
      end else if (8'h34 == _T_19[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_1;
      end else if (8'h34 == _T_15[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_53 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h35 == _T_37[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_7;
      end else if (8'h35 == _T_34[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_6;
      end else if (8'h35 == _T_31[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_5;
      end else if (8'h35 == _T_28[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_4;
      end else if (8'h35 == _T_25[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_3;
      end else if (8'h35 == _T_22[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_2;
      end else if (8'h35 == _T_19[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_1;
      end else if (8'h35 == _T_15[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_54 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h36 == _T_37[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_7;
      end else if (8'h36 == _T_34[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_6;
      end else if (8'h36 == _T_31[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_5;
      end else if (8'h36 == _T_28[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_4;
      end else if (8'h36 == _T_25[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_3;
      end else if (8'h36 == _T_22[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_2;
      end else if (8'h36 == _T_19[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_1;
      end else if (8'h36 == _T_15[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_55 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h37 == _T_37[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_7;
      end else if (8'h37 == _T_34[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_6;
      end else if (8'h37 == _T_31[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_5;
      end else if (8'h37 == _T_28[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_4;
      end else if (8'h37 == _T_25[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_3;
      end else if (8'h37 == _T_22[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_2;
      end else if (8'h37 == _T_19[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_1;
      end else if (8'h37 == _T_15[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_56 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h38 == _T_37[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_7;
      end else if (8'h38 == _T_34[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_6;
      end else if (8'h38 == _T_31[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_5;
      end else if (8'h38 == _T_28[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_4;
      end else if (8'h38 == _T_25[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_3;
      end else if (8'h38 == _T_22[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_2;
      end else if (8'h38 == _T_19[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_1;
      end else if (8'h38 == _T_15[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_57 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h39 == _T_37[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_7;
      end else if (8'h39 == _T_34[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_6;
      end else if (8'h39 == _T_31[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_5;
      end else if (8'h39 == _T_28[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_4;
      end else if (8'h39 == _T_25[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_3;
      end else if (8'h39 == _T_22[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_2;
      end else if (8'h39 == _T_19[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_1;
      end else if (8'h39 == _T_15[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_58 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3a == _T_37[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_7;
      end else if (8'h3a == _T_34[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_6;
      end else if (8'h3a == _T_31[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_5;
      end else if (8'h3a == _T_28[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_4;
      end else if (8'h3a == _T_25[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_3;
      end else if (8'h3a == _T_22[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_2;
      end else if (8'h3a == _T_19[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_1;
      end else if (8'h3a == _T_15[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_59 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3b == _T_37[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_7;
      end else if (8'h3b == _T_34[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_6;
      end else if (8'h3b == _T_31[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_5;
      end else if (8'h3b == _T_28[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_4;
      end else if (8'h3b == _T_25[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_3;
      end else if (8'h3b == _T_22[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_2;
      end else if (8'h3b == _T_19[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_1;
      end else if (8'h3b == _T_15[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_60 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3c == _T_37[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_7;
      end else if (8'h3c == _T_34[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_6;
      end else if (8'h3c == _T_31[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_5;
      end else if (8'h3c == _T_28[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_4;
      end else if (8'h3c == _T_25[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_3;
      end else if (8'h3c == _T_22[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_2;
      end else if (8'h3c == _T_19[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_1;
      end else if (8'h3c == _T_15[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_61 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3d == _T_37[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_7;
      end else if (8'h3d == _T_34[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_6;
      end else if (8'h3d == _T_31[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_5;
      end else if (8'h3d == _T_28[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_4;
      end else if (8'h3d == _T_25[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_3;
      end else if (8'h3d == _T_22[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_2;
      end else if (8'h3d == _T_19[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_1;
      end else if (8'h3d == _T_15[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_62 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3e == _T_37[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_7;
      end else if (8'h3e == _T_34[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_6;
      end else if (8'h3e == _T_31[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_5;
      end else if (8'h3e == _T_28[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_4;
      end else if (8'h3e == _T_25[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_3;
      end else if (8'h3e == _T_22[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_2;
      end else if (8'h3e == _T_19[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_1;
      end else if (8'h3e == _T_15[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_63 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3f == _T_37[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_7;
      end else if (8'h3f == _T_34[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_6;
      end else if (8'h3f == _T_31[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_5;
      end else if (8'h3f == _T_28[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_4;
      end else if (8'h3f == _T_25[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_3;
      end else if (8'h3f == _T_22[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_2;
      end else if (8'h3f == _T_19[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_1;
      end else if (8'h3f == _T_15[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_64 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h40 == _T_37[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_7;
      end else if (8'h40 == _T_34[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_6;
      end else if (8'h40 == _T_31[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_5;
      end else if (8'h40 == _T_28[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_4;
      end else if (8'h40 == _T_25[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_3;
      end else if (8'h40 == _T_22[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_2;
      end else if (8'h40 == _T_19[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_1;
      end else if (8'h40 == _T_15[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_65 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h41 == _T_37[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_7;
      end else if (8'h41 == _T_34[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_6;
      end else if (8'h41 == _T_31[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_5;
      end else if (8'h41 == _T_28[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_4;
      end else if (8'h41 == _T_25[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_3;
      end else if (8'h41 == _T_22[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_2;
      end else if (8'h41 == _T_19[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_1;
      end else if (8'h41 == _T_15[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_66 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h42 == _T_37[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_7;
      end else if (8'h42 == _T_34[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_6;
      end else if (8'h42 == _T_31[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_5;
      end else if (8'h42 == _T_28[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_4;
      end else if (8'h42 == _T_25[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_3;
      end else if (8'h42 == _T_22[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_2;
      end else if (8'h42 == _T_19[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_1;
      end else if (8'h42 == _T_15[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_67 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h43 == _T_37[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_7;
      end else if (8'h43 == _T_34[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_6;
      end else if (8'h43 == _T_31[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_5;
      end else if (8'h43 == _T_28[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_4;
      end else if (8'h43 == _T_25[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_3;
      end else if (8'h43 == _T_22[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_2;
      end else if (8'h43 == _T_19[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_1;
      end else if (8'h43 == _T_15[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_68 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h44 == _T_37[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_7;
      end else if (8'h44 == _T_34[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_6;
      end else if (8'h44 == _T_31[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_5;
      end else if (8'h44 == _T_28[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_4;
      end else if (8'h44 == _T_25[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_3;
      end else if (8'h44 == _T_22[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_2;
      end else if (8'h44 == _T_19[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_1;
      end else if (8'h44 == _T_15[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_69 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h45 == _T_37[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_7;
      end else if (8'h45 == _T_34[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_6;
      end else if (8'h45 == _T_31[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_5;
      end else if (8'h45 == _T_28[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_4;
      end else if (8'h45 == _T_25[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_3;
      end else if (8'h45 == _T_22[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_2;
      end else if (8'h45 == _T_19[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_1;
      end else if (8'h45 == _T_15[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_70 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h46 == _T_37[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_7;
      end else if (8'h46 == _T_34[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_6;
      end else if (8'h46 == _T_31[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_5;
      end else if (8'h46 == _T_28[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_4;
      end else if (8'h46 == _T_25[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_3;
      end else if (8'h46 == _T_22[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_2;
      end else if (8'h46 == _T_19[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_1;
      end else if (8'h46 == _T_15[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_71 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h47 == _T_37[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_7;
      end else if (8'h47 == _T_34[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_6;
      end else if (8'h47 == _T_31[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_5;
      end else if (8'h47 == _T_28[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_4;
      end else if (8'h47 == _T_25[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_3;
      end else if (8'h47 == _T_22[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_2;
      end else if (8'h47 == _T_19[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_1;
      end else if (8'h47 == _T_15[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_72 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h48 == _T_37[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_7;
      end else if (8'h48 == _T_34[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_6;
      end else if (8'h48 == _T_31[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_5;
      end else if (8'h48 == _T_28[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_4;
      end else if (8'h48 == _T_25[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_3;
      end else if (8'h48 == _T_22[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_2;
      end else if (8'h48 == _T_19[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_1;
      end else if (8'h48 == _T_15[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_73 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h49 == _T_37[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_7;
      end else if (8'h49 == _T_34[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_6;
      end else if (8'h49 == _T_31[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_5;
      end else if (8'h49 == _T_28[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_4;
      end else if (8'h49 == _T_25[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_3;
      end else if (8'h49 == _T_22[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_2;
      end else if (8'h49 == _T_19[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_1;
      end else if (8'h49 == _T_15[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_74 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4a == _T_37[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_7;
      end else if (8'h4a == _T_34[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_6;
      end else if (8'h4a == _T_31[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_5;
      end else if (8'h4a == _T_28[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_4;
      end else if (8'h4a == _T_25[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_3;
      end else if (8'h4a == _T_22[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_2;
      end else if (8'h4a == _T_19[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_1;
      end else if (8'h4a == _T_15[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_75 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4b == _T_37[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_7;
      end else if (8'h4b == _T_34[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_6;
      end else if (8'h4b == _T_31[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_5;
      end else if (8'h4b == _T_28[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_4;
      end else if (8'h4b == _T_25[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_3;
      end else if (8'h4b == _T_22[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_2;
      end else if (8'h4b == _T_19[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_1;
      end else if (8'h4b == _T_15[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_76 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4c == _T_37[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_7;
      end else if (8'h4c == _T_34[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_6;
      end else if (8'h4c == _T_31[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_5;
      end else if (8'h4c == _T_28[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_4;
      end else if (8'h4c == _T_25[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_3;
      end else if (8'h4c == _T_22[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_2;
      end else if (8'h4c == _T_19[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_1;
      end else if (8'h4c == _T_15[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_77 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4d == _T_37[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_7;
      end else if (8'h4d == _T_34[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_6;
      end else if (8'h4d == _T_31[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_5;
      end else if (8'h4d == _T_28[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_4;
      end else if (8'h4d == _T_25[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_3;
      end else if (8'h4d == _T_22[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_2;
      end else if (8'h4d == _T_19[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_1;
      end else if (8'h4d == _T_15[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_78 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4e == _T_37[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_7;
      end else if (8'h4e == _T_34[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_6;
      end else if (8'h4e == _T_31[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_5;
      end else if (8'h4e == _T_28[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_4;
      end else if (8'h4e == _T_25[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_3;
      end else if (8'h4e == _T_22[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_2;
      end else if (8'h4e == _T_19[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_1;
      end else if (8'h4e == _T_15[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_79 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4f == _T_37[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_7;
      end else if (8'h4f == _T_34[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_6;
      end else if (8'h4f == _T_31[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_5;
      end else if (8'h4f == _T_28[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_4;
      end else if (8'h4f == _T_25[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_3;
      end else if (8'h4f == _T_22[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_2;
      end else if (8'h4f == _T_19[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_1;
      end else if (8'h4f == _T_15[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_80 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h50 == _T_37[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_7;
      end else if (8'h50 == _T_34[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_6;
      end else if (8'h50 == _T_31[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_5;
      end else if (8'h50 == _T_28[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_4;
      end else if (8'h50 == _T_25[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_3;
      end else if (8'h50 == _T_22[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_2;
      end else if (8'h50 == _T_19[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_1;
      end else if (8'h50 == _T_15[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_81 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h51 == _T_37[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_7;
      end else if (8'h51 == _T_34[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_6;
      end else if (8'h51 == _T_31[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_5;
      end else if (8'h51 == _T_28[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_4;
      end else if (8'h51 == _T_25[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_3;
      end else if (8'h51 == _T_22[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_2;
      end else if (8'h51 == _T_19[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_1;
      end else if (8'h51 == _T_15[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_82 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h52 == _T_37[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_7;
      end else if (8'h52 == _T_34[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_6;
      end else if (8'h52 == _T_31[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_5;
      end else if (8'h52 == _T_28[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_4;
      end else if (8'h52 == _T_25[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_3;
      end else if (8'h52 == _T_22[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_2;
      end else if (8'h52 == _T_19[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_1;
      end else if (8'h52 == _T_15[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_83 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h53 == _T_37[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_7;
      end else if (8'h53 == _T_34[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_6;
      end else if (8'h53 == _T_31[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_5;
      end else if (8'h53 == _T_28[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_4;
      end else if (8'h53 == _T_25[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_3;
      end else if (8'h53 == _T_22[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_2;
      end else if (8'h53 == _T_19[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_1;
      end else if (8'h53 == _T_15[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_84 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h54 == _T_37[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_7;
      end else if (8'h54 == _T_34[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_6;
      end else if (8'h54 == _T_31[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_5;
      end else if (8'h54 == _T_28[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_4;
      end else if (8'h54 == _T_25[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_3;
      end else if (8'h54 == _T_22[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_2;
      end else if (8'h54 == _T_19[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_1;
      end else if (8'h54 == _T_15[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_85 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h55 == _T_37[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_7;
      end else if (8'h55 == _T_34[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_6;
      end else if (8'h55 == _T_31[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_5;
      end else if (8'h55 == _T_28[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_4;
      end else if (8'h55 == _T_25[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_3;
      end else if (8'h55 == _T_22[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_2;
      end else if (8'h55 == _T_19[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_1;
      end else if (8'h55 == _T_15[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_86 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h56 == _T_37[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_7;
      end else if (8'h56 == _T_34[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_6;
      end else if (8'h56 == _T_31[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_5;
      end else if (8'h56 == _T_28[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_4;
      end else if (8'h56 == _T_25[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_3;
      end else if (8'h56 == _T_22[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_2;
      end else if (8'h56 == _T_19[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_1;
      end else if (8'h56 == _T_15[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_87 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h57 == _T_37[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_7;
      end else if (8'h57 == _T_34[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_6;
      end else if (8'h57 == _T_31[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_5;
      end else if (8'h57 == _T_28[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_4;
      end else if (8'h57 == _T_25[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_3;
      end else if (8'h57 == _T_22[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_2;
      end else if (8'h57 == _T_19[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_1;
      end else if (8'h57 == _T_15[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_88 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h58 == _T_37[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_7;
      end else if (8'h58 == _T_34[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_6;
      end else if (8'h58 == _T_31[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_5;
      end else if (8'h58 == _T_28[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_4;
      end else if (8'h58 == _T_25[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_3;
      end else if (8'h58 == _T_22[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_2;
      end else if (8'h58 == _T_19[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_1;
      end else if (8'h58 == _T_15[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_89 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h59 == _T_37[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_7;
      end else if (8'h59 == _T_34[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_6;
      end else if (8'h59 == _T_31[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_5;
      end else if (8'h59 == _T_28[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_4;
      end else if (8'h59 == _T_25[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_3;
      end else if (8'h59 == _T_22[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_2;
      end else if (8'h59 == _T_19[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_1;
      end else if (8'h59 == _T_15[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_90 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5a == _T_37[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_7;
      end else if (8'h5a == _T_34[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_6;
      end else if (8'h5a == _T_31[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_5;
      end else if (8'h5a == _T_28[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_4;
      end else if (8'h5a == _T_25[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_3;
      end else if (8'h5a == _T_22[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_2;
      end else if (8'h5a == _T_19[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_1;
      end else if (8'h5a == _T_15[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_91 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5b == _T_37[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_7;
      end else if (8'h5b == _T_34[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_6;
      end else if (8'h5b == _T_31[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_5;
      end else if (8'h5b == _T_28[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_4;
      end else if (8'h5b == _T_25[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_3;
      end else if (8'h5b == _T_22[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_2;
      end else if (8'h5b == _T_19[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_1;
      end else if (8'h5b == _T_15[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_92 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5c == _T_37[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_7;
      end else if (8'h5c == _T_34[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_6;
      end else if (8'h5c == _T_31[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_5;
      end else if (8'h5c == _T_28[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_4;
      end else if (8'h5c == _T_25[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_3;
      end else if (8'h5c == _T_22[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_2;
      end else if (8'h5c == _T_19[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_1;
      end else if (8'h5c == _T_15[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_93 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5d == _T_37[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_7;
      end else if (8'h5d == _T_34[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_6;
      end else if (8'h5d == _T_31[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_5;
      end else if (8'h5d == _T_28[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_4;
      end else if (8'h5d == _T_25[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_3;
      end else if (8'h5d == _T_22[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_2;
      end else if (8'h5d == _T_19[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_1;
      end else if (8'h5d == _T_15[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_94 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5e == _T_37[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_7;
      end else if (8'h5e == _T_34[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_6;
      end else if (8'h5e == _T_31[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_5;
      end else if (8'h5e == _T_28[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_4;
      end else if (8'h5e == _T_25[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_3;
      end else if (8'h5e == _T_22[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_2;
      end else if (8'h5e == _T_19[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_1;
      end else if (8'h5e == _T_15[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_95 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5f == _T_37[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_7;
      end else if (8'h5f == _T_34[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_6;
      end else if (8'h5f == _T_31[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_5;
      end else if (8'h5f == _T_28[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_4;
      end else if (8'h5f == _T_25[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_3;
      end else if (8'h5f == _T_22[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_2;
      end else if (8'h5f == _T_19[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_1;
      end else if (8'h5f == _T_15[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_96 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h60 == _T_37[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_7;
      end else if (8'h60 == _T_34[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_6;
      end else if (8'h60 == _T_31[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_5;
      end else if (8'h60 == _T_28[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_4;
      end else if (8'h60 == _T_25[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_3;
      end else if (8'h60 == _T_22[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_2;
      end else if (8'h60 == _T_19[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_1;
      end else if (8'h60 == _T_15[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_97 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h61 == _T_37[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_7;
      end else if (8'h61 == _T_34[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_6;
      end else if (8'h61 == _T_31[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_5;
      end else if (8'h61 == _T_28[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_4;
      end else if (8'h61 == _T_25[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_3;
      end else if (8'h61 == _T_22[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_2;
      end else if (8'h61 == _T_19[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_1;
      end else if (8'h61 == _T_15[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_98 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h62 == _T_37[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_7;
      end else if (8'h62 == _T_34[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_6;
      end else if (8'h62 == _T_31[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_5;
      end else if (8'h62 == _T_28[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_4;
      end else if (8'h62 == _T_25[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_3;
      end else if (8'h62 == _T_22[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_2;
      end else if (8'h62 == _T_19[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_1;
      end else if (8'h62 == _T_15[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_99 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h63 == _T_37[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_7;
      end else if (8'h63 == _T_34[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_6;
      end else if (8'h63 == _T_31[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_5;
      end else if (8'h63 == _T_28[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_4;
      end else if (8'h63 == _T_25[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_3;
      end else if (8'h63 == _T_22[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_2;
      end else if (8'h63 == _T_19[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_1;
      end else if (8'h63 == _T_15[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_100 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h64 == _T_37[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_7;
      end else if (8'h64 == _T_34[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_6;
      end else if (8'h64 == _T_31[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_5;
      end else if (8'h64 == _T_28[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_4;
      end else if (8'h64 == _T_25[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_3;
      end else if (8'h64 == _T_22[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_2;
      end else if (8'h64 == _T_19[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_1;
      end else if (8'h64 == _T_15[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_101 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h65 == _T_37[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_7;
      end else if (8'h65 == _T_34[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_6;
      end else if (8'h65 == _T_31[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_5;
      end else if (8'h65 == _T_28[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_4;
      end else if (8'h65 == _T_25[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_3;
      end else if (8'h65 == _T_22[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_2;
      end else if (8'h65 == _T_19[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_1;
      end else if (8'h65 == _T_15[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_102 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h66 == _T_37[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_7;
      end else if (8'h66 == _T_34[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_6;
      end else if (8'h66 == _T_31[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_5;
      end else if (8'h66 == _T_28[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_4;
      end else if (8'h66 == _T_25[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_3;
      end else if (8'h66 == _T_22[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_2;
      end else if (8'h66 == _T_19[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_1;
      end else if (8'h66 == _T_15[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_103 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h67 == _T_37[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_7;
      end else if (8'h67 == _T_34[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_6;
      end else if (8'h67 == _T_31[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_5;
      end else if (8'h67 == _T_28[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_4;
      end else if (8'h67 == _T_25[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_3;
      end else if (8'h67 == _T_22[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_2;
      end else if (8'h67 == _T_19[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_1;
      end else if (8'h67 == _T_15[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_104 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h68 == _T_37[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_7;
      end else if (8'h68 == _T_34[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_6;
      end else if (8'h68 == _T_31[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_5;
      end else if (8'h68 == _T_28[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_4;
      end else if (8'h68 == _T_25[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_3;
      end else if (8'h68 == _T_22[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_2;
      end else if (8'h68 == _T_19[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_1;
      end else if (8'h68 == _T_15[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_105 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h69 == _T_37[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_7;
      end else if (8'h69 == _T_34[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_6;
      end else if (8'h69 == _T_31[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_5;
      end else if (8'h69 == _T_28[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_4;
      end else if (8'h69 == _T_25[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_3;
      end else if (8'h69 == _T_22[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_2;
      end else if (8'h69 == _T_19[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_1;
      end else if (8'h69 == _T_15[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_106 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6a == _T_37[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_7;
      end else if (8'h6a == _T_34[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_6;
      end else if (8'h6a == _T_31[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_5;
      end else if (8'h6a == _T_28[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_4;
      end else if (8'h6a == _T_25[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_3;
      end else if (8'h6a == _T_22[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_2;
      end else if (8'h6a == _T_19[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_1;
      end else if (8'h6a == _T_15[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_107 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6b == _T_37[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_7;
      end else if (8'h6b == _T_34[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_6;
      end else if (8'h6b == _T_31[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_5;
      end else if (8'h6b == _T_28[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_4;
      end else if (8'h6b == _T_25[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_3;
      end else if (8'h6b == _T_22[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_2;
      end else if (8'h6b == _T_19[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_1;
      end else if (8'h6b == _T_15[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_108 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6c == _T_37[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_7;
      end else if (8'h6c == _T_34[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_6;
      end else if (8'h6c == _T_31[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_5;
      end else if (8'h6c == _T_28[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_4;
      end else if (8'h6c == _T_25[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_3;
      end else if (8'h6c == _T_22[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_2;
      end else if (8'h6c == _T_19[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_1;
      end else if (8'h6c == _T_15[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_109 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6d == _T_37[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_7;
      end else if (8'h6d == _T_34[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_6;
      end else if (8'h6d == _T_31[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_5;
      end else if (8'h6d == _T_28[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_4;
      end else if (8'h6d == _T_25[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_3;
      end else if (8'h6d == _T_22[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_2;
      end else if (8'h6d == _T_19[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_1;
      end else if (8'h6d == _T_15[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_110 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6e == _T_37[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_7;
      end else if (8'h6e == _T_34[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_6;
      end else if (8'h6e == _T_31[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_5;
      end else if (8'h6e == _T_28[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_4;
      end else if (8'h6e == _T_25[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_3;
      end else if (8'h6e == _T_22[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_2;
      end else if (8'h6e == _T_19[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_1;
      end else if (8'h6e == _T_15[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_111 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6f == _T_37[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_7;
      end else if (8'h6f == _T_34[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_6;
      end else if (8'h6f == _T_31[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_5;
      end else if (8'h6f == _T_28[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_4;
      end else if (8'h6f == _T_25[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_3;
      end else if (8'h6f == _T_22[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_2;
      end else if (8'h6f == _T_19[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_1;
      end else if (8'h6f == _T_15[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_112 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h70 == _T_37[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_7;
      end else if (8'h70 == _T_34[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_6;
      end else if (8'h70 == _T_31[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_5;
      end else if (8'h70 == _T_28[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_4;
      end else if (8'h70 == _T_25[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_3;
      end else if (8'h70 == _T_22[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_2;
      end else if (8'h70 == _T_19[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_1;
      end else if (8'h70 == _T_15[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_113 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h71 == _T_37[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_7;
      end else if (8'h71 == _T_34[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_6;
      end else if (8'h71 == _T_31[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_5;
      end else if (8'h71 == _T_28[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_4;
      end else if (8'h71 == _T_25[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_3;
      end else if (8'h71 == _T_22[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_2;
      end else if (8'h71 == _T_19[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_1;
      end else if (8'h71 == _T_15[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_114 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h72 == _T_37[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_7;
      end else if (8'h72 == _T_34[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_6;
      end else if (8'h72 == _T_31[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_5;
      end else if (8'h72 == _T_28[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_4;
      end else if (8'h72 == _T_25[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_3;
      end else if (8'h72 == _T_22[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_2;
      end else if (8'h72 == _T_19[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_1;
      end else if (8'h72 == _T_15[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_115 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h73 == _T_37[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_7;
      end else if (8'h73 == _T_34[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_6;
      end else if (8'h73 == _T_31[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_5;
      end else if (8'h73 == _T_28[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_4;
      end else if (8'h73 == _T_25[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_3;
      end else if (8'h73 == _T_22[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_2;
      end else if (8'h73 == _T_19[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_1;
      end else if (8'h73 == _T_15[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_116 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h74 == _T_37[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_7;
      end else if (8'h74 == _T_34[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_6;
      end else if (8'h74 == _T_31[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_5;
      end else if (8'h74 == _T_28[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_4;
      end else if (8'h74 == _T_25[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_3;
      end else if (8'h74 == _T_22[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_2;
      end else if (8'h74 == _T_19[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_1;
      end else if (8'h74 == _T_15[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_117 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h75 == _T_37[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_7;
      end else if (8'h75 == _T_34[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_6;
      end else if (8'h75 == _T_31[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_5;
      end else if (8'h75 == _T_28[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_4;
      end else if (8'h75 == _T_25[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_3;
      end else if (8'h75 == _T_22[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_2;
      end else if (8'h75 == _T_19[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_1;
      end else if (8'h75 == _T_15[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_118 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h76 == _T_37[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_7;
      end else if (8'h76 == _T_34[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_6;
      end else if (8'h76 == _T_31[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_5;
      end else if (8'h76 == _T_28[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_4;
      end else if (8'h76 == _T_25[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_3;
      end else if (8'h76 == _T_22[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_2;
      end else if (8'h76 == _T_19[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_1;
      end else if (8'h76 == _T_15[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_119 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h77 == _T_37[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_7;
      end else if (8'h77 == _T_34[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_6;
      end else if (8'h77 == _T_31[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_5;
      end else if (8'h77 == _T_28[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_4;
      end else if (8'h77 == _T_25[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_3;
      end else if (8'h77 == _T_22[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_2;
      end else if (8'h77 == _T_19[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_1;
      end else if (8'h77 == _T_15[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_120 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h78 == _T_37[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_7;
      end else if (8'h78 == _T_34[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_6;
      end else if (8'h78 == _T_31[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_5;
      end else if (8'h78 == _T_28[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_4;
      end else if (8'h78 == _T_25[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_3;
      end else if (8'h78 == _T_22[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_2;
      end else if (8'h78 == _T_19[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_1;
      end else if (8'h78 == _T_15[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_121 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h79 == _T_37[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_7;
      end else if (8'h79 == _T_34[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_6;
      end else if (8'h79 == _T_31[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_5;
      end else if (8'h79 == _T_28[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_4;
      end else if (8'h79 == _T_25[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_3;
      end else if (8'h79 == _T_22[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_2;
      end else if (8'h79 == _T_19[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_1;
      end else if (8'h79 == _T_15[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_122 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7a == _T_37[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_7;
      end else if (8'h7a == _T_34[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_6;
      end else if (8'h7a == _T_31[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_5;
      end else if (8'h7a == _T_28[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_4;
      end else if (8'h7a == _T_25[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_3;
      end else if (8'h7a == _T_22[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_2;
      end else if (8'h7a == _T_19[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_1;
      end else if (8'h7a == _T_15[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_123 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7b == _T_37[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_7;
      end else if (8'h7b == _T_34[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_6;
      end else if (8'h7b == _T_31[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_5;
      end else if (8'h7b == _T_28[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_4;
      end else if (8'h7b == _T_25[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_3;
      end else if (8'h7b == _T_22[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_2;
      end else if (8'h7b == _T_19[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_1;
      end else if (8'h7b == _T_15[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_124 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7c == _T_37[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_7;
      end else if (8'h7c == _T_34[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_6;
      end else if (8'h7c == _T_31[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_5;
      end else if (8'h7c == _T_28[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_4;
      end else if (8'h7c == _T_25[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_3;
      end else if (8'h7c == _T_22[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_2;
      end else if (8'h7c == _T_19[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_1;
      end else if (8'h7c == _T_15[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_125 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7d == _T_37[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_7;
      end else if (8'h7d == _T_34[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_6;
      end else if (8'h7d == _T_31[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_5;
      end else if (8'h7d == _T_28[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_4;
      end else if (8'h7d == _T_25[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_3;
      end else if (8'h7d == _T_22[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_2;
      end else if (8'h7d == _T_19[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_1;
      end else if (8'h7d == _T_15[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_126 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7e == _T_37[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_7;
      end else if (8'h7e == _T_34[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_6;
      end else if (8'h7e == _T_31[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_5;
      end else if (8'h7e == _T_28[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_4;
      end else if (8'h7e == _T_25[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_3;
      end else if (8'h7e == _T_22[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_2;
      end else if (8'h7e == _T_19[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_1;
      end else if (8'h7e == _T_15[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_127 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7f == _T_37[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_7;
      end else if (8'h7f == _T_34[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_6;
      end else if (8'h7f == _T_31[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_5;
      end else if (8'h7f == _T_28[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_4;
      end else if (8'h7f == _T_25[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_3;
      end else if (8'h7f == _T_22[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_2;
      end else if (8'h7f == _T_19[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_1;
      end else if (8'h7f == _T_15[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_128 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h80 == _T_37[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_7;
      end else if (8'h80 == _T_34[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_6;
      end else if (8'h80 == _T_31[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_5;
      end else if (8'h80 == _T_28[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_4;
      end else if (8'h80 == _T_25[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_3;
      end else if (8'h80 == _T_22[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_2;
      end else if (8'h80 == _T_19[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_1;
      end else if (8'h80 == _T_15[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_129 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h81 == _T_37[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_7;
      end else if (8'h81 == _T_34[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_6;
      end else if (8'h81 == _T_31[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_5;
      end else if (8'h81 == _T_28[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_4;
      end else if (8'h81 == _T_25[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_3;
      end else if (8'h81 == _T_22[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_2;
      end else if (8'h81 == _T_19[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_1;
      end else if (8'h81 == _T_15[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_130 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h82 == _T_37[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_7;
      end else if (8'h82 == _T_34[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_6;
      end else if (8'h82 == _T_31[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_5;
      end else if (8'h82 == _T_28[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_4;
      end else if (8'h82 == _T_25[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_3;
      end else if (8'h82 == _T_22[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_2;
      end else if (8'h82 == _T_19[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_1;
      end else if (8'h82 == _T_15[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_131 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h83 == _T_37[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_7;
      end else if (8'h83 == _T_34[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_6;
      end else if (8'h83 == _T_31[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_5;
      end else if (8'h83 == _T_28[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_4;
      end else if (8'h83 == _T_25[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_3;
      end else if (8'h83 == _T_22[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_2;
      end else if (8'h83 == _T_19[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_1;
      end else if (8'h83 == _T_15[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_132 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h84 == _T_37[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_7;
      end else if (8'h84 == _T_34[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_6;
      end else if (8'h84 == _T_31[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_5;
      end else if (8'h84 == _T_28[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_4;
      end else if (8'h84 == _T_25[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_3;
      end else if (8'h84 == _T_22[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_2;
      end else if (8'h84 == _T_19[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_1;
      end else if (8'h84 == _T_15[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_133 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h85 == _T_37[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_7;
      end else if (8'h85 == _T_34[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_6;
      end else if (8'h85 == _T_31[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_5;
      end else if (8'h85 == _T_28[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_4;
      end else if (8'h85 == _T_25[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_3;
      end else if (8'h85 == _T_22[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_2;
      end else if (8'h85 == _T_19[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_1;
      end else if (8'h85 == _T_15[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_134 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h86 == _T_37[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_7;
      end else if (8'h86 == _T_34[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_6;
      end else if (8'h86 == _T_31[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_5;
      end else if (8'h86 == _T_28[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_4;
      end else if (8'h86 == _T_25[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_3;
      end else if (8'h86 == _T_22[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_2;
      end else if (8'h86 == _T_19[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_1;
      end else if (8'h86 == _T_15[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_135 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h87 == _T_37[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_7;
      end else if (8'h87 == _T_34[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_6;
      end else if (8'h87 == _T_31[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_5;
      end else if (8'h87 == _T_28[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_4;
      end else if (8'h87 == _T_25[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_3;
      end else if (8'h87 == _T_22[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_2;
      end else if (8'h87 == _T_19[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_1;
      end else if (8'h87 == _T_15[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_136 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h88 == _T_37[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_7;
      end else if (8'h88 == _T_34[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_6;
      end else if (8'h88 == _T_31[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_5;
      end else if (8'h88 == _T_28[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_4;
      end else if (8'h88 == _T_25[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_3;
      end else if (8'h88 == _T_22[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_2;
      end else if (8'h88 == _T_19[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_1;
      end else if (8'h88 == _T_15[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_137 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h89 == _T_37[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_7;
      end else if (8'h89 == _T_34[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_6;
      end else if (8'h89 == _T_31[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_5;
      end else if (8'h89 == _T_28[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_4;
      end else if (8'h89 == _T_25[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_3;
      end else if (8'h89 == _T_22[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_2;
      end else if (8'h89 == _T_19[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_1;
      end else if (8'h89 == _T_15[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_138 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8a == _T_37[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_7;
      end else if (8'h8a == _T_34[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_6;
      end else if (8'h8a == _T_31[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_5;
      end else if (8'h8a == _T_28[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_4;
      end else if (8'h8a == _T_25[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_3;
      end else if (8'h8a == _T_22[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_2;
      end else if (8'h8a == _T_19[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_1;
      end else if (8'h8a == _T_15[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_139 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8b == _T_37[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_7;
      end else if (8'h8b == _T_34[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_6;
      end else if (8'h8b == _T_31[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_5;
      end else if (8'h8b == _T_28[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_4;
      end else if (8'h8b == _T_25[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_3;
      end else if (8'h8b == _T_22[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_2;
      end else if (8'h8b == _T_19[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_1;
      end else if (8'h8b == _T_15[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_140 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8c == _T_37[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_7;
      end else if (8'h8c == _T_34[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_6;
      end else if (8'h8c == _T_31[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_5;
      end else if (8'h8c == _T_28[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_4;
      end else if (8'h8c == _T_25[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_3;
      end else if (8'h8c == _T_22[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_2;
      end else if (8'h8c == _T_19[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_1;
      end else if (8'h8c == _T_15[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_141 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8d == _T_37[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_7;
      end else if (8'h8d == _T_34[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_6;
      end else if (8'h8d == _T_31[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_5;
      end else if (8'h8d == _T_28[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_4;
      end else if (8'h8d == _T_25[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_3;
      end else if (8'h8d == _T_22[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_2;
      end else if (8'h8d == _T_19[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_1;
      end else if (8'h8d == _T_15[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_142 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8e == _T_37[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_7;
      end else if (8'h8e == _T_34[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_6;
      end else if (8'h8e == _T_31[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_5;
      end else if (8'h8e == _T_28[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_4;
      end else if (8'h8e == _T_25[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_3;
      end else if (8'h8e == _T_22[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_2;
      end else if (8'h8e == _T_19[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_1;
      end else if (8'h8e == _T_15[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_143 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8f == _T_37[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_7;
      end else if (8'h8f == _T_34[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_6;
      end else if (8'h8f == _T_31[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_5;
      end else if (8'h8f == _T_28[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_4;
      end else if (8'h8f == _T_25[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_3;
      end else if (8'h8f == _T_22[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_2;
      end else if (8'h8f == _T_19[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_1;
      end else if (8'h8f == _T_15[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_144 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h90 == _T_37[7:0]) begin
        image_1_144 <= io_pixelVal_in_1_7;
      end else if (8'h90 == _T_34[7:0]) begin
        image_1_144 <= io_pixelVal_in_1_6;
      end else if (8'h90 == _T_31[7:0]) begin
        image_1_144 <= io_pixelVal_in_1_5;
      end else if (8'h90 == _T_28[7:0]) begin
        image_1_144 <= io_pixelVal_in_1_4;
      end else if (8'h90 == _T_25[7:0]) begin
        image_1_144 <= io_pixelVal_in_1_3;
      end else if (8'h90 == _T_22[7:0]) begin
        image_1_144 <= io_pixelVal_in_1_2;
      end else if (8'h90 == _T_19[7:0]) begin
        image_1_144 <= io_pixelVal_in_1_1;
      end else if (8'h90 == _T_15[7:0]) begin
        image_1_144 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_145 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h91 == _T_37[7:0]) begin
        image_1_145 <= io_pixelVal_in_1_7;
      end else if (8'h91 == _T_34[7:0]) begin
        image_1_145 <= io_pixelVal_in_1_6;
      end else if (8'h91 == _T_31[7:0]) begin
        image_1_145 <= io_pixelVal_in_1_5;
      end else if (8'h91 == _T_28[7:0]) begin
        image_1_145 <= io_pixelVal_in_1_4;
      end else if (8'h91 == _T_25[7:0]) begin
        image_1_145 <= io_pixelVal_in_1_3;
      end else if (8'h91 == _T_22[7:0]) begin
        image_1_145 <= io_pixelVal_in_1_2;
      end else if (8'h91 == _T_19[7:0]) begin
        image_1_145 <= io_pixelVal_in_1_1;
      end else if (8'h91 == _T_15[7:0]) begin
        image_1_145 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_146 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h92 == _T_37[7:0]) begin
        image_1_146 <= io_pixelVal_in_1_7;
      end else if (8'h92 == _T_34[7:0]) begin
        image_1_146 <= io_pixelVal_in_1_6;
      end else if (8'h92 == _T_31[7:0]) begin
        image_1_146 <= io_pixelVal_in_1_5;
      end else if (8'h92 == _T_28[7:0]) begin
        image_1_146 <= io_pixelVal_in_1_4;
      end else if (8'h92 == _T_25[7:0]) begin
        image_1_146 <= io_pixelVal_in_1_3;
      end else if (8'h92 == _T_22[7:0]) begin
        image_1_146 <= io_pixelVal_in_1_2;
      end else if (8'h92 == _T_19[7:0]) begin
        image_1_146 <= io_pixelVal_in_1_1;
      end else if (8'h92 == _T_15[7:0]) begin
        image_1_146 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_147 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h93 == _T_37[7:0]) begin
        image_1_147 <= io_pixelVal_in_1_7;
      end else if (8'h93 == _T_34[7:0]) begin
        image_1_147 <= io_pixelVal_in_1_6;
      end else if (8'h93 == _T_31[7:0]) begin
        image_1_147 <= io_pixelVal_in_1_5;
      end else if (8'h93 == _T_28[7:0]) begin
        image_1_147 <= io_pixelVal_in_1_4;
      end else if (8'h93 == _T_25[7:0]) begin
        image_1_147 <= io_pixelVal_in_1_3;
      end else if (8'h93 == _T_22[7:0]) begin
        image_1_147 <= io_pixelVal_in_1_2;
      end else if (8'h93 == _T_19[7:0]) begin
        image_1_147 <= io_pixelVal_in_1_1;
      end else if (8'h93 == _T_15[7:0]) begin
        image_1_147 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_148 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h94 == _T_37[7:0]) begin
        image_1_148 <= io_pixelVal_in_1_7;
      end else if (8'h94 == _T_34[7:0]) begin
        image_1_148 <= io_pixelVal_in_1_6;
      end else if (8'h94 == _T_31[7:0]) begin
        image_1_148 <= io_pixelVal_in_1_5;
      end else if (8'h94 == _T_28[7:0]) begin
        image_1_148 <= io_pixelVal_in_1_4;
      end else if (8'h94 == _T_25[7:0]) begin
        image_1_148 <= io_pixelVal_in_1_3;
      end else if (8'h94 == _T_22[7:0]) begin
        image_1_148 <= io_pixelVal_in_1_2;
      end else if (8'h94 == _T_19[7:0]) begin
        image_1_148 <= io_pixelVal_in_1_1;
      end else if (8'h94 == _T_15[7:0]) begin
        image_1_148 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_149 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h95 == _T_37[7:0]) begin
        image_1_149 <= io_pixelVal_in_1_7;
      end else if (8'h95 == _T_34[7:0]) begin
        image_1_149 <= io_pixelVal_in_1_6;
      end else if (8'h95 == _T_31[7:0]) begin
        image_1_149 <= io_pixelVal_in_1_5;
      end else if (8'h95 == _T_28[7:0]) begin
        image_1_149 <= io_pixelVal_in_1_4;
      end else if (8'h95 == _T_25[7:0]) begin
        image_1_149 <= io_pixelVal_in_1_3;
      end else if (8'h95 == _T_22[7:0]) begin
        image_1_149 <= io_pixelVal_in_1_2;
      end else if (8'h95 == _T_19[7:0]) begin
        image_1_149 <= io_pixelVal_in_1_1;
      end else if (8'h95 == _T_15[7:0]) begin
        image_1_149 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_150 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h96 == _T_37[7:0]) begin
        image_1_150 <= io_pixelVal_in_1_7;
      end else if (8'h96 == _T_34[7:0]) begin
        image_1_150 <= io_pixelVal_in_1_6;
      end else if (8'h96 == _T_31[7:0]) begin
        image_1_150 <= io_pixelVal_in_1_5;
      end else if (8'h96 == _T_28[7:0]) begin
        image_1_150 <= io_pixelVal_in_1_4;
      end else if (8'h96 == _T_25[7:0]) begin
        image_1_150 <= io_pixelVal_in_1_3;
      end else if (8'h96 == _T_22[7:0]) begin
        image_1_150 <= io_pixelVal_in_1_2;
      end else if (8'h96 == _T_19[7:0]) begin
        image_1_150 <= io_pixelVal_in_1_1;
      end else if (8'h96 == _T_15[7:0]) begin
        image_1_150 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_151 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h97 == _T_37[7:0]) begin
        image_1_151 <= io_pixelVal_in_1_7;
      end else if (8'h97 == _T_34[7:0]) begin
        image_1_151 <= io_pixelVal_in_1_6;
      end else if (8'h97 == _T_31[7:0]) begin
        image_1_151 <= io_pixelVal_in_1_5;
      end else if (8'h97 == _T_28[7:0]) begin
        image_1_151 <= io_pixelVal_in_1_4;
      end else if (8'h97 == _T_25[7:0]) begin
        image_1_151 <= io_pixelVal_in_1_3;
      end else if (8'h97 == _T_22[7:0]) begin
        image_1_151 <= io_pixelVal_in_1_2;
      end else if (8'h97 == _T_19[7:0]) begin
        image_1_151 <= io_pixelVal_in_1_1;
      end else if (8'h97 == _T_15[7:0]) begin
        image_1_151 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_152 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h98 == _T_37[7:0]) begin
        image_1_152 <= io_pixelVal_in_1_7;
      end else if (8'h98 == _T_34[7:0]) begin
        image_1_152 <= io_pixelVal_in_1_6;
      end else if (8'h98 == _T_31[7:0]) begin
        image_1_152 <= io_pixelVal_in_1_5;
      end else if (8'h98 == _T_28[7:0]) begin
        image_1_152 <= io_pixelVal_in_1_4;
      end else if (8'h98 == _T_25[7:0]) begin
        image_1_152 <= io_pixelVal_in_1_3;
      end else if (8'h98 == _T_22[7:0]) begin
        image_1_152 <= io_pixelVal_in_1_2;
      end else if (8'h98 == _T_19[7:0]) begin
        image_1_152 <= io_pixelVal_in_1_1;
      end else if (8'h98 == _T_15[7:0]) begin
        image_1_152 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_153 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h99 == _T_37[7:0]) begin
        image_1_153 <= io_pixelVal_in_1_7;
      end else if (8'h99 == _T_34[7:0]) begin
        image_1_153 <= io_pixelVal_in_1_6;
      end else if (8'h99 == _T_31[7:0]) begin
        image_1_153 <= io_pixelVal_in_1_5;
      end else if (8'h99 == _T_28[7:0]) begin
        image_1_153 <= io_pixelVal_in_1_4;
      end else if (8'h99 == _T_25[7:0]) begin
        image_1_153 <= io_pixelVal_in_1_3;
      end else if (8'h99 == _T_22[7:0]) begin
        image_1_153 <= io_pixelVal_in_1_2;
      end else if (8'h99 == _T_19[7:0]) begin
        image_1_153 <= io_pixelVal_in_1_1;
      end else if (8'h99 == _T_15[7:0]) begin
        image_1_153 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_154 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9a == _T_37[7:0]) begin
        image_1_154 <= io_pixelVal_in_1_7;
      end else if (8'h9a == _T_34[7:0]) begin
        image_1_154 <= io_pixelVal_in_1_6;
      end else if (8'h9a == _T_31[7:0]) begin
        image_1_154 <= io_pixelVal_in_1_5;
      end else if (8'h9a == _T_28[7:0]) begin
        image_1_154 <= io_pixelVal_in_1_4;
      end else if (8'h9a == _T_25[7:0]) begin
        image_1_154 <= io_pixelVal_in_1_3;
      end else if (8'h9a == _T_22[7:0]) begin
        image_1_154 <= io_pixelVal_in_1_2;
      end else if (8'h9a == _T_19[7:0]) begin
        image_1_154 <= io_pixelVal_in_1_1;
      end else if (8'h9a == _T_15[7:0]) begin
        image_1_154 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_155 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9b == _T_37[7:0]) begin
        image_1_155 <= io_pixelVal_in_1_7;
      end else if (8'h9b == _T_34[7:0]) begin
        image_1_155 <= io_pixelVal_in_1_6;
      end else if (8'h9b == _T_31[7:0]) begin
        image_1_155 <= io_pixelVal_in_1_5;
      end else if (8'h9b == _T_28[7:0]) begin
        image_1_155 <= io_pixelVal_in_1_4;
      end else if (8'h9b == _T_25[7:0]) begin
        image_1_155 <= io_pixelVal_in_1_3;
      end else if (8'h9b == _T_22[7:0]) begin
        image_1_155 <= io_pixelVal_in_1_2;
      end else if (8'h9b == _T_19[7:0]) begin
        image_1_155 <= io_pixelVal_in_1_1;
      end else if (8'h9b == _T_15[7:0]) begin
        image_1_155 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_156 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9c == _T_37[7:0]) begin
        image_1_156 <= io_pixelVal_in_1_7;
      end else if (8'h9c == _T_34[7:0]) begin
        image_1_156 <= io_pixelVal_in_1_6;
      end else if (8'h9c == _T_31[7:0]) begin
        image_1_156 <= io_pixelVal_in_1_5;
      end else if (8'h9c == _T_28[7:0]) begin
        image_1_156 <= io_pixelVal_in_1_4;
      end else if (8'h9c == _T_25[7:0]) begin
        image_1_156 <= io_pixelVal_in_1_3;
      end else if (8'h9c == _T_22[7:0]) begin
        image_1_156 <= io_pixelVal_in_1_2;
      end else if (8'h9c == _T_19[7:0]) begin
        image_1_156 <= io_pixelVal_in_1_1;
      end else if (8'h9c == _T_15[7:0]) begin
        image_1_156 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_157 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9d == _T_37[7:0]) begin
        image_1_157 <= io_pixelVal_in_1_7;
      end else if (8'h9d == _T_34[7:0]) begin
        image_1_157 <= io_pixelVal_in_1_6;
      end else if (8'h9d == _T_31[7:0]) begin
        image_1_157 <= io_pixelVal_in_1_5;
      end else if (8'h9d == _T_28[7:0]) begin
        image_1_157 <= io_pixelVal_in_1_4;
      end else if (8'h9d == _T_25[7:0]) begin
        image_1_157 <= io_pixelVal_in_1_3;
      end else if (8'h9d == _T_22[7:0]) begin
        image_1_157 <= io_pixelVal_in_1_2;
      end else if (8'h9d == _T_19[7:0]) begin
        image_1_157 <= io_pixelVal_in_1_1;
      end else if (8'h9d == _T_15[7:0]) begin
        image_1_157 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_158 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9e == _T_37[7:0]) begin
        image_1_158 <= io_pixelVal_in_1_7;
      end else if (8'h9e == _T_34[7:0]) begin
        image_1_158 <= io_pixelVal_in_1_6;
      end else if (8'h9e == _T_31[7:0]) begin
        image_1_158 <= io_pixelVal_in_1_5;
      end else if (8'h9e == _T_28[7:0]) begin
        image_1_158 <= io_pixelVal_in_1_4;
      end else if (8'h9e == _T_25[7:0]) begin
        image_1_158 <= io_pixelVal_in_1_3;
      end else if (8'h9e == _T_22[7:0]) begin
        image_1_158 <= io_pixelVal_in_1_2;
      end else if (8'h9e == _T_19[7:0]) begin
        image_1_158 <= io_pixelVal_in_1_1;
      end else if (8'h9e == _T_15[7:0]) begin
        image_1_158 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_159 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9f == _T_37[7:0]) begin
        image_1_159 <= io_pixelVal_in_1_7;
      end else if (8'h9f == _T_34[7:0]) begin
        image_1_159 <= io_pixelVal_in_1_6;
      end else if (8'h9f == _T_31[7:0]) begin
        image_1_159 <= io_pixelVal_in_1_5;
      end else if (8'h9f == _T_28[7:0]) begin
        image_1_159 <= io_pixelVal_in_1_4;
      end else if (8'h9f == _T_25[7:0]) begin
        image_1_159 <= io_pixelVal_in_1_3;
      end else if (8'h9f == _T_22[7:0]) begin
        image_1_159 <= io_pixelVal_in_1_2;
      end else if (8'h9f == _T_19[7:0]) begin
        image_1_159 <= io_pixelVal_in_1_1;
      end else if (8'h9f == _T_15[7:0]) begin
        image_1_159 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_160 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha0 == _T_37[7:0]) begin
        image_1_160 <= io_pixelVal_in_1_7;
      end else if (8'ha0 == _T_34[7:0]) begin
        image_1_160 <= io_pixelVal_in_1_6;
      end else if (8'ha0 == _T_31[7:0]) begin
        image_1_160 <= io_pixelVal_in_1_5;
      end else if (8'ha0 == _T_28[7:0]) begin
        image_1_160 <= io_pixelVal_in_1_4;
      end else if (8'ha0 == _T_25[7:0]) begin
        image_1_160 <= io_pixelVal_in_1_3;
      end else if (8'ha0 == _T_22[7:0]) begin
        image_1_160 <= io_pixelVal_in_1_2;
      end else if (8'ha0 == _T_19[7:0]) begin
        image_1_160 <= io_pixelVal_in_1_1;
      end else if (8'ha0 == _T_15[7:0]) begin
        image_1_160 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_161 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha1 == _T_37[7:0]) begin
        image_1_161 <= io_pixelVal_in_1_7;
      end else if (8'ha1 == _T_34[7:0]) begin
        image_1_161 <= io_pixelVal_in_1_6;
      end else if (8'ha1 == _T_31[7:0]) begin
        image_1_161 <= io_pixelVal_in_1_5;
      end else if (8'ha1 == _T_28[7:0]) begin
        image_1_161 <= io_pixelVal_in_1_4;
      end else if (8'ha1 == _T_25[7:0]) begin
        image_1_161 <= io_pixelVal_in_1_3;
      end else if (8'ha1 == _T_22[7:0]) begin
        image_1_161 <= io_pixelVal_in_1_2;
      end else if (8'ha1 == _T_19[7:0]) begin
        image_1_161 <= io_pixelVal_in_1_1;
      end else if (8'ha1 == _T_15[7:0]) begin
        image_1_161 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_162 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha2 == _T_37[7:0]) begin
        image_1_162 <= io_pixelVal_in_1_7;
      end else if (8'ha2 == _T_34[7:0]) begin
        image_1_162 <= io_pixelVal_in_1_6;
      end else if (8'ha2 == _T_31[7:0]) begin
        image_1_162 <= io_pixelVal_in_1_5;
      end else if (8'ha2 == _T_28[7:0]) begin
        image_1_162 <= io_pixelVal_in_1_4;
      end else if (8'ha2 == _T_25[7:0]) begin
        image_1_162 <= io_pixelVal_in_1_3;
      end else if (8'ha2 == _T_22[7:0]) begin
        image_1_162 <= io_pixelVal_in_1_2;
      end else if (8'ha2 == _T_19[7:0]) begin
        image_1_162 <= io_pixelVal_in_1_1;
      end else if (8'ha2 == _T_15[7:0]) begin
        image_1_162 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_163 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha3 == _T_37[7:0]) begin
        image_1_163 <= io_pixelVal_in_1_7;
      end else if (8'ha3 == _T_34[7:0]) begin
        image_1_163 <= io_pixelVal_in_1_6;
      end else if (8'ha3 == _T_31[7:0]) begin
        image_1_163 <= io_pixelVal_in_1_5;
      end else if (8'ha3 == _T_28[7:0]) begin
        image_1_163 <= io_pixelVal_in_1_4;
      end else if (8'ha3 == _T_25[7:0]) begin
        image_1_163 <= io_pixelVal_in_1_3;
      end else if (8'ha3 == _T_22[7:0]) begin
        image_1_163 <= io_pixelVal_in_1_2;
      end else if (8'ha3 == _T_19[7:0]) begin
        image_1_163 <= io_pixelVal_in_1_1;
      end else if (8'ha3 == _T_15[7:0]) begin
        image_1_163 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_164 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha4 == _T_37[7:0]) begin
        image_1_164 <= io_pixelVal_in_1_7;
      end else if (8'ha4 == _T_34[7:0]) begin
        image_1_164 <= io_pixelVal_in_1_6;
      end else if (8'ha4 == _T_31[7:0]) begin
        image_1_164 <= io_pixelVal_in_1_5;
      end else if (8'ha4 == _T_28[7:0]) begin
        image_1_164 <= io_pixelVal_in_1_4;
      end else if (8'ha4 == _T_25[7:0]) begin
        image_1_164 <= io_pixelVal_in_1_3;
      end else if (8'ha4 == _T_22[7:0]) begin
        image_1_164 <= io_pixelVal_in_1_2;
      end else if (8'ha4 == _T_19[7:0]) begin
        image_1_164 <= io_pixelVal_in_1_1;
      end else if (8'ha4 == _T_15[7:0]) begin
        image_1_164 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_165 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha5 == _T_37[7:0]) begin
        image_1_165 <= io_pixelVal_in_1_7;
      end else if (8'ha5 == _T_34[7:0]) begin
        image_1_165 <= io_pixelVal_in_1_6;
      end else if (8'ha5 == _T_31[7:0]) begin
        image_1_165 <= io_pixelVal_in_1_5;
      end else if (8'ha5 == _T_28[7:0]) begin
        image_1_165 <= io_pixelVal_in_1_4;
      end else if (8'ha5 == _T_25[7:0]) begin
        image_1_165 <= io_pixelVal_in_1_3;
      end else if (8'ha5 == _T_22[7:0]) begin
        image_1_165 <= io_pixelVal_in_1_2;
      end else if (8'ha5 == _T_19[7:0]) begin
        image_1_165 <= io_pixelVal_in_1_1;
      end else if (8'ha5 == _T_15[7:0]) begin
        image_1_165 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_166 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha6 == _T_37[7:0]) begin
        image_1_166 <= io_pixelVal_in_1_7;
      end else if (8'ha6 == _T_34[7:0]) begin
        image_1_166 <= io_pixelVal_in_1_6;
      end else if (8'ha6 == _T_31[7:0]) begin
        image_1_166 <= io_pixelVal_in_1_5;
      end else if (8'ha6 == _T_28[7:0]) begin
        image_1_166 <= io_pixelVal_in_1_4;
      end else if (8'ha6 == _T_25[7:0]) begin
        image_1_166 <= io_pixelVal_in_1_3;
      end else if (8'ha6 == _T_22[7:0]) begin
        image_1_166 <= io_pixelVal_in_1_2;
      end else if (8'ha6 == _T_19[7:0]) begin
        image_1_166 <= io_pixelVal_in_1_1;
      end else if (8'ha6 == _T_15[7:0]) begin
        image_1_166 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_167 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha7 == _T_37[7:0]) begin
        image_1_167 <= io_pixelVal_in_1_7;
      end else if (8'ha7 == _T_34[7:0]) begin
        image_1_167 <= io_pixelVal_in_1_6;
      end else if (8'ha7 == _T_31[7:0]) begin
        image_1_167 <= io_pixelVal_in_1_5;
      end else if (8'ha7 == _T_28[7:0]) begin
        image_1_167 <= io_pixelVal_in_1_4;
      end else if (8'ha7 == _T_25[7:0]) begin
        image_1_167 <= io_pixelVal_in_1_3;
      end else if (8'ha7 == _T_22[7:0]) begin
        image_1_167 <= io_pixelVal_in_1_2;
      end else if (8'ha7 == _T_19[7:0]) begin
        image_1_167 <= io_pixelVal_in_1_1;
      end else if (8'ha7 == _T_15[7:0]) begin
        image_1_167 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_168 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha8 == _T_37[7:0]) begin
        image_1_168 <= io_pixelVal_in_1_7;
      end else if (8'ha8 == _T_34[7:0]) begin
        image_1_168 <= io_pixelVal_in_1_6;
      end else if (8'ha8 == _T_31[7:0]) begin
        image_1_168 <= io_pixelVal_in_1_5;
      end else if (8'ha8 == _T_28[7:0]) begin
        image_1_168 <= io_pixelVal_in_1_4;
      end else if (8'ha8 == _T_25[7:0]) begin
        image_1_168 <= io_pixelVal_in_1_3;
      end else if (8'ha8 == _T_22[7:0]) begin
        image_1_168 <= io_pixelVal_in_1_2;
      end else if (8'ha8 == _T_19[7:0]) begin
        image_1_168 <= io_pixelVal_in_1_1;
      end else if (8'ha8 == _T_15[7:0]) begin
        image_1_168 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_169 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha9 == _T_37[7:0]) begin
        image_1_169 <= io_pixelVal_in_1_7;
      end else if (8'ha9 == _T_34[7:0]) begin
        image_1_169 <= io_pixelVal_in_1_6;
      end else if (8'ha9 == _T_31[7:0]) begin
        image_1_169 <= io_pixelVal_in_1_5;
      end else if (8'ha9 == _T_28[7:0]) begin
        image_1_169 <= io_pixelVal_in_1_4;
      end else if (8'ha9 == _T_25[7:0]) begin
        image_1_169 <= io_pixelVal_in_1_3;
      end else if (8'ha9 == _T_22[7:0]) begin
        image_1_169 <= io_pixelVal_in_1_2;
      end else if (8'ha9 == _T_19[7:0]) begin
        image_1_169 <= io_pixelVal_in_1_1;
      end else if (8'ha9 == _T_15[7:0]) begin
        image_1_169 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_170 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'haa == _T_37[7:0]) begin
        image_1_170 <= io_pixelVal_in_1_7;
      end else if (8'haa == _T_34[7:0]) begin
        image_1_170 <= io_pixelVal_in_1_6;
      end else if (8'haa == _T_31[7:0]) begin
        image_1_170 <= io_pixelVal_in_1_5;
      end else if (8'haa == _T_28[7:0]) begin
        image_1_170 <= io_pixelVal_in_1_4;
      end else if (8'haa == _T_25[7:0]) begin
        image_1_170 <= io_pixelVal_in_1_3;
      end else if (8'haa == _T_22[7:0]) begin
        image_1_170 <= io_pixelVal_in_1_2;
      end else if (8'haa == _T_19[7:0]) begin
        image_1_170 <= io_pixelVal_in_1_1;
      end else if (8'haa == _T_15[7:0]) begin
        image_1_170 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_171 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hab == _T_37[7:0]) begin
        image_1_171 <= io_pixelVal_in_1_7;
      end else if (8'hab == _T_34[7:0]) begin
        image_1_171 <= io_pixelVal_in_1_6;
      end else if (8'hab == _T_31[7:0]) begin
        image_1_171 <= io_pixelVal_in_1_5;
      end else if (8'hab == _T_28[7:0]) begin
        image_1_171 <= io_pixelVal_in_1_4;
      end else if (8'hab == _T_25[7:0]) begin
        image_1_171 <= io_pixelVal_in_1_3;
      end else if (8'hab == _T_22[7:0]) begin
        image_1_171 <= io_pixelVal_in_1_2;
      end else if (8'hab == _T_19[7:0]) begin
        image_1_171 <= io_pixelVal_in_1_1;
      end else if (8'hab == _T_15[7:0]) begin
        image_1_171 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_172 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hac == _T_37[7:0]) begin
        image_1_172 <= io_pixelVal_in_1_7;
      end else if (8'hac == _T_34[7:0]) begin
        image_1_172 <= io_pixelVal_in_1_6;
      end else if (8'hac == _T_31[7:0]) begin
        image_1_172 <= io_pixelVal_in_1_5;
      end else if (8'hac == _T_28[7:0]) begin
        image_1_172 <= io_pixelVal_in_1_4;
      end else if (8'hac == _T_25[7:0]) begin
        image_1_172 <= io_pixelVal_in_1_3;
      end else if (8'hac == _T_22[7:0]) begin
        image_1_172 <= io_pixelVal_in_1_2;
      end else if (8'hac == _T_19[7:0]) begin
        image_1_172 <= io_pixelVal_in_1_1;
      end else if (8'hac == _T_15[7:0]) begin
        image_1_172 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_173 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'had == _T_37[7:0]) begin
        image_1_173 <= io_pixelVal_in_1_7;
      end else if (8'had == _T_34[7:0]) begin
        image_1_173 <= io_pixelVal_in_1_6;
      end else if (8'had == _T_31[7:0]) begin
        image_1_173 <= io_pixelVal_in_1_5;
      end else if (8'had == _T_28[7:0]) begin
        image_1_173 <= io_pixelVal_in_1_4;
      end else if (8'had == _T_25[7:0]) begin
        image_1_173 <= io_pixelVal_in_1_3;
      end else if (8'had == _T_22[7:0]) begin
        image_1_173 <= io_pixelVal_in_1_2;
      end else if (8'had == _T_19[7:0]) begin
        image_1_173 <= io_pixelVal_in_1_1;
      end else if (8'had == _T_15[7:0]) begin
        image_1_173 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_174 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hae == _T_37[7:0]) begin
        image_1_174 <= io_pixelVal_in_1_7;
      end else if (8'hae == _T_34[7:0]) begin
        image_1_174 <= io_pixelVal_in_1_6;
      end else if (8'hae == _T_31[7:0]) begin
        image_1_174 <= io_pixelVal_in_1_5;
      end else if (8'hae == _T_28[7:0]) begin
        image_1_174 <= io_pixelVal_in_1_4;
      end else if (8'hae == _T_25[7:0]) begin
        image_1_174 <= io_pixelVal_in_1_3;
      end else if (8'hae == _T_22[7:0]) begin
        image_1_174 <= io_pixelVal_in_1_2;
      end else if (8'hae == _T_19[7:0]) begin
        image_1_174 <= io_pixelVal_in_1_1;
      end else if (8'hae == _T_15[7:0]) begin
        image_1_174 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_175 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'haf == _T_37[7:0]) begin
        image_1_175 <= io_pixelVal_in_1_7;
      end else if (8'haf == _T_34[7:0]) begin
        image_1_175 <= io_pixelVal_in_1_6;
      end else if (8'haf == _T_31[7:0]) begin
        image_1_175 <= io_pixelVal_in_1_5;
      end else if (8'haf == _T_28[7:0]) begin
        image_1_175 <= io_pixelVal_in_1_4;
      end else if (8'haf == _T_25[7:0]) begin
        image_1_175 <= io_pixelVal_in_1_3;
      end else if (8'haf == _T_22[7:0]) begin
        image_1_175 <= io_pixelVal_in_1_2;
      end else if (8'haf == _T_19[7:0]) begin
        image_1_175 <= io_pixelVal_in_1_1;
      end else if (8'haf == _T_15[7:0]) begin
        image_1_175 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_176 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb0 == _T_37[7:0]) begin
        image_1_176 <= io_pixelVal_in_1_7;
      end else if (8'hb0 == _T_34[7:0]) begin
        image_1_176 <= io_pixelVal_in_1_6;
      end else if (8'hb0 == _T_31[7:0]) begin
        image_1_176 <= io_pixelVal_in_1_5;
      end else if (8'hb0 == _T_28[7:0]) begin
        image_1_176 <= io_pixelVal_in_1_4;
      end else if (8'hb0 == _T_25[7:0]) begin
        image_1_176 <= io_pixelVal_in_1_3;
      end else if (8'hb0 == _T_22[7:0]) begin
        image_1_176 <= io_pixelVal_in_1_2;
      end else if (8'hb0 == _T_19[7:0]) begin
        image_1_176 <= io_pixelVal_in_1_1;
      end else if (8'hb0 == _T_15[7:0]) begin
        image_1_176 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_177 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb1 == _T_37[7:0]) begin
        image_1_177 <= io_pixelVal_in_1_7;
      end else if (8'hb1 == _T_34[7:0]) begin
        image_1_177 <= io_pixelVal_in_1_6;
      end else if (8'hb1 == _T_31[7:0]) begin
        image_1_177 <= io_pixelVal_in_1_5;
      end else if (8'hb1 == _T_28[7:0]) begin
        image_1_177 <= io_pixelVal_in_1_4;
      end else if (8'hb1 == _T_25[7:0]) begin
        image_1_177 <= io_pixelVal_in_1_3;
      end else if (8'hb1 == _T_22[7:0]) begin
        image_1_177 <= io_pixelVal_in_1_2;
      end else if (8'hb1 == _T_19[7:0]) begin
        image_1_177 <= io_pixelVal_in_1_1;
      end else if (8'hb1 == _T_15[7:0]) begin
        image_1_177 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_178 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb2 == _T_37[7:0]) begin
        image_1_178 <= io_pixelVal_in_1_7;
      end else if (8'hb2 == _T_34[7:0]) begin
        image_1_178 <= io_pixelVal_in_1_6;
      end else if (8'hb2 == _T_31[7:0]) begin
        image_1_178 <= io_pixelVal_in_1_5;
      end else if (8'hb2 == _T_28[7:0]) begin
        image_1_178 <= io_pixelVal_in_1_4;
      end else if (8'hb2 == _T_25[7:0]) begin
        image_1_178 <= io_pixelVal_in_1_3;
      end else if (8'hb2 == _T_22[7:0]) begin
        image_1_178 <= io_pixelVal_in_1_2;
      end else if (8'hb2 == _T_19[7:0]) begin
        image_1_178 <= io_pixelVal_in_1_1;
      end else if (8'hb2 == _T_15[7:0]) begin
        image_1_178 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_179 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb3 == _T_37[7:0]) begin
        image_1_179 <= io_pixelVal_in_1_7;
      end else if (8'hb3 == _T_34[7:0]) begin
        image_1_179 <= io_pixelVal_in_1_6;
      end else if (8'hb3 == _T_31[7:0]) begin
        image_1_179 <= io_pixelVal_in_1_5;
      end else if (8'hb3 == _T_28[7:0]) begin
        image_1_179 <= io_pixelVal_in_1_4;
      end else if (8'hb3 == _T_25[7:0]) begin
        image_1_179 <= io_pixelVal_in_1_3;
      end else if (8'hb3 == _T_22[7:0]) begin
        image_1_179 <= io_pixelVal_in_1_2;
      end else if (8'hb3 == _T_19[7:0]) begin
        image_1_179 <= io_pixelVal_in_1_1;
      end else if (8'hb3 == _T_15[7:0]) begin
        image_1_179 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_180 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb4 == _T_37[7:0]) begin
        image_1_180 <= io_pixelVal_in_1_7;
      end else if (8'hb4 == _T_34[7:0]) begin
        image_1_180 <= io_pixelVal_in_1_6;
      end else if (8'hb4 == _T_31[7:0]) begin
        image_1_180 <= io_pixelVal_in_1_5;
      end else if (8'hb4 == _T_28[7:0]) begin
        image_1_180 <= io_pixelVal_in_1_4;
      end else if (8'hb4 == _T_25[7:0]) begin
        image_1_180 <= io_pixelVal_in_1_3;
      end else if (8'hb4 == _T_22[7:0]) begin
        image_1_180 <= io_pixelVal_in_1_2;
      end else if (8'hb4 == _T_19[7:0]) begin
        image_1_180 <= io_pixelVal_in_1_1;
      end else if (8'hb4 == _T_15[7:0]) begin
        image_1_180 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_181 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb5 == _T_37[7:0]) begin
        image_1_181 <= io_pixelVal_in_1_7;
      end else if (8'hb5 == _T_34[7:0]) begin
        image_1_181 <= io_pixelVal_in_1_6;
      end else if (8'hb5 == _T_31[7:0]) begin
        image_1_181 <= io_pixelVal_in_1_5;
      end else if (8'hb5 == _T_28[7:0]) begin
        image_1_181 <= io_pixelVal_in_1_4;
      end else if (8'hb5 == _T_25[7:0]) begin
        image_1_181 <= io_pixelVal_in_1_3;
      end else if (8'hb5 == _T_22[7:0]) begin
        image_1_181 <= io_pixelVal_in_1_2;
      end else if (8'hb5 == _T_19[7:0]) begin
        image_1_181 <= io_pixelVal_in_1_1;
      end else if (8'hb5 == _T_15[7:0]) begin
        image_1_181 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_182 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb6 == _T_37[7:0]) begin
        image_1_182 <= io_pixelVal_in_1_7;
      end else if (8'hb6 == _T_34[7:0]) begin
        image_1_182 <= io_pixelVal_in_1_6;
      end else if (8'hb6 == _T_31[7:0]) begin
        image_1_182 <= io_pixelVal_in_1_5;
      end else if (8'hb6 == _T_28[7:0]) begin
        image_1_182 <= io_pixelVal_in_1_4;
      end else if (8'hb6 == _T_25[7:0]) begin
        image_1_182 <= io_pixelVal_in_1_3;
      end else if (8'hb6 == _T_22[7:0]) begin
        image_1_182 <= io_pixelVal_in_1_2;
      end else if (8'hb6 == _T_19[7:0]) begin
        image_1_182 <= io_pixelVal_in_1_1;
      end else if (8'hb6 == _T_15[7:0]) begin
        image_1_182 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_183 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb7 == _T_37[7:0]) begin
        image_1_183 <= io_pixelVal_in_1_7;
      end else if (8'hb7 == _T_34[7:0]) begin
        image_1_183 <= io_pixelVal_in_1_6;
      end else if (8'hb7 == _T_31[7:0]) begin
        image_1_183 <= io_pixelVal_in_1_5;
      end else if (8'hb7 == _T_28[7:0]) begin
        image_1_183 <= io_pixelVal_in_1_4;
      end else if (8'hb7 == _T_25[7:0]) begin
        image_1_183 <= io_pixelVal_in_1_3;
      end else if (8'hb7 == _T_22[7:0]) begin
        image_1_183 <= io_pixelVal_in_1_2;
      end else if (8'hb7 == _T_19[7:0]) begin
        image_1_183 <= io_pixelVal_in_1_1;
      end else if (8'hb7 == _T_15[7:0]) begin
        image_1_183 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_184 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb8 == _T_37[7:0]) begin
        image_1_184 <= io_pixelVal_in_1_7;
      end else if (8'hb8 == _T_34[7:0]) begin
        image_1_184 <= io_pixelVal_in_1_6;
      end else if (8'hb8 == _T_31[7:0]) begin
        image_1_184 <= io_pixelVal_in_1_5;
      end else if (8'hb8 == _T_28[7:0]) begin
        image_1_184 <= io_pixelVal_in_1_4;
      end else if (8'hb8 == _T_25[7:0]) begin
        image_1_184 <= io_pixelVal_in_1_3;
      end else if (8'hb8 == _T_22[7:0]) begin
        image_1_184 <= io_pixelVal_in_1_2;
      end else if (8'hb8 == _T_19[7:0]) begin
        image_1_184 <= io_pixelVal_in_1_1;
      end else if (8'hb8 == _T_15[7:0]) begin
        image_1_184 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_185 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb9 == _T_37[7:0]) begin
        image_1_185 <= io_pixelVal_in_1_7;
      end else if (8'hb9 == _T_34[7:0]) begin
        image_1_185 <= io_pixelVal_in_1_6;
      end else if (8'hb9 == _T_31[7:0]) begin
        image_1_185 <= io_pixelVal_in_1_5;
      end else if (8'hb9 == _T_28[7:0]) begin
        image_1_185 <= io_pixelVal_in_1_4;
      end else if (8'hb9 == _T_25[7:0]) begin
        image_1_185 <= io_pixelVal_in_1_3;
      end else if (8'hb9 == _T_22[7:0]) begin
        image_1_185 <= io_pixelVal_in_1_2;
      end else if (8'hb9 == _T_19[7:0]) begin
        image_1_185 <= io_pixelVal_in_1_1;
      end else if (8'hb9 == _T_15[7:0]) begin
        image_1_185 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_186 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hba == _T_37[7:0]) begin
        image_1_186 <= io_pixelVal_in_1_7;
      end else if (8'hba == _T_34[7:0]) begin
        image_1_186 <= io_pixelVal_in_1_6;
      end else if (8'hba == _T_31[7:0]) begin
        image_1_186 <= io_pixelVal_in_1_5;
      end else if (8'hba == _T_28[7:0]) begin
        image_1_186 <= io_pixelVal_in_1_4;
      end else if (8'hba == _T_25[7:0]) begin
        image_1_186 <= io_pixelVal_in_1_3;
      end else if (8'hba == _T_22[7:0]) begin
        image_1_186 <= io_pixelVal_in_1_2;
      end else if (8'hba == _T_19[7:0]) begin
        image_1_186 <= io_pixelVal_in_1_1;
      end else if (8'hba == _T_15[7:0]) begin
        image_1_186 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_187 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbb == _T_37[7:0]) begin
        image_1_187 <= io_pixelVal_in_1_7;
      end else if (8'hbb == _T_34[7:0]) begin
        image_1_187 <= io_pixelVal_in_1_6;
      end else if (8'hbb == _T_31[7:0]) begin
        image_1_187 <= io_pixelVal_in_1_5;
      end else if (8'hbb == _T_28[7:0]) begin
        image_1_187 <= io_pixelVal_in_1_4;
      end else if (8'hbb == _T_25[7:0]) begin
        image_1_187 <= io_pixelVal_in_1_3;
      end else if (8'hbb == _T_22[7:0]) begin
        image_1_187 <= io_pixelVal_in_1_2;
      end else if (8'hbb == _T_19[7:0]) begin
        image_1_187 <= io_pixelVal_in_1_1;
      end else if (8'hbb == _T_15[7:0]) begin
        image_1_187 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_188 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbc == _T_37[7:0]) begin
        image_1_188 <= io_pixelVal_in_1_7;
      end else if (8'hbc == _T_34[7:0]) begin
        image_1_188 <= io_pixelVal_in_1_6;
      end else if (8'hbc == _T_31[7:0]) begin
        image_1_188 <= io_pixelVal_in_1_5;
      end else if (8'hbc == _T_28[7:0]) begin
        image_1_188 <= io_pixelVal_in_1_4;
      end else if (8'hbc == _T_25[7:0]) begin
        image_1_188 <= io_pixelVal_in_1_3;
      end else if (8'hbc == _T_22[7:0]) begin
        image_1_188 <= io_pixelVal_in_1_2;
      end else if (8'hbc == _T_19[7:0]) begin
        image_1_188 <= io_pixelVal_in_1_1;
      end else if (8'hbc == _T_15[7:0]) begin
        image_1_188 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_189 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbd == _T_37[7:0]) begin
        image_1_189 <= io_pixelVal_in_1_7;
      end else if (8'hbd == _T_34[7:0]) begin
        image_1_189 <= io_pixelVal_in_1_6;
      end else if (8'hbd == _T_31[7:0]) begin
        image_1_189 <= io_pixelVal_in_1_5;
      end else if (8'hbd == _T_28[7:0]) begin
        image_1_189 <= io_pixelVal_in_1_4;
      end else if (8'hbd == _T_25[7:0]) begin
        image_1_189 <= io_pixelVal_in_1_3;
      end else if (8'hbd == _T_22[7:0]) begin
        image_1_189 <= io_pixelVal_in_1_2;
      end else if (8'hbd == _T_19[7:0]) begin
        image_1_189 <= io_pixelVal_in_1_1;
      end else if (8'hbd == _T_15[7:0]) begin
        image_1_189 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_190 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbe == _T_37[7:0]) begin
        image_1_190 <= io_pixelVal_in_1_7;
      end else if (8'hbe == _T_34[7:0]) begin
        image_1_190 <= io_pixelVal_in_1_6;
      end else if (8'hbe == _T_31[7:0]) begin
        image_1_190 <= io_pixelVal_in_1_5;
      end else if (8'hbe == _T_28[7:0]) begin
        image_1_190 <= io_pixelVal_in_1_4;
      end else if (8'hbe == _T_25[7:0]) begin
        image_1_190 <= io_pixelVal_in_1_3;
      end else if (8'hbe == _T_22[7:0]) begin
        image_1_190 <= io_pixelVal_in_1_2;
      end else if (8'hbe == _T_19[7:0]) begin
        image_1_190 <= io_pixelVal_in_1_1;
      end else if (8'hbe == _T_15[7:0]) begin
        image_1_190 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_191 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbf == _T_37[7:0]) begin
        image_1_191 <= io_pixelVal_in_1_7;
      end else if (8'hbf == _T_34[7:0]) begin
        image_1_191 <= io_pixelVal_in_1_6;
      end else if (8'hbf == _T_31[7:0]) begin
        image_1_191 <= io_pixelVal_in_1_5;
      end else if (8'hbf == _T_28[7:0]) begin
        image_1_191 <= io_pixelVal_in_1_4;
      end else if (8'hbf == _T_25[7:0]) begin
        image_1_191 <= io_pixelVal_in_1_3;
      end else if (8'hbf == _T_22[7:0]) begin
        image_1_191 <= io_pixelVal_in_1_2;
      end else if (8'hbf == _T_19[7:0]) begin
        image_1_191 <= io_pixelVal_in_1_1;
      end else if (8'hbf == _T_15[7:0]) begin
        image_1_191 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_2_0 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h0 == _T_37[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_7;
      end else if (8'h0 == _T_34[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_6;
      end else if (8'h0 == _T_31[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_5;
      end else if (8'h0 == _T_28[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_4;
      end else if (8'h0 == _T_25[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_3;
      end else if (8'h0 == _T_22[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_2;
      end else if (8'h0 == _T_19[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_1;
      end else if (8'h0 == _T_15[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_1 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1 == _T_37[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_7;
      end else if (8'h1 == _T_34[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_6;
      end else if (8'h1 == _T_31[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_5;
      end else if (8'h1 == _T_28[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_4;
      end else if (8'h1 == _T_25[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_3;
      end else if (8'h1 == _T_22[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_2;
      end else if (8'h1 == _T_19[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_1;
      end else if (8'h1 == _T_15[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_2 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2 == _T_37[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_7;
      end else if (8'h2 == _T_34[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_6;
      end else if (8'h2 == _T_31[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_5;
      end else if (8'h2 == _T_28[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_4;
      end else if (8'h2 == _T_25[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_3;
      end else if (8'h2 == _T_22[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_2;
      end else if (8'h2 == _T_19[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_1;
      end else if (8'h2 == _T_15[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_3 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3 == _T_37[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_7;
      end else if (8'h3 == _T_34[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_6;
      end else if (8'h3 == _T_31[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_5;
      end else if (8'h3 == _T_28[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_4;
      end else if (8'h3 == _T_25[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_3;
      end else if (8'h3 == _T_22[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_2;
      end else if (8'h3 == _T_19[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_1;
      end else if (8'h3 == _T_15[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_4 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4 == _T_37[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_7;
      end else if (8'h4 == _T_34[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_6;
      end else if (8'h4 == _T_31[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_5;
      end else if (8'h4 == _T_28[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_4;
      end else if (8'h4 == _T_25[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_3;
      end else if (8'h4 == _T_22[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_2;
      end else if (8'h4 == _T_19[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_1;
      end else if (8'h4 == _T_15[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_5 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5 == _T_37[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_7;
      end else if (8'h5 == _T_34[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_6;
      end else if (8'h5 == _T_31[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_5;
      end else if (8'h5 == _T_28[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_4;
      end else if (8'h5 == _T_25[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_3;
      end else if (8'h5 == _T_22[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_2;
      end else if (8'h5 == _T_19[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_1;
      end else if (8'h5 == _T_15[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_6 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6 == _T_37[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_7;
      end else if (8'h6 == _T_34[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_6;
      end else if (8'h6 == _T_31[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_5;
      end else if (8'h6 == _T_28[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_4;
      end else if (8'h6 == _T_25[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_3;
      end else if (8'h6 == _T_22[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_2;
      end else if (8'h6 == _T_19[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_1;
      end else if (8'h6 == _T_15[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_7 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7 == _T_37[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_7;
      end else if (8'h7 == _T_34[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_6;
      end else if (8'h7 == _T_31[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_5;
      end else if (8'h7 == _T_28[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_4;
      end else if (8'h7 == _T_25[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_3;
      end else if (8'h7 == _T_22[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_2;
      end else if (8'h7 == _T_19[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_1;
      end else if (8'h7 == _T_15[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_8 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8 == _T_37[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_7;
      end else if (8'h8 == _T_34[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_6;
      end else if (8'h8 == _T_31[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_5;
      end else if (8'h8 == _T_28[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_4;
      end else if (8'h8 == _T_25[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_3;
      end else if (8'h8 == _T_22[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_2;
      end else if (8'h8 == _T_19[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_1;
      end else if (8'h8 == _T_15[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_9 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9 == _T_37[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_7;
      end else if (8'h9 == _T_34[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_6;
      end else if (8'h9 == _T_31[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_5;
      end else if (8'h9 == _T_28[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_4;
      end else if (8'h9 == _T_25[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_3;
      end else if (8'h9 == _T_22[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_2;
      end else if (8'h9 == _T_19[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_1;
      end else if (8'h9 == _T_15[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_10 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha == _T_37[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_7;
      end else if (8'ha == _T_34[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_6;
      end else if (8'ha == _T_31[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_5;
      end else if (8'ha == _T_28[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_4;
      end else if (8'ha == _T_25[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_3;
      end else if (8'ha == _T_22[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_2;
      end else if (8'ha == _T_19[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_1;
      end else if (8'ha == _T_15[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_11 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb == _T_37[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_7;
      end else if (8'hb == _T_34[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_6;
      end else if (8'hb == _T_31[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_5;
      end else if (8'hb == _T_28[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_4;
      end else if (8'hb == _T_25[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_3;
      end else if (8'hb == _T_22[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_2;
      end else if (8'hb == _T_19[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_1;
      end else if (8'hb == _T_15[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_12 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc == _T_37[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_7;
      end else if (8'hc == _T_34[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_6;
      end else if (8'hc == _T_31[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_5;
      end else if (8'hc == _T_28[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_4;
      end else if (8'hc == _T_25[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_3;
      end else if (8'hc == _T_22[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_2;
      end else if (8'hc == _T_19[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_1;
      end else if (8'hc == _T_15[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_13 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd == _T_37[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_7;
      end else if (8'hd == _T_34[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_6;
      end else if (8'hd == _T_31[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_5;
      end else if (8'hd == _T_28[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_4;
      end else if (8'hd == _T_25[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_3;
      end else if (8'hd == _T_22[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_2;
      end else if (8'hd == _T_19[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_1;
      end else if (8'hd == _T_15[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_14 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he == _T_37[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_7;
      end else if (8'he == _T_34[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_6;
      end else if (8'he == _T_31[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_5;
      end else if (8'he == _T_28[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_4;
      end else if (8'he == _T_25[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_3;
      end else if (8'he == _T_22[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_2;
      end else if (8'he == _T_19[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_1;
      end else if (8'he == _T_15[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_15 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf == _T_37[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_7;
      end else if (8'hf == _T_34[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_6;
      end else if (8'hf == _T_31[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_5;
      end else if (8'hf == _T_28[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_4;
      end else if (8'hf == _T_25[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_3;
      end else if (8'hf == _T_22[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_2;
      end else if (8'hf == _T_19[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_1;
      end else if (8'hf == _T_15[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_16 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h10 == _T_37[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_7;
      end else if (8'h10 == _T_34[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_6;
      end else if (8'h10 == _T_31[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_5;
      end else if (8'h10 == _T_28[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_4;
      end else if (8'h10 == _T_25[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_3;
      end else if (8'h10 == _T_22[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_2;
      end else if (8'h10 == _T_19[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_1;
      end else if (8'h10 == _T_15[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_17 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h11 == _T_37[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_7;
      end else if (8'h11 == _T_34[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_6;
      end else if (8'h11 == _T_31[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_5;
      end else if (8'h11 == _T_28[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_4;
      end else if (8'h11 == _T_25[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_3;
      end else if (8'h11 == _T_22[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_2;
      end else if (8'h11 == _T_19[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_1;
      end else if (8'h11 == _T_15[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_18 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h12 == _T_37[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_7;
      end else if (8'h12 == _T_34[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_6;
      end else if (8'h12 == _T_31[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_5;
      end else if (8'h12 == _T_28[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_4;
      end else if (8'h12 == _T_25[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_3;
      end else if (8'h12 == _T_22[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_2;
      end else if (8'h12 == _T_19[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_1;
      end else if (8'h12 == _T_15[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_19 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h13 == _T_37[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_7;
      end else if (8'h13 == _T_34[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_6;
      end else if (8'h13 == _T_31[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_5;
      end else if (8'h13 == _T_28[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_4;
      end else if (8'h13 == _T_25[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_3;
      end else if (8'h13 == _T_22[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_2;
      end else if (8'h13 == _T_19[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_1;
      end else if (8'h13 == _T_15[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_20 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h14 == _T_37[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_7;
      end else if (8'h14 == _T_34[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_6;
      end else if (8'h14 == _T_31[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_5;
      end else if (8'h14 == _T_28[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_4;
      end else if (8'h14 == _T_25[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_3;
      end else if (8'h14 == _T_22[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_2;
      end else if (8'h14 == _T_19[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_1;
      end else if (8'h14 == _T_15[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_21 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h15 == _T_37[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_7;
      end else if (8'h15 == _T_34[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_6;
      end else if (8'h15 == _T_31[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_5;
      end else if (8'h15 == _T_28[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_4;
      end else if (8'h15 == _T_25[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_3;
      end else if (8'h15 == _T_22[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_2;
      end else if (8'h15 == _T_19[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_1;
      end else if (8'h15 == _T_15[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_22 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h16 == _T_37[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_7;
      end else if (8'h16 == _T_34[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_6;
      end else if (8'h16 == _T_31[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_5;
      end else if (8'h16 == _T_28[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_4;
      end else if (8'h16 == _T_25[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_3;
      end else if (8'h16 == _T_22[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_2;
      end else if (8'h16 == _T_19[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_1;
      end else if (8'h16 == _T_15[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_23 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h17 == _T_37[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_7;
      end else if (8'h17 == _T_34[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_6;
      end else if (8'h17 == _T_31[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_5;
      end else if (8'h17 == _T_28[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_4;
      end else if (8'h17 == _T_25[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_3;
      end else if (8'h17 == _T_22[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_2;
      end else if (8'h17 == _T_19[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_1;
      end else if (8'h17 == _T_15[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_24 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h18 == _T_37[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_7;
      end else if (8'h18 == _T_34[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_6;
      end else if (8'h18 == _T_31[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_5;
      end else if (8'h18 == _T_28[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_4;
      end else if (8'h18 == _T_25[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_3;
      end else if (8'h18 == _T_22[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_2;
      end else if (8'h18 == _T_19[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_1;
      end else if (8'h18 == _T_15[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_25 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h19 == _T_37[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_7;
      end else if (8'h19 == _T_34[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_6;
      end else if (8'h19 == _T_31[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_5;
      end else if (8'h19 == _T_28[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_4;
      end else if (8'h19 == _T_25[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_3;
      end else if (8'h19 == _T_22[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_2;
      end else if (8'h19 == _T_19[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_1;
      end else if (8'h19 == _T_15[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_26 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1a == _T_37[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_7;
      end else if (8'h1a == _T_34[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_6;
      end else if (8'h1a == _T_31[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_5;
      end else if (8'h1a == _T_28[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_4;
      end else if (8'h1a == _T_25[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_3;
      end else if (8'h1a == _T_22[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_2;
      end else if (8'h1a == _T_19[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_1;
      end else if (8'h1a == _T_15[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_27 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1b == _T_37[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_7;
      end else if (8'h1b == _T_34[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_6;
      end else if (8'h1b == _T_31[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_5;
      end else if (8'h1b == _T_28[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_4;
      end else if (8'h1b == _T_25[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_3;
      end else if (8'h1b == _T_22[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_2;
      end else if (8'h1b == _T_19[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_1;
      end else if (8'h1b == _T_15[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_28 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1c == _T_37[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_7;
      end else if (8'h1c == _T_34[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_6;
      end else if (8'h1c == _T_31[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_5;
      end else if (8'h1c == _T_28[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_4;
      end else if (8'h1c == _T_25[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_3;
      end else if (8'h1c == _T_22[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_2;
      end else if (8'h1c == _T_19[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_1;
      end else if (8'h1c == _T_15[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_29 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1d == _T_37[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_7;
      end else if (8'h1d == _T_34[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_6;
      end else if (8'h1d == _T_31[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_5;
      end else if (8'h1d == _T_28[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_4;
      end else if (8'h1d == _T_25[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_3;
      end else if (8'h1d == _T_22[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_2;
      end else if (8'h1d == _T_19[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_1;
      end else if (8'h1d == _T_15[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_30 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1e == _T_37[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_7;
      end else if (8'h1e == _T_34[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_6;
      end else if (8'h1e == _T_31[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_5;
      end else if (8'h1e == _T_28[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_4;
      end else if (8'h1e == _T_25[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_3;
      end else if (8'h1e == _T_22[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_2;
      end else if (8'h1e == _T_19[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_1;
      end else if (8'h1e == _T_15[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_31 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1f == _T_37[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_7;
      end else if (8'h1f == _T_34[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_6;
      end else if (8'h1f == _T_31[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_5;
      end else if (8'h1f == _T_28[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_4;
      end else if (8'h1f == _T_25[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_3;
      end else if (8'h1f == _T_22[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_2;
      end else if (8'h1f == _T_19[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_1;
      end else if (8'h1f == _T_15[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_32 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h20 == _T_37[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_7;
      end else if (8'h20 == _T_34[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_6;
      end else if (8'h20 == _T_31[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_5;
      end else if (8'h20 == _T_28[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_4;
      end else if (8'h20 == _T_25[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_3;
      end else if (8'h20 == _T_22[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_2;
      end else if (8'h20 == _T_19[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_1;
      end else if (8'h20 == _T_15[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_33 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h21 == _T_37[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_7;
      end else if (8'h21 == _T_34[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_6;
      end else if (8'h21 == _T_31[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_5;
      end else if (8'h21 == _T_28[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_4;
      end else if (8'h21 == _T_25[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_3;
      end else if (8'h21 == _T_22[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_2;
      end else if (8'h21 == _T_19[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_1;
      end else if (8'h21 == _T_15[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_34 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h22 == _T_37[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_7;
      end else if (8'h22 == _T_34[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_6;
      end else if (8'h22 == _T_31[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_5;
      end else if (8'h22 == _T_28[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_4;
      end else if (8'h22 == _T_25[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_3;
      end else if (8'h22 == _T_22[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_2;
      end else if (8'h22 == _T_19[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_1;
      end else if (8'h22 == _T_15[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_35 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h23 == _T_37[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_7;
      end else if (8'h23 == _T_34[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_6;
      end else if (8'h23 == _T_31[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_5;
      end else if (8'h23 == _T_28[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_4;
      end else if (8'h23 == _T_25[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_3;
      end else if (8'h23 == _T_22[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_2;
      end else if (8'h23 == _T_19[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_1;
      end else if (8'h23 == _T_15[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_36 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h24 == _T_37[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_7;
      end else if (8'h24 == _T_34[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_6;
      end else if (8'h24 == _T_31[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_5;
      end else if (8'h24 == _T_28[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_4;
      end else if (8'h24 == _T_25[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_3;
      end else if (8'h24 == _T_22[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_2;
      end else if (8'h24 == _T_19[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_1;
      end else if (8'h24 == _T_15[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_37 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h25 == _T_37[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_7;
      end else if (8'h25 == _T_34[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_6;
      end else if (8'h25 == _T_31[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_5;
      end else if (8'h25 == _T_28[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_4;
      end else if (8'h25 == _T_25[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_3;
      end else if (8'h25 == _T_22[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_2;
      end else if (8'h25 == _T_19[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_1;
      end else if (8'h25 == _T_15[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_38 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h26 == _T_37[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_7;
      end else if (8'h26 == _T_34[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_6;
      end else if (8'h26 == _T_31[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_5;
      end else if (8'h26 == _T_28[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_4;
      end else if (8'h26 == _T_25[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_3;
      end else if (8'h26 == _T_22[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_2;
      end else if (8'h26 == _T_19[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_1;
      end else if (8'h26 == _T_15[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_39 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h27 == _T_37[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_7;
      end else if (8'h27 == _T_34[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_6;
      end else if (8'h27 == _T_31[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_5;
      end else if (8'h27 == _T_28[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_4;
      end else if (8'h27 == _T_25[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_3;
      end else if (8'h27 == _T_22[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_2;
      end else if (8'h27 == _T_19[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_1;
      end else if (8'h27 == _T_15[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_40 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h28 == _T_37[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_7;
      end else if (8'h28 == _T_34[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_6;
      end else if (8'h28 == _T_31[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_5;
      end else if (8'h28 == _T_28[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_4;
      end else if (8'h28 == _T_25[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_3;
      end else if (8'h28 == _T_22[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_2;
      end else if (8'h28 == _T_19[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_1;
      end else if (8'h28 == _T_15[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_41 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h29 == _T_37[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_7;
      end else if (8'h29 == _T_34[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_6;
      end else if (8'h29 == _T_31[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_5;
      end else if (8'h29 == _T_28[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_4;
      end else if (8'h29 == _T_25[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_3;
      end else if (8'h29 == _T_22[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_2;
      end else if (8'h29 == _T_19[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_1;
      end else if (8'h29 == _T_15[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_42 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2a == _T_37[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_7;
      end else if (8'h2a == _T_34[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_6;
      end else if (8'h2a == _T_31[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_5;
      end else if (8'h2a == _T_28[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_4;
      end else if (8'h2a == _T_25[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_3;
      end else if (8'h2a == _T_22[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_2;
      end else if (8'h2a == _T_19[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_1;
      end else if (8'h2a == _T_15[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_43 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2b == _T_37[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_7;
      end else if (8'h2b == _T_34[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_6;
      end else if (8'h2b == _T_31[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_5;
      end else if (8'h2b == _T_28[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_4;
      end else if (8'h2b == _T_25[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_3;
      end else if (8'h2b == _T_22[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_2;
      end else if (8'h2b == _T_19[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_1;
      end else if (8'h2b == _T_15[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_44 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2c == _T_37[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_7;
      end else if (8'h2c == _T_34[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_6;
      end else if (8'h2c == _T_31[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_5;
      end else if (8'h2c == _T_28[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_4;
      end else if (8'h2c == _T_25[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_3;
      end else if (8'h2c == _T_22[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_2;
      end else if (8'h2c == _T_19[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_1;
      end else if (8'h2c == _T_15[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_45 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2d == _T_37[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_7;
      end else if (8'h2d == _T_34[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_6;
      end else if (8'h2d == _T_31[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_5;
      end else if (8'h2d == _T_28[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_4;
      end else if (8'h2d == _T_25[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_3;
      end else if (8'h2d == _T_22[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_2;
      end else if (8'h2d == _T_19[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_1;
      end else if (8'h2d == _T_15[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_46 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2e == _T_37[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_7;
      end else if (8'h2e == _T_34[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_6;
      end else if (8'h2e == _T_31[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_5;
      end else if (8'h2e == _T_28[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_4;
      end else if (8'h2e == _T_25[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_3;
      end else if (8'h2e == _T_22[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_2;
      end else if (8'h2e == _T_19[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_1;
      end else if (8'h2e == _T_15[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_47 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2f == _T_37[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_7;
      end else if (8'h2f == _T_34[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_6;
      end else if (8'h2f == _T_31[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_5;
      end else if (8'h2f == _T_28[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_4;
      end else if (8'h2f == _T_25[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_3;
      end else if (8'h2f == _T_22[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_2;
      end else if (8'h2f == _T_19[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_1;
      end else if (8'h2f == _T_15[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_48 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h30 == _T_37[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_7;
      end else if (8'h30 == _T_34[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_6;
      end else if (8'h30 == _T_31[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_5;
      end else if (8'h30 == _T_28[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_4;
      end else if (8'h30 == _T_25[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_3;
      end else if (8'h30 == _T_22[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_2;
      end else if (8'h30 == _T_19[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_1;
      end else if (8'h30 == _T_15[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_49 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h31 == _T_37[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_7;
      end else if (8'h31 == _T_34[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_6;
      end else if (8'h31 == _T_31[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_5;
      end else if (8'h31 == _T_28[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_4;
      end else if (8'h31 == _T_25[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_3;
      end else if (8'h31 == _T_22[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_2;
      end else if (8'h31 == _T_19[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_1;
      end else if (8'h31 == _T_15[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_50 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h32 == _T_37[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_7;
      end else if (8'h32 == _T_34[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_6;
      end else if (8'h32 == _T_31[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_5;
      end else if (8'h32 == _T_28[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_4;
      end else if (8'h32 == _T_25[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_3;
      end else if (8'h32 == _T_22[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_2;
      end else if (8'h32 == _T_19[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_1;
      end else if (8'h32 == _T_15[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_51 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h33 == _T_37[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_7;
      end else if (8'h33 == _T_34[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_6;
      end else if (8'h33 == _T_31[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_5;
      end else if (8'h33 == _T_28[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_4;
      end else if (8'h33 == _T_25[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_3;
      end else if (8'h33 == _T_22[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_2;
      end else if (8'h33 == _T_19[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_1;
      end else if (8'h33 == _T_15[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_52 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h34 == _T_37[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_7;
      end else if (8'h34 == _T_34[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_6;
      end else if (8'h34 == _T_31[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_5;
      end else if (8'h34 == _T_28[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_4;
      end else if (8'h34 == _T_25[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_3;
      end else if (8'h34 == _T_22[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_2;
      end else if (8'h34 == _T_19[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_1;
      end else if (8'h34 == _T_15[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_53 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h35 == _T_37[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_7;
      end else if (8'h35 == _T_34[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_6;
      end else if (8'h35 == _T_31[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_5;
      end else if (8'h35 == _T_28[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_4;
      end else if (8'h35 == _T_25[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_3;
      end else if (8'h35 == _T_22[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_2;
      end else if (8'h35 == _T_19[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_1;
      end else if (8'h35 == _T_15[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_54 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h36 == _T_37[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_7;
      end else if (8'h36 == _T_34[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_6;
      end else if (8'h36 == _T_31[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_5;
      end else if (8'h36 == _T_28[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_4;
      end else if (8'h36 == _T_25[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_3;
      end else if (8'h36 == _T_22[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_2;
      end else if (8'h36 == _T_19[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_1;
      end else if (8'h36 == _T_15[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_55 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h37 == _T_37[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_7;
      end else if (8'h37 == _T_34[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_6;
      end else if (8'h37 == _T_31[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_5;
      end else if (8'h37 == _T_28[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_4;
      end else if (8'h37 == _T_25[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_3;
      end else if (8'h37 == _T_22[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_2;
      end else if (8'h37 == _T_19[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_1;
      end else if (8'h37 == _T_15[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_56 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h38 == _T_37[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_7;
      end else if (8'h38 == _T_34[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_6;
      end else if (8'h38 == _T_31[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_5;
      end else if (8'h38 == _T_28[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_4;
      end else if (8'h38 == _T_25[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_3;
      end else if (8'h38 == _T_22[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_2;
      end else if (8'h38 == _T_19[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_1;
      end else if (8'h38 == _T_15[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_57 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h39 == _T_37[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_7;
      end else if (8'h39 == _T_34[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_6;
      end else if (8'h39 == _T_31[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_5;
      end else if (8'h39 == _T_28[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_4;
      end else if (8'h39 == _T_25[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_3;
      end else if (8'h39 == _T_22[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_2;
      end else if (8'h39 == _T_19[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_1;
      end else if (8'h39 == _T_15[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_58 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3a == _T_37[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_7;
      end else if (8'h3a == _T_34[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_6;
      end else if (8'h3a == _T_31[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_5;
      end else if (8'h3a == _T_28[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_4;
      end else if (8'h3a == _T_25[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_3;
      end else if (8'h3a == _T_22[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_2;
      end else if (8'h3a == _T_19[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_1;
      end else if (8'h3a == _T_15[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_59 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3b == _T_37[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_7;
      end else if (8'h3b == _T_34[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_6;
      end else if (8'h3b == _T_31[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_5;
      end else if (8'h3b == _T_28[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_4;
      end else if (8'h3b == _T_25[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_3;
      end else if (8'h3b == _T_22[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_2;
      end else if (8'h3b == _T_19[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_1;
      end else if (8'h3b == _T_15[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_60 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3c == _T_37[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_7;
      end else if (8'h3c == _T_34[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_6;
      end else if (8'h3c == _T_31[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_5;
      end else if (8'h3c == _T_28[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_4;
      end else if (8'h3c == _T_25[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_3;
      end else if (8'h3c == _T_22[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_2;
      end else if (8'h3c == _T_19[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_1;
      end else if (8'h3c == _T_15[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_61 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3d == _T_37[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_7;
      end else if (8'h3d == _T_34[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_6;
      end else if (8'h3d == _T_31[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_5;
      end else if (8'h3d == _T_28[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_4;
      end else if (8'h3d == _T_25[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_3;
      end else if (8'h3d == _T_22[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_2;
      end else if (8'h3d == _T_19[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_1;
      end else if (8'h3d == _T_15[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_62 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3e == _T_37[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_7;
      end else if (8'h3e == _T_34[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_6;
      end else if (8'h3e == _T_31[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_5;
      end else if (8'h3e == _T_28[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_4;
      end else if (8'h3e == _T_25[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_3;
      end else if (8'h3e == _T_22[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_2;
      end else if (8'h3e == _T_19[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_1;
      end else if (8'h3e == _T_15[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_63 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3f == _T_37[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_7;
      end else if (8'h3f == _T_34[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_6;
      end else if (8'h3f == _T_31[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_5;
      end else if (8'h3f == _T_28[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_4;
      end else if (8'h3f == _T_25[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_3;
      end else if (8'h3f == _T_22[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_2;
      end else if (8'h3f == _T_19[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_1;
      end else if (8'h3f == _T_15[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_64 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h40 == _T_37[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_7;
      end else if (8'h40 == _T_34[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_6;
      end else if (8'h40 == _T_31[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_5;
      end else if (8'h40 == _T_28[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_4;
      end else if (8'h40 == _T_25[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_3;
      end else if (8'h40 == _T_22[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_2;
      end else if (8'h40 == _T_19[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_1;
      end else if (8'h40 == _T_15[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_65 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h41 == _T_37[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_7;
      end else if (8'h41 == _T_34[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_6;
      end else if (8'h41 == _T_31[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_5;
      end else if (8'h41 == _T_28[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_4;
      end else if (8'h41 == _T_25[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_3;
      end else if (8'h41 == _T_22[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_2;
      end else if (8'h41 == _T_19[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_1;
      end else if (8'h41 == _T_15[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_66 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h42 == _T_37[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_7;
      end else if (8'h42 == _T_34[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_6;
      end else if (8'h42 == _T_31[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_5;
      end else if (8'h42 == _T_28[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_4;
      end else if (8'h42 == _T_25[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_3;
      end else if (8'h42 == _T_22[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_2;
      end else if (8'h42 == _T_19[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_1;
      end else if (8'h42 == _T_15[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_67 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h43 == _T_37[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_7;
      end else if (8'h43 == _T_34[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_6;
      end else if (8'h43 == _T_31[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_5;
      end else if (8'h43 == _T_28[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_4;
      end else if (8'h43 == _T_25[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_3;
      end else if (8'h43 == _T_22[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_2;
      end else if (8'h43 == _T_19[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_1;
      end else if (8'h43 == _T_15[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_68 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h44 == _T_37[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_7;
      end else if (8'h44 == _T_34[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_6;
      end else if (8'h44 == _T_31[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_5;
      end else if (8'h44 == _T_28[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_4;
      end else if (8'h44 == _T_25[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_3;
      end else if (8'h44 == _T_22[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_2;
      end else if (8'h44 == _T_19[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_1;
      end else if (8'h44 == _T_15[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_69 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h45 == _T_37[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_7;
      end else if (8'h45 == _T_34[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_6;
      end else if (8'h45 == _T_31[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_5;
      end else if (8'h45 == _T_28[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_4;
      end else if (8'h45 == _T_25[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_3;
      end else if (8'h45 == _T_22[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_2;
      end else if (8'h45 == _T_19[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_1;
      end else if (8'h45 == _T_15[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_70 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h46 == _T_37[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_7;
      end else if (8'h46 == _T_34[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_6;
      end else if (8'h46 == _T_31[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_5;
      end else if (8'h46 == _T_28[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_4;
      end else if (8'h46 == _T_25[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_3;
      end else if (8'h46 == _T_22[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_2;
      end else if (8'h46 == _T_19[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_1;
      end else if (8'h46 == _T_15[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_71 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h47 == _T_37[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_7;
      end else if (8'h47 == _T_34[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_6;
      end else if (8'h47 == _T_31[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_5;
      end else if (8'h47 == _T_28[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_4;
      end else if (8'h47 == _T_25[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_3;
      end else if (8'h47 == _T_22[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_2;
      end else if (8'h47 == _T_19[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_1;
      end else if (8'h47 == _T_15[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_72 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h48 == _T_37[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_7;
      end else if (8'h48 == _T_34[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_6;
      end else if (8'h48 == _T_31[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_5;
      end else if (8'h48 == _T_28[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_4;
      end else if (8'h48 == _T_25[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_3;
      end else if (8'h48 == _T_22[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_2;
      end else if (8'h48 == _T_19[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_1;
      end else if (8'h48 == _T_15[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_73 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h49 == _T_37[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_7;
      end else if (8'h49 == _T_34[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_6;
      end else if (8'h49 == _T_31[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_5;
      end else if (8'h49 == _T_28[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_4;
      end else if (8'h49 == _T_25[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_3;
      end else if (8'h49 == _T_22[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_2;
      end else if (8'h49 == _T_19[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_1;
      end else if (8'h49 == _T_15[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_74 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4a == _T_37[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_7;
      end else if (8'h4a == _T_34[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_6;
      end else if (8'h4a == _T_31[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_5;
      end else if (8'h4a == _T_28[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_4;
      end else if (8'h4a == _T_25[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_3;
      end else if (8'h4a == _T_22[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_2;
      end else if (8'h4a == _T_19[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_1;
      end else if (8'h4a == _T_15[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_75 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4b == _T_37[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_7;
      end else if (8'h4b == _T_34[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_6;
      end else if (8'h4b == _T_31[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_5;
      end else if (8'h4b == _T_28[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_4;
      end else if (8'h4b == _T_25[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_3;
      end else if (8'h4b == _T_22[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_2;
      end else if (8'h4b == _T_19[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_1;
      end else if (8'h4b == _T_15[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_76 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4c == _T_37[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_7;
      end else if (8'h4c == _T_34[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_6;
      end else if (8'h4c == _T_31[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_5;
      end else if (8'h4c == _T_28[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_4;
      end else if (8'h4c == _T_25[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_3;
      end else if (8'h4c == _T_22[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_2;
      end else if (8'h4c == _T_19[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_1;
      end else if (8'h4c == _T_15[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_77 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4d == _T_37[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_7;
      end else if (8'h4d == _T_34[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_6;
      end else if (8'h4d == _T_31[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_5;
      end else if (8'h4d == _T_28[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_4;
      end else if (8'h4d == _T_25[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_3;
      end else if (8'h4d == _T_22[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_2;
      end else if (8'h4d == _T_19[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_1;
      end else if (8'h4d == _T_15[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_78 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4e == _T_37[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_7;
      end else if (8'h4e == _T_34[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_6;
      end else if (8'h4e == _T_31[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_5;
      end else if (8'h4e == _T_28[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_4;
      end else if (8'h4e == _T_25[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_3;
      end else if (8'h4e == _T_22[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_2;
      end else if (8'h4e == _T_19[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_1;
      end else if (8'h4e == _T_15[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_79 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4f == _T_37[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_7;
      end else if (8'h4f == _T_34[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_6;
      end else if (8'h4f == _T_31[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_5;
      end else if (8'h4f == _T_28[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_4;
      end else if (8'h4f == _T_25[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_3;
      end else if (8'h4f == _T_22[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_2;
      end else if (8'h4f == _T_19[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_1;
      end else if (8'h4f == _T_15[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_80 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h50 == _T_37[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_7;
      end else if (8'h50 == _T_34[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_6;
      end else if (8'h50 == _T_31[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_5;
      end else if (8'h50 == _T_28[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_4;
      end else if (8'h50 == _T_25[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_3;
      end else if (8'h50 == _T_22[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_2;
      end else if (8'h50 == _T_19[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_1;
      end else if (8'h50 == _T_15[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_81 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h51 == _T_37[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_7;
      end else if (8'h51 == _T_34[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_6;
      end else if (8'h51 == _T_31[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_5;
      end else if (8'h51 == _T_28[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_4;
      end else if (8'h51 == _T_25[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_3;
      end else if (8'h51 == _T_22[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_2;
      end else if (8'h51 == _T_19[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_1;
      end else if (8'h51 == _T_15[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_82 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h52 == _T_37[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_7;
      end else if (8'h52 == _T_34[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_6;
      end else if (8'h52 == _T_31[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_5;
      end else if (8'h52 == _T_28[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_4;
      end else if (8'h52 == _T_25[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_3;
      end else if (8'h52 == _T_22[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_2;
      end else if (8'h52 == _T_19[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_1;
      end else if (8'h52 == _T_15[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_83 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h53 == _T_37[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_7;
      end else if (8'h53 == _T_34[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_6;
      end else if (8'h53 == _T_31[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_5;
      end else if (8'h53 == _T_28[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_4;
      end else if (8'h53 == _T_25[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_3;
      end else if (8'h53 == _T_22[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_2;
      end else if (8'h53 == _T_19[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_1;
      end else if (8'h53 == _T_15[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_84 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h54 == _T_37[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_7;
      end else if (8'h54 == _T_34[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_6;
      end else if (8'h54 == _T_31[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_5;
      end else if (8'h54 == _T_28[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_4;
      end else if (8'h54 == _T_25[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_3;
      end else if (8'h54 == _T_22[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_2;
      end else if (8'h54 == _T_19[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_1;
      end else if (8'h54 == _T_15[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_85 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h55 == _T_37[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_7;
      end else if (8'h55 == _T_34[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_6;
      end else if (8'h55 == _T_31[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_5;
      end else if (8'h55 == _T_28[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_4;
      end else if (8'h55 == _T_25[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_3;
      end else if (8'h55 == _T_22[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_2;
      end else if (8'h55 == _T_19[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_1;
      end else if (8'h55 == _T_15[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_86 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h56 == _T_37[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_7;
      end else if (8'h56 == _T_34[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_6;
      end else if (8'h56 == _T_31[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_5;
      end else if (8'h56 == _T_28[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_4;
      end else if (8'h56 == _T_25[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_3;
      end else if (8'h56 == _T_22[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_2;
      end else if (8'h56 == _T_19[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_1;
      end else if (8'h56 == _T_15[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_87 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h57 == _T_37[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_7;
      end else if (8'h57 == _T_34[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_6;
      end else if (8'h57 == _T_31[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_5;
      end else if (8'h57 == _T_28[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_4;
      end else if (8'h57 == _T_25[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_3;
      end else if (8'h57 == _T_22[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_2;
      end else if (8'h57 == _T_19[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_1;
      end else if (8'h57 == _T_15[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_88 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h58 == _T_37[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_7;
      end else if (8'h58 == _T_34[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_6;
      end else if (8'h58 == _T_31[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_5;
      end else if (8'h58 == _T_28[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_4;
      end else if (8'h58 == _T_25[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_3;
      end else if (8'h58 == _T_22[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_2;
      end else if (8'h58 == _T_19[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_1;
      end else if (8'h58 == _T_15[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_89 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h59 == _T_37[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_7;
      end else if (8'h59 == _T_34[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_6;
      end else if (8'h59 == _T_31[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_5;
      end else if (8'h59 == _T_28[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_4;
      end else if (8'h59 == _T_25[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_3;
      end else if (8'h59 == _T_22[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_2;
      end else if (8'h59 == _T_19[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_1;
      end else if (8'h59 == _T_15[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_90 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5a == _T_37[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_7;
      end else if (8'h5a == _T_34[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_6;
      end else if (8'h5a == _T_31[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_5;
      end else if (8'h5a == _T_28[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_4;
      end else if (8'h5a == _T_25[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_3;
      end else if (8'h5a == _T_22[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_2;
      end else if (8'h5a == _T_19[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_1;
      end else if (8'h5a == _T_15[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_91 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5b == _T_37[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_7;
      end else if (8'h5b == _T_34[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_6;
      end else if (8'h5b == _T_31[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_5;
      end else if (8'h5b == _T_28[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_4;
      end else if (8'h5b == _T_25[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_3;
      end else if (8'h5b == _T_22[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_2;
      end else if (8'h5b == _T_19[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_1;
      end else if (8'h5b == _T_15[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_92 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5c == _T_37[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_7;
      end else if (8'h5c == _T_34[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_6;
      end else if (8'h5c == _T_31[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_5;
      end else if (8'h5c == _T_28[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_4;
      end else if (8'h5c == _T_25[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_3;
      end else if (8'h5c == _T_22[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_2;
      end else if (8'h5c == _T_19[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_1;
      end else if (8'h5c == _T_15[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_93 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5d == _T_37[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_7;
      end else if (8'h5d == _T_34[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_6;
      end else if (8'h5d == _T_31[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_5;
      end else if (8'h5d == _T_28[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_4;
      end else if (8'h5d == _T_25[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_3;
      end else if (8'h5d == _T_22[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_2;
      end else if (8'h5d == _T_19[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_1;
      end else if (8'h5d == _T_15[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_94 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5e == _T_37[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_7;
      end else if (8'h5e == _T_34[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_6;
      end else if (8'h5e == _T_31[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_5;
      end else if (8'h5e == _T_28[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_4;
      end else if (8'h5e == _T_25[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_3;
      end else if (8'h5e == _T_22[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_2;
      end else if (8'h5e == _T_19[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_1;
      end else if (8'h5e == _T_15[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_95 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5f == _T_37[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_7;
      end else if (8'h5f == _T_34[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_6;
      end else if (8'h5f == _T_31[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_5;
      end else if (8'h5f == _T_28[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_4;
      end else if (8'h5f == _T_25[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_3;
      end else if (8'h5f == _T_22[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_2;
      end else if (8'h5f == _T_19[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_1;
      end else if (8'h5f == _T_15[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_96 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h60 == _T_37[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_7;
      end else if (8'h60 == _T_34[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_6;
      end else if (8'h60 == _T_31[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_5;
      end else if (8'h60 == _T_28[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_4;
      end else if (8'h60 == _T_25[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_3;
      end else if (8'h60 == _T_22[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_2;
      end else if (8'h60 == _T_19[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_1;
      end else if (8'h60 == _T_15[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_97 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h61 == _T_37[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_7;
      end else if (8'h61 == _T_34[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_6;
      end else if (8'h61 == _T_31[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_5;
      end else if (8'h61 == _T_28[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_4;
      end else if (8'h61 == _T_25[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_3;
      end else if (8'h61 == _T_22[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_2;
      end else if (8'h61 == _T_19[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_1;
      end else if (8'h61 == _T_15[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_98 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h62 == _T_37[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_7;
      end else if (8'h62 == _T_34[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_6;
      end else if (8'h62 == _T_31[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_5;
      end else if (8'h62 == _T_28[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_4;
      end else if (8'h62 == _T_25[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_3;
      end else if (8'h62 == _T_22[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_2;
      end else if (8'h62 == _T_19[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_1;
      end else if (8'h62 == _T_15[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_99 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h63 == _T_37[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_7;
      end else if (8'h63 == _T_34[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_6;
      end else if (8'h63 == _T_31[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_5;
      end else if (8'h63 == _T_28[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_4;
      end else if (8'h63 == _T_25[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_3;
      end else if (8'h63 == _T_22[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_2;
      end else if (8'h63 == _T_19[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_1;
      end else if (8'h63 == _T_15[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_100 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h64 == _T_37[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_7;
      end else if (8'h64 == _T_34[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_6;
      end else if (8'h64 == _T_31[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_5;
      end else if (8'h64 == _T_28[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_4;
      end else if (8'h64 == _T_25[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_3;
      end else if (8'h64 == _T_22[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_2;
      end else if (8'h64 == _T_19[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_1;
      end else if (8'h64 == _T_15[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_101 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h65 == _T_37[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_7;
      end else if (8'h65 == _T_34[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_6;
      end else if (8'h65 == _T_31[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_5;
      end else if (8'h65 == _T_28[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_4;
      end else if (8'h65 == _T_25[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_3;
      end else if (8'h65 == _T_22[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_2;
      end else if (8'h65 == _T_19[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_1;
      end else if (8'h65 == _T_15[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_102 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h66 == _T_37[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_7;
      end else if (8'h66 == _T_34[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_6;
      end else if (8'h66 == _T_31[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_5;
      end else if (8'h66 == _T_28[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_4;
      end else if (8'h66 == _T_25[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_3;
      end else if (8'h66 == _T_22[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_2;
      end else if (8'h66 == _T_19[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_1;
      end else if (8'h66 == _T_15[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_103 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h67 == _T_37[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_7;
      end else if (8'h67 == _T_34[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_6;
      end else if (8'h67 == _T_31[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_5;
      end else if (8'h67 == _T_28[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_4;
      end else if (8'h67 == _T_25[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_3;
      end else if (8'h67 == _T_22[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_2;
      end else if (8'h67 == _T_19[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_1;
      end else if (8'h67 == _T_15[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_104 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h68 == _T_37[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_7;
      end else if (8'h68 == _T_34[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_6;
      end else if (8'h68 == _T_31[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_5;
      end else if (8'h68 == _T_28[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_4;
      end else if (8'h68 == _T_25[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_3;
      end else if (8'h68 == _T_22[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_2;
      end else if (8'h68 == _T_19[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_1;
      end else if (8'h68 == _T_15[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_105 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h69 == _T_37[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_7;
      end else if (8'h69 == _T_34[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_6;
      end else if (8'h69 == _T_31[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_5;
      end else if (8'h69 == _T_28[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_4;
      end else if (8'h69 == _T_25[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_3;
      end else if (8'h69 == _T_22[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_2;
      end else if (8'h69 == _T_19[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_1;
      end else if (8'h69 == _T_15[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_106 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6a == _T_37[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_7;
      end else if (8'h6a == _T_34[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_6;
      end else if (8'h6a == _T_31[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_5;
      end else if (8'h6a == _T_28[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_4;
      end else if (8'h6a == _T_25[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_3;
      end else if (8'h6a == _T_22[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_2;
      end else if (8'h6a == _T_19[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_1;
      end else if (8'h6a == _T_15[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_107 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6b == _T_37[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_7;
      end else if (8'h6b == _T_34[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_6;
      end else if (8'h6b == _T_31[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_5;
      end else if (8'h6b == _T_28[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_4;
      end else if (8'h6b == _T_25[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_3;
      end else if (8'h6b == _T_22[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_2;
      end else if (8'h6b == _T_19[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_1;
      end else if (8'h6b == _T_15[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_108 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6c == _T_37[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_7;
      end else if (8'h6c == _T_34[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_6;
      end else if (8'h6c == _T_31[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_5;
      end else if (8'h6c == _T_28[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_4;
      end else if (8'h6c == _T_25[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_3;
      end else if (8'h6c == _T_22[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_2;
      end else if (8'h6c == _T_19[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_1;
      end else if (8'h6c == _T_15[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_109 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6d == _T_37[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_7;
      end else if (8'h6d == _T_34[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_6;
      end else if (8'h6d == _T_31[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_5;
      end else if (8'h6d == _T_28[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_4;
      end else if (8'h6d == _T_25[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_3;
      end else if (8'h6d == _T_22[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_2;
      end else if (8'h6d == _T_19[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_1;
      end else if (8'h6d == _T_15[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_110 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6e == _T_37[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_7;
      end else if (8'h6e == _T_34[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_6;
      end else if (8'h6e == _T_31[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_5;
      end else if (8'h6e == _T_28[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_4;
      end else if (8'h6e == _T_25[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_3;
      end else if (8'h6e == _T_22[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_2;
      end else if (8'h6e == _T_19[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_1;
      end else if (8'h6e == _T_15[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_111 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6f == _T_37[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_7;
      end else if (8'h6f == _T_34[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_6;
      end else if (8'h6f == _T_31[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_5;
      end else if (8'h6f == _T_28[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_4;
      end else if (8'h6f == _T_25[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_3;
      end else if (8'h6f == _T_22[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_2;
      end else if (8'h6f == _T_19[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_1;
      end else if (8'h6f == _T_15[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_112 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h70 == _T_37[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_7;
      end else if (8'h70 == _T_34[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_6;
      end else if (8'h70 == _T_31[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_5;
      end else if (8'h70 == _T_28[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_4;
      end else if (8'h70 == _T_25[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_3;
      end else if (8'h70 == _T_22[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_2;
      end else if (8'h70 == _T_19[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_1;
      end else if (8'h70 == _T_15[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_113 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h71 == _T_37[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_7;
      end else if (8'h71 == _T_34[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_6;
      end else if (8'h71 == _T_31[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_5;
      end else if (8'h71 == _T_28[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_4;
      end else if (8'h71 == _T_25[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_3;
      end else if (8'h71 == _T_22[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_2;
      end else if (8'h71 == _T_19[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_1;
      end else if (8'h71 == _T_15[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_114 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h72 == _T_37[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_7;
      end else if (8'h72 == _T_34[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_6;
      end else if (8'h72 == _T_31[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_5;
      end else if (8'h72 == _T_28[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_4;
      end else if (8'h72 == _T_25[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_3;
      end else if (8'h72 == _T_22[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_2;
      end else if (8'h72 == _T_19[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_1;
      end else if (8'h72 == _T_15[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_115 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h73 == _T_37[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_7;
      end else if (8'h73 == _T_34[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_6;
      end else if (8'h73 == _T_31[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_5;
      end else if (8'h73 == _T_28[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_4;
      end else if (8'h73 == _T_25[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_3;
      end else if (8'h73 == _T_22[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_2;
      end else if (8'h73 == _T_19[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_1;
      end else if (8'h73 == _T_15[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_116 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h74 == _T_37[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_7;
      end else if (8'h74 == _T_34[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_6;
      end else if (8'h74 == _T_31[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_5;
      end else if (8'h74 == _T_28[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_4;
      end else if (8'h74 == _T_25[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_3;
      end else if (8'h74 == _T_22[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_2;
      end else if (8'h74 == _T_19[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_1;
      end else if (8'h74 == _T_15[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_117 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h75 == _T_37[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_7;
      end else if (8'h75 == _T_34[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_6;
      end else if (8'h75 == _T_31[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_5;
      end else if (8'h75 == _T_28[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_4;
      end else if (8'h75 == _T_25[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_3;
      end else if (8'h75 == _T_22[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_2;
      end else if (8'h75 == _T_19[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_1;
      end else if (8'h75 == _T_15[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_118 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h76 == _T_37[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_7;
      end else if (8'h76 == _T_34[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_6;
      end else if (8'h76 == _T_31[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_5;
      end else if (8'h76 == _T_28[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_4;
      end else if (8'h76 == _T_25[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_3;
      end else if (8'h76 == _T_22[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_2;
      end else if (8'h76 == _T_19[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_1;
      end else if (8'h76 == _T_15[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_119 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h77 == _T_37[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_7;
      end else if (8'h77 == _T_34[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_6;
      end else if (8'h77 == _T_31[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_5;
      end else if (8'h77 == _T_28[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_4;
      end else if (8'h77 == _T_25[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_3;
      end else if (8'h77 == _T_22[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_2;
      end else if (8'h77 == _T_19[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_1;
      end else if (8'h77 == _T_15[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_120 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h78 == _T_37[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_7;
      end else if (8'h78 == _T_34[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_6;
      end else if (8'h78 == _T_31[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_5;
      end else if (8'h78 == _T_28[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_4;
      end else if (8'h78 == _T_25[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_3;
      end else if (8'h78 == _T_22[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_2;
      end else if (8'h78 == _T_19[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_1;
      end else if (8'h78 == _T_15[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_121 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h79 == _T_37[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_7;
      end else if (8'h79 == _T_34[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_6;
      end else if (8'h79 == _T_31[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_5;
      end else if (8'h79 == _T_28[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_4;
      end else if (8'h79 == _T_25[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_3;
      end else if (8'h79 == _T_22[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_2;
      end else if (8'h79 == _T_19[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_1;
      end else if (8'h79 == _T_15[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_122 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7a == _T_37[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_7;
      end else if (8'h7a == _T_34[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_6;
      end else if (8'h7a == _T_31[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_5;
      end else if (8'h7a == _T_28[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_4;
      end else if (8'h7a == _T_25[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_3;
      end else if (8'h7a == _T_22[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_2;
      end else if (8'h7a == _T_19[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_1;
      end else if (8'h7a == _T_15[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_123 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7b == _T_37[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_7;
      end else if (8'h7b == _T_34[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_6;
      end else if (8'h7b == _T_31[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_5;
      end else if (8'h7b == _T_28[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_4;
      end else if (8'h7b == _T_25[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_3;
      end else if (8'h7b == _T_22[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_2;
      end else if (8'h7b == _T_19[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_1;
      end else if (8'h7b == _T_15[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_124 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7c == _T_37[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_7;
      end else if (8'h7c == _T_34[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_6;
      end else if (8'h7c == _T_31[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_5;
      end else if (8'h7c == _T_28[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_4;
      end else if (8'h7c == _T_25[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_3;
      end else if (8'h7c == _T_22[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_2;
      end else if (8'h7c == _T_19[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_1;
      end else if (8'h7c == _T_15[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_125 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7d == _T_37[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_7;
      end else if (8'h7d == _T_34[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_6;
      end else if (8'h7d == _T_31[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_5;
      end else if (8'h7d == _T_28[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_4;
      end else if (8'h7d == _T_25[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_3;
      end else if (8'h7d == _T_22[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_2;
      end else if (8'h7d == _T_19[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_1;
      end else if (8'h7d == _T_15[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_126 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7e == _T_37[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_7;
      end else if (8'h7e == _T_34[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_6;
      end else if (8'h7e == _T_31[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_5;
      end else if (8'h7e == _T_28[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_4;
      end else if (8'h7e == _T_25[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_3;
      end else if (8'h7e == _T_22[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_2;
      end else if (8'h7e == _T_19[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_1;
      end else if (8'h7e == _T_15[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_127 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7f == _T_37[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_7;
      end else if (8'h7f == _T_34[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_6;
      end else if (8'h7f == _T_31[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_5;
      end else if (8'h7f == _T_28[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_4;
      end else if (8'h7f == _T_25[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_3;
      end else if (8'h7f == _T_22[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_2;
      end else if (8'h7f == _T_19[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_1;
      end else if (8'h7f == _T_15[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_128 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h80 == _T_37[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_7;
      end else if (8'h80 == _T_34[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_6;
      end else if (8'h80 == _T_31[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_5;
      end else if (8'h80 == _T_28[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_4;
      end else if (8'h80 == _T_25[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_3;
      end else if (8'h80 == _T_22[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_2;
      end else if (8'h80 == _T_19[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_1;
      end else if (8'h80 == _T_15[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_129 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h81 == _T_37[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_7;
      end else if (8'h81 == _T_34[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_6;
      end else if (8'h81 == _T_31[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_5;
      end else if (8'h81 == _T_28[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_4;
      end else if (8'h81 == _T_25[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_3;
      end else if (8'h81 == _T_22[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_2;
      end else if (8'h81 == _T_19[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_1;
      end else if (8'h81 == _T_15[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_130 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h82 == _T_37[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_7;
      end else if (8'h82 == _T_34[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_6;
      end else if (8'h82 == _T_31[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_5;
      end else if (8'h82 == _T_28[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_4;
      end else if (8'h82 == _T_25[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_3;
      end else if (8'h82 == _T_22[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_2;
      end else if (8'h82 == _T_19[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_1;
      end else if (8'h82 == _T_15[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_131 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h83 == _T_37[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_7;
      end else if (8'h83 == _T_34[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_6;
      end else if (8'h83 == _T_31[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_5;
      end else if (8'h83 == _T_28[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_4;
      end else if (8'h83 == _T_25[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_3;
      end else if (8'h83 == _T_22[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_2;
      end else if (8'h83 == _T_19[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_1;
      end else if (8'h83 == _T_15[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_132 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h84 == _T_37[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_7;
      end else if (8'h84 == _T_34[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_6;
      end else if (8'h84 == _T_31[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_5;
      end else if (8'h84 == _T_28[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_4;
      end else if (8'h84 == _T_25[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_3;
      end else if (8'h84 == _T_22[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_2;
      end else if (8'h84 == _T_19[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_1;
      end else if (8'h84 == _T_15[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_133 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h85 == _T_37[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_7;
      end else if (8'h85 == _T_34[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_6;
      end else if (8'h85 == _T_31[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_5;
      end else if (8'h85 == _T_28[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_4;
      end else if (8'h85 == _T_25[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_3;
      end else if (8'h85 == _T_22[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_2;
      end else if (8'h85 == _T_19[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_1;
      end else if (8'h85 == _T_15[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_134 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h86 == _T_37[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_7;
      end else if (8'h86 == _T_34[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_6;
      end else if (8'h86 == _T_31[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_5;
      end else if (8'h86 == _T_28[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_4;
      end else if (8'h86 == _T_25[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_3;
      end else if (8'h86 == _T_22[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_2;
      end else if (8'h86 == _T_19[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_1;
      end else if (8'h86 == _T_15[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_135 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h87 == _T_37[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_7;
      end else if (8'h87 == _T_34[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_6;
      end else if (8'h87 == _T_31[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_5;
      end else if (8'h87 == _T_28[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_4;
      end else if (8'h87 == _T_25[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_3;
      end else if (8'h87 == _T_22[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_2;
      end else if (8'h87 == _T_19[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_1;
      end else if (8'h87 == _T_15[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_136 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h88 == _T_37[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_7;
      end else if (8'h88 == _T_34[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_6;
      end else if (8'h88 == _T_31[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_5;
      end else if (8'h88 == _T_28[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_4;
      end else if (8'h88 == _T_25[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_3;
      end else if (8'h88 == _T_22[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_2;
      end else if (8'h88 == _T_19[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_1;
      end else if (8'h88 == _T_15[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_137 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h89 == _T_37[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_7;
      end else if (8'h89 == _T_34[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_6;
      end else if (8'h89 == _T_31[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_5;
      end else if (8'h89 == _T_28[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_4;
      end else if (8'h89 == _T_25[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_3;
      end else if (8'h89 == _T_22[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_2;
      end else if (8'h89 == _T_19[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_1;
      end else if (8'h89 == _T_15[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_138 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8a == _T_37[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_7;
      end else if (8'h8a == _T_34[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_6;
      end else if (8'h8a == _T_31[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_5;
      end else if (8'h8a == _T_28[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_4;
      end else if (8'h8a == _T_25[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_3;
      end else if (8'h8a == _T_22[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_2;
      end else if (8'h8a == _T_19[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_1;
      end else if (8'h8a == _T_15[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_139 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8b == _T_37[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_7;
      end else if (8'h8b == _T_34[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_6;
      end else if (8'h8b == _T_31[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_5;
      end else if (8'h8b == _T_28[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_4;
      end else if (8'h8b == _T_25[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_3;
      end else if (8'h8b == _T_22[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_2;
      end else if (8'h8b == _T_19[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_1;
      end else if (8'h8b == _T_15[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_140 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8c == _T_37[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_7;
      end else if (8'h8c == _T_34[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_6;
      end else if (8'h8c == _T_31[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_5;
      end else if (8'h8c == _T_28[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_4;
      end else if (8'h8c == _T_25[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_3;
      end else if (8'h8c == _T_22[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_2;
      end else if (8'h8c == _T_19[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_1;
      end else if (8'h8c == _T_15[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_141 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8d == _T_37[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_7;
      end else if (8'h8d == _T_34[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_6;
      end else if (8'h8d == _T_31[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_5;
      end else if (8'h8d == _T_28[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_4;
      end else if (8'h8d == _T_25[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_3;
      end else if (8'h8d == _T_22[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_2;
      end else if (8'h8d == _T_19[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_1;
      end else if (8'h8d == _T_15[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_142 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8e == _T_37[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_7;
      end else if (8'h8e == _T_34[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_6;
      end else if (8'h8e == _T_31[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_5;
      end else if (8'h8e == _T_28[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_4;
      end else if (8'h8e == _T_25[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_3;
      end else if (8'h8e == _T_22[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_2;
      end else if (8'h8e == _T_19[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_1;
      end else if (8'h8e == _T_15[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_143 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8f == _T_37[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_7;
      end else if (8'h8f == _T_34[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_6;
      end else if (8'h8f == _T_31[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_5;
      end else if (8'h8f == _T_28[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_4;
      end else if (8'h8f == _T_25[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_3;
      end else if (8'h8f == _T_22[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_2;
      end else if (8'h8f == _T_19[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_1;
      end else if (8'h8f == _T_15[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_144 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h90 == _T_37[7:0]) begin
        image_2_144 <= io_pixelVal_in_2_7;
      end else if (8'h90 == _T_34[7:0]) begin
        image_2_144 <= io_pixelVal_in_2_6;
      end else if (8'h90 == _T_31[7:0]) begin
        image_2_144 <= io_pixelVal_in_2_5;
      end else if (8'h90 == _T_28[7:0]) begin
        image_2_144 <= io_pixelVal_in_2_4;
      end else if (8'h90 == _T_25[7:0]) begin
        image_2_144 <= io_pixelVal_in_2_3;
      end else if (8'h90 == _T_22[7:0]) begin
        image_2_144 <= io_pixelVal_in_2_2;
      end else if (8'h90 == _T_19[7:0]) begin
        image_2_144 <= io_pixelVal_in_2_1;
      end else if (8'h90 == _T_15[7:0]) begin
        image_2_144 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_145 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h91 == _T_37[7:0]) begin
        image_2_145 <= io_pixelVal_in_2_7;
      end else if (8'h91 == _T_34[7:0]) begin
        image_2_145 <= io_pixelVal_in_2_6;
      end else if (8'h91 == _T_31[7:0]) begin
        image_2_145 <= io_pixelVal_in_2_5;
      end else if (8'h91 == _T_28[7:0]) begin
        image_2_145 <= io_pixelVal_in_2_4;
      end else if (8'h91 == _T_25[7:0]) begin
        image_2_145 <= io_pixelVal_in_2_3;
      end else if (8'h91 == _T_22[7:0]) begin
        image_2_145 <= io_pixelVal_in_2_2;
      end else if (8'h91 == _T_19[7:0]) begin
        image_2_145 <= io_pixelVal_in_2_1;
      end else if (8'h91 == _T_15[7:0]) begin
        image_2_145 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_146 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h92 == _T_37[7:0]) begin
        image_2_146 <= io_pixelVal_in_2_7;
      end else if (8'h92 == _T_34[7:0]) begin
        image_2_146 <= io_pixelVal_in_2_6;
      end else if (8'h92 == _T_31[7:0]) begin
        image_2_146 <= io_pixelVal_in_2_5;
      end else if (8'h92 == _T_28[7:0]) begin
        image_2_146 <= io_pixelVal_in_2_4;
      end else if (8'h92 == _T_25[7:0]) begin
        image_2_146 <= io_pixelVal_in_2_3;
      end else if (8'h92 == _T_22[7:0]) begin
        image_2_146 <= io_pixelVal_in_2_2;
      end else if (8'h92 == _T_19[7:0]) begin
        image_2_146 <= io_pixelVal_in_2_1;
      end else if (8'h92 == _T_15[7:0]) begin
        image_2_146 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_147 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h93 == _T_37[7:0]) begin
        image_2_147 <= io_pixelVal_in_2_7;
      end else if (8'h93 == _T_34[7:0]) begin
        image_2_147 <= io_pixelVal_in_2_6;
      end else if (8'h93 == _T_31[7:0]) begin
        image_2_147 <= io_pixelVal_in_2_5;
      end else if (8'h93 == _T_28[7:0]) begin
        image_2_147 <= io_pixelVal_in_2_4;
      end else if (8'h93 == _T_25[7:0]) begin
        image_2_147 <= io_pixelVal_in_2_3;
      end else if (8'h93 == _T_22[7:0]) begin
        image_2_147 <= io_pixelVal_in_2_2;
      end else if (8'h93 == _T_19[7:0]) begin
        image_2_147 <= io_pixelVal_in_2_1;
      end else if (8'h93 == _T_15[7:0]) begin
        image_2_147 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_148 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h94 == _T_37[7:0]) begin
        image_2_148 <= io_pixelVal_in_2_7;
      end else if (8'h94 == _T_34[7:0]) begin
        image_2_148 <= io_pixelVal_in_2_6;
      end else if (8'h94 == _T_31[7:0]) begin
        image_2_148 <= io_pixelVal_in_2_5;
      end else if (8'h94 == _T_28[7:0]) begin
        image_2_148 <= io_pixelVal_in_2_4;
      end else if (8'h94 == _T_25[7:0]) begin
        image_2_148 <= io_pixelVal_in_2_3;
      end else if (8'h94 == _T_22[7:0]) begin
        image_2_148 <= io_pixelVal_in_2_2;
      end else if (8'h94 == _T_19[7:0]) begin
        image_2_148 <= io_pixelVal_in_2_1;
      end else if (8'h94 == _T_15[7:0]) begin
        image_2_148 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_149 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h95 == _T_37[7:0]) begin
        image_2_149 <= io_pixelVal_in_2_7;
      end else if (8'h95 == _T_34[7:0]) begin
        image_2_149 <= io_pixelVal_in_2_6;
      end else if (8'h95 == _T_31[7:0]) begin
        image_2_149 <= io_pixelVal_in_2_5;
      end else if (8'h95 == _T_28[7:0]) begin
        image_2_149 <= io_pixelVal_in_2_4;
      end else if (8'h95 == _T_25[7:0]) begin
        image_2_149 <= io_pixelVal_in_2_3;
      end else if (8'h95 == _T_22[7:0]) begin
        image_2_149 <= io_pixelVal_in_2_2;
      end else if (8'h95 == _T_19[7:0]) begin
        image_2_149 <= io_pixelVal_in_2_1;
      end else if (8'h95 == _T_15[7:0]) begin
        image_2_149 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_150 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h96 == _T_37[7:0]) begin
        image_2_150 <= io_pixelVal_in_2_7;
      end else if (8'h96 == _T_34[7:0]) begin
        image_2_150 <= io_pixelVal_in_2_6;
      end else if (8'h96 == _T_31[7:0]) begin
        image_2_150 <= io_pixelVal_in_2_5;
      end else if (8'h96 == _T_28[7:0]) begin
        image_2_150 <= io_pixelVal_in_2_4;
      end else if (8'h96 == _T_25[7:0]) begin
        image_2_150 <= io_pixelVal_in_2_3;
      end else if (8'h96 == _T_22[7:0]) begin
        image_2_150 <= io_pixelVal_in_2_2;
      end else if (8'h96 == _T_19[7:0]) begin
        image_2_150 <= io_pixelVal_in_2_1;
      end else if (8'h96 == _T_15[7:0]) begin
        image_2_150 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_151 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h97 == _T_37[7:0]) begin
        image_2_151 <= io_pixelVal_in_2_7;
      end else if (8'h97 == _T_34[7:0]) begin
        image_2_151 <= io_pixelVal_in_2_6;
      end else if (8'h97 == _T_31[7:0]) begin
        image_2_151 <= io_pixelVal_in_2_5;
      end else if (8'h97 == _T_28[7:0]) begin
        image_2_151 <= io_pixelVal_in_2_4;
      end else if (8'h97 == _T_25[7:0]) begin
        image_2_151 <= io_pixelVal_in_2_3;
      end else if (8'h97 == _T_22[7:0]) begin
        image_2_151 <= io_pixelVal_in_2_2;
      end else if (8'h97 == _T_19[7:0]) begin
        image_2_151 <= io_pixelVal_in_2_1;
      end else if (8'h97 == _T_15[7:0]) begin
        image_2_151 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_152 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h98 == _T_37[7:0]) begin
        image_2_152 <= io_pixelVal_in_2_7;
      end else if (8'h98 == _T_34[7:0]) begin
        image_2_152 <= io_pixelVal_in_2_6;
      end else if (8'h98 == _T_31[7:0]) begin
        image_2_152 <= io_pixelVal_in_2_5;
      end else if (8'h98 == _T_28[7:0]) begin
        image_2_152 <= io_pixelVal_in_2_4;
      end else if (8'h98 == _T_25[7:0]) begin
        image_2_152 <= io_pixelVal_in_2_3;
      end else if (8'h98 == _T_22[7:0]) begin
        image_2_152 <= io_pixelVal_in_2_2;
      end else if (8'h98 == _T_19[7:0]) begin
        image_2_152 <= io_pixelVal_in_2_1;
      end else if (8'h98 == _T_15[7:0]) begin
        image_2_152 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_153 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h99 == _T_37[7:0]) begin
        image_2_153 <= io_pixelVal_in_2_7;
      end else if (8'h99 == _T_34[7:0]) begin
        image_2_153 <= io_pixelVal_in_2_6;
      end else if (8'h99 == _T_31[7:0]) begin
        image_2_153 <= io_pixelVal_in_2_5;
      end else if (8'h99 == _T_28[7:0]) begin
        image_2_153 <= io_pixelVal_in_2_4;
      end else if (8'h99 == _T_25[7:0]) begin
        image_2_153 <= io_pixelVal_in_2_3;
      end else if (8'h99 == _T_22[7:0]) begin
        image_2_153 <= io_pixelVal_in_2_2;
      end else if (8'h99 == _T_19[7:0]) begin
        image_2_153 <= io_pixelVal_in_2_1;
      end else if (8'h99 == _T_15[7:0]) begin
        image_2_153 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_154 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9a == _T_37[7:0]) begin
        image_2_154 <= io_pixelVal_in_2_7;
      end else if (8'h9a == _T_34[7:0]) begin
        image_2_154 <= io_pixelVal_in_2_6;
      end else if (8'h9a == _T_31[7:0]) begin
        image_2_154 <= io_pixelVal_in_2_5;
      end else if (8'h9a == _T_28[7:0]) begin
        image_2_154 <= io_pixelVal_in_2_4;
      end else if (8'h9a == _T_25[7:0]) begin
        image_2_154 <= io_pixelVal_in_2_3;
      end else if (8'h9a == _T_22[7:0]) begin
        image_2_154 <= io_pixelVal_in_2_2;
      end else if (8'h9a == _T_19[7:0]) begin
        image_2_154 <= io_pixelVal_in_2_1;
      end else if (8'h9a == _T_15[7:0]) begin
        image_2_154 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_155 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9b == _T_37[7:0]) begin
        image_2_155 <= io_pixelVal_in_2_7;
      end else if (8'h9b == _T_34[7:0]) begin
        image_2_155 <= io_pixelVal_in_2_6;
      end else if (8'h9b == _T_31[7:0]) begin
        image_2_155 <= io_pixelVal_in_2_5;
      end else if (8'h9b == _T_28[7:0]) begin
        image_2_155 <= io_pixelVal_in_2_4;
      end else if (8'h9b == _T_25[7:0]) begin
        image_2_155 <= io_pixelVal_in_2_3;
      end else if (8'h9b == _T_22[7:0]) begin
        image_2_155 <= io_pixelVal_in_2_2;
      end else if (8'h9b == _T_19[7:0]) begin
        image_2_155 <= io_pixelVal_in_2_1;
      end else if (8'h9b == _T_15[7:0]) begin
        image_2_155 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_156 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9c == _T_37[7:0]) begin
        image_2_156 <= io_pixelVal_in_2_7;
      end else if (8'h9c == _T_34[7:0]) begin
        image_2_156 <= io_pixelVal_in_2_6;
      end else if (8'h9c == _T_31[7:0]) begin
        image_2_156 <= io_pixelVal_in_2_5;
      end else if (8'h9c == _T_28[7:0]) begin
        image_2_156 <= io_pixelVal_in_2_4;
      end else if (8'h9c == _T_25[7:0]) begin
        image_2_156 <= io_pixelVal_in_2_3;
      end else if (8'h9c == _T_22[7:0]) begin
        image_2_156 <= io_pixelVal_in_2_2;
      end else if (8'h9c == _T_19[7:0]) begin
        image_2_156 <= io_pixelVal_in_2_1;
      end else if (8'h9c == _T_15[7:0]) begin
        image_2_156 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_157 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9d == _T_37[7:0]) begin
        image_2_157 <= io_pixelVal_in_2_7;
      end else if (8'h9d == _T_34[7:0]) begin
        image_2_157 <= io_pixelVal_in_2_6;
      end else if (8'h9d == _T_31[7:0]) begin
        image_2_157 <= io_pixelVal_in_2_5;
      end else if (8'h9d == _T_28[7:0]) begin
        image_2_157 <= io_pixelVal_in_2_4;
      end else if (8'h9d == _T_25[7:0]) begin
        image_2_157 <= io_pixelVal_in_2_3;
      end else if (8'h9d == _T_22[7:0]) begin
        image_2_157 <= io_pixelVal_in_2_2;
      end else if (8'h9d == _T_19[7:0]) begin
        image_2_157 <= io_pixelVal_in_2_1;
      end else if (8'h9d == _T_15[7:0]) begin
        image_2_157 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_158 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9e == _T_37[7:0]) begin
        image_2_158 <= io_pixelVal_in_2_7;
      end else if (8'h9e == _T_34[7:0]) begin
        image_2_158 <= io_pixelVal_in_2_6;
      end else if (8'h9e == _T_31[7:0]) begin
        image_2_158 <= io_pixelVal_in_2_5;
      end else if (8'h9e == _T_28[7:0]) begin
        image_2_158 <= io_pixelVal_in_2_4;
      end else if (8'h9e == _T_25[7:0]) begin
        image_2_158 <= io_pixelVal_in_2_3;
      end else if (8'h9e == _T_22[7:0]) begin
        image_2_158 <= io_pixelVal_in_2_2;
      end else if (8'h9e == _T_19[7:0]) begin
        image_2_158 <= io_pixelVal_in_2_1;
      end else if (8'h9e == _T_15[7:0]) begin
        image_2_158 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_159 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9f == _T_37[7:0]) begin
        image_2_159 <= io_pixelVal_in_2_7;
      end else if (8'h9f == _T_34[7:0]) begin
        image_2_159 <= io_pixelVal_in_2_6;
      end else if (8'h9f == _T_31[7:0]) begin
        image_2_159 <= io_pixelVal_in_2_5;
      end else if (8'h9f == _T_28[7:0]) begin
        image_2_159 <= io_pixelVal_in_2_4;
      end else if (8'h9f == _T_25[7:0]) begin
        image_2_159 <= io_pixelVal_in_2_3;
      end else if (8'h9f == _T_22[7:0]) begin
        image_2_159 <= io_pixelVal_in_2_2;
      end else if (8'h9f == _T_19[7:0]) begin
        image_2_159 <= io_pixelVal_in_2_1;
      end else if (8'h9f == _T_15[7:0]) begin
        image_2_159 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_160 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha0 == _T_37[7:0]) begin
        image_2_160 <= io_pixelVal_in_2_7;
      end else if (8'ha0 == _T_34[7:0]) begin
        image_2_160 <= io_pixelVal_in_2_6;
      end else if (8'ha0 == _T_31[7:0]) begin
        image_2_160 <= io_pixelVal_in_2_5;
      end else if (8'ha0 == _T_28[7:0]) begin
        image_2_160 <= io_pixelVal_in_2_4;
      end else if (8'ha0 == _T_25[7:0]) begin
        image_2_160 <= io_pixelVal_in_2_3;
      end else if (8'ha0 == _T_22[7:0]) begin
        image_2_160 <= io_pixelVal_in_2_2;
      end else if (8'ha0 == _T_19[7:0]) begin
        image_2_160 <= io_pixelVal_in_2_1;
      end else if (8'ha0 == _T_15[7:0]) begin
        image_2_160 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_161 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha1 == _T_37[7:0]) begin
        image_2_161 <= io_pixelVal_in_2_7;
      end else if (8'ha1 == _T_34[7:0]) begin
        image_2_161 <= io_pixelVal_in_2_6;
      end else if (8'ha1 == _T_31[7:0]) begin
        image_2_161 <= io_pixelVal_in_2_5;
      end else if (8'ha1 == _T_28[7:0]) begin
        image_2_161 <= io_pixelVal_in_2_4;
      end else if (8'ha1 == _T_25[7:0]) begin
        image_2_161 <= io_pixelVal_in_2_3;
      end else if (8'ha1 == _T_22[7:0]) begin
        image_2_161 <= io_pixelVal_in_2_2;
      end else if (8'ha1 == _T_19[7:0]) begin
        image_2_161 <= io_pixelVal_in_2_1;
      end else if (8'ha1 == _T_15[7:0]) begin
        image_2_161 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_162 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha2 == _T_37[7:0]) begin
        image_2_162 <= io_pixelVal_in_2_7;
      end else if (8'ha2 == _T_34[7:0]) begin
        image_2_162 <= io_pixelVal_in_2_6;
      end else if (8'ha2 == _T_31[7:0]) begin
        image_2_162 <= io_pixelVal_in_2_5;
      end else if (8'ha2 == _T_28[7:0]) begin
        image_2_162 <= io_pixelVal_in_2_4;
      end else if (8'ha2 == _T_25[7:0]) begin
        image_2_162 <= io_pixelVal_in_2_3;
      end else if (8'ha2 == _T_22[7:0]) begin
        image_2_162 <= io_pixelVal_in_2_2;
      end else if (8'ha2 == _T_19[7:0]) begin
        image_2_162 <= io_pixelVal_in_2_1;
      end else if (8'ha2 == _T_15[7:0]) begin
        image_2_162 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_163 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha3 == _T_37[7:0]) begin
        image_2_163 <= io_pixelVal_in_2_7;
      end else if (8'ha3 == _T_34[7:0]) begin
        image_2_163 <= io_pixelVal_in_2_6;
      end else if (8'ha3 == _T_31[7:0]) begin
        image_2_163 <= io_pixelVal_in_2_5;
      end else if (8'ha3 == _T_28[7:0]) begin
        image_2_163 <= io_pixelVal_in_2_4;
      end else if (8'ha3 == _T_25[7:0]) begin
        image_2_163 <= io_pixelVal_in_2_3;
      end else if (8'ha3 == _T_22[7:0]) begin
        image_2_163 <= io_pixelVal_in_2_2;
      end else if (8'ha3 == _T_19[7:0]) begin
        image_2_163 <= io_pixelVal_in_2_1;
      end else if (8'ha3 == _T_15[7:0]) begin
        image_2_163 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_164 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha4 == _T_37[7:0]) begin
        image_2_164 <= io_pixelVal_in_2_7;
      end else if (8'ha4 == _T_34[7:0]) begin
        image_2_164 <= io_pixelVal_in_2_6;
      end else if (8'ha4 == _T_31[7:0]) begin
        image_2_164 <= io_pixelVal_in_2_5;
      end else if (8'ha4 == _T_28[7:0]) begin
        image_2_164 <= io_pixelVal_in_2_4;
      end else if (8'ha4 == _T_25[7:0]) begin
        image_2_164 <= io_pixelVal_in_2_3;
      end else if (8'ha4 == _T_22[7:0]) begin
        image_2_164 <= io_pixelVal_in_2_2;
      end else if (8'ha4 == _T_19[7:0]) begin
        image_2_164 <= io_pixelVal_in_2_1;
      end else if (8'ha4 == _T_15[7:0]) begin
        image_2_164 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_165 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha5 == _T_37[7:0]) begin
        image_2_165 <= io_pixelVal_in_2_7;
      end else if (8'ha5 == _T_34[7:0]) begin
        image_2_165 <= io_pixelVal_in_2_6;
      end else if (8'ha5 == _T_31[7:0]) begin
        image_2_165 <= io_pixelVal_in_2_5;
      end else if (8'ha5 == _T_28[7:0]) begin
        image_2_165 <= io_pixelVal_in_2_4;
      end else if (8'ha5 == _T_25[7:0]) begin
        image_2_165 <= io_pixelVal_in_2_3;
      end else if (8'ha5 == _T_22[7:0]) begin
        image_2_165 <= io_pixelVal_in_2_2;
      end else if (8'ha5 == _T_19[7:0]) begin
        image_2_165 <= io_pixelVal_in_2_1;
      end else if (8'ha5 == _T_15[7:0]) begin
        image_2_165 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_166 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha6 == _T_37[7:0]) begin
        image_2_166 <= io_pixelVal_in_2_7;
      end else if (8'ha6 == _T_34[7:0]) begin
        image_2_166 <= io_pixelVal_in_2_6;
      end else if (8'ha6 == _T_31[7:0]) begin
        image_2_166 <= io_pixelVal_in_2_5;
      end else if (8'ha6 == _T_28[7:0]) begin
        image_2_166 <= io_pixelVal_in_2_4;
      end else if (8'ha6 == _T_25[7:0]) begin
        image_2_166 <= io_pixelVal_in_2_3;
      end else if (8'ha6 == _T_22[7:0]) begin
        image_2_166 <= io_pixelVal_in_2_2;
      end else if (8'ha6 == _T_19[7:0]) begin
        image_2_166 <= io_pixelVal_in_2_1;
      end else if (8'ha6 == _T_15[7:0]) begin
        image_2_166 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_167 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha7 == _T_37[7:0]) begin
        image_2_167 <= io_pixelVal_in_2_7;
      end else if (8'ha7 == _T_34[7:0]) begin
        image_2_167 <= io_pixelVal_in_2_6;
      end else if (8'ha7 == _T_31[7:0]) begin
        image_2_167 <= io_pixelVal_in_2_5;
      end else if (8'ha7 == _T_28[7:0]) begin
        image_2_167 <= io_pixelVal_in_2_4;
      end else if (8'ha7 == _T_25[7:0]) begin
        image_2_167 <= io_pixelVal_in_2_3;
      end else if (8'ha7 == _T_22[7:0]) begin
        image_2_167 <= io_pixelVal_in_2_2;
      end else if (8'ha7 == _T_19[7:0]) begin
        image_2_167 <= io_pixelVal_in_2_1;
      end else if (8'ha7 == _T_15[7:0]) begin
        image_2_167 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_168 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha8 == _T_37[7:0]) begin
        image_2_168 <= io_pixelVal_in_2_7;
      end else if (8'ha8 == _T_34[7:0]) begin
        image_2_168 <= io_pixelVal_in_2_6;
      end else if (8'ha8 == _T_31[7:0]) begin
        image_2_168 <= io_pixelVal_in_2_5;
      end else if (8'ha8 == _T_28[7:0]) begin
        image_2_168 <= io_pixelVal_in_2_4;
      end else if (8'ha8 == _T_25[7:0]) begin
        image_2_168 <= io_pixelVal_in_2_3;
      end else if (8'ha8 == _T_22[7:0]) begin
        image_2_168 <= io_pixelVal_in_2_2;
      end else if (8'ha8 == _T_19[7:0]) begin
        image_2_168 <= io_pixelVal_in_2_1;
      end else if (8'ha8 == _T_15[7:0]) begin
        image_2_168 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_169 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha9 == _T_37[7:0]) begin
        image_2_169 <= io_pixelVal_in_2_7;
      end else if (8'ha9 == _T_34[7:0]) begin
        image_2_169 <= io_pixelVal_in_2_6;
      end else if (8'ha9 == _T_31[7:0]) begin
        image_2_169 <= io_pixelVal_in_2_5;
      end else if (8'ha9 == _T_28[7:0]) begin
        image_2_169 <= io_pixelVal_in_2_4;
      end else if (8'ha9 == _T_25[7:0]) begin
        image_2_169 <= io_pixelVal_in_2_3;
      end else if (8'ha9 == _T_22[7:0]) begin
        image_2_169 <= io_pixelVal_in_2_2;
      end else if (8'ha9 == _T_19[7:0]) begin
        image_2_169 <= io_pixelVal_in_2_1;
      end else if (8'ha9 == _T_15[7:0]) begin
        image_2_169 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_170 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'haa == _T_37[7:0]) begin
        image_2_170 <= io_pixelVal_in_2_7;
      end else if (8'haa == _T_34[7:0]) begin
        image_2_170 <= io_pixelVal_in_2_6;
      end else if (8'haa == _T_31[7:0]) begin
        image_2_170 <= io_pixelVal_in_2_5;
      end else if (8'haa == _T_28[7:0]) begin
        image_2_170 <= io_pixelVal_in_2_4;
      end else if (8'haa == _T_25[7:0]) begin
        image_2_170 <= io_pixelVal_in_2_3;
      end else if (8'haa == _T_22[7:0]) begin
        image_2_170 <= io_pixelVal_in_2_2;
      end else if (8'haa == _T_19[7:0]) begin
        image_2_170 <= io_pixelVal_in_2_1;
      end else if (8'haa == _T_15[7:0]) begin
        image_2_170 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_171 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hab == _T_37[7:0]) begin
        image_2_171 <= io_pixelVal_in_2_7;
      end else if (8'hab == _T_34[7:0]) begin
        image_2_171 <= io_pixelVal_in_2_6;
      end else if (8'hab == _T_31[7:0]) begin
        image_2_171 <= io_pixelVal_in_2_5;
      end else if (8'hab == _T_28[7:0]) begin
        image_2_171 <= io_pixelVal_in_2_4;
      end else if (8'hab == _T_25[7:0]) begin
        image_2_171 <= io_pixelVal_in_2_3;
      end else if (8'hab == _T_22[7:0]) begin
        image_2_171 <= io_pixelVal_in_2_2;
      end else if (8'hab == _T_19[7:0]) begin
        image_2_171 <= io_pixelVal_in_2_1;
      end else if (8'hab == _T_15[7:0]) begin
        image_2_171 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_172 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hac == _T_37[7:0]) begin
        image_2_172 <= io_pixelVal_in_2_7;
      end else if (8'hac == _T_34[7:0]) begin
        image_2_172 <= io_pixelVal_in_2_6;
      end else if (8'hac == _T_31[7:0]) begin
        image_2_172 <= io_pixelVal_in_2_5;
      end else if (8'hac == _T_28[7:0]) begin
        image_2_172 <= io_pixelVal_in_2_4;
      end else if (8'hac == _T_25[7:0]) begin
        image_2_172 <= io_pixelVal_in_2_3;
      end else if (8'hac == _T_22[7:0]) begin
        image_2_172 <= io_pixelVal_in_2_2;
      end else if (8'hac == _T_19[7:0]) begin
        image_2_172 <= io_pixelVal_in_2_1;
      end else if (8'hac == _T_15[7:0]) begin
        image_2_172 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_173 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'had == _T_37[7:0]) begin
        image_2_173 <= io_pixelVal_in_2_7;
      end else if (8'had == _T_34[7:0]) begin
        image_2_173 <= io_pixelVal_in_2_6;
      end else if (8'had == _T_31[7:0]) begin
        image_2_173 <= io_pixelVal_in_2_5;
      end else if (8'had == _T_28[7:0]) begin
        image_2_173 <= io_pixelVal_in_2_4;
      end else if (8'had == _T_25[7:0]) begin
        image_2_173 <= io_pixelVal_in_2_3;
      end else if (8'had == _T_22[7:0]) begin
        image_2_173 <= io_pixelVal_in_2_2;
      end else if (8'had == _T_19[7:0]) begin
        image_2_173 <= io_pixelVal_in_2_1;
      end else if (8'had == _T_15[7:0]) begin
        image_2_173 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_174 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hae == _T_37[7:0]) begin
        image_2_174 <= io_pixelVal_in_2_7;
      end else if (8'hae == _T_34[7:0]) begin
        image_2_174 <= io_pixelVal_in_2_6;
      end else if (8'hae == _T_31[7:0]) begin
        image_2_174 <= io_pixelVal_in_2_5;
      end else if (8'hae == _T_28[7:0]) begin
        image_2_174 <= io_pixelVal_in_2_4;
      end else if (8'hae == _T_25[7:0]) begin
        image_2_174 <= io_pixelVal_in_2_3;
      end else if (8'hae == _T_22[7:0]) begin
        image_2_174 <= io_pixelVal_in_2_2;
      end else if (8'hae == _T_19[7:0]) begin
        image_2_174 <= io_pixelVal_in_2_1;
      end else if (8'hae == _T_15[7:0]) begin
        image_2_174 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_175 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'haf == _T_37[7:0]) begin
        image_2_175 <= io_pixelVal_in_2_7;
      end else if (8'haf == _T_34[7:0]) begin
        image_2_175 <= io_pixelVal_in_2_6;
      end else if (8'haf == _T_31[7:0]) begin
        image_2_175 <= io_pixelVal_in_2_5;
      end else if (8'haf == _T_28[7:0]) begin
        image_2_175 <= io_pixelVal_in_2_4;
      end else if (8'haf == _T_25[7:0]) begin
        image_2_175 <= io_pixelVal_in_2_3;
      end else if (8'haf == _T_22[7:0]) begin
        image_2_175 <= io_pixelVal_in_2_2;
      end else if (8'haf == _T_19[7:0]) begin
        image_2_175 <= io_pixelVal_in_2_1;
      end else if (8'haf == _T_15[7:0]) begin
        image_2_175 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_176 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb0 == _T_37[7:0]) begin
        image_2_176 <= io_pixelVal_in_2_7;
      end else if (8'hb0 == _T_34[7:0]) begin
        image_2_176 <= io_pixelVal_in_2_6;
      end else if (8'hb0 == _T_31[7:0]) begin
        image_2_176 <= io_pixelVal_in_2_5;
      end else if (8'hb0 == _T_28[7:0]) begin
        image_2_176 <= io_pixelVal_in_2_4;
      end else if (8'hb0 == _T_25[7:0]) begin
        image_2_176 <= io_pixelVal_in_2_3;
      end else if (8'hb0 == _T_22[7:0]) begin
        image_2_176 <= io_pixelVal_in_2_2;
      end else if (8'hb0 == _T_19[7:0]) begin
        image_2_176 <= io_pixelVal_in_2_1;
      end else if (8'hb0 == _T_15[7:0]) begin
        image_2_176 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_177 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb1 == _T_37[7:0]) begin
        image_2_177 <= io_pixelVal_in_2_7;
      end else if (8'hb1 == _T_34[7:0]) begin
        image_2_177 <= io_pixelVal_in_2_6;
      end else if (8'hb1 == _T_31[7:0]) begin
        image_2_177 <= io_pixelVal_in_2_5;
      end else if (8'hb1 == _T_28[7:0]) begin
        image_2_177 <= io_pixelVal_in_2_4;
      end else if (8'hb1 == _T_25[7:0]) begin
        image_2_177 <= io_pixelVal_in_2_3;
      end else if (8'hb1 == _T_22[7:0]) begin
        image_2_177 <= io_pixelVal_in_2_2;
      end else if (8'hb1 == _T_19[7:0]) begin
        image_2_177 <= io_pixelVal_in_2_1;
      end else if (8'hb1 == _T_15[7:0]) begin
        image_2_177 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_178 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb2 == _T_37[7:0]) begin
        image_2_178 <= io_pixelVal_in_2_7;
      end else if (8'hb2 == _T_34[7:0]) begin
        image_2_178 <= io_pixelVal_in_2_6;
      end else if (8'hb2 == _T_31[7:0]) begin
        image_2_178 <= io_pixelVal_in_2_5;
      end else if (8'hb2 == _T_28[7:0]) begin
        image_2_178 <= io_pixelVal_in_2_4;
      end else if (8'hb2 == _T_25[7:0]) begin
        image_2_178 <= io_pixelVal_in_2_3;
      end else if (8'hb2 == _T_22[7:0]) begin
        image_2_178 <= io_pixelVal_in_2_2;
      end else if (8'hb2 == _T_19[7:0]) begin
        image_2_178 <= io_pixelVal_in_2_1;
      end else if (8'hb2 == _T_15[7:0]) begin
        image_2_178 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_179 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb3 == _T_37[7:0]) begin
        image_2_179 <= io_pixelVal_in_2_7;
      end else if (8'hb3 == _T_34[7:0]) begin
        image_2_179 <= io_pixelVal_in_2_6;
      end else if (8'hb3 == _T_31[7:0]) begin
        image_2_179 <= io_pixelVal_in_2_5;
      end else if (8'hb3 == _T_28[7:0]) begin
        image_2_179 <= io_pixelVal_in_2_4;
      end else if (8'hb3 == _T_25[7:0]) begin
        image_2_179 <= io_pixelVal_in_2_3;
      end else if (8'hb3 == _T_22[7:0]) begin
        image_2_179 <= io_pixelVal_in_2_2;
      end else if (8'hb3 == _T_19[7:0]) begin
        image_2_179 <= io_pixelVal_in_2_1;
      end else if (8'hb3 == _T_15[7:0]) begin
        image_2_179 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_180 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb4 == _T_37[7:0]) begin
        image_2_180 <= io_pixelVal_in_2_7;
      end else if (8'hb4 == _T_34[7:0]) begin
        image_2_180 <= io_pixelVal_in_2_6;
      end else if (8'hb4 == _T_31[7:0]) begin
        image_2_180 <= io_pixelVal_in_2_5;
      end else if (8'hb4 == _T_28[7:0]) begin
        image_2_180 <= io_pixelVal_in_2_4;
      end else if (8'hb4 == _T_25[7:0]) begin
        image_2_180 <= io_pixelVal_in_2_3;
      end else if (8'hb4 == _T_22[7:0]) begin
        image_2_180 <= io_pixelVal_in_2_2;
      end else if (8'hb4 == _T_19[7:0]) begin
        image_2_180 <= io_pixelVal_in_2_1;
      end else if (8'hb4 == _T_15[7:0]) begin
        image_2_180 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_181 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb5 == _T_37[7:0]) begin
        image_2_181 <= io_pixelVal_in_2_7;
      end else if (8'hb5 == _T_34[7:0]) begin
        image_2_181 <= io_pixelVal_in_2_6;
      end else if (8'hb5 == _T_31[7:0]) begin
        image_2_181 <= io_pixelVal_in_2_5;
      end else if (8'hb5 == _T_28[7:0]) begin
        image_2_181 <= io_pixelVal_in_2_4;
      end else if (8'hb5 == _T_25[7:0]) begin
        image_2_181 <= io_pixelVal_in_2_3;
      end else if (8'hb5 == _T_22[7:0]) begin
        image_2_181 <= io_pixelVal_in_2_2;
      end else if (8'hb5 == _T_19[7:0]) begin
        image_2_181 <= io_pixelVal_in_2_1;
      end else if (8'hb5 == _T_15[7:0]) begin
        image_2_181 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_182 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb6 == _T_37[7:0]) begin
        image_2_182 <= io_pixelVal_in_2_7;
      end else if (8'hb6 == _T_34[7:0]) begin
        image_2_182 <= io_pixelVal_in_2_6;
      end else if (8'hb6 == _T_31[7:0]) begin
        image_2_182 <= io_pixelVal_in_2_5;
      end else if (8'hb6 == _T_28[7:0]) begin
        image_2_182 <= io_pixelVal_in_2_4;
      end else if (8'hb6 == _T_25[7:0]) begin
        image_2_182 <= io_pixelVal_in_2_3;
      end else if (8'hb6 == _T_22[7:0]) begin
        image_2_182 <= io_pixelVal_in_2_2;
      end else if (8'hb6 == _T_19[7:0]) begin
        image_2_182 <= io_pixelVal_in_2_1;
      end else if (8'hb6 == _T_15[7:0]) begin
        image_2_182 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_183 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb7 == _T_37[7:0]) begin
        image_2_183 <= io_pixelVal_in_2_7;
      end else if (8'hb7 == _T_34[7:0]) begin
        image_2_183 <= io_pixelVal_in_2_6;
      end else if (8'hb7 == _T_31[7:0]) begin
        image_2_183 <= io_pixelVal_in_2_5;
      end else if (8'hb7 == _T_28[7:0]) begin
        image_2_183 <= io_pixelVal_in_2_4;
      end else if (8'hb7 == _T_25[7:0]) begin
        image_2_183 <= io_pixelVal_in_2_3;
      end else if (8'hb7 == _T_22[7:0]) begin
        image_2_183 <= io_pixelVal_in_2_2;
      end else if (8'hb7 == _T_19[7:0]) begin
        image_2_183 <= io_pixelVal_in_2_1;
      end else if (8'hb7 == _T_15[7:0]) begin
        image_2_183 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_184 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb8 == _T_37[7:0]) begin
        image_2_184 <= io_pixelVal_in_2_7;
      end else if (8'hb8 == _T_34[7:0]) begin
        image_2_184 <= io_pixelVal_in_2_6;
      end else if (8'hb8 == _T_31[7:0]) begin
        image_2_184 <= io_pixelVal_in_2_5;
      end else if (8'hb8 == _T_28[7:0]) begin
        image_2_184 <= io_pixelVal_in_2_4;
      end else if (8'hb8 == _T_25[7:0]) begin
        image_2_184 <= io_pixelVal_in_2_3;
      end else if (8'hb8 == _T_22[7:0]) begin
        image_2_184 <= io_pixelVal_in_2_2;
      end else if (8'hb8 == _T_19[7:0]) begin
        image_2_184 <= io_pixelVal_in_2_1;
      end else if (8'hb8 == _T_15[7:0]) begin
        image_2_184 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_185 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb9 == _T_37[7:0]) begin
        image_2_185 <= io_pixelVal_in_2_7;
      end else if (8'hb9 == _T_34[7:0]) begin
        image_2_185 <= io_pixelVal_in_2_6;
      end else if (8'hb9 == _T_31[7:0]) begin
        image_2_185 <= io_pixelVal_in_2_5;
      end else if (8'hb9 == _T_28[7:0]) begin
        image_2_185 <= io_pixelVal_in_2_4;
      end else if (8'hb9 == _T_25[7:0]) begin
        image_2_185 <= io_pixelVal_in_2_3;
      end else if (8'hb9 == _T_22[7:0]) begin
        image_2_185 <= io_pixelVal_in_2_2;
      end else if (8'hb9 == _T_19[7:0]) begin
        image_2_185 <= io_pixelVal_in_2_1;
      end else if (8'hb9 == _T_15[7:0]) begin
        image_2_185 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_186 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hba == _T_37[7:0]) begin
        image_2_186 <= io_pixelVal_in_2_7;
      end else if (8'hba == _T_34[7:0]) begin
        image_2_186 <= io_pixelVal_in_2_6;
      end else if (8'hba == _T_31[7:0]) begin
        image_2_186 <= io_pixelVal_in_2_5;
      end else if (8'hba == _T_28[7:0]) begin
        image_2_186 <= io_pixelVal_in_2_4;
      end else if (8'hba == _T_25[7:0]) begin
        image_2_186 <= io_pixelVal_in_2_3;
      end else if (8'hba == _T_22[7:0]) begin
        image_2_186 <= io_pixelVal_in_2_2;
      end else if (8'hba == _T_19[7:0]) begin
        image_2_186 <= io_pixelVal_in_2_1;
      end else if (8'hba == _T_15[7:0]) begin
        image_2_186 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_187 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbb == _T_37[7:0]) begin
        image_2_187 <= io_pixelVal_in_2_7;
      end else if (8'hbb == _T_34[7:0]) begin
        image_2_187 <= io_pixelVal_in_2_6;
      end else if (8'hbb == _T_31[7:0]) begin
        image_2_187 <= io_pixelVal_in_2_5;
      end else if (8'hbb == _T_28[7:0]) begin
        image_2_187 <= io_pixelVal_in_2_4;
      end else if (8'hbb == _T_25[7:0]) begin
        image_2_187 <= io_pixelVal_in_2_3;
      end else if (8'hbb == _T_22[7:0]) begin
        image_2_187 <= io_pixelVal_in_2_2;
      end else if (8'hbb == _T_19[7:0]) begin
        image_2_187 <= io_pixelVal_in_2_1;
      end else if (8'hbb == _T_15[7:0]) begin
        image_2_187 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_188 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbc == _T_37[7:0]) begin
        image_2_188 <= io_pixelVal_in_2_7;
      end else if (8'hbc == _T_34[7:0]) begin
        image_2_188 <= io_pixelVal_in_2_6;
      end else if (8'hbc == _T_31[7:0]) begin
        image_2_188 <= io_pixelVal_in_2_5;
      end else if (8'hbc == _T_28[7:0]) begin
        image_2_188 <= io_pixelVal_in_2_4;
      end else if (8'hbc == _T_25[7:0]) begin
        image_2_188 <= io_pixelVal_in_2_3;
      end else if (8'hbc == _T_22[7:0]) begin
        image_2_188 <= io_pixelVal_in_2_2;
      end else if (8'hbc == _T_19[7:0]) begin
        image_2_188 <= io_pixelVal_in_2_1;
      end else if (8'hbc == _T_15[7:0]) begin
        image_2_188 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_189 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbd == _T_37[7:0]) begin
        image_2_189 <= io_pixelVal_in_2_7;
      end else if (8'hbd == _T_34[7:0]) begin
        image_2_189 <= io_pixelVal_in_2_6;
      end else if (8'hbd == _T_31[7:0]) begin
        image_2_189 <= io_pixelVal_in_2_5;
      end else if (8'hbd == _T_28[7:0]) begin
        image_2_189 <= io_pixelVal_in_2_4;
      end else if (8'hbd == _T_25[7:0]) begin
        image_2_189 <= io_pixelVal_in_2_3;
      end else if (8'hbd == _T_22[7:0]) begin
        image_2_189 <= io_pixelVal_in_2_2;
      end else if (8'hbd == _T_19[7:0]) begin
        image_2_189 <= io_pixelVal_in_2_1;
      end else if (8'hbd == _T_15[7:0]) begin
        image_2_189 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_190 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbe == _T_37[7:0]) begin
        image_2_190 <= io_pixelVal_in_2_7;
      end else if (8'hbe == _T_34[7:0]) begin
        image_2_190 <= io_pixelVal_in_2_6;
      end else if (8'hbe == _T_31[7:0]) begin
        image_2_190 <= io_pixelVal_in_2_5;
      end else if (8'hbe == _T_28[7:0]) begin
        image_2_190 <= io_pixelVal_in_2_4;
      end else if (8'hbe == _T_25[7:0]) begin
        image_2_190 <= io_pixelVal_in_2_3;
      end else if (8'hbe == _T_22[7:0]) begin
        image_2_190 <= io_pixelVal_in_2_2;
      end else if (8'hbe == _T_19[7:0]) begin
        image_2_190 <= io_pixelVal_in_2_1;
      end else if (8'hbe == _T_15[7:0]) begin
        image_2_190 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_191 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbf == _T_37[7:0]) begin
        image_2_191 <= io_pixelVal_in_2_7;
      end else if (8'hbf == _T_34[7:0]) begin
        image_2_191 <= io_pixelVal_in_2_6;
      end else if (8'hbf == _T_31[7:0]) begin
        image_2_191 <= io_pixelVal_in_2_5;
      end else if (8'hbf == _T_28[7:0]) begin
        image_2_191 <= io_pixelVal_in_2_4;
      end else if (8'hbf == _T_25[7:0]) begin
        image_2_191 <= io_pixelVal_in_2_3;
      end else if (8'hbf == _T_22[7:0]) begin
        image_2_191 <= io_pixelVal_in_2_2;
      end else if (8'hbf == _T_19[7:0]) begin
        image_2_191 <= io_pixelVal_in_2_1;
      end else if (8'hbf == _T_15[7:0]) begin
        image_2_191 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      pixelIndex <= 32'h0;
    end else if (io_valid_in) begin
      if (_T_90) begin
        pixelIndex <= 32'h0;
      end else begin
        pixelIndex <= _T_88;
      end
    end
  end
endmodule
module ImageProcessing(
  input         clock,
  input         reset,
  input  [5:0]  io_SPI_filterIndex,
  input         io_SPI_invert,
  input         io_SPI_distort,
  input  [10:0] io_rowIndex,
  input  [10:0] io_colIndex,
  output [3:0]  io_pixelVal_out_0,
  output [3:0]  io_pixelVal_out_1,
  output [3:0]  io_pixelVal_out_2
);
  wire  filter_clock; // @[ImageProcessing.scala 23:22]
  wire  filter_reset; // @[ImageProcessing.scala 23:22]
  wire [5:0] filter_io_SPI_filterIndex; // @[ImageProcessing.scala 23:22]
  wire  filter_io_SPI_distort; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_0; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_1; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_2; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_3; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_4; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_5; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_6; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_7; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_0; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_1; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_2; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_3; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_4; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_5; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_6; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_7; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_0; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_1; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_2; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_3; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_4; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_5; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_6; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_7; // @[ImageProcessing.scala 23:22]
  wire  filter_io_valid_out; // @[ImageProcessing.scala 23:22]
  wire  videoBuffer_clock; // @[ImageProcessing.scala 24:27]
  wire  videoBuffer_reset; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_0; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_1; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_2; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_3; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_4; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_5; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_6; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_7; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_0; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_1; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_2; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_3; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_4; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_5; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_6; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_7; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_0; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_1; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_2; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_3; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_4; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_5; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_6; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_7; // @[ImageProcessing.scala 24:27]
  wire  videoBuffer_io_valid_in; // @[ImageProcessing.scala 24:27]
  wire [10:0] videoBuffer_io_rowIndex; // @[ImageProcessing.scala 24:27]
  wire [10:0] videoBuffer_io_colIndex; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_out_0; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_out_1; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_out_2; // @[ImageProcessing.scala 24:27]
  Filter filter ( // @[ImageProcessing.scala 23:22]
    .clock(filter_clock),
    .reset(filter_reset),
    .io_SPI_filterIndex(filter_io_SPI_filterIndex),
    .io_SPI_distort(filter_io_SPI_distort),
    .io_pixelVal_out_0_0(filter_io_pixelVal_out_0_0),
    .io_pixelVal_out_0_1(filter_io_pixelVal_out_0_1),
    .io_pixelVal_out_0_2(filter_io_pixelVal_out_0_2),
    .io_pixelVal_out_0_3(filter_io_pixelVal_out_0_3),
    .io_pixelVal_out_0_4(filter_io_pixelVal_out_0_4),
    .io_pixelVal_out_0_5(filter_io_pixelVal_out_0_5),
    .io_pixelVal_out_0_6(filter_io_pixelVal_out_0_6),
    .io_pixelVal_out_0_7(filter_io_pixelVal_out_0_7),
    .io_pixelVal_out_1_0(filter_io_pixelVal_out_1_0),
    .io_pixelVal_out_1_1(filter_io_pixelVal_out_1_1),
    .io_pixelVal_out_1_2(filter_io_pixelVal_out_1_2),
    .io_pixelVal_out_1_3(filter_io_pixelVal_out_1_3),
    .io_pixelVal_out_1_4(filter_io_pixelVal_out_1_4),
    .io_pixelVal_out_1_5(filter_io_pixelVal_out_1_5),
    .io_pixelVal_out_1_6(filter_io_pixelVal_out_1_6),
    .io_pixelVal_out_1_7(filter_io_pixelVal_out_1_7),
    .io_pixelVal_out_2_0(filter_io_pixelVal_out_2_0),
    .io_pixelVal_out_2_1(filter_io_pixelVal_out_2_1),
    .io_pixelVal_out_2_2(filter_io_pixelVal_out_2_2),
    .io_pixelVal_out_2_3(filter_io_pixelVal_out_2_3),
    .io_pixelVal_out_2_4(filter_io_pixelVal_out_2_4),
    .io_pixelVal_out_2_5(filter_io_pixelVal_out_2_5),
    .io_pixelVal_out_2_6(filter_io_pixelVal_out_2_6),
    .io_pixelVal_out_2_7(filter_io_pixelVal_out_2_7),
    .io_valid_out(filter_io_valid_out)
  );
  VideoBuffer videoBuffer ( // @[ImageProcessing.scala 24:27]
    .clock(videoBuffer_clock),
    .reset(videoBuffer_reset),
    .io_pixelVal_in_0_0(videoBuffer_io_pixelVal_in_0_0),
    .io_pixelVal_in_0_1(videoBuffer_io_pixelVal_in_0_1),
    .io_pixelVal_in_0_2(videoBuffer_io_pixelVal_in_0_2),
    .io_pixelVal_in_0_3(videoBuffer_io_pixelVal_in_0_3),
    .io_pixelVal_in_0_4(videoBuffer_io_pixelVal_in_0_4),
    .io_pixelVal_in_0_5(videoBuffer_io_pixelVal_in_0_5),
    .io_pixelVal_in_0_6(videoBuffer_io_pixelVal_in_0_6),
    .io_pixelVal_in_0_7(videoBuffer_io_pixelVal_in_0_7),
    .io_pixelVal_in_1_0(videoBuffer_io_pixelVal_in_1_0),
    .io_pixelVal_in_1_1(videoBuffer_io_pixelVal_in_1_1),
    .io_pixelVal_in_1_2(videoBuffer_io_pixelVal_in_1_2),
    .io_pixelVal_in_1_3(videoBuffer_io_pixelVal_in_1_3),
    .io_pixelVal_in_1_4(videoBuffer_io_pixelVal_in_1_4),
    .io_pixelVal_in_1_5(videoBuffer_io_pixelVal_in_1_5),
    .io_pixelVal_in_1_6(videoBuffer_io_pixelVal_in_1_6),
    .io_pixelVal_in_1_7(videoBuffer_io_pixelVal_in_1_7),
    .io_pixelVal_in_2_0(videoBuffer_io_pixelVal_in_2_0),
    .io_pixelVal_in_2_1(videoBuffer_io_pixelVal_in_2_1),
    .io_pixelVal_in_2_2(videoBuffer_io_pixelVal_in_2_2),
    .io_pixelVal_in_2_3(videoBuffer_io_pixelVal_in_2_3),
    .io_pixelVal_in_2_4(videoBuffer_io_pixelVal_in_2_4),
    .io_pixelVal_in_2_5(videoBuffer_io_pixelVal_in_2_5),
    .io_pixelVal_in_2_6(videoBuffer_io_pixelVal_in_2_6),
    .io_pixelVal_in_2_7(videoBuffer_io_pixelVal_in_2_7),
    .io_valid_in(videoBuffer_io_valid_in),
    .io_rowIndex(videoBuffer_io_rowIndex),
    .io_colIndex(videoBuffer_io_colIndex),
    .io_pixelVal_out_0(videoBuffer_io_pixelVal_out_0),
    .io_pixelVal_out_1(videoBuffer_io_pixelVal_out_1),
    .io_pixelVal_out_2(videoBuffer_io_pixelVal_out_2)
  );
  assign io_pixelVal_out_0 = videoBuffer_io_pixelVal_out_0; // @[ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25]
  assign io_pixelVal_out_1 = videoBuffer_io_pixelVal_out_1; // @[ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25]
  assign io_pixelVal_out_2 = videoBuffer_io_pixelVal_out_2; // @[ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25]
  assign filter_clock = clock;
  assign filter_reset = reset;
  assign filter_io_SPI_filterIndex = io_SPI_filterIndex; // @[ImageProcessing.scala 29:29]
  assign filter_io_SPI_distort = io_SPI_distort; // @[ImageProcessing.scala 31:29]
  assign videoBuffer_clock = clock;
  assign videoBuffer_reset = reset;
  assign videoBuffer_io_pixelVal_in_0_0 = filter_io_pixelVal_out_0_0; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_1 = filter_io_pixelVal_out_0_1; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_2 = filter_io_pixelVal_out_0_2; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_3 = filter_io_pixelVal_out_0_3; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_4 = filter_io_pixelVal_out_0_4; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_5 = filter_io_pixelVal_out_0_5; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_6 = filter_io_pixelVal_out_0_6; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_7 = filter_io_pixelVal_out_0_7; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_0 = filter_io_pixelVal_out_1_0; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_1 = filter_io_pixelVal_out_1_1; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_2 = filter_io_pixelVal_out_1_2; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_3 = filter_io_pixelVal_out_1_3; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_4 = filter_io_pixelVal_out_1_4; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_5 = filter_io_pixelVal_out_1_5; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_6 = filter_io_pixelVal_out_1_6; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_7 = filter_io_pixelVal_out_1_7; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_0 = filter_io_pixelVal_out_2_0; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_1 = filter_io_pixelVal_out_2_1; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_2 = filter_io_pixelVal_out_2_2; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_3 = filter_io_pixelVal_out_2_3; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_4 = filter_io_pixelVal_out_2_4; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_5 = filter_io_pixelVal_out_2_5; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_6 = filter_io_pixelVal_out_2_6; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_7 = filter_io_pixelVal_out_2_7; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_valid_in = filter_io_valid_out; // @[ImageProcessing.scala 39:27]
  assign videoBuffer_io_rowIndex = io_rowIndex; // @[ImageProcessing.scala 26:27]
  assign videoBuffer_io_colIndex = io_colIndex; // @[ImageProcessing.scala 27:27]
endmodule
