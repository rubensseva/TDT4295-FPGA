module DotProd(
  input        clock,
  input        reset,
  input  [7:0] io_dataInA,
  input  [7:0] io_dataInB,
  output [8:0] io_dataOut,
  output       io_outputValid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] countVal; // @[Counter.scala 29:33]
  wire  countReset = countVal == 4'h8; // @[Counter.scala 38:24]
  wire [3:0] _T_2 = countVal + 4'h1; // @[Counter.scala 39:22]
  reg [8:0] accumulator; // @[DotProd.scala 19:28]
  wire [15:0] product = $signed(io_dataInA) * $signed(io_dataInB); // @[DotProd.scala 20:35]
  wire [15:0] _GEN_5 = {{7{accumulator[8]}},accumulator}; // @[DotProd.scala 21:30]
  wire [15:0] _T_6 = $signed(_GEN_5) + $signed(product); // @[DotProd.scala 21:30]
  wire [15:0] _GEN_4 = countReset ? $signed(16'sh0) : $signed(_T_6); // @[DotProd.scala 25:20]
  assign io_dataOut = _T_6[8:0]; // @[DotProd.scala 23:14]
  assign io_outputValid = countVal == 4'h8; // @[DotProd.scala 26:20 DotProd.scala 29:20]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  countVal = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  accumulator = _RAND_1[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      countVal <= 4'h0;
    end else if (countReset) begin
      countVal <= 4'h0;
    end else begin
      countVal <= _T_2;
    end
    if (reset) begin
      accumulator <= 9'sh0;
    end else begin
      accumulator <= _GEN_4[8:0];
    end
  end
endmodule
module KernelConvolution(
  input        clock,
  input        reset,
  input  [4:0] io_kernelVal_in,
  input  [3:0] io_pixelVal_in_0,
  input  [3:0] io_pixelVal_in_1,
  input  [3:0] io_pixelVal_in_2,
  input  [3:0] io_pixelVal_in_3,
  input  [3:0] io_pixelVal_in_4,
  input  [3:0] io_pixelVal_in_5,
  input  [3:0] io_pixelVal_in_6,
  input  [3:0] io_pixelVal_in_7,
  output [8:0] io_pixelVal_out_0,
  output [8:0] io_pixelVal_out_1,
  output [8:0] io_pixelVal_out_2,
  output [8:0] io_pixelVal_out_3,
  output [8:0] io_pixelVal_out_4,
  output [8:0] io_pixelVal_out_5,
  output [8:0] io_pixelVal_out_6,
  output [8:0] io_pixelVal_out_7,
  output       io_valid_out
);
  wire  DotProd_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_1_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_1_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_1_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_1_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_1_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_1_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_2_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_2_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_2_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_2_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_2_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_2_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_3_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_3_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_3_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_3_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_3_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_3_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_4_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_4_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_4_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_4_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_4_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_4_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_5_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_5_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_5_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_5_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_5_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_5_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_6_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_6_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_6_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_6_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_6_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_6_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_7_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_7_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_7_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_7_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_7_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_7_io_outputValid; // @[KernelConvolution.scala 21:58]
  DotProd DotProd ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_clock),
    .reset(DotProd_reset),
    .io_dataInA(DotProd_io_dataInA),
    .io_dataInB(DotProd_io_dataInB),
    .io_dataOut(DotProd_io_dataOut),
    .io_outputValid(DotProd_io_outputValid)
  );
  DotProd DotProd_1 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_1_clock),
    .reset(DotProd_1_reset),
    .io_dataInA(DotProd_1_io_dataInA),
    .io_dataInB(DotProd_1_io_dataInB),
    .io_dataOut(DotProd_1_io_dataOut),
    .io_outputValid(DotProd_1_io_outputValid)
  );
  DotProd DotProd_2 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_2_clock),
    .reset(DotProd_2_reset),
    .io_dataInA(DotProd_2_io_dataInA),
    .io_dataInB(DotProd_2_io_dataInB),
    .io_dataOut(DotProd_2_io_dataOut),
    .io_outputValid(DotProd_2_io_outputValid)
  );
  DotProd DotProd_3 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_3_clock),
    .reset(DotProd_3_reset),
    .io_dataInA(DotProd_3_io_dataInA),
    .io_dataInB(DotProd_3_io_dataInB),
    .io_dataOut(DotProd_3_io_dataOut),
    .io_outputValid(DotProd_3_io_outputValid)
  );
  DotProd DotProd_4 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_4_clock),
    .reset(DotProd_4_reset),
    .io_dataInA(DotProd_4_io_dataInA),
    .io_dataInB(DotProd_4_io_dataInB),
    .io_dataOut(DotProd_4_io_dataOut),
    .io_outputValid(DotProd_4_io_outputValid)
  );
  DotProd DotProd_5 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_5_clock),
    .reset(DotProd_5_reset),
    .io_dataInA(DotProd_5_io_dataInA),
    .io_dataInB(DotProd_5_io_dataInB),
    .io_dataOut(DotProd_5_io_dataOut),
    .io_outputValid(DotProd_5_io_outputValid)
  );
  DotProd DotProd_6 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_6_clock),
    .reset(DotProd_6_reset),
    .io_dataInA(DotProd_6_io_dataInA),
    .io_dataInB(DotProd_6_io_dataInB),
    .io_dataOut(DotProd_6_io_dataOut),
    .io_outputValid(DotProd_6_io_outputValid)
  );
  DotProd DotProd_7 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_7_clock),
    .reset(DotProd_7_reset),
    .io_dataInA(DotProd_7_io_dataInA),
    .io_dataInB(DotProd_7_io_dataInB),
    .io_dataOut(DotProd_7_io_dataOut),
    .io_outputValid(DotProd_7_io_outputValid)
  );
  assign io_pixelVal_out_0 = DotProd_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_1 = DotProd_1_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_2 = DotProd_2_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_3 = DotProd_3_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_4 = DotProd_4_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_5 = DotProd_5_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_6 = DotProd_6_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_7 = DotProd_7_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_valid_out = DotProd_io_outputValid; // @[KernelConvolution.scala 35:30]
  assign DotProd_clock = clock;
  assign DotProd_reset = reset;
  assign DotProd_io_dataInA = {{4'd0}, io_pixelVal_in_0}; // @[KernelConvolution.scala 21:32]
  assign DotProd_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_1_clock = clock;
  assign DotProd_1_reset = reset;
  assign DotProd_1_io_dataInA = {{4'd0}, io_pixelVal_in_1}; // @[KernelConvolution.scala 21:32]
  assign DotProd_1_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_2_clock = clock;
  assign DotProd_2_reset = reset;
  assign DotProd_2_io_dataInA = {{4'd0}, io_pixelVal_in_2}; // @[KernelConvolution.scala 21:32]
  assign DotProd_2_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_3_clock = clock;
  assign DotProd_3_reset = reset;
  assign DotProd_3_io_dataInA = {{4'd0}, io_pixelVal_in_3}; // @[KernelConvolution.scala 21:32]
  assign DotProd_3_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_4_clock = clock;
  assign DotProd_4_reset = reset;
  assign DotProd_4_io_dataInA = {{4'd0}, io_pixelVal_in_4}; // @[KernelConvolution.scala 21:32]
  assign DotProd_4_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_5_clock = clock;
  assign DotProd_5_reset = reset;
  assign DotProd_5_io_dataInA = {{4'd0}, io_pixelVal_in_5}; // @[KernelConvolution.scala 21:32]
  assign DotProd_5_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_6_clock = clock;
  assign DotProd_6_reset = reset;
  assign DotProd_6_io_dataInA = {{4'd0}, io_pixelVal_in_6}; // @[KernelConvolution.scala 21:32]
  assign DotProd_6_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_7_clock = clock;
  assign DotProd_7_reset = reset;
  assign DotProd_7_io_dataInA = {{4'd0}, io_pixelVal_in_7}; // @[KernelConvolution.scala 21:32]
  assign DotProd_7_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
endmodule
module Filter(
  input        clock,
  input        reset,
  input  [5:0] io_SPI_filterIndex,
  input        io_SPI_distort,
  output [3:0] io_pixelVal_out_0_0,
  output [3:0] io_pixelVal_out_0_1,
  output [3:0] io_pixelVal_out_0_2,
  output [3:0] io_pixelVal_out_0_3,
  output [3:0] io_pixelVal_out_0_4,
  output [3:0] io_pixelVal_out_0_5,
  output [3:0] io_pixelVal_out_0_6,
  output [3:0] io_pixelVal_out_0_7,
  output [3:0] io_pixelVal_out_1_0,
  output [3:0] io_pixelVal_out_1_1,
  output [3:0] io_pixelVal_out_1_2,
  output [3:0] io_pixelVal_out_1_3,
  output [3:0] io_pixelVal_out_1_4,
  output [3:0] io_pixelVal_out_1_5,
  output [3:0] io_pixelVal_out_1_6,
  output [3:0] io_pixelVal_out_1_7,
  output [3:0] io_pixelVal_out_2_0,
  output [3:0] io_pixelVal_out_2_1,
  output [3:0] io_pixelVal_out_2_2,
  output [3:0] io_pixelVal_out_2_3,
  output [3:0] io_pixelVal_out_2_4,
  output [3:0] io_pixelVal_out_2_5,
  output [3:0] io_pixelVal_out_2_6,
  output [3:0] io_pixelVal_out_2_7,
  output       io_valid_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
`endif // RANDOMIZE_REG_INIT
  wire  KernelConvolution_clock; // @[Filter.scala 212:36]
  wire  KernelConvolution_reset; // @[Filter.scala 212:36]
  wire [4:0] KernelConvolution_io_kernelVal_in; // @[Filter.scala 212:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_0; // @[Filter.scala 212:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_1; // @[Filter.scala 212:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_2; // @[Filter.scala 212:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_3; // @[Filter.scala 212:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_4; // @[Filter.scala 212:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_5; // @[Filter.scala 212:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_6; // @[Filter.scala 212:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_7; // @[Filter.scala 212:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_0; // @[Filter.scala 212:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_1; // @[Filter.scala 212:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_2; // @[Filter.scala 212:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_3; // @[Filter.scala 212:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_4; // @[Filter.scala 212:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_5; // @[Filter.scala 212:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_6; // @[Filter.scala 212:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_7; // @[Filter.scala 212:36]
  wire  KernelConvolution_io_valid_out; // @[Filter.scala 212:36]
  wire  KernelConvolution_1_clock; // @[Filter.scala 213:36]
  wire  KernelConvolution_1_reset; // @[Filter.scala 213:36]
  wire [4:0] KernelConvolution_1_io_kernelVal_in; // @[Filter.scala 213:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_0; // @[Filter.scala 213:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_1; // @[Filter.scala 213:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_2; // @[Filter.scala 213:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_3; // @[Filter.scala 213:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_4; // @[Filter.scala 213:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_5; // @[Filter.scala 213:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_6; // @[Filter.scala 213:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_7; // @[Filter.scala 213:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_0; // @[Filter.scala 213:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_1; // @[Filter.scala 213:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_2; // @[Filter.scala 213:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_3; // @[Filter.scala 213:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_4; // @[Filter.scala 213:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_5; // @[Filter.scala 213:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_6; // @[Filter.scala 213:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_7; // @[Filter.scala 213:36]
  wire  KernelConvolution_1_io_valid_out; // @[Filter.scala 213:36]
  wire  KernelConvolution_2_clock; // @[Filter.scala 214:36]
  wire  KernelConvolution_2_reset; // @[Filter.scala 214:36]
  wire [4:0] KernelConvolution_2_io_kernelVal_in; // @[Filter.scala 214:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_0; // @[Filter.scala 214:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_1; // @[Filter.scala 214:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_2; // @[Filter.scala 214:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_3; // @[Filter.scala 214:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_4; // @[Filter.scala 214:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_5; // @[Filter.scala 214:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_6; // @[Filter.scala 214:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_7; // @[Filter.scala 214:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_0; // @[Filter.scala 214:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_1; // @[Filter.scala 214:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_2; // @[Filter.scala 214:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_3; // @[Filter.scala 214:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_4; // @[Filter.scala 214:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_5; // @[Filter.scala 214:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_6; // @[Filter.scala 214:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_7; // @[Filter.scala 214:36]
  wire  KernelConvolution_2_io_valid_out; // @[Filter.scala 214:36]
  reg [3:0] kernelCounter; // @[Counter.scala 29:33]
  wire  kernelCountReset = kernelCounter == 4'h8; // @[Counter.scala 38:24]
  wire [3:0] _T_14 = kernelCounter + 4'h1; // @[Counter.scala 39:22]
  wire  _GEN_38651 = 3'h0 == io_SPI_filterIndex[2:0]; // @[Filter.scala 220:41]
  wire  _GEN_38652 = 4'h4 == kernelCounter; // @[Filter.scala 220:41]
  wire [4:0] _GEN_7 = _GEN_38651 & _GEN_38652 ? $signed(5'sh1) : $signed(5'sh0); // @[Filter.scala 220:41]
  wire  _GEN_38654 = 4'h5 == kernelCounter; // @[Filter.scala 220:41]
  wire [4:0] _GEN_8 = _GEN_38651 & _GEN_38654 ? $signed(5'sh0) : $signed(_GEN_7); // @[Filter.scala 220:41]
  wire  _GEN_38656 = 4'h6 == kernelCounter; // @[Filter.scala 220:41]
  wire [4:0] _GEN_9 = _GEN_38651 & _GEN_38656 ? $signed(5'sh0) : $signed(_GEN_8); // @[Filter.scala 220:41]
  wire  _GEN_38658 = 4'h7 == kernelCounter; // @[Filter.scala 220:41]
  wire [4:0] _GEN_10 = _GEN_38651 & _GEN_38658 ? $signed(5'sh0) : $signed(_GEN_9); // @[Filter.scala 220:41]
  wire  _GEN_38660 = 4'h8 == kernelCounter; // @[Filter.scala 220:41]
  wire [4:0] _GEN_11 = _GEN_38651 & _GEN_38660 ? $signed(5'sh0) : $signed(_GEN_10); // @[Filter.scala 220:41]
  wire  _GEN_38661 = 3'h1 == io_SPI_filterIndex[2:0]; // @[Filter.scala 220:41]
  wire  _GEN_38662 = 4'h0 == kernelCounter; // @[Filter.scala 220:41]
  wire [4:0] _GEN_12 = _GEN_38661 & _GEN_38662 ? $signed(5'sh1) : $signed(_GEN_11); // @[Filter.scala 220:41]
  wire  _GEN_38664 = 4'h1 == kernelCounter; // @[Filter.scala 220:41]
  wire [4:0] _GEN_13 = _GEN_38661 & _GEN_38664 ? $signed(5'sh1) : $signed(_GEN_12); // @[Filter.scala 220:41]
  wire  _GEN_38666 = 4'h2 == kernelCounter; // @[Filter.scala 220:41]
  wire [4:0] _GEN_14 = _GEN_38661 & _GEN_38666 ? $signed(5'sh1) : $signed(_GEN_13); // @[Filter.scala 220:41]
  wire  _GEN_38668 = 4'h3 == kernelCounter; // @[Filter.scala 220:41]
  wire [4:0] _GEN_15 = _GEN_38661 & _GEN_38668 ? $signed(5'sh1) : $signed(_GEN_14); // @[Filter.scala 220:41]
  wire [4:0] _GEN_16 = _GEN_38661 & _GEN_38652 ? $signed(5'sh1) : $signed(_GEN_15); // @[Filter.scala 220:41]
  wire [4:0] _GEN_17 = _GEN_38661 & _GEN_38654 ? $signed(5'sh1) : $signed(_GEN_16); // @[Filter.scala 220:41]
  wire [4:0] _GEN_18 = _GEN_38661 & _GEN_38656 ? $signed(5'sh1) : $signed(_GEN_17); // @[Filter.scala 220:41]
  wire [4:0] _GEN_19 = _GEN_38661 & _GEN_38658 ? $signed(5'sh1) : $signed(_GEN_18); // @[Filter.scala 220:41]
  wire [4:0] _GEN_20 = _GEN_38661 & _GEN_38660 ? $signed(5'sh1) : $signed(_GEN_19); // @[Filter.scala 220:41]
  wire  _GEN_38679 = 3'h2 == io_SPI_filterIndex[2:0]; // @[Filter.scala 220:41]
  wire [4:0] _GEN_21 = _GEN_38679 & _GEN_38662 ? $signed(5'sh1) : $signed(_GEN_20); // @[Filter.scala 220:41]
  wire [4:0] _GEN_22 = _GEN_38679 & _GEN_38664 ? $signed(5'sh2) : $signed(_GEN_21); // @[Filter.scala 220:41]
  wire [4:0] _GEN_23 = _GEN_38679 & _GEN_38666 ? $signed(5'sh1) : $signed(_GEN_22); // @[Filter.scala 220:41]
  wire [4:0] _GEN_24 = _GEN_38679 & _GEN_38668 ? $signed(5'sh2) : $signed(_GEN_23); // @[Filter.scala 220:41]
  wire [4:0] _GEN_25 = _GEN_38679 & _GEN_38652 ? $signed(5'sh4) : $signed(_GEN_24); // @[Filter.scala 220:41]
  wire [4:0] _GEN_26 = _GEN_38679 & _GEN_38654 ? $signed(5'sh2) : $signed(_GEN_25); // @[Filter.scala 220:41]
  wire [4:0] _GEN_27 = _GEN_38679 & _GEN_38656 ? $signed(5'sh1) : $signed(_GEN_26); // @[Filter.scala 220:41]
  wire [4:0] _GEN_28 = _GEN_38679 & _GEN_38658 ? $signed(5'sh2) : $signed(_GEN_27); // @[Filter.scala 220:41]
  wire [4:0] _GEN_29 = _GEN_38679 & _GEN_38660 ? $signed(5'sh1) : $signed(_GEN_28); // @[Filter.scala 220:41]
  wire  _GEN_38697 = 3'h3 == io_SPI_filterIndex[2:0]; // @[Filter.scala 220:41]
  wire [4:0] _GEN_30 = _GEN_38697 & _GEN_38662 ? $signed(5'sh0) : $signed(_GEN_29); // @[Filter.scala 220:41]
  wire [4:0] _GEN_31 = _GEN_38697 & _GEN_38664 ? $signed(-5'sh1) : $signed(_GEN_30); // @[Filter.scala 220:41]
  wire [4:0] _GEN_32 = _GEN_38697 & _GEN_38666 ? $signed(5'sh0) : $signed(_GEN_31); // @[Filter.scala 220:41]
  wire [4:0] _GEN_33 = _GEN_38697 & _GEN_38668 ? $signed(-5'sh1) : $signed(_GEN_32); // @[Filter.scala 220:41]
  wire [4:0] _GEN_34 = _GEN_38697 & _GEN_38652 ? $signed(5'sh4) : $signed(_GEN_33); // @[Filter.scala 220:41]
  wire [4:0] _GEN_35 = _GEN_38697 & _GEN_38654 ? $signed(-5'sh1) : $signed(_GEN_34); // @[Filter.scala 220:41]
  wire [4:0] _GEN_36 = _GEN_38697 & _GEN_38656 ? $signed(5'sh0) : $signed(_GEN_35); // @[Filter.scala 220:41]
  wire [4:0] _GEN_37 = _GEN_38697 & _GEN_38658 ? $signed(-5'sh1) : $signed(_GEN_36); // @[Filter.scala 220:41]
  wire [4:0] _GEN_38 = _GEN_38697 & _GEN_38660 ? $signed(5'sh0) : $signed(_GEN_37); // @[Filter.scala 220:41]
  wire  _GEN_38715 = 3'h4 == io_SPI_filterIndex[2:0]; // @[Filter.scala 220:41]
  wire [4:0] _GEN_39 = _GEN_38715 & _GEN_38662 ? $signed(-5'sh1) : $signed(_GEN_38); // @[Filter.scala 220:41]
  wire [4:0] _GEN_40 = _GEN_38715 & _GEN_38664 ? $signed(-5'sh1) : $signed(_GEN_39); // @[Filter.scala 220:41]
  wire [4:0] _GEN_41 = _GEN_38715 & _GEN_38666 ? $signed(-5'sh1) : $signed(_GEN_40); // @[Filter.scala 220:41]
  wire [4:0] _GEN_42 = _GEN_38715 & _GEN_38668 ? $signed(-5'sh1) : $signed(_GEN_41); // @[Filter.scala 220:41]
  wire [4:0] _GEN_43 = _GEN_38715 & _GEN_38652 ? $signed(5'sh8) : $signed(_GEN_42); // @[Filter.scala 220:41]
  wire [4:0] _GEN_44 = _GEN_38715 & _GEN_38654 ? $signed(-5'sh1) : $signed(_GEN_43); // @[Filter.scala 220:41]
  wire [4:0] _GEN_45 = _GEN_38715 & _GEN_38656 ? $signed(-5'sh1) : $signed(_GEN_44); // @[Filter.scala 220:41]
  wire [4:0] _GEN_46 = _GEN_38715 & _GEN_38658 ? $signed(-5'sh1) : $signed(_GEN_45); // @[Filter.scala 220:41]
  wire [4:0] _GEN_47 = _GEN_38715 & _GEN_38660 ? $signed(-5'sh1) : $signed(_GEN_46); // @[Filter.scala 220:41]
  wire  _GEN_38733 = 3'h5 == io_SPI_filterIndex[2:0]; // @[Filter.scala 220:41]
  wire [4:0] _GEN_48 = _GEN_38733 & _GEN_38662 ? $signed(5'sh0) : $signed(_GEN_47); // @[Filter.scala 220:41]
  wire [4:0] _GEN_49 = _GEN_38733 & _GEN_38664 ? $signed(-5'sh1) : $signed(_GEN_48); // @[Filter.scala 220:41]
  wire [4:0] _GEN_50 = _GEN_38733 & _GEN_38666 ? $signed(5'sh0) : $signed(_GEN_49); // @[Filter.scala 220:41]
  wire [4:0] _GEN_51 = _GEN_38733 & _GEN_38668 ? $signed(-5'sh1) : $signed(_GEN_50); // @[Filter.scala 220:41]
  wire [4:0] _GEN_52 = _GEN_38733 & _GEN_38652 ? $signed(5'sh5) : $signed(_GEN_51); // @[Filter.scala 220:41]
  wire [4:0] _GEN_53 = _GEN_38733 & _GEN_38654 ? $signed(-5'sh1) : $signed(_GEN_52); // @[Filter.scala 220:41]
  wire [4:0] _GEN_54 = _GEN_38733 & _GEN_38656 ? $signed(5'sh0) : $signed(_GEN_53); // @[Filter.scala 220:41]
  wire [4:0] _GEN_55 = _GEN_38733 & _GEN_38658 ? $signed(-5'sh1) : $signed(_GEN_54); // @[Filter.scala 220:41]
  reg [1:0] imageCounterX; // @[Counter.scala 29:33]
  wire  imageCounterXReset = imageCounterX == 2'h2; // @[Counter.scala 38:24]
  wire [1:0] _T_20 = imageCounterX + 2'h1; // @[Counter.scala 39:22]
  reg [1:0] imageCounterY; // @[Counter.scala 29:33]
  wire  _T_21 = imageCounterY == 2'h2; // @[Counter.scala 38:24]
  wire [1:0] _T_23 = imageCounterY + 2'h1; // @[Counter.scala 39:22]
  reg [31:0] pixelIndex; // @[Filter.scala 225:31]
  wire [32:0] _T_24 = {{1'd0}, pixelIndex}; // @[Filter.scala 228:31]
  wire [31:0] _GEN_0 = _T_24[31:0] % 32'h20; // @[Filter.scala 228:38]
  wire [5:0] _T_26 = _GEN_0[5:0]; // @[Filter.scala 228:38]
  wire [5:0] _GEN_38951 = {{4'd0}, imageCounterX}; // @[Filter.scala 228:53]
  wire [5:0] _T_28 = _T_26 + _GEN_38951; // @[Filter.scala 228:53]
  wire [5:0] _T_30 = _T_28 - 6'h1; // @[Filter.scala 228:69]
  wire [31:0] _T_33 = _T_24[31:0] / 32'h20; // @[Filter.scala 229:38]
  wire [31:0] _GEN_38952 = {{30'd0}, imageCounterY}; // @[Filter.scala 229:53]
  wire [31:0] _T_35 = _T_33 + _GEN_38952; // @[Filter.scala 229:53]
  wire [31:0] _T_37 = _T_35 - 32'h1; // @[Filter.scala 229:69]
  wire [37:0] _T_38 = _T_37 * 32'h20; // @[Filter.scala 230:42]
  wire [37:0] _GEN_38953 = {{32'd0}, _T_30}; // @[Filter.scala 230:57]
  wire [37:0] _T_40 = _T_38 + _GEN_38953; // @[Filter.scala 230:57]
  wire [3:0] _GEN_193 = 10'h16 == _T_40[9:0] ? 4'h9 : 4'ha; // @[Filter.scala 230:62]
  wire [3:0] _GEN_194 = 10'h17 == _T_40[9:0] ? 4'h3 : _GEN_193; // @[Filter.scala 230:62]
  wire [3:0] _GEN_195 = 10'h18 == _T_40[9:0] ? 4'h6 : _GEN_194; // @[Filter.scala 230:62]
  wire [3:0] _GEN_196 = 10'h19 == _T_40[9:0] ? 4'ha : _GEN_195; // @[Filter.scala 230:62]
  wire [3:0] _GEN_197 = 10'h1a == _T_40[9:0] ? 4'ha : _GEN_196; // @[Filter.scala 230:62]
  wire [3:0] _GEN_198 = 10'h1b == _T_40[9:0] ? 4'ha : _GEN_197; // @[Filter.scala 230:62]
  wire [3:0] _GEN_199 = 10'h1c == _T_40[9:0] ? 4'ha : _GEN_198; // @[Filter.scala 230:62]
  wire [3:0] _GEN_200 = 10'h1d == _T_40[9:0] ? 4'ha : _GEN_199; // @[Filter.scala 230:62]
  wire [3:0] _GEN_201 = 10'h1e == _T_40[9:0] ? 4'ha : _GEN_200; // @[Filter.scala 230:62]
  wire [3:0] _GEN_202 = 10'h1f == _T_40[9:0] ? 4'ha : _GEN_201; // @[Filter.scala 230:62]
  wire [3:0] _GEN_203 = 10'h20 == _T_40[9:0] ? 4'ha : _GEN_202; // @[Filter.scala 230:62]
  wire [3:0] _GEN_204 = 10'h21 == _T_40[9:0] ? 4'ha : _GEN_203; // @[Filter.scala 230:62]
  wire [3:0] _GEN_205 = 10'h22 == _T_40[9:0] ? 4'ha : _GEN_204; // @[Filter.scala 230:62]
  wire [3:0] _GEN_206 = 10'h23 == _T_40[9:0] ? 4'ha : _GEN_205; // @[Filter.scala 230:62]
  wire [3:0] _GEN_207 = 10'h24 == _T_40[9:0] ? 4'ha : _GEN_206; // @[Filter.scala 230:62]
  wire [3:0] _GEN_208 = 10'h25 == _T_40[9:0] ? 4'ha : _GEN_207; // @[Filter.scala 230:62]
  wire [3:0] _GEN_209 = 10'h26 == _T_40[9:0] ? 4'ha : _GEN_208; // @[Filter.scala 230:62]
  wire [3:0] _GEN_210 = 10'h27 == _T_40[9:0] ? 4'ha : _GEN_209; // @[Filter.scala 230:62]
  wire [3:0] _GEN_211 = 10'h28 == _T_40[9:0] ? 4'ha : _GEN_210; // @[Filter.scala 230:62]
  wire [3:0] _GEN_212 = 10'h29 == _T_40[9:0] ? 4'ha : _GEN_211; // @[Filter.scala 230:62]
  wire [3:0] _GEN_213 = 10'h2a == _T_40[9:0] ? 4'ha : _GEN_212; // @[Filter.scala 230:62]
  wire [3:0] _GEN_214 = 10'h2b == _T_40[9:0] ? 4'ha : _GEN_213; // @[Filter.scala 230:62]
  wire [3:0] _GEN_215 = 10'h2c == _T_40[9:0] ? 4'ha : _GEN_214; // @[Filter.scala 230:62]
  wire [3:0] _GEN_216 = 10'h2d == _T_40[9:0] ? 4'ha : _GEN_215; // @[Filter.scala 230:62]
  wire [3:0] _GEN_217 = 10'h2e == _T_40[9:0] ? 4'ha : _GEN_216; // @[Filter.scala 230:62]
  wire [3:0] _GEN_218 = 10'h2f == _T_40[9:0] ? 4'ha : _GEN_217; // @[Filter.scala 230:62]
  wire [3:0] _GEN_219 = 10'h30 == _T_40[9:0] ? 4'ha : _GEN_218; // @[Filter.scala 230:62]
  wire [3:0] _GEN_220 = 10'h31 == _T_40[9:0] ? 4'ha : _GEN_219; // @[Filter.scala 230:62]
  wire [3:0] _GEN_221 = 10'h32 == _T_40[9:0] ? 4'ha : _GEN_220; // @[Filter.scala 230:62]
  wire [3:0] _GEN_222 = 10'h33 == _T_40[9:0] ? 4'ha : _GEN_221; // @[Filter.scala 230:62]
  wire [3:0] _GEN_223 = 10'h34 == _T_40[9:0] ? 4'ha : _GEN_222; // @[Filter.scala 230:62]
  wire [3:0] _GEN_224 = 10'h35 == _T_40[9:0] ? 4'ha : _GEN_223; // @[Filter.scala 230:62]
  wire [3:0] _GEN_225 = 10'h36 == _T_40[9:0] ? 4'ha : _GEN_224; // @[Filter.scala 230:62]
  wire [3:0] _GEN_226 = 10'h37 == _T_40[9:0] ? 4'ha : _GEN_225; // @[Filter.scala 230:62]
  wire [3:0] _GEN_227 = 10'h38 == _T_40[9:0] ? 4'ha : _GEN_226; // @[Filter.scala 230:62]
  wire [3:0] _GEN_228 = 10'h39 == _T_40[9:0] ? 4'ha : _GEN_227; // @[Filter.scala 230:62]
  wire [3:0] _GEN_229 = 10'h3a == _T_40[9:0] ? 4'ha : _GEN_228; // @[Filter.scala 230:62]
  wire [3:0] _GEN_230 = 10'h3b == _T_40[9:0] ? 4'h9 : _GEN_229; // @[Filter.scala 230:62]
  wire [3:0] _GEN_231 = 10'h3c == _T_40[9:0] ? 4'h4 : _GEN_230; // @[Filter.scala 230:62]
  wire [3:0] _GEN_232 = 10'h3d == _T_40[9:0] ? 4'h3 : _GEN_231; // @[Filter.scala 230:62]
  wire [3:0] _GEN_233 = 10'h3e == _T_40[9:0] ? 4'h4 : _GEN_232; // @[Filter.scala 230:62]
  wire [3:0] _GEN_234 = 10'h3f == _T_40[9:0] ? 4'ha : _GEN_233; // @[Filter.scala 230:62]
  wire [3:0] _GEN_235 = 10'h40 == _T_40[9:0] ? 4'ha : _GEN_234; // @[Filter.scala 230:62]
  wire [3:0] _GEN_236 = 10'h41 == _T_40[9:0] ? 4'ha : _GEN_235; // @[Filter.scala 230:62]
  wire [3:0] _GEN_237 = 10'h42 == _T_40[9:0] ? 4'ha : _GEN_236; // @[Filter.scala 230:62]
  wire [3:0] _GEN_238 = 10'h43 == _T_40[9:0] ? 4'ha : _GEN_237; // @[Filter.scala 230:62]
  wire [3:0] _GEN_239 = 10'h44 == _T_40[9:0] ? 4'ha : _GEN_238; // @[Filter.scala 230:62]
  wire [3:0] _GEN_240 = 10'h45 == _T_40[9:0] ? 4'ha : _GEN_239; // @[Filter.scala 230:62]
  wire [3:0] _GEN_241 = 10'h46 == _T_40[9:0] ? 4'ha : _GEN_240; // @[Filter.scala 230:62]
  wire [3:0] _GEN_242 = 10'h47 == _T_40[9:0] ? 4'ha : _GEN_241; // @[Filter.scala 230:62]
  wire [3:0] _GEN_243 = 10'h48 == _T_40[9:0] ? 4'ha : _GEN_242; // @[Filter.scala 230:62]
  wire [3:0] _GEN_244 = 10'h49 == _T_40[9:0] ? 4'ha : _GEN_243; // @[Filter.scala 230:62]
  wire [3:0] _GEN_245 = 10'h4a == _T_40[9:0] ? 4'ha : _GEN_244; // @[Filter.scala 230:62]
  wire [3:0] _GEN_246 = 10'h4b == _T_40[9:0] ? 4'ha : _GEN_245; // @[Filter.scala 230:62]
  wire [3:0] _GEN_247 = 10'h4c == _T_40[9:0] ? 4'ha : _GEN_246; // @[Filter.scala 230:62]
  wire [3:0] _GEN_248 = 10'h4d == _T_40[9:0] ? 4'ha : _GEN_247; // @[Filter.scala 230:62]
  wire [3:0] _GEN_249 = 10'h4e == _T_40[9:0] ? 4'ha : _GEN_248; // @[Filter.scala 230:62]
  wire [3:0] _GEN_250 = 10'h4f == _T_40[9:0] ? 4'ha : _GEN_249; // @[Filter.scala 230:62]
  wire [3:0] _GEN_251 = 10'h50 == _T_40[9:0] ? 4'ha : _GEN_250; // @[Filter.scala 230:62]
  wire [3:0] _GEN_252 = 10'h51 == _T_40[9:0] ? 4'ha : _GEN_251; // @[Filter.scala 230:62]
  wire [3:0] _GEN_253 = 10'h52 == _T_40[9:0] ? 4'ha : _GEN_252; // @[Filter.scala 230:62]
  wire [3:0] _GEN_254 = 10'h53 == _T_40[9:0] ? 4'ha : _GEN_253; // @[Filter.scala 230:62]
  wire [3:0] _GEN_255 = 10'h54 == _T_40[9:0] ? 4'ha : _GEN_254; // @[Filter.scala 230:62]
  wire [3:0] _GEN_256 = 10'h55 == _T_40[9:0] ? 4'ha : _GEN_255; // @[Filter.scala 230:62]
  wire [3:0] _GEN_257 = 10'h56 == _T_40[9:0] ? 4'ha : _GEN_256; // @[Filter.scala 230:62]
  wire [3:0] _GEN_258 = 10'h57 == _T_40[9:0] ? 4'ha : _GEN_257; // @[Filter.scala 230:62]
  wire [3:0] _GEN_259 = 10'h58 == _T_40[9:0] ? 4'ha : _GEN_258; // @[Filter.scala 230:62]
  wire [3:0] _GEN_260 = 10'h59 == _T_40[9:0] ? 4'ha : _GEN_259; // @[Filter.scala 230:62]
  wire [3:0] _GEN_261 = 10'h5a == _T_40[9:0] ? 4'h7 : _GEN_260; // @[Filter.scala 230:62]
  wire [3:0] _GEN_262 = 10'h5b == _T_40[9:0] ? 4'h7 : _GEN_261; // @[Filter.scala 230:62]
  wire [3:0] _GEN_263 = 10'h5c == _T_40[9:0] ? 4'ha : _GEN_262; // @[Filter.scala 230:62]
  wire [3:0] _GEN_264 = 10'h5d == _T_40[9:0] ? 4'ha : _GEN_263; // @[Filter.scala 230:62]
  wire [3:0] _GEN_265 = 10'h5e == _T_40[9:0] ? 4'ha : _GEN_264; // @[Filter.scala 230:62]
  wire [3:0] _GEN_266 = 10'h5f == _T_40[9:0] ? 4'ha : _GEN_265; // @[Filter.scala 230:62]
  wire [3:0] _GEN_267 = 10'h60 == _T_40[9:0] ? 4'ha : _GEN_266; // @[Filter.scala 230:62]
  wire [3:0] _GEN_268 = 10'h61 == _T_40[9:0] ? 4'h8 : _GEN_267; // @[Filter.scala 230:62]
  wire [3:0] _GEN_269 = 10'h62 == _T_40[9:0] ? 4'h3 : _GEN_268; // @[Filter.scala 230:62]
  wire [3:0] _GEN_270 = 10'h63 == _T_40[9:0] ? 4'h3 : _GEN_269; // @[Filter.scala 230:62]
  wire [3:0] _GEN_271 = 10'h64 == _T_40[9:0] ? 4'h3 : _GEN_270; // @[Filter.scala 230:62]
  wire [3:0] _GEN_272 = 10'h65 == _T_40[9:0] ? 4'h9 : _GEN_271; // @[Filter.scala 230:62]
  wire [3:0] _GEN_273 = 10'h66 == _T_40[9:0] ? 4'ha : _GEN_272; // @[Filter.scala 230:62]
  wire [3:0] _GEN_274 = 10'h67 == _T_40[9:0] ? 4'ha : _GEN_273; // @[Filter.scala 230:62]
  wire [3:0] _GEN_275 = 10'h68 == _T_40[9:0] ? 4'ha : _GEN_274; // @[Filter.scala 230:62]
  wire [3:0] _GEN_276 = 10'h69 == _T_40[9:0] ? 4'ha : _GEN_275; // @[Filter.scala 230:62]
  wire [3:0] _GEN_277 = 10'h6a == _T_40[9:0] ? 4'ha : _GEN_276; // @[Filter.scala 230:62]
  wire [3:0] _GEN_278 = 10'h6b == _T_40[9:0] ? 4'h8 : _GEN_277; // @[Filter.scala 230:62]
  wire [3:0] _GEN_279 = 10'h6c == _T_40[9:0] ? 4'h5 : _GEN_278; // @[Filter.scala 230:62]
  wire [3:0] _GEN_280 = 10'h6d == _T_40[9:0] ? 4'h8 : _GEN_279; // @[Filter.scala 230:62]
  wire [3:0] _GEN_281 = 10'h6e == _T_40[9:0] ? 4'ha : _GEN_280; // @[Filter.scala 230:62]
  wire [3:0] _GEN_282 = 10'h6f == _T_40[9:0] ? 4'ha : _GEN_281; // @[Filter.scala 230:62]
  wire [3:0] _GEN_283 = 10'h70 == _T_40[9:0] ? 4'ha : _GEN_282; // @[Filter.scala 230:62]
  wire [3:0] _GEN_284 = 10'h71 == _T_40[9:0] ? 4'ha : _GEN_283; // @[Filter.scala 230:62]
  wire [3:0] _GEN_285 = 10'h72 == _T_40[9:0] ? 4'ha : _GEN_284; // @[Filter.scala 230:62]
  wire [3:0] _GEN_286 = 10'h73 == _T_40[9:0] ? 4'ha : _GEN_285; // @[Filter.scala 230:62]
  wire [3:0] _GEN_287 = 10'h74 == _T_40[9:0] ? 4'ha : _GEN_286; // @[Filter.scala 230:62]
  wire [3:0] _GEN_288 = 10'h75 == _T_40[9:0] ? 4'ha : _GEN_287; // @[Filter.scala 230:62]
  wire [3:0] _GEN_289 = 10'h76 == _T_40[9:0] ? 4'ha : _GEN_288; // @[Filter.scala 230:62]
  wire [3:0] _GEN_290 = 10'h77 == _T_40[9:0] ? 4'ha : _GEN_289; // @[Filter.scala 230:62]
  wire [3:0] _GEN_291 = 10'h78 == _T_40[9:0] ? 4'ha : _GEN_290; // @[Filter.scala 230:62]
  wire [3:0] _GEN_292 = 10'h79 == _T_40[9:0] ? 4'ha : _GEN_291; // @[Filter.scala 230:62]
  wire [3:0] _GEN_293 = 10'h7a == _T_40[9:0] ? 4'ha : _GEN_292; // @[Filter.scala 230:62]
  wire [3:0] _GEN_294 = 10'h7b == _T_40[9:0] ? 4'ha : _GEN_293; // @[Filter.scala 230:62]
  wire [3:0] _GEN_295 = 10'h7c == _T_40[9:0] ? 4'ha : _GEN_294; // @[Filter.scala 230:62]
  wire [3:0] _GEN_296 = 10'h7d == _T_40[9:0] ? 4'ha : _GEN_295; // @[Filter.scala 230:62]
  wire [3:0] _GEN_297 = 10'h7e == _T_40[9:0] ? 4'ha : _GEN_296; // @[Filter.scala 230:62]
  wire [3:0] _GEN_298 = 10'h7f == _T_40[9:0] ? 4'ha : _GEN_297; // @[Filter.scala 230:62]
  wire [3:0] _GEN_299 = 10'h80 == _T_40[9:0] ? 4'ha : _GEN_298; // @[Filter.scala 230:62]
  wire [3:0] _GEN_300 = 10'h81 == _T_40[9:0] ? 4'h5 : _GEN_299; // @[Filter.scala 230:62]
  wire [3:0] _GEN_301 = 10'h82 == _T_40[9:0] ? 4'h5 : _GEN_300; // @[Filter.scala 230:62]
  wire [3:0] _GEN_302 = 10'h83 == _T_40[9:0] ? 4'h7 : _GEN_301; // @[Filter.scala 230:62]
  wire [3:0] _GEN_303 = 10'h84 == _T_40[9:0] ? 4'ha : _GEN_302; // @[Filter.scala 230:62]
  wire [3:0] _GEN_304 = 10'h85 == _T_40[9:0] ? 4'ha : _GEN_303; // @[Filter.scala 230:62]
  wire [3:0] _GEN_305 = 10'h86 == _T_40[9:0] ? 4'ha : _GEN_304; // @[Filter.scala 230:62]
  wire [3:0] _GEN_306 = 10'h87 == _T_40[9:0] ? 4'h5 : _GEN_305; // @[Filter.scala 230:62]
  wire [3:0] _GEN_307 = 10'h88 == _T_40[9:0] ? 4'h3 : _GEN_306; // @[Filter.scala 230:62]
  wire [3:0] _GEN_308 = 10'h89 == _T_40[9:0] ? 4'h3 : _GEN_307; // @[Filter.scala 230:62]
  wire [3:0] _GEN_309 = 10'h8a == _T_40[9:0] ? 4'h4 : _GEN_308; // @[Filter.scala 230:62]
  wire [3:0] _GEN_310 = 10'h8b == _T_40[9:0] ? 4'h9 : _GEN_309; // @[Filter.scala 230:62]
  wire [3:0] _GEN_311 = 10'h8c == _T_40[9:0] ? 4'ha : _GEN_310; // @[Filter.scala 230:62]
  wire [3:0] _GEN_312 = 10'h8d == _T_40[9:0] ? 4'ha : _GEN_311; // @[Filter.scala 230:62]
  wire [3:0] _GEN_313 = 10'h8e == _T_40[9:0] ? 4'ha : _GEN_312; // @[Filter.scala 230:62]
  wire [3:0] _GEN_314 = 10'h8f == _T_40[9:0] ? 4'h6 : _GEN_313; // @[Filter.scala 230:62]
  wire [3:0] _GEN_315 = 10'h90 == _T_40[9:0] ? 4'h4 : _GEN_314; // @[Filter.scala 230:62]
  wire [3:0] _GEN_316 = 10'h91 == _T_40[9:0] ? 4'h3 : _GEN_315; // @[Filter.scala 230:62]
  wire [3:0] _GEN_317 = 10'h92 == _T_40[9:0] ? 4'h7 : _GEN_316; // @[Filter.scala 230:62]
  wire [3:0] _GEN_318 = 10'h93 == _T_40[9:0] ? 4'ha : _GEN_317; // @[Filter.scala 230:62]
  wire [3:0] _GEN_319 = 10'h94 == _T_40[9:0] ? 4'ha : _GEN_318; // @[Filter.scala 230:62]
  wire [3:0] _GEN_320 = 10'h95 == _T_40[9:0] ? 4'ha : _GEN_319; // @[Filter.scala 230:62]
  wire [3:0] _GEN_321 = 10'h96 == _T_40[9:0] ? 4'ha : _GEN_320; // @[Filter.scala 230:62]
  wire [3:0] _GEN_322 = 10'h97 == _T_40[9:0] ? 4'ha : _GEN_321; // @[Filter.scala 230:62]
  wire [3:0] _GEN_323 = 10'h98 == _T_40[9:0] ? 4'ha : _GEN_322; // @[Filter.scala 230:62]
  wire [3:0] _GEN_324 = 10'h99 == _T_40[9:0] ? 4'ha : _GEN_323; // @[Filter.scala 230:62]
  wire [3:0] _GEN_325 = 10'h9a == _T_40[9:0] ? 4'ha : _GEN_324; // @[Filter.scala 230:62]
  wire [3:0] _GEN_326 = 10'h9b == _T_40[9:0] ? 4'ha : _GEN_325; // @[Filter.scala 230:62]
  wire [3:0] _GEN_327 = 10'h9c == _T_40[9:0] ? 4'ha : _GEN_326; // @[Filter.scala 230:62]
  wire [3:0] _GEN_328 = 10'h9d == _T_40[9:0] ? 4'ha : _GEN_327; // @[Filter.scala 230:62]
  wire [3:0] _GEN_329 = 10'h9e == _T_40[9:0] ? 4'ha : _GEN_328; // @[Filter.scala 230:62]
  wire [3:0] _GEN_330 = 10'h9f == _T_40[9:0] ? 4'ha : _GEN_329; // @[Filter.scala 230:62]
  wire [3:0] _GEN_331 = 10'ha0 == _T_40[9:0] ? 4'ha : _GEN_330; // @[Filter.scala 230:62]
  wire [3:0] _GEN_332 = 10'ha1 == _T_40[9:0] ? 4'ha : _GEN_331; // @[Filter.scala 230:62]
  wire [3:0] _GEN_333 = 10'ha2 == _T_40[9:0] ? 4'ha : _GEN_332; // @[Filter.scala 230:62]
  wire [3:0] _GEN_334 = 10'ha3 == _T_40[9:0] ? 4'ha : _GEN_333; // @[Filter.scala 230:62]
  wire [3:0] _GEN_335 = 10'ha4 == _T_40[9:0] ? 4'ha : _GEN_334; // @[Filter.scala 230:62]
  wire [3:0] _GEN_336 = 10'ha5 == _T_40[9:0] ? 4'ha : _GEN_335; // @[Filter.scala 230:62]
  wire [3:0] _GEN_337 = 10'ha6 == _T_40[9:0] ? 4'ha : _GEN_336; // @[Filter.scala 230:62]
  wire [3:0] _GEN_338 = 10'ha7 == _T_40[9:0] ? 4'h9 : _GEN_337; // @[Filter.scala 230:62]
  wire [3:0] _GEN_339 = 10'ha8 == _T_40[9:0] ? 4'h4 : _GEN_338; // @[Filter.scala 230:62]
  wire [3:0] _GEN_340 = 10'ha9 == _T_40[9:0] ? 4'h3 : _GEN_339; // @[Filter.scala 230:62]
  wire [3:0] _GEN_341 = 10'haa == _T_40[9:0] ? 4'h4 : _GEN_340; // @[Filter.scala 230:62]
  wire [3:0] _GEN_342 = 10'hab == _T_40[9:0] ? 4'h7 : _GEN_341; // @[Filter.scala 230:62]
  wire [3:0] _GEN_343 = 10'hac == _T_40[9:0] ? 4'h8 : _GEN_342; // @[Filter.scala 230:62]
  wire [3:0] _GEN_344 = 10'had == _T_40[9:0] ? 4'h3 : _GEN_343; // @[Filter.scala 230:62]
  wire [3:0] _GEN_345 = 10'hae == _T_40[9:0] ? 4'h3 : _GEN_344; // @[Filter.scala 230:62]
  wire [3:0] _GEN_346 = 10'haf == _T_40[9:0] ? 4'h3 : _GEN_345; // @[Filter.scala 230:62]
  wire [3:0] _GEN_347 = 10'hb0 == _T_40[9:0] ? 4'h3 : _GEN_346; // @[Filter.scala 230:62]
  wire [3:0] _GEN_348 = 10'hb1 == _T_40[9:0] ? 4'h7 : _GEN_347; // @[Filter.scala 230:62]
  wire [3:0] _GEN_349 = 10'hb2 == _T_40[9:0] ? 4'h9 : _GEN_348; // @[Filter.scala 230:62]
  wire [3:0] _GEN_350 = 10'hb3 == _T_40[9:0] ? 4'h6 : _GEN_349; // @[Filter.scala 230:62]
  wire [3:0] _GEN_351 = 10'hb4 == _T_40[9:0] ? 4'h4 : _GEN_350; // @[Filter.scala 230:62]
  wire [3:0] _GEN_352 = 10'hb5 == _T_40[9:0] ? 4'h3 : _GEN_351; // @[Filter.scala 230:62]
  wire [3:0] _GEN_353 = 10'hb6 == _T_40[9:0] ? 4'h3 : _GEN_352; // @[Filter.scala 230:62]
  wire [3:0] _GEN_354 = 10'hb7 == _T_40[9:0] ? 4'h6 : _GEN_353; // @[Filter.scala 230:62]
  wire [3:0] _GEN_355 = 10'hb8 == _T_40[9:0] ? 4'ha : _GEN_354; // @[Filter.scala 230:62]
  wire [3:0] _GEN_356 = 10'hb9 == _T_40[9:0] ? 4'ha : _GEN_355; // @[Filter.scala 230:62]
  wire [3:0] _GEN_357 = 10'hba == _T_40[9:0] ? 4'ha : _GEN_356; // @[Filter.scala 230:62]
  wire [3:0] _GEN_358 = 10'hbb == _T_40[9:0] ? 4'ha : _GEN_357; // @[Filter.scala 230:62]
  wire [3:0] _GEN_359 = 10'hbc == _T_40[9:0] ? 4'ha : _GEN_358; // @[Filter.scala 230:62]
  wire [3:0] _GEN_360 = 10'hbd == _T_40[9:0] ? 4'h9 : _GEN_359; // @[Filter.scala 230:62]
  wire [3:0] _GEN_361 = 10'hbe == _T_40[9:0] ? 4'ha : _GEN_360; // @[Filter.scala 230:62]
  wire [3:0] _GEN_362 = 10'hbf == _T_40[9:0] ? 4'ha : _GEN_361; // @[Filter.scala 230:62]
  wire [3:0] _GEN_363 = 10'hc0 == _T_40[9:0] ? 4'ha : _GEN_362; // @[Filter.scala 230:62]
  wire [3:0] _GEN_364 = 10'hc1 == _T_40[9:0] ? 4'ha : _GEN_363; // @[Filter.scala 230:62]
  wire [3:0] _GEN_365 = 10'hc2 == _T_40[9:0] ? 4'ha : _GEN_364; // @[Filter.scala 230:62]
  wire [3:0] _GEN_366 = 10'hc3 == _T_40[9:0] ? 4'ha : _GEN_365; // @[Filter.scala 230:62]
  wire [3:0] _GEN_367 = 10'hc4 == _T_40[9:0] ? 4'ha : _GEN_366; // @[Filter.scala 230:62]
  wire [3:0] _GEN_368 = 10'hc5 == _T_40[9:0] ? 4'ha : _GEN_367; // @[Filter.scala 230:62]
  wire [3:0] _GEN_369 = 10'hc6 == _T_40[9:0] ? 4'ha : _GEN_368; // @[Filter.scala 230:62]
  wire [3:0] _GEN_370 = 10'hc7 == _T_40[9:0] ? 4'h9 : _GEN_369; // @[Filter.scala 230:62]
  wire [3:0] _GEN_371 = 10'hc8 == _T_40[9:0] ? 4'h8 : _GEN_370; // @[Filter.scala 230:62]
  wire [3:0] _GEN_372 = 10'hc9 == _T_40[9:0] ? 4'h8 : _GEN_371; // @[Filter.scala 230:62]
  wire [3:0] _GEN_373 = 10'hca == _T_40[9:0] ? 4'h9 : _GEN_372; // @[Filter.scala 230:62]
  wire [3:0] _GEN_374 = 10'hcb == _T_40[9:0] ? 4'ha : _GEN_373; // @[Filter.scala 230:62]
  wire [3:0] _GEN_375 = 10'hcc == _T_40[9:0] ? 4'ha : _GEN_374; // @[Filter.scala 230:62]
  wire [3:0] _GEN_376 = 10'hcd == _T_40[9:0] ? 4'ha : _GEN_375; // @[Filter.scala 230:62]
  wire [3:0] _GEN_377 = 10'hce == _T_40[9:0] ? 4'h8 : _GEN_376; // @[Filter.scala 230:62]
  wire [3:0] _GEN_378 = 10'hcf == _T_40[9:0] ? 4'h3 : _GEN_377; // @[Filter.scala 230:62]
  wire [3:0] _GEN_379 = 10'hd0 == _T_40[9:0] ? 4'h3 : _GEN_378; // @[Filter.scala 230:62]
  wire [3:0] _GEN_380 = 10'hd1 == _T_40[9:0] ? 4'h3 : _GEN_379; // @[Filter.scala 230:62]
  wire [3:0] _GEN_381 = 10'hd2 == _T_40[9:0] ? 4'h4 : _GEN_380; // @[Filter.scala 230:62]
  wire [3:0] _GEN_382 = 10'hd3 == _T_40[9:0] ? 4'h3 : _GEN_381; // @[Filter.scala 230:62]
  wire [3:0] _GEN_383 = 10'hd4 == _T_40[9:0] ? 4'h3 : _GEN_382; // @[Filter.scala 230:62]
  wire [3:0] _GEN_384 = 10'hd5 == _T_40[9:0] ? 4'h3 : _GEN_383; // @[Filter.scala 230:62]
  wire [3:0] _GEN_385 = 10'hd6 == _T_40[9:0] ? 4'h3 : _GEN_384; // @[Filter.scala 230:62]
  wire [3:0] _GEN_386 = 10'hd7 == _T_40[9:0] ? 4'h5 : _GEN_385; // @[Filter.scala 230:62]
  wire [3:0] _GEN_387 = 10'hd8 == _T_40[9:0] ? 4'h4 : _GEN_386; // @[Filter.scala 230:62]
  wire [3:0] _GEN_388 = 10'hd9 == _T_40[9:0] ? 4'h3 : _GEN_387; // @[Filter.scala 230:62]
  wire [3:0] _GEN_389 = 10'hda == _T_40[9:0] ? 4'h3 : _GEN_388; // @[Filter.scala 230:62]
  wire [3:0] _GEN_390 = 10'hdb == _T_40[9:0] ? 4'h3 : _GEN_389; // @[Filter.scala 230:62]
  wire [3:0] _GEN_391 = 10'hdc == _T_40[9:0] ? 4'h4 : _GEN_390; // @[Filter.scala 230:62]
  wire [3:0] _GEN_392 = 10'hdd == _T_40[9:0] ? 4'ha : _GEN_391; // @[Filter.scala 230:62]
  wire [3:0] _GEN_393 = 10'hde == _T_40[9:0] ? 4'ha : _GEN_392; // @[Filter.scala 230:62]
  wire [3:0] _GEN_394 = 10'hdf == _T_40[9:0] ? 4'ha : _GEN_393; // @[Filter.scala 230:62]
  wire [3:0] _GEN_395 = 10'he0 == _T_40[9:0] ? 4'ha : _GEN_394; // @[Filter.scala 230:62]
  wire [3:0] _GEN_396 = 10'he1 == _T_40[9:0] ? 4'ha : _GEN_395; // @[Filter.scala 230:62]
  wire [3:0] _GEN_397 = 10'he2 == _T_40[9:0] ? 4'ha : _GEN_396; // @[Filter.scala 230:62]
  wire [3:0] _GEN_398 = 10'he3 == _T_40[9:0] ? 4'h5 : _GEN_397; // @[Filter.scala 230:62]
  wire [3:0] _GEN_399 = 10'he4 == _T_40[9:0] ? 4'ha : _GEN_398; // @[Filter.scala 230:62]
  wire [3:0] _GEN_400 = 10'he5 == _T_40[9:0] ? 4'ha : _GEN_399; // @[Filter.scala 230:62]
  wire [3:0] _GEN_401 = 10'he6 == _T_40[9:0] ? 4'ha : _GEN_400; // @[Filter.scala 230:62]
  wire [3:0] _GEN_402 = 10'he7 == _T_40[9:0] ? 4'ha : _GEN_401; // @[Filter.scala 230:62]
  wire [3:0] _GEN_403 = 10'he8 == _T_40[9:0] ? 4'ha : _GEN_402; // @[Filter.scala 230:62]
  wire [3:0] _GEN_404 = 10'he9 == _T_40[9:0] ? 4'ha : _GEN_403; // @[Filter.scala 230:62]
  wire [3:0] _GEN_405 = 10'hea == _T_40[9:0] ? 4'ha : _GEN_404; // @[Filter.scala 230:62]
  wire [3:0] _GEN_406 = 10'heb == _T_40[9:0] ? 4'h9 : _GEN_405; // @[Filter.scala 230:62]
  wire [3:0] _GEN_407 = 10'hec == _T_40[9:0] ? 4'h7 : _GEN_406; // @[Filter.scala 230:62]
  wire [3:0] _GEN_408 = 10'hed == _T_40[9:0] ? 4'h3 : _GEN_407; // @[Filter.scala 230:62]
  wire [3:0] _GEN_409 = 10'hee == _T_40[9:0] ? 4'h3 : _GEN_408; // @[Filter.scala 230:62]
  wire [3:0] _GEN_410 = 10'hef == _T_40[9:0] ? 4'h3 : _GEN_409; // @[Filter.scala 230:62]
  wire [3:0] _GEN_411 = 10'hf0 == _T_40[9:0] ? 4'h4 : _GEN_410; // @[Filter.scala 230:62]
  wire [3:0] _GEN_412 = 10'hf1 == _T_40[9:0] ? 4'h7 : _GEN_411; // @[Filter.scala 230:62]
  wire [3:0] _GEN_413 = 10'hf2 == _T_40[9:0] ? 4'ha : _GEN_412; // @[Filter.scala 230:62]
  wire [3:0] _GEN_414 = 10'hf3 == _T_40[9:0] ? 4'ha : _GEN_413; // @[Filter.scala 230:62]
  wire [3:0] _GEN_415 = 10'hf4 == _T_40[9:0] ? 4'ha : _GEN_414; // @[Filter.scala 230:62]
  wire [3:0] _GEN_416 = 10'hf5 == _T_40[9:0] ? 4'h7 : _GEN_415; // @[Filter.scala 230:62]
  wire [3:0] _GEN_417 = 10'hf6 == _T_40[9:0] ? 4'h3 : _GEN_416; // @[Filter.scala 230:62]
  wire [3:0] _GEN_418 = 10'hf7 == _T_40[9:0] ? 4'h3 : _GEN_417; // @[Filter.scala 230:62]
  wire [3:0] _GEN_419 = 10'hf8 == _T_40[9:0] ? 4'h3 : _GEN_418; // @[Filter.scala 230:62]
  wire [3:0] _GEN_420 = 10'hf9 == _T_40[9:0] ? 4'h3 : _GEN_419; // @[Filter.scala 230:62]
  wire [3:0] _GEN_421 = 10'hfa == _T_40[9:0] ? 4'h3 : _GEN_420; // @[Filter.scala 230:62]
  wire [3:0] _GEN_422 = 10'hfb == _T_40[9:0] ? 4'h3 : _GEN_421; // @[Filter.scala 230:62]
  wire [3:0] _GEN_423 = 10'hfc == _T_40[9:0] ? 4'h3 : _GEN_422; // @[Filter.scala 230:62]
  wire [3:0] _GEN_424 = 10'hfd == _T_40[9:0] ? 4'h3 : _GEN_423; // @[Filter.scala 230:62]
  wire [3:0] _GEN_425 = 10'hfe == _T_40[9:0] ? 4'h3 : _GEN_424; // @[Filter.scala 230:62]
  wire [3:0] _GEN_426 = 10'hff == _T_40[9:0] ? 4'h3 : _GEN_425; // @[Filter.scala 230:62]
  wire [3:0] _GEN_427 = 10'h100 == _T_40[9:0] ? 4'h3 : _GEN_426; // @[Filter.scala 230:62]
  wire [3:0] _GEN_428 = 10'h101 == _T_40[9:0] ? 4'h4 : _GEN_427; // @[Filter.scala 230:62]
  wire [3:0] _GEN_429 = 10'h102 == _T_40[9:0] ? 4'h6 : _GEN_428; // @[Filter.scala 230:62]
  wire [3:0] _GEN_430 = 10'h103 == _T_40[9:0] ? 4'ha : _GEN_429; // @[Filter.scala 230:62]
  wire [3:0] _GEN_431 = 10'h104 == _T_40[9:0] ? 4'ha : _GEN_430; // @[Filter.scala 230:62]
  wire [3:0] _GEN_432 = 10'h105 == _T_40[9:0] ? 4'h9 : _GEN_431; // @[Filter.scala 230:62]
  wire [3:0] _GEN_433 = 10'h106 == _T_40[9:0] ? 4'h9 : _GEN_432; // @[Filter.scala 230:62]
  wire [3:0] _GEN_434 = 10'h107 == _T_40[9:0] ? 4'h9 : _GEN_433; // @[Filter.scala 230:62]
  wire [3:0] _GEN_435 = 10'h108 == _T_40[9:0] ? 4'h9 : _GEN_434; // @[Filter.scala 230:62]
  wire [3:0] _GEN_436 = 10'h109 == _T_40[9:0] ? 4'h3 : _GEN_435; // @[Filter.scala 230:62]
  wire [3:0] _GEN_437 = 10'h10a == _T_40[9:0] ? 4'ha : _GEN_436; // @[Filter.scala 230:62]
  wire [3:0] _GEN_438 = 10'h10b == _T_40[9:0] ? 4'ha : _GEN_437; // @[Filter.scala 230:62]
  wire [3:0] _GEN_439 = 10'h10c == _T_40[9:0] ? 4'ha : _GEN_438; // @[Filter.scala 230:62]
  wire [3:0] _GEN_440 = 10'h10d == _T_40[9:0] ? 4'ha : _GEN_439; // @[Filter.scala 230:62]
  wire [3:0] _GEN_441 = 10'h10e == _T_40[9:0] ? 4'ha : _GEN_440; // @[Filter.scala 230:62]
  wire [3:0] _GEN_442 = 10'h10f == _T_40[9:0] ? 4'h9 : _GEN_441; // @[Filter.scala 230:62]
  wire [3:0] _GEN_443 = 10'h110 == _T_40[9:0] ? 4'h9 : _GEN_442; // @[Filter.scala 230:62]
  wire [3:0] _GEN_444 = 10'h111 == _T_40[9:0] ? 4'h4 : _GEN_443; // @[Filter.scala 230:62]
  wire [3:0] _GEN_445 = 10'h112 == _T_40[9:0] ? 4'h8 : _GEN_444; // @[Filter.scala 230:62]
  wire [3:0] _GEN_446 = 10'h113 == _T_40[9:0] ? 4'h3 : _GEN_445; // @[Filter.scala 230:62]
  wire [3:0] _GEN_447 = 10'h114 == _T_40[9:0] ? 4'h3 : _GEN_446; // @[Filter.scala 230:62]
  wire [3:0] _GEN_448 = 10'h115 == _T_40[9:0] ? 4'h4 : _GEN_447; // @[Filter.scala 230:62]
  wire [3:0] _GEN_449 = 10'h116 == _T_40[9:0] ? 4'h4 : _GEN_448; // @[Filter.scala 230:62]
  wire [3:0] _GEN_450 = 10'h117 == _T_40[9:0] ? 4'h3 : _GEN_449; // @[Filter.scala 230:62]
  wire [3:0] _GEN_451 = 10'h118 == _T_40[9:0] ? 4'h8 : _GEN_450; // @[Filter.scala 230:62]
  wire [3:0] _GEN_452 = 10'h119 == _T_40[9:0] ? 4'ha : _GEN_451; // @[Filter.scala 230:62]
  wire [3:0] _GEN_453 = 10'h11a == _T_40[9:0] ? 4'ha : _GEN_452; // @[Filter.scala 230:62]
  wire [3:0] _GEN_454 = 10'h11b == _T_40[9:0] ? 4'ha : _GEN_453; // @[Filter.scala 230:62]
  wire [3:0] _GEN_455 = 10'h11c == _T_40[9:0] ? 4'h6 : _GEN_454; // @[Filter.scala 230:62]
  wire [3:0] _GEN_456 = 10'h11d == _T_40[9:0] ? 4'h3 : _GEN_455; // @[Filter.scala 230:62]
  wire [3:0] _GEN_457 = 10'h11e == _T_40[9:0] ? 4'h3 : _GEN_456; // @[Filter.scala 230:62]
  wire [3:0] _GEN_458 = 10'h11f == _T_40[9:0] ? 4'h3 : _GEN_457; // @[Filter.scala 230:62]
  wire [3:0] _GEN_459 = 10'h120 == _T_40[9:0] ? 4'h3 : _GEN_458; // @[Filter.scala 230:62]
  wire [3:0] _GEN_460 = 10'h121 == _T_40[9:0] ? 4'h3 : _GEN_459; // @[Filter.scala 230:62]
  wire [3:0] _GEN_461 = 10'h122 == _T_40[9:0] ? 4'h3 : _GEN_460; // @[Filter.scala 230:62]
  wire [3:0] _GEN_462 = 10'h123 == _T_40[9:0] ? 4'h3 : _GEN_461; // @[Filter.scala 230:62]
  wire [3:0] _GEN_463 = 10'h124 == _T_40[9:0] ? 4'h3 : _GEN_462; // @[Filter.scala 230:62]
  wire [3:0] _GEN_464 = 10'h125 == _T_40[9:0] ? 4'h3 : _GEN_463; // @[Filter.scala 230:62]
  wire [3:0] _GEN_465 = 10'h126 == _T_40[9:0] ? 4'h4 : _GEN_464; // @[Filter.scala 230:62]
  wire [3:0] _GEN_466 = 10'h127 == _T_40[9:0] ? 4'h6 : _GEN_465; // @[Filter.scala 230:62]
  wire [3:0] _GEN_467 = 10'h128 == _T_40[9:0] ? 4'h5 : _GEN_466; // @[Filter.scala 230:62]
  wire [3:0] _GEN_468 = 10'h129 == _T_40[9:0] ? 4'h8 : _GEN_467; // @[Filter.scala 230:62]
  wire [3:0] _GEN_469 = 10'h12a == _T_40[9:0] ? 4'h5 : _GEN_468; // @[Filter.scala 230:62]
  wire [3:0] _GEN_470 = 10'h12b == _T_40[9:0] ? 4'h3 : _GEN_469; // @[Filter.scala 230:62]
  wire [3:0] _GEN_471 = 10'h12c == _T_40[9:0] ? 4'h3 : _GEN_470; // @[Filter.scala 230:62]
  wire [3:0] _GEN_472 = 10'h12d == _T_40[9:0] ? 4'h3 : _GEN_471; // @[Filter.scala 230:62]
  wire [3:0] _GEN_473 = 10'h12e == _T_40[9:0] ? 4'h4 : _GEN_472; // @[Filter.scala 230:62]
  wire [3:0] _GEN_474 = 10'h12f == _T_40[9:0] ? 4'h4 : _GEN_473; // @[Filter.scala 230:62]
  wire [3:0] _GEN_475 = 10'h130 == _T_40[9:0] ? 4'ha : _GEN_474; // @[Filter.scala 230:62]
  wire [3:0] _GEN_476 = 10'h131 == _T_40[9:0] ? 4'h9 : _GEN_475; // @[Filter.scala 230:62]
  wire [3:0] _GEN_477 = 10'h132 == _T_40[9:0] ? 4'h9 : _GEN_476; // @[Filter.scala 230:62]
  wire [3:0] _GEN_478 = 10'h133 == _T_40[9:0] ? 4'h8 : _GEN_477; // @[Filter.scala 230:62]
  wire [3:0] _GEN_479 = 10'h134 == _T_40[9:0] ? 4'h9 : _GEN_478; // @[Filter.scala 230:62]
  wire [3:0] _GEN_480 = 10'h135 == _T_40[9:0] ? 4'h8 : _GEN_479; // @[Filter.scala 230:62]
  wire [3:0] _GEN_481 = 10'h136 == _T_40[9:0] ? 4'h7 : _GEN_480; // @[Filter.scala 230:62]
  wire [3:0] _GEN_482 = 10'h137 == _T_40[9:0] ? 4'h6 : _GEN_481; // @[Filter.scala 230:62]
  wire [3:0] _GEN_483 = 10'h138 == _T_40[9:0] ? 4'h8 : _GEN_482; // @[Filter.scala 230:62]
  wire [3:0] _GEN_484 = 10'h139 == _T_40[9:0] ? 4'h3 : _GEN_483; // @[Filter.scala 230:62]
  wire [3:0] _GEN_485 = 10'h13a == _T_40[9:0] ? 4'h3 : _GEN_484; // @[Filter.scala 230:62]
  wire [3:0] _GEN_486 = 10'h13b == _T_40[9:0] ? 4'h4 : _GEN_485; // @[Filter.scala 230:62]
  wire [3:0] _GEN_487 = 10'h13c == _T_40[9:0] ? 4'h4 : _GEN_486; // @[Filter.scala 230:62]
  wire [3:0] _GEN_488 = 10'h13d == _T_40[9:0] ? 4'h3 : _GEN_487; // @[Filter.scala 230:62]
  wire [3:0] _GEN_489 = 10'h13e == _T_40[9:0] ? 4'h5 : _GEN_488; // @[Filter.scala 230:62]
  wire [3:0] _GEN_490 = 10'h13f == _T_40[9:0] ? 4'h9 : _GEN_489; // @[Filter.scala 230:62]
  wire [3:0] _GEN_491 = 10'h140 == _T_40[9:0] ? 4'ha : _GEN_490; // @[Filter.scala 230:62]
  wire [3:0] _GEN_492 = 10'h141 == _T_40[9:0] ? 4'ha : _GEN_491; // @[Filter.scala 230:62]
  wire [3:0] _GEN_493 = 10'h142 == _T_40[9:0] ? 4'ha : _GEN_492; // @[Filter.scala 230:62]
  wire [3:0] _GEN_494 = 10'h143 == _T_40[9:0] ? 4'h5 : _GEN_493; // @[Filter.scala 230:62]
  wire [3:0] _GEN_495 = 10'h144 == _T_40[9:0] ? 4'h3 : _GEN_494; // @[Filter.scala 230:62]
  wire [3:0] _GEN_496 = 10'h145 == _T_40[9:0] ? 4'h3 : _GEN_495; // @[Filter.scala 230:62]
  wire [3:0] _GEN_497 = 10'h146 == _T_40[9:0] ? 4'h3 : _GEN_496; // @[Filter.scala 230:62]
  wire [3:0] _GEN_498 = 10'h147 == _T_40[9:0] ? 4'h4 : _GEN_497; // @[Filter.scala 230:62]
  wire [3:0] _GEN_499 = 10'h148 == _T_40[9:0] ? 4'h3 : _GEN_498; // @[Filter.scala 230:62]
  wire [3:0] _GEN_500 = 10'h149 == _T_40[9:0] ? 4'h3 : _GEN_499; // @[Filter.scala 230:62]
  wire [3:0] _GEN_501 = 10'h14a == _T_40[9:0] ? 4'h3 : _GEN_500; // @[Filter.scala 230:62]
  wire [3:0] _GEN_502 = 10'h14b == _T_40[9:0] ? 4'h6 : _GEN_501; // @[Filter.scala 230:62]
  wire [3:0] _GEN_503 = 10'h14c == _T_40[9:0] ? 4'h8 : _GEN_502; // @[Filter.scala 230:62]
  wire [3:0] _GEN_504 = 10'h14d == _T_40[9:0] ? 4'h5 : _GEN_503; // @[Filter.scala 230:62]
  wire [3:0] _GEN_505 = 10'h14e == _T_40[9:0] ? 4'h4 : _GEN_504; // @[Filter.scala 230:62]
  wire [3:0] _GEN_506 = 10'h14f == _T_40[9:0] ? 4'h3 : _GEN_505; // @[Filter.scala 230:62]
  wire [3:0] _GEN_507 = 10'h150 == _T_40[9:0] ? 4'h3 : _GEN_506; // @[Filter.scala 230:62]
  wire [3:0] _GEN_508 = 10'h151 == _T_40[9:0] ? 4'h3 : _GEN_507; // @[Filter.scala 230:62]
  wire [3:0] _GEN_509 = 10'h152 == _T_40[9:0] ? 4'h3 : _GEN_508; // @[Filter.scala 230:62]
  wire [3:0] _GEN_510 = 10'h153 == _T_40[9:0] ? 4'h3 : _GEN_509; // @[Filter.scala 230:62]
  wire [3:0] _GEN_511 = 10'h154 == _T_40[9:0] ? 4'h3 : _GEN_510; // @[Filter.scala 230:62]
  wire [3:0] _GEN_512 = 10'h155 == _T_40[9:0] ? 4'h4 : _GEN_511; // @[Filter.scala 230:62]
  wire [3:0] _GEN_513 = 10'h156 == _T_40[9:0] ? 4'h9 : _GEN_512; // @[Filter.scala 230:62]
  wire [3:0] _GEN_514 = 10'h157 == _T_40[9:0] ? 4'h8 : _GEN_513; // @[Filter.scala 230:62]
  wire [3:0] _GEN_515 = 10'h158 == _T_40[9:0] ? 4'h8 : _GEN_514; // @[Filter.scala 230:62]
  wire [3:0] _GEN_516 = 10'h159 == _T_40[9:0] ? 4'h8 : _GEN_515; // @[Filter.scala 230:62]
  wire [3:0] _GEN_517 = 10'h15a == _T_40[9:0] ? 4'h8 : _GEN_516; // @[Filter.scala 230:62]
  wire [3:0] _GEN_518 = 10'h15b == _T_40[9:0] ? 4'h8 : _GEN_517; // @[Filter.scala 230:62]
  wire [3:0] _GEN_519 = 10'h15c == _T_40[9:0] ? 4'h7 : _GEN_518; // @[Filter.scala 230:62]
  wire [3:0] _GEN_520 = 10'h15d == _T_40[9:0] ? 4'h7 : _GEN_519; // @[Filter.scala 230:62]
  wire [3:0] _GEN_521 = 10'h15e == _T_40[9:0] ? 4'h8 : _GEN_520; // @[Filter.scala 230:62]
  wire [3:0] _GEN_522 = 10'h15f == _T_40[9:0] ? 4'h3 : _GEN_521; // @[Filter.scala 230:62]
  wire [3:0] _GEN_523 = 10'h160 == _T_40[9:0] ? 4'h4 : _GEN_522; // @[Filter.scala 230:62]
  wire [3:0] _GEN_524 = 10'h161 == _T_40[9:0] ? 4'h4 : _GEN_523; // @[Filter.scala 230:62]
  wire [3:0] _GEN_525 = 10'h162 == _T_40[9:0] ? 4'h4 : _GEN_524; // @[Filter.scala 230:62]
  wire [3:0] _GEN_526 = 10'h163 == _T_40[9:0] ? 4'h4 : _GEN_525; // @[Filter.scala 230:62]
  wire [3:0] _GEN_527 = 10'h164 == _T_40[9:0] ? 4'h5 : _GEN_526; // @[Filter.scala 230:62]
  wire [3:0] _GEN_528 = 10'h165 == _T_40[9:0] ? 4'ha : _GEN_527; // @[Filter.scala 230:62]
  wire [3:0] _GEN_529 = 10'h166 == _T_40[9:0] ? 4'h9 : _GEN_528; // @[Filter.scala 230:62]
  wire [3:0] _GEN_530 = 10'h167 == _T_40[9:0] ? 4'ha : _GEN_529; // @[Filter.scala 230:62]
  wire [3:0] _GEN_531 = 10'h168 == _T_40[9:0] ? 4'ha : _GEN_530; // @[Filter.scala 230:62]
  wire [3:0] _GEN_532 = 10'h169 == _T_40[9:0] ? 4'h6 : _GEN_531; // @[Filter.scala 230:62]
  wire [3:0] _GEN_533 = 10'h16a == _T_40[9:0] ? 4'h3 : _GEN_532; // @[Filter.scala 230:62]
  wire [3:0] _GEN_534 = 10'h16b == _T_40[9:0] ? 4'h3 : _GEN_533; // @[Filter.scala 230:62]
  wire [3:0] _GEN_535 = 10'h16c == _T_40[9:0] ? 4'h3 : _GEN_534; // @[Filter.scala 230:62]
  wire [3:0] _GEN_536 = 10'h16d == _T_40[9:0] ? 4'h4 : _GEN_535; // @[Filter.scala 230:62]
  wire [3:0] _GEN_537 = 10'h16e == _T_40[9:0] ? 4'h3 : _GEN_536; // @[Filter.scala 230:62]
  wire [3:0] _GEN_538 = 10'h16f == _T_40[9:0] ? 4'h3 : _GEN_537; // @[Filter.scala 230:62]
  wire [3:0] _GEN_539 = 10'h170 == _T_40[9:0] ? 4'h3 : _GEN_538; // @[Filter.scala 230:62]
  wire [3:0] _GEN_540 = 10'h171 == _T_40[9:0] ? 4'h7 : _GEN_539; // @[Filter.scala 230:62]
  wire [3:0] _GEN_541 = 10'h172 == _T_40[9:0] ? 4'ha : _GEN_540; // @[Filter.scala 230:62]
  wire [3:0] _GEN_542 = 10'h173 == _T_40[9:0] ? 4'h5 : _GEN_541; // @[Filter.scala 230:62]
  wire [3:0] _GEN_543 = 10'h174 == _T_40[9:0] ? 4'h3 : _GEN_542; // @[Filter.scala 230:62]
  wire [3:0] _GEN_544 = 10'h175 == _T_40[9:0] ? 4'h4 : _GEN_543; // @[Filter.scala 230:62]
  wire [3:0] _GEN_545 = 10'h176 == _T_40[9:0] ? 4'h4 : _GEN_544; // @[Filter.scala 230:62]
  wire [3:0] _GEN_546 = 10'h177 == _T_40[9:0] ? 4'h4 : _GEN_545; // @[Filter.scala 230:62]
  wire [3:0] _GEN_547 = 10'h178 == _T_40[9:0] ? 4'h4 : _GEN_546; // @[Filter.scala 230:62]
  wire [3:0] _GEN_548 = 10'h179 == _T_40[9:0] ? 4'h3 : _GEN_547; // @[Filter.scala 230:62]
  wire [3:0] _GEN_549 = 10'h17a == _T_40[9:0] ? 4'h3 : _GEN_548; // @[Filter.scala 230:62]
  wire [3:0] _GEN_550 = 10'h17b == _T_40[9:0] ? 4'h3 : _GEN_549; // @[Filter.scala 230:62]
  wire [3:0] _GEN_551 = 10'h17c == _T_40[9:0] ? 4'h8 : _GEN_550; // @[Filter.scala 230:62]
  wire [3:0] _GEN_552 = 10'h17d == _T_40[9:0] ? 4'h8 : _GEN_551; // @[Filter.scala 230:62]
  wire [3:0] _GEN_553 = 10'h17e == _T_40[9:0] ? 4'h8 : _GEN_552; // @[Filter.scala 230:62]
  wire [3:0] _GEN_554 = 10'h17f == _T_40[9:0] ? 4'h8 : _GEN_553; // @[Filter.scala 230:62]
  wire [3:0] _GEN_555 = 10'h180 == _T_40[9:0] ? 4'h8 : _GEN_554; // @[Filter.scala 230:62]
  wire [3:0] _GEN_556 = 10'h181 == _T_40[9:0] ? 4'h8 : _GEN_555; // @[Filter.scala 230:62]
  wire [3:0] _GEN_557 = 10'h182 == _T_40[9:0] ? 4'h8 : _GEN_556; // @[Filter.scala 230:62]
  wire [3:0] _GEN_558 = 10'h183 == _T_40[9:0] ? 4'h8 : _GEN_557; // @[Filter.scala 230:62]
  wire [3:0] _GEN_559 = 10'h184 == _T_40[9:0] ? 4'h8 : _GEN_558; // @[Filter.scala 230:62]
  wire [3:0] _GEN_560 = 10'h185 == _T_40[9:0] ? 4'h5 : _GEN_559; // @[Filter.scala 230:62]
  wire [3:0] _GEN_561 = 10'h186 == _T_40[9:0] ? 4'h3 : _GEN_560; // @[Filter.scala 230:62]
  wire [3:0] _GEN_562 = 10'h187 == _T_40[9:0] ? 4'h4 : _GEN_561; // @[Filter.scala 230:62]
  wire [3:0] _GEN_563 = 10'h188 == _T_40[9:0] ? 4'h4 : _GEN_562; // @[Filter.scala 230:62]
  wire [3:0] _GEN_564 = 10'h189 == _T_40[9:0] ? 4'h4 : _GEN_563; // @[Filter.scala 230:62]
  wire [3:0] _GEN_565 = 10'h18a == _T_40[9:0] ? 4'h5 : _GEN_564; // @[Filter.scala 230:62]
  wire [3:0] _GEN_566 = 10'h18b == _T_40[9:0] ? 4'ha : _GEN_565; // @[Filter.scala 230:62]
  wire [3:0] _GEN_567 = 10'h18c == _T_40[9:0] ? 4'ha : _GEN_566; // @[Filter.scala 230:62]
  wire [3:0] _GEN_568 = 10'h18d == _T_40[9:0] ? 4'h9 : _GEN_567; // @[Filter.scala 230:62]
  wire [3:0] _GEN_569 = 10'h18e == _T_40[9:0] ? 4'ha : _GEN_568; // @[Filter.scala 230:62]
  wire [3:0] _GEN_570 = 10'h18f == _T_40[9:0] ? 4'h4 : _GEN_569; // @[Filter.scala 230:62]
  wire [3:0] _GEN_571 = 10'h190 == _T_40[9:0] ? 4'h3 : _GEN_570; // @[Filter.scala 230:62]
  wire [3:0] _GEN_572 = 10'h191 == _T_40[9:0] ? 4'h3 : _GEN_571; // @[Filter.scala 230:62]
  wire [3:0] _GEN_573 = 10'h192 == _T_40[9:0] ? 4'h5 : _GEN_572; // @[Filter.scala 230:62]
  wire [3:0] _GEN_574 = 10'h193 == _T_40[9:0] ? 4'h6 : _GEN_573; // @[Filter.scala 230:62]
  wire [3:0] _GEN_575 = 10'h194 == _T_40[9:0] ? 4'h5 : _GEN_574; // @[Filter.scala 230:62]
  wire [3:0] _GEN_576 = 10'h195 == _T_40[9:0] ? 4'h3 : _GEN_575; // @[Filter.scala 230:62]
  wire [3:0] _GEN_577 = 10'h196 == _T_40[9:0] ? 4'h3 : _GEN_576; // @[Filter.scala 230:62]
  wire [3:0] _GEN_578 = 10'h197 == _T_40[9:0] ? 4'h5 : _GEN_577; // @[Filter.scala 230:62]
  wire [3:0] _GEN_579 = 10'h198 == _T_40[9:0] ? 4'ha : _GEN_578; // @[Filter.scala 230:62]
  wire [3:0] _GEN_580 = 10'h199 == _T_40[9:0] ? 4'h3 : _GEN_579; // @[Filter.scala 230:62]
  wire [3:0] _GEN_581 = 10'h19a == _T_40[9:0] ? 4'h1 : _GEN_580; // @[Filter.scala 230:62]
  wire [3:0] _GEN_582 = 10'h19b == _T_40[9:0] ? 4'h2 : _GEN_581; // @[Filter.scala 230:62]
  wire [3:0] _GEN_583 = 10'h19c == _T_40[9:0] ? 4'h4 : _GEN_582; // @[Filter.scala 230:62]
  wire [3:0] _GEN_584 = 10'h19d == _T_40[9:0] ? 4'h3 : _GEN_583; // @[Filter.scala 230:62]
  wire [3:0] _GEN_585 = 10'h19e == _T_40[9:0] ? 4'h1 : _GEN_584; // @[Filter.scala 230:62]
  wire [3:0] _GEN_586 = 10'h19f == _T_40[9:0] ? 4'h2 : _GEN_585; // @[Filter.scala 230:62]
  wire [3:0] _GEN_587 = 10'h1a0 == _T_40[9:0] ? 4'h3 : _GEN_586; // @[Filter.scala 230:62]
  wire [3:0] _GEN_588 = 10'h1a1 == _T_40[9:0] ? 4'h4 : _GEN_587; // @[Filter.scala 230:62]
  wire [3:0] _GEN_589 = 10'h1a2 == _T_40[9:0] ? 4'h8 : _GEN_588; // @[Filter.scala 230:62]
  wire [3:0] _GEN_590 = 10'h1a3 == _T_40[9:0] ? 4'h8 : _GEN_589; // @[Filter.scala 230:62]
  wire [3:0] _GEN_591 = 10'h1a4 == _T_40[9:0] ? 4'h8 : _GEN_590; // @[Filter.scala 230:62]
  wire [3:0] _GEN_592 = 10'h1a5 == _T_40[9:0] ? 4'h8 : _GEN_591; // @[Filter.scala 230:62]
  wire [3:0] _GEN_593 = 10'h1a6 == _T_40[9:0] ? 4'h7 : _GEN_592; // @[Filter.scala 230:62]
  wire [3:0] _GEN_594 = 10'h1a7 == _T_40[9:0] ? 4'h8 : _GEN_593; // @[Filter.scala 230:62]
  wire [3:0] _GEN_595 = 10'h1a8 == _T_40[9:0] ? 4'h8 : _GEN_594; // @[Filter.scala 230:62]
  wire [3:0] _GEN_596 = 10'h1a9 == _T_40[9:0] ? 4'h8 : _GEN_595; // @[Filter.scala 230:62]
  wire [3:0] _GEN_597 = 10'h1aa == _T_40[9:0] ? 4'h7 : _GEN_596; // @[Filter.scala 230:62]
  wire [3:0] _GEN_598 = 10'h1ab == _T_40[9:0] ? 4'h4 : _GEN_597; // @[Filter.scala 230:62]
  wire [3:0] _GEN_599 = 10'h1ac == _T_40[9:0] ? 4'h4 : _GEN_598; // @[Filter.scala 230:62]
  wire [3:0] _GEN_600 = 10'h1ad == _T_40[9:0] ? 4'h3 : _GEN_599; // @[Filter.scala 230:62]
  wire [3:0] _GEN_601 = 10'h1ae == _T_40[9:0] ? 4'h3 : _GEN_600; // @[Filter.scala 230:62]
  wire [3:0] _GEN_602 = 10'h1af == _T_40[9:0] ? 4'h4 : _GEN_601; // @[Filter.scala 230:62]
  wire [3:0] _GEN_603 = 10'h1b0 == _T_40[9:0] ? 4'h6 : _GEN_602; // @[Filter.scala 230:62]
  wire [3:0] _GEN_604 = 10'h1b1 == _T_40[9:0] ? 4'ha : _GEN_603; // @[Filter.scala 230:62]
  wire [3:0] _GEN_605 = 10'h1b2 == _T_40[9:0] ? 4'ha : _GEN_604; // @[Filter.scala 230:62]
  wire [3:0] _GEN_606 = 10'h1b3 == _T_40[9:0] ? 4'h9 : _GEN_605; // @[Filter.scala 230:62]
  wire [3:0] _GEN_607 = 10'h1b4 == _T_40[9:0] ? 4'h9 : _GEN_606; // @[Filter.scala 230:62]
  wire [3:0] _GEN_608 = 10'h1b5 == _T_40[9:0] ? 4'h3 : _GEN_607; // @[Filter.scala 230:62]
  wire [3:0] _GEN_609 = 10'h1b6 == _T_40[9:0] ? 4'h3 : _GEN_608; // @[Filter.scala 230:62]
  wire [3:0] _GEN_610 = 10'h1b7 == _T_40[9:0] ? 4'h4 : _GEN_609; // @[Filter.scala 230:62]
  wire [3:0] _GEN_611 = 10'h1b8 == _T_40[9:0] ? 4'h5 : _GEN_610; // @[Filter.scala 230:62]
  wire [3:0] _GEN_612 = 10'h1b9 == _T_40[9:0] ? 4'h6 : _GEN_611; // @[Filter.scala 230:62]
  wire [3:0] _GEN_613 = 10'h1ba == _T_40[9:0] ? 4'h4 : _GEN_612; // @[Filter.scala 230:62]
  wire [3:0] _GEN_614 = 10'h1bb == _T_40[9:0] ? 4'h3 : _GEN_613; // @[Filter.scala 230:62]
  wire [3:0] _GEN_615 = 10'h1bc == _T_40[9:0] ? 4'h3 : _GEN_614; // @[Filter.scala 230:62]
  wire [3:0] _GEN_616 = 10'h1bd == _T_40[9:0] ? 4'h4 : _GEN_615; // @[Filter.scala 230:62]
  wire [3:0] _GEN_617 = 10'h1be == _T_40[9:0] ? 4'ha : _GEN_616; // @[Filter.scala 230:62]
  wire [3:0] _GEN_618 = 10'h1bf == _T_40[9:0] ? 4'h4 : _GEN_617; // @[Filter.scala 230:62]
  wire [3:0] _GEN_619 = 10'h1c0 == _T_40[9:0] ? 4'h5 : _GEN_618; // @[Filter.scala 230:62]
  wire [3:0] _GEN_620 = 10'h1c1 == _T_40[9:0] ? 4'h5 : _GEN_619; // @[Filter.scala 230:62]
  wire [3:0] _GEN_621 = 10'h1c2 == _T_40[9:0] ? 4'h4 : _GEN_620; // @[Filter.scala 230:62]
  wire [3:0] _GEN_622 = 10'h1c3 == _T_40[9:0] ? 4'h5 : _GEN_621; // @[Filter.scala 230:62]
  wire [3:0] _GEN_623 = 10'h1c4 == _T_40[9:0] ? 4'h4 : _GEN_622; // @[Filter.scala 230:62]
  wire [3:0] _GEN_624 = 10'h1c5 == _T_40[9:0] ? 4'h3 : _GEN_623; // @[Filter.scala 230:62]
  wire [3:0] _GEN_625 = 10'h1c6 == _T_40[9:0] ? 4'h4 : _GEN_624; // @[Filter.scala 230:62]
  wire [3:0] _GEN_626 = 10'h1c7 == _T_40[9:0] ? 4'h3 : _GEN_625; // @[Filter.scala 230:62]
  wire [3:0] _GEN_627 = 10'h1c8 == _T_40[9:0] ? 4'h8 : _GEN_626; // @[Filter.scala 230:62]
  wire [3:0] _GEN_628 = 10'h1c9 == _T_40[9:0] ? 4'h8 : _GEN_627; // @[Filter.scala 230:62]
  wire [3:0] _GEN_629 = 10'h1ca == _T_40[9:0] ? 4'h8 : _GEN_628; // @[Filter.scala 230:62]
  wire [3:0] _GEN_630 = 10'h1cb == _T_40[9:0] ? 4'h8 : _GEN_629; // @[Filter.scala 230:62]
  wire [3:0] _GEN_631 = 10'h1cc == _T_40[9:0] ? 4'h8 : _GEN_630; // @[Filter.scala 230:62]
  wire [3:0] _GEN_632 = 10'h1cd == _T_40[9:0] ? 4'h8 : _GEN_631; // @[Filter.scala 230:62]
  wire [3:0] _GEN_633 = 10'h1ce == _T_40[9:0] ? 4'h8 : _GEN_632; // @[Filter.scala 230:62]
  wire [3:0] _GEN_634 = 10'h1cf == _T_40[9:0] ? 4'h8 : _GEN_633; // @[Filter.scala 230:62]
  wire [3:0] _GEN_635 = 10'h1d0 == _T_40[9:0] ? 4'h5 : _GEN_634; // @[Filter.scala 230:62]
  wire [3:0] _GEN_636 = 10'h1d1 == _T_40[9:0] ? 4'h4 : _GEN_635; // @[Filter.scala 230:62]
  wire [3:0] _GEN_637 = 10'h1d2 == _T_40[9:0] ? 4'h6 : _GEN_636; // @[Filter.scala 230:62]
  wire [3:0] _GEN_638 = 10'h1d3 == _T_40[9:0] ? 4'h6 : _GEN_637; // @[Filter.scala 230:62]
  wire [3:0] _GEN_639 = 10'h1d4 == _T_40[9:0] ? 4'h6 : _GEN_638; // @[Filter.scala 230:62]
  wire [3:0] _GEN_640 = 10'h1d5 == _T_40[9:0] ? 4'h5 : _GEN_639; // @[Filter.scala 230:62]
  wire [3:0] _GEN_641 = 10'h1d6 == _T_40[9:0] ? 4'h8 : _GEN_640; // @[Filter.scala 230:62]
  wire [3:0] _GEN_642 = 10'h1d7 == _T_40[9:0] ? 4'ha : _GEN_641; // @[Filter.scala 230:62]
  wire [3:0] _GEN_643 = 10'h1d8 == _T_40[9:0] ? 4'ha : _GEN_642; // @[Filter.scala 230:62]
  wire [3:0] _GEN_644 = 10'h1d9 == _T_40[9:0] ? 4'ha : _GEN_643; // @[Filter.scala 230:62]
  wire [3:0] _GEN_645 = 10'h1da == _T_40[9:0] ? 4'h6 : _GEN_644; // @[Filter.scala 230:62]
  wire [3:0] _GEN_646 = 10'h1db == _T_40[9:0] ? 4'h3 : _GEN_645; // @[Filter.scala 230:62]
  wire [3:0] _GEN_647 = 10'h1dc == _T_40[9:0] ? 4'h5 : _GEN_646; // @[Filter.scala 230:62]
  wire [3:0] _GEN_648 = 10'h1dd == _T_40[9:0] ? 4'h2 : _GEN_647; // @[Filter.scala 230:62]
  wire [3:0] _GEN_649 = 10'h1de == _T_40[9:0] ? 4'h5 : _GEN_648; // @[Filter.scala 230:62]
  wire [3:0] _GEN_650 = 10'h1df == _T_40[9:0] ? 4'h5 : _GEN_649; // @[Filter.scala 230:62]
  wire [3:0] _GEN_651 = 10'h1e0 == _T_40[9:0] ? 4'h5 : _GEN_650; // @[Filter.scala 230:62]
  wire [3:0] _GEN_652 = 10'h1e1 == _T_40[9:0] ? 4'h3 : _GEN_651; // @[Filter.scala 230:62]
  wire [3:0] _GEN_653 = 10'h1e2 == _T_40[9:0] ? 4'h3 : _GEN_652; // @[Filter.scala 230:62]
  wire [3:0] _GEN_654 = 10'h1e3 == _T_40[9:0] ? 4'h3 : _GEN_653; // @[Filter.scala 230:62]
  wire [3:0] _GEN_655 = 10'h1e4 == _T_40[9:0] ? 4'h9 : _GEN_654; // @[Filter.scala 230:62]
  wire [3:0] _GEN_656 = 10'h1e5 == _T_40[9:0] ? 4'h4 : _GEN_655; // @[Filter.scala 230:62]
  wire [3:0] _GEN_657 = 10'h1e6 == _T_40[9:0] ? 4'h4 : _GEN_656; // @[Filter.scala 230:62]
  wire [3:0] _GEN_658 = 10'h1e7 == _T_40[9:0] ? 4'h4 : _GEN_657; // @[Filter.scala 230:62]
  wire [3:0] _GEN_659 = 10'h1e8 == _T_40[9:0] ? 4'h4 : _GEN_658; // @[Filter.scala 230:62]
  wire [3:0] _GEN_660 = 10'h1e9 == _T_40[9:0] ? 4'h4 : _GEN_659; // @[Filter.scala 230:62]
  wire [3:0] _GEN_661 = 10'h1ea == _T_40[9:0] ? 4'h4 : _GEN_660; // @[Filter.scala 230:62]
  wire [3:0] _GEN_662 = 10'h1eb == _T_40[9:0] ? 4'h4 : _GEN_661; // @[Filter.scala 230:62]
  wire [3:0] _GEN_663 = 10'h1ec == _T_40[9:0] ? 4'h4 : _GEN_662; // @[Filter.scala 230:62]
  wire [3:0] _GEN_664 = 10'h1ed == _T_40[9:0] ? 4'h4 : _GEN_663; // @[Filter.scala 230:62]
  wire [3:0] _GEN_665 = 10'h1ee == _T_40[9:0] ? 4'h8 : _GEN_664; // @[Filter.scala 230:62]
  wire [3:0] _GEN_666 = 10'h1ef == _T_40[9:0] ? 4'h8 : _GEN_665; // @[Filter.scala 230:62]
  wire [3:0] _GEN_667 = 10'h1f0 == _T_40[9:0] ? 4'h8 : _GEN_666; // @[Filter.scala 230:62]
  wire [3:0] _GEN_668 = 10'h1f1 == _T_40[9:0] ? 4'h8 : _GEN_667; // @[Filter.scala 230:62]
  wire [3:0] _GEN_669 = 10'h1f2 == _T_40[9:0] ? 4'h8 : _GEN_668; // @[Filter.scala 230:62]
  wire [3:0] _GEN_670 = 10'h1f3 == _T_40[9:0] ? 4'h8 : _GEN_669; // @[Filter.scala 230:62]
  wire [3:0] _GEN_671 = 10'h1f4 == _T_40[9:0] ? 4'h9 : _GEN_670; // @[Filter.scala 230:62]
  wire [3:0] _GEN_672 = 10'h1f5 == _T_40[9:0] ? 4'h9 : _GEN_671; // @[Filter.scala 230:62]
  wire [3:0] _GEN_673 = 10'h1f6 == _T_40[9:0] ? 4'ha : _GEN_672; // @[Filter.scala 230:62]
  wire [3:0] _GEN_674 = 10'h1f7 == _T_40[9:0] ? 4'h5 : _GEN_673; // @[Filter.scala 230:62]
  wire [3:0] _GEN_675 = 10'h1f8 == _T_40[9:0] ? 4'h5 : _GEN_674; // @[Filter.scala 230:62]
  wire [3:0] _GEN_676 = 10'h1f9 == _T_40[9:0] ? 4'h7 : _GEN_675; // @[Filter.scala 230:62]
  wire [3:0] _GEN_677 = 10'h1fa == _T_40[9:0] ? 4'h7 : _GEN_676; // @[Filter.scala 230:62]
  wire [3:0] _GEN_678 = 10'h1fb == _T_40[9:0] ? 4'h5 : _GEN_677; // @[Filter.scala 230:62]
  wire [3:0] _GEN_679 = 10'h1fc == _T_40[9:0] ? 4'ha : _GEN_678; // @[Filter.scala 230:62]
  wire [3:0] _GEN_680 = 10'h1fd == _T_40[9:0] ? 4'hb : _GEN_679; // @[Filter.scala 230:62]
  wire [3:0] _GEN_681 = 10'h1fe == _T_40[9:0] ? 4'hb : _GEN_680; // @[Filter.scala 230:62]
  wire [3:0] _GEN_682 = 10'h1ff == _T_40[9:0] ? 4'ha : _GEN_681; // @[Filter.scala 230:62]
  wire [3:0] _GEN_683 = 10'h200 == _T_40[9:0] ? 4'h4 : _GEN_682; // @[Filter.scala 230:62]
  wire [3:0] _GEN_684 = 10'h201 == _T_40[9:0] ? 4'h3 : _GEN_683; // @[Filter.scala 230:62]
  wire [3:0] _GEN_685 = 10'h202 == _T_40[9:0] ? 4'h2 : _GEN_684; // @[Filter.scala 230:62]
  wire [3:0] _GEN_686 = 10'h203 == _T_40[9:0] ? 4'h2 : _GEN_685; // @[Filter.scala 230:62]
  wire [3:0] _GEN_687 = 10'h204 == _T_40[9:0] ? 4'h2 : _GEN_686; // @[Filter.scala 230:62]
  wire [3:0] _GEN_688 = 10'h205 == _T_40[9:0] ? 4'h2 : _GEN_687; // @[Filter.scala 230:62]
  wire [3:0] _GEN_689 = 10'h206 == _T_40[9:0] ? 4'h2 : _GEN_688; // @[Filter.scala 230:62]
  wire [3:0] _GEN_690 = 10'h207 == _T_40[9:0] ? 4'h2 : _GEN_689; // @[Filter.scala 230:62]
  wire [3:0] _GEN_691 = 10'h208 == _T_40[9:0] ? 4'h3 : _GEN_690; // @[Filter.scala 230:62]
  wire [3:0] _GEN_692 = 10'h209 == _T_40[9:0] ? 4'h3 : _GEN_691; // @[Filter.scala 230:62]
  wire [3:0] _GEN_693 = 10'h20a == _T_40[9:0] ? 4'h8 : _GEN_692; // @[Filter.scala 230:62]
  wire [3:0] _GEN_694 = 10'h20b == _T_40[9:0] ? 4'h4 : _GEN_693; // @[Filter.scala 230:62]
  wire [3:0] _GEN_695 = 10'h20c == _T_40[9:0] ? 4'h4 : _GEN_694; // @[Filter.scala 230:62]
  wire [3:0] _GEN_696 = 10'h20d == _T_40[9:0] ? 4'h4 : _GEN_695; // @[Filter.scala 230:62]
  wire [3:0] _GEN_697 = 10'h20e == _T_40[9:0] ? 4'h4 : _GEN_696; // @[Filter.scala 230:62]
  wire [3:0] _GEN_698 = 10'h20f == _T_40[9:0] ? 4'h4 : _GEN_697; // @[Filter.scala 230:62]
  wire [3:0] _GEN_699 = 10'h210 == _T_40[9:0] ? 4'h4 : _GEN_698; // @[Filter.scala 230:62]
  wire [3:0] _GEN_700 = 10'h211 == _T_40[9:0] ? 4'h4 : _GEN_699; // @[Filter.scala 230:62]
  wire [3:0] _GEN_701 = 10'h212 == _T_40[9:0] ? 4'h4 : _GEN_700; // @[Filter.scala 230:62]
  wire [3:0] _GEN_702 = 10'h213 == _T_40[9:0] ? 4'h6 : _GEN_701; // @[Filter.scala 230:62]
  wire [3:0] _GEN_703 = 10'h214 == _T_40[9:0] ? 4'h7 : _GEN_702; // @[Filter.scala 230:62]
  wire [3:0] _GEN_704 = 10'h215 == _T_40[9:0] ? 4'h8 : _GEN_703; // @[Filter.scala 230:62]
  wire [3:0] _GEN_705 = 10'h216 == _T_40[9:0] ? 4'h8 : _GEN_704; // @[Filter.scala 230:62]
  wire [3:0] _GEN_706 = 10'h217 == _T_40[9:0] ? 4'h8 : _GEN_705; // @[Filter.scala 230:62]
  wire [3:0] _GEN_707 = 10'h218 == _T_40[9:0] ? 4'h8 : _GEN_706; // @[Filter.scala 230:62]
  wire [3:0] _GEN_708 = 10'h219 == _T_40[9:0] ? 4'h8 : _GEN_707; // @[Filter.scala 230:62]
  wire [3:0] _GEN_709 = 10'h21a == _T_40[9:0] ? 4'h8 : _GEN_708; // @[Filter.scala 230:62]
  wire [3:0] _GEN_710 = 10'h21b == _T_40[9:0] ? 4'h8 : _GEN_709; // @[Filter.scala 230:62]
  wire [3:0] _GEN_711 = 10'h21c == _T_40[9:0] ? 4'ha : _GEN_710; // @[Filter.scala 230:62]
  wire [3:0] _GEN_712 = 10'h21d == _T_40[9:0] ? 4'h9 : _GEN_711; // @[Filter.scala 230:62]
  wire [3:0] _GEN_713 = 10'h21e == _T_40[9:0] ? 4'h6 : _GEN_712; // @[Filter.scala 230:62]
  wire [3:0] _GEN_714 = 10'h21f == _T_40[9:0] ? 4'h4 : _GEN_713; // @[Filter.scala 230:62]
  wire [3:0] _GEN_715 = 10'h220 == _T_40[9:0] ? 4'h4 : _GEN_714; // @[Filter.scala 230:62]
  wire [3:0] _GEN_716 = 10'h221 == _T_40[9:0] ? 4'h5 : _GEN_715; // @[Filter.scala 230:62]
  wire [3:0] _GEN_717 = 10'h222 == _T_40[9:0] ? 4'ha : _GEN_716; // @[Filter.scala 230:62]
  wire [3:0] _GEN_718 = 10'h223 == _T_40[9:0] ? 4'ha : _GEN_717; // @[Filter.scala 230:62]
  wire [3:0] _GEN_719 = 10'h224 == _T_40[9:0] ? 4'ha : _GEN_718; // @[Filter.scala 230:62]
  wire [3:0] _GEN_720 = 10'h225 == _T_40[9:0] ? 4'h8 : _GEN_719; // @[Filter.scala 230:62]
  wire [3:0] _GEN_721 = 10'h226 == _T_40[9:0] ? 4'h4 : _GEN_720; // @[Filter.scala 230:62]
  wire [3:0] _GEN_722 = 10'h227 == _T_40[9:0] ? 4'h2 : _GEN_721; // @[Filter.scala 230:62]
  wire [3:0] _GEN_723 = 10'h228 == _T_40[9:0] ? 4'h2 : _GEN_722; // @[Filter.scala 230:62]
  wire [3:0] _GEN_724 = 10'h229 == _T_40[9:0] ? 4'h2 : _GEN_723; // @[Filter.scala 230:62]
  wire [3:0] _GEN_725 = 10'h22a == _T_40[9:0] ? 4'h2 : _GEN_724; // @[Filter.scala 230:62]
  wire [3:0] _GEN_726 = 10'h22b == _T_40[9:0] ? 4'h2 : _GEN_725; // @[Filter.scala 230:62]
  wire [3:0] _GEN_727 = 10'h22c == _T_40[9:0] ? 4'h2 : _GEN_726; // @[Filter.scala 230:62]
  wire [3:0] _GEN_728 = 10'h22d == _T_40[9:0] ? 4'h2 : _GEN_727; // @[Filter.scala 230:62]
  wire [3:0] _GEN_729 = 10'h22e == _T_40[9:0] ? 4'h2 : _GEN_728; // @[Filter.scala 230:62]
  wire [3:0] _GEN_730 = 10'h22f == _T_40[9:0] ? 4'h3 : _GEN_729; // @[Filter.scala 230:62]
  wire [3:0] _GEN_731 = 10'h230 == _T_40[9:0] ? 4'h3 : _GEN_730; // @[Filter.scala 230:62]
  wire [3:0] _GEN_732 = 10'h231 == _T_40[9:0] ? 4'h3 : _GEN_731; // @[Filter.scala 230:62]
  wire [3:0] _GEN_733 = 10'h232 == _T_40[9:0] ? 4'h4 : _GEN_732; // @[Filter.scala 230:62]
  wire [3:0] _GEN_734 = 10'h233 == _T_40[9:0] ? 4'h6 : _GEN_733; // @[Filter.scala 230:62]
  wire [3:0] _GEN_735 = 10'h234 == _T_40[9:0] ? 4'h6 : _GEN_734; // @[Filter.scala 230:62]
  wire [3:0] _GEN_736 = 10'h235 == _T_40[9:0] ? 4'h4 : _GEN_735; // @[Filter.scala 230:62]
  wire [3:0] _GEN_737 = 10'h236 == _T_40[9:0] ? 4'h4 : _GEN_736; // @[Filter.scala 230:62]
  wire [3:0] _GEN_738 = 10'h237 == _T_40[9:0] ? 4'h4 : _GEN_737; // @[Filter.scala 230:62]
  wire [3:0] _GEN_739 = 10'h238 == _T_40[9:0] ? 4'h4 : _GEN_738; // @[Filter.scala 230:62]
  wire [3:0] _GEN_740 = 10'h239 == _T_40[9:0] ? 4'h3 : _GEN_739; // @[Filter.scala 230:62]
  wire [3:0] _GEN_741 = 10'h23a == _T_40[9:0] ? 4'h7 : _GEN_740; // @[Filter.scala 230:62]
  wire [3:0] _GEN_742 = 10'h23b == _T_40[9:0] ? 4'h7 : _GEN_741; // @[Filter.scala 230:62]
  wire [3:0] _GEN_743 = 10'h23c == _T_40[9:0] ? 4'h7 : _GEN_742; // @[Filter.scala 230:62]
  wire [3:0] _GEN_744 = 10'h23d == _T_40[9:0] ? 4'h7 : _GEN_743; // @[Filter.scala 230:62]
  wire [3:0] _GEN_745 = 10'h23e == _T_40[9:0] ? 4'h7 : _GEN_744; // @[Filter.scala 230:62]
  wire [3:0] _GEN_746 = 10'h23f == _T_40[9:0] ? 4'h7 : _GEN_745; // @[Filter.scala 230:62]
  wire [3:0] _GEN_747 = 10'h240 == _T_40[9:0] ? 4'h7 : _GEN_746; // @[Filter.scala 230:62]
  wire [3:0] _GEN_748 = 10'h241 == _T_40[9:0] ? 4'h8 : _GEN_747; // @[Filter.scala 230:62]
  wire [3:0] _GEN_749 = 10'h242 == _T_40[9:0] ? 4'ha : _GEN_748; // @[Filter.scala 230:62]
  wire [3:0] _GEN_750 = 10'h243 == _T_40[9:0] ? 4'ha : _GEN_749; // @[Filter.scala 230:62]
  wire [3:0] _GEN_751 = 10'h244 == _T_40[9:0] ? 4'ha : _GEN_750; // @[Filter.scala 230:62]
  wire [3:0] _GEN_752 = 10'h245 == _T_40[9:0] ? 4'h8 : _GEN_751; // @[Filter.scala 230:62]
  wire [3:0] _GEN_753 = 10'h246 == _T_40[9:0] ? 4'h7 : _GEN_752; // @[Filter.scala 230:62]
  wire [3:0] _GEN_754 = 10'h247 == _T_40[9:0] ? 4'h8 : _GEN_753; // @[Filter.scala 230:62]
  wire [3:0] _GEN_755 = 10'h248 == _T_40[9:0] ? 4'ha : _GEN_754; // @[Filter.scala 230:62]
  wire [3:0] _GEN_756 = 10'h249 == _T_40[9:0] ? 4'ha : _GEN_755; // @[Filter.scala 230:62]
  wire [3:0] _GEN_757 = 10'h24a == _T_40[9:0] ? 4'ha : _GEN_756; // @[Filter.scala 230:62]
  wire [3:0] _GEN_758 = 10'h24b == _T_40[9:0] ? 4'h4 : _GEN_757; // @[Filter.scala 230:62]
  wire [3:0] _GEN_759 = 10'h24c == _T_40[9:0] ? 4'h4 : _GEN_758; // @[Filter.scala 230:62]
  wire [3:0] _GEN_760 = 10'h24d == _T_40[9:0] ? 4'h2 : _GEN_759; // @[Filter.scala 230:62]
  wire [3:0] _GEN_761 = 10'h24e == _T_40[9:0] ? 4'h2 : _GEN_760; // @[Filter.scala 230:62]
  wire [3:0] _GEN_762 = 10'h24f == _T_40[9:0] ? 4'h2 : _GEN_761; // @[Filter.scala 230:62]
  wire [3:0] _GEN_763 = 10'h250 == _T_40[9:0] ? 4'h2 : _GEN_762; // @[Filter.scala 230:62]
  wire [3:0] _GEN_764 = 10'h251 == _T_40[9:0] ? 4'h2 : _GEN_763; // @[Filter.scala 230:62]
  wire [3:0] _GEN_765 = 10'h252 == _T_40[9:0] ? 4'h2 : _GEN_764; // @[Filter.scala 230:62]
  wire [3:0] _GEN_766 = 10'h253 == _T_40[9:0] ? 4'h2 : _GEN_765; // @[Filter.scala 230:62]
  wire [3:0] _GEN_767 = 10'h254 == _T_40[9:0] ? 4'h2 : _GEN_766; // @[Filter.scala 230:62]
  wire [3:0] _GEN_768 = 10'h255 == _T_40[9:0] ? 4'h3 : _GEN_767; // @[Filter.scala 230:62]
  wire [3:0] _GEN_769 = 10'h256 == _T_40[9:0] ? 4'h4 : _GEN_768; // @[Filter.scala 230:62]
  wire [3:0] _GEN_770 = 10'h257 == _T_40[9:0] ? 4'h3 : _GEN_769; // @[Filter.scala 230:62]
  wire [3:0] _GEN_771 = 10'h258 == _T_40[9:0] ? 4'h4 : _GEN_770; // @[Filter.scala 230:62]
  wire [3:0] _GEN_772 = 10'h259 == _T_40[9:0] ? 4'h4 : _GEN_771; // @[Filter.scala 230:62]
  wire [3:0] _GEN_773 = 10'h25a == _T_40[9:0] ? 4'h4 : _GEN_772; // @[Filter.scala 230:62]
  wire [3:0] _GEN_774 = 10'h25b == _T_40[9:0] ? 4'h3 : _GEN_773; // @[Filter.scala 230:62]
  wire [3:0] _GEN_775 = 10'h25c == _T_40[9:0] ? 4'h4 : _GEN_774; // @[Filter.scala 230:62]
  wire [3:0] _GEN_776 = 10'h25d == _T_40[9:0] ? 4'h4 : _GEN_775; // @[Filter.scala 230:62]
  wire [3:0] _GEN_777 = 10'h25e == _T_40[9:0] ? 4'h3 : _GEN_776; // @[Filter.scala 230:62]
  wire [3:0] _GEN_778 = 10'h25f == _T_40[9:0] ? 4'h3 : _GEN_777; // @[Filter.scala 230:62]
  wire [3:0] _GEN_779 = 10'h260 == _T_40[9:0] ? 4'h8 : _GEN_778; // @[Filter.scala 230:62]
  wire [3:0] _GEN_780 = 10'h261 == _T_40[9:0] ? 4'h7 : _GEN_779; // @[Filter.scala 230:62]
  wire [3:0] _GEN_781 = 10'h262 == _T_40[9:0] ? 4'h6 : _GEN_780; // @[Filter.scala 230:62]
  wire [3:0] _GEN_782 = 10'h263 == _T_40[9:0] ? 4'h5 : _GEN_781; // @[Filter.scala 230:62]
  wire [3:0] _GEN_783 = 10'h264 == _T_40[9:0] ? 4'h6 : _GEN_782; // @[Filter.scala 230:62]
  wire [3:0] _GEN_784 = 10'h265 == _T_40[9:0] ? 4'h5 : _GEN_783; // @[Filter.scala 230:62]
  wire [3:0] _GEN_785 = 10'h266 == _T_40[9:0] ? 4'h5 : _GEN_784; // @[Filter.scala 230:62]
  wire [3:0] _GEN_786 = 10'h267 == _T_40[9:0] ? 4'h7 : _GEN_785; // @[Filter.scala 230:62]
  wire [3:0] _GEN_787 = 10'h268 == _T_40[9:0] ? 4'ha : _GEN_786; // @[Filter.scala 230:62]
  wire [3:0] _GEN_788 = 10'h269 == _T_40[9:0] ? 4'ha : _GEN_787; // @[Filter.scala 230:62]
  wire [3:0] _GEN_789 = 10'h26a == _T_40[9:0] ? 4'ha : _GEN_788; // @[Filter.scala 230:62]
  wire [3:0] _GEN_790 = 10'h26b == _T_40[9:0] ? 4'ha : _GEN_789; // @[Filter.scala 230:62]
  wire [3:0] _GEN_791 = 10'h26c == _T_40[9:0] ? 4'ha : _GEN_790; // @[Filter.scala 230:62]
  wire [3:0] _GEN_792 = 10'h26d == _T_40[9:0] ? 4'ha : _GEN_791; // @[Filter.scala 230:62]
  wire [3:0] _GEN_793 = 10'h26e == _T_40[9:0] ? 4'ha : _GEN_792; // @[Filter.scala 230:62]
  wire [3:0] _GEN_794 = 10'h26f == _T_40[9:0] ? 4'ha : _GEN_793; // @[Filter.scala 230:62]
  wire [3:0] _GEN_795 = 10'h270 == _T_40[9:0] ? 4'h5 : _GEN_794; // @[Filter.scala 230:62]
  wire [3:0] _GEN_796 = 10'h271 == _T_40[9:0] ? 4'h4 : _GEN_795; // @[Filter.scala 230:62]
  wire [3:0] _GEN_797 = 10'h272 == _T_40[9:0] ? 4'h3 : _GEN_796; // @[Filter.scala 230:62]
  wire [3:0] _GEN_798 = 10'h273 == _T_40[9:0] ? 4'h2 : _GEN_797; // @[Filter.scala 230:62]
  wire [3:0] _GEN_799 = 10'h274 == _T_40[9:0] ? 4'h2 : _GEN_798; // @[Filter.scala 230:62]
  wire [3:0] _GEN_800 = 10'h275 == _T_40[9:0] ? 4'h2 : _GEN_799; // @[Filter.scala 230:62]
  wire [3:0] _GEN_801 = 10'h276 == _T_40[9:0] ? 4'h2 : _GEN_800; // @[Filter.scala 230:62]
  wire [3:0] _GEN_802 = 10'h277 == _T_40[9:0] ? 4'h2 : _GEN_801; // @[Filter.scala 230:62]
  wire [3:0] _GEN_803 = 10'h278 == _T_40[9:0] ? 4'h2 : _GEN_802; // @[Filter.scala 230:62]
  wire [3:0] _GEN_804 = 10'h279 == _T_40[9:0] ? 4'h2 : _GEN_803; // @[Filter.scala 230:62]
  wire [3:0] _GEN_805 = 10'h27a == _T_40[9:0] ? 4'h2 : _GEN_804; // @[Filter.scala 230:62]
  wire [3:0] _GEN_806 = 10'h27b == _T_40[9:0] ? 4'h4 : _GEN_805; // @[Filter.scala 230:62]
  wire [3:0] _GEN_807 = 10'h27c == _T_40[9:0] ? 4'h3 : _GEN_806; // @[Filter.scala 230:62]
  wire [3:0] _GEN_808 = 10'h27d == _T_40[9:0] ? 4'h4 : _GEN_807; // @[Filter.scala 230:62]
  wire [3:0] _GEN_809 = 10'h27e == _T_40[9:0] ? 4'h5 : _GEN_808; // @[Filter.scala 230:62]
  wire [3:0] _GEN_810 = 10'h27f == _T_40[9:0] ? 4'h4 : _GEN_809; // @[Filter.scala 230:62]
  wire [3:0] _GEN_811 = 10'h280 == _T_40[9:0] ? 4'h4 : _GEN_810; // @[Filter.scala 230:62]
  wire [3:0] _GEN_812 = 10'h281 == _T_40[9:0] ? 4'h4 : _GEN_811; // @[Filter.scala 230:62]
  wire [3:0] _GEN_813 = 10'h282 == _T_40[9:0] ? 4'h4 : _GEN_812; // @[Filter.scala 230:62]
  wire [3:0] _GEN_814 = 10'h283 == _T_40[9:0] ? 4'h3 : _GEN_813; // @[Filter.scala 230:62]
  wire [3:0] _GEN_815 = 10'h284 == _T_40[9:0] ? 4'h3 : _GEN_814; // @[Filter.scala 230:62]
  wire [3:0] _GEN_816 = 10'h285 == _T_40[9:0] ? 4'h3 : _GEN_815; // @[Filter.scala 230:62]
  wire [3:0] _GEN_817 = 10'h286 == _T_40[9:0] ? 4'h8 : _GEN_816; // @[Filter.scala 230:62]
  wire [3:0] _GEN_818 = 10'h287 == _T_40[9:0] ? 4'h6 : _GEN_817; // @[Filter.scala 230:62]
  wire [3:0] _GEN_819 = 10'h288 == _T_40[9:0] ? 4'h6 : _GEN_818; // @[Filter.scala 230:62]
  wire [3:0] _GEN_820 = 10'h289 == _T_40[9:0] ? 4'h6 : _GEN_819; // @[Filter.scala 230:62]
  wire [3:0] _GEN_821 = 10'h28a == _T_40[9:0] ? 4'h7 : _GEN_820; // @[Filter.scala 230:62]
  wire [3:0] _GEN_822 = 10'h28b == _T_40[9:0] ? 4'h7 : _GEN_821; // @[Filter.scala 230:62]
  wire [3:0] _GEN_823 = 10'h28c == _T_40[9:0] ? 4'h6 : _GEN_822; // @[Filter.scala 230:62]
  wire [3:0] _GEN_824 = 10'h28d == _T_40[9:0] ? 4'h6 : _GEN_823; // @[Filter.scala 230:62]
  wire [3:0] _GEN_825 = 10'h28e == _T_40[9:0] ? 4'h4 : _GEN_824; // @[Filter.scala 230:62]
  wire [3:0] _GEN_826 = 10'h28f == _T_40[9:0] ? 4'h7 : _GEN_825; // @[Filter.scala 230:62]
  wire [3:0] _GEN_827 = 10'h290 == _T_40[9:0] ? 4'h9 : _GEN_826; // @[Filter.scala 230:62]
  wire [3:0] _GEN_828 = 10'h291 == _T_40[9:0] ? 4'ha : _GEN_827; // @[Filter.scala 230:62]
  wire [3:0] _GEN_829 = 10'h292 == _T_40[9:0] ? 4'ha : _GEN_828; // @[Filter.scala 230:62]
  wire [3:0] _GEN_830 = 10'h293 == _T_40[9:0] ? 4'ha : _GEN_829; // @[Filter.scala 230:62]
  wire [3:0] _GEN_831 = 10'h294 == _T_40[9:0] ? 4'h9 : _GEN_830; // @[Filter.scala 230:62]
  wire [3:0] _GEN_832 = 10'h295 == _T_40[9:0] ? 4'h5 : _GEN_831; // @[Filter.scala 230:62]
  wire [3:0] _GEN_833 = 10'h296 == _T_40[9:0] ? 4'h4 : _GEN_832; // @[Filter.scala 230:62]
  wire [3:0] _GEN_834 = 10'h297 == _T_40[9:0] ? 4'h4 : _GEN_833; // @[Filter.scala 230:62]
  wire [3:0] _GEN_835 = 10'h298 == _T_40[9:0] ? 4'h3 : _GEN_834; // @[Filter.scala 230:62]
  wire [3:0] _GEN_836 = 10'h299 == _T_40[9:0] ? 4'h3 : _GEN_835; // @[Filter.scala 230:62]
  wire [3:0] _GEN_837 = 10'h29a == _T_40[9:0] ? 4'h2 : _GEN_836; // @[Filter.scala 230:62]
  wire [3:0] _GEN_838 = 10'h29b == _T_40[9:0] ? 4'h2 : _GEN_837; // @[Filter.scala 230:62]
  wire [3:0] _GEN_839 = 10'h29c == _T_40[9:0] ? 4'h2 : _GEN_838; // @[Filter.scala 230:62]
  wire [3:0] _GEN_840 = 10'h29d == _T_40[9:0] ? 4'h2 : _GEN_839; // @[Filter.scala 230:62]
  wire [3:0] _GEN_841 = 10'h29e == _T_40[9:0] ? 4'h2 : _GEN_840; // @[Filter.scala 230:62]
  wire [3:0] _GEN_842 = 10'h29f == _T_40[9:0] ? 4'h2 : _GEN_841; // @[Filter.scala 230:62]
  wire [3:0] _GEN_843 = 10'h2a0 == _T_40[9:0] ? 4'h2 : _GEN_842; // @[Filter.scala 230:62]
  wire [3:0] _GEN_844 = 10'h2a1 == _T_40[9:0] ? 4'h4 : _GEN_843; // @[Filter.scala 230:62]
  wire [3:0] _GEN_845 = 10'h2a2 == _T_40[9:0] ? 4'h3 : _GEN_844; // @[Filter.scala 230:62]
  wire [3:0] _GEN_846 = 10'h2a3 == _T_40[9:0] ? 4'h4 : _GEN_845; // @[Filter.scala 230:62]
  wire [3:0] _GEN_847 = 10'h2a4 == _T_40[9:0] ? 4'h5 : _GEN_846; // @[Filter.scala 230:62]
  wire [3:0] _GEN_848 = 10'h2a5 == _T_40[9:0] ? 4'h4 : _GEN_847; // @[Filter.scala 230:62]
  wire [3:0] _GEN_849 = 10'h2a6 == _T_40[9:0] ? 4'h4 : _GEN_848; // @[Filter.scala 230:62]
  wire [3:0] _GEN_850 = 10'h2a7 == _T_40[9:0] ? 4'h4 : _GEN_849; // @[Filter.scala 230:62]
  wire [3:0] _GEN_851 = 10'h2a8 == _T_40[9:0] ? 4'h3 : _GEN_850; // @[Filter.scala 230:62]
  wire [3:0] _GEN_852 = 10'h2a9 == _T_40[9:0] ? 4'h3 : _GEN_851; // @[Filter.scala 230:62]
  wire [3:0] _GEN_853 = 10'h2aa == _T_40[9:0] ? 4'h3 : _GEN_852; // @[Filter.scala 230:62]
  wire [3:0] _GEN_854 = 10'h2ab == _T_40[9:0] ? 4'h3 : _GEN_853; // @[Filter.scala 230:62]
  wire [3:0] _GEN_855 = 10'h2ac == _T_40[9:0] ? 4'h8 : _GEN_854; // @[Filter.scala 230:62]
  wire [3:0] _GEN_856 = 10'h2ad == _T_40[9:0] ? 4'h7 : _GEN_855; // @[Filter.scala 230:62]
  wire [3:0] _GEN_857 = 10'h2ae == _T_40[9:0] ? 4'h5 : _GEN_856; // @[Filter.scala 230:62]
  wire [3:0] _GEN_858 = 10'h2af == _T_40[9:0] ? 4'h6 : _GEN_857; // @[Filter.scala 230:62]
  wire [3:0] _GEN_859 = 10'h2b0 == _T_40[9:0] ? 4'h7 : _GEN_858; // @[Filter.scala 230:62]
  wire [3:0] _GEN_860 = 10'h2b1 == _T_40[9:0] ? 4'h6 : _GEN_859; // @[Filter.scala 230:62]
  wire [3:0] _GEN_861 = 10'h2b2 == _T_40[9:0] ? 4'h6 : _GEN_860; // @[Filter.scala 230:62]
  wire [3:0] _GEN_862 = 10'h2b3 == _T_40[9:0] ? 4'h6 : _GEN_861; // @[Filter.scala 230:62]
  wire [3:0] _GEN_863 = 10'h2b4 == _T_40[9:0] ? 4'h3 : _GEN_862; // @[Filter.scala 230:62]
  wire [3:0] _GEN_864 = 10'h2b5 == _T_40[9:0] ? 4'h3 : _GEN_863; // @[Filter.scala 230:62]
  wire [3:0] _GEN_865 = 10'h2b6 == _T_40[9:0] ? 4'h3 : _GEN_864; // @[Filter.scala 230:62]
  wire [3:0] _GEN_866 = 10'h2b7 == _T_40[9:0] ? 4'h4 : _GEN_865; // @[Filter.scala 230:62]
  wire [3:0] _GEN_867 = 10'h2b8 == _T_40[9:0] ? 4'h6 : _GEN_866; // @[Filter.scala 230:62]
  wire [3:0] _GEN_868 = 10'h2b9 == _T_40[9:0] ? 4'h9 : _GEN_867; // @[Filter.scala 230:62]
  wire [3:0] _GEN_869 = 10'h2ba == _T_40[9:0] ? 4'h4 : _GEN_868; // @[Filter.scala 230:62]
  wire [3:0] _GEN_870 = 10'h2bb == _T_40[9:0] ? 4'h3 : _GEN_869; // @[Filter.scala 230:62]
  wire [3:0] _GEN_871 = 10'h2bc == _T_40[9:0] ? 4'h4 : _GEN_870; // @[Filter.scala 230:62]
  wire [3:0] _GEN_872 = 10'h2bd == _T_40[9:0] ? 4'h3 : _GEN_871; // @[Filter.scala 230:62]
  wire [3:0] _GEN_873 = 10'h2be == _T_40[9:0] ? 4'h3 : _GEN_872; // @[Filter.scala 230:62]
  wire [3:0] _GEN_874 = 10'h2bf == _T_40[9:0] ? 4'h3 : _GEN_873; // @[Filter.scala 230:62]
  wire [3:0] _GEN_875 = 10'h2c0 == _T_40[9:0] ? 4'h2 : _GEN_874; // @[Filter.scala 230:62]
  wire [3:0] _GEN_876 = 10'h2c1 == _T_40[9:0] ? 4'h2 : _GEN_875; // @[Filter.scala 230:62]
  wire [3:0] _GEN_877 = 10'h2c2 == _T_40[9:0] ? 4'h2 : _GEN_876; // @[Filter.scala 230:62]
  wire [3:0] _GEN_878 = 10'h2c3 == _T_40[9:0] ? 4'h2 : _GEN_877; // @[Filter.scala 230:62]
  wire [3:0] _GEN_879 = 10'h2c4 == _T_40[9:0] ? 4'h2 : _GEN_878; // @[Filter.scala 230:62]
  wire [3:0] _GEN_880 = 10'h2c5 == _T_40[9:0] ? 4'h2 : _GEN_879; // @[Filter.scala 230:62]
  wire [3:0] _GEN_881 = 10'h2c6 == _T_40[9:0] ? 4'h2 : _GEN_880; // @[Filter.scala 230:62]
  wire [3:0] _GEN_882 = 10'h2c7 == _T_40[9:0] ? 4'h4 : _GEN_881; // @[Filter.scala 230:62]
  wire [3:0] _GEN_883 = 10'h2c8 == _T_40[9:0] ? 4'h3 : _GEN_882; // @[Filter.scala 230:62]
  wire [3:0] _GEN_884 = 10'h2c9 == _T_40[9:0] ? 4'h4 : _GEN_883; // @[Filter.scala 230:62]
  wire [3:0] _GEN_885 = 10'h2ca == _T_40[9:0] ? 4'h5 : _GEN_884; // @[Filter.scala 230:62]
  wire [3:0] _GEN_886 = 10'h2cb == _T_40[9:0] ? 4'h3 : _GEN_885; // @[Filter.scala 230:62]
  wire [3:0] _GEN_887 = 10'h2cc == _T_40[9:0] ? 4'h3 : _GEN_886; // @[Filter.scala 230:62]
  wire [3:0] _GEN_888 = 10'h2cd == _T_40[9:0] ? 4'h3 : _GEN_887; // @[Filter.scala 230:62]
  wire [3:0] _GEN_889 = 10'h2ce == _T_40[9:0] ? 4'h3 : _GEN_888; // @[Filter.scala 230:62]
  wire [3:0] _GEN_890 = 10'h2cf == _T_40[9:0] ? 4'h3 : _GEN_889; // @[Filter.scala 230:62]
  wire [3:0] _GEN_891 = 10'h2d0 == _T_40[9:0] ? 4'h3 : _GEN_890; // @[Filter.scala 230:62]
  wire [3:0] _GEN_892 = 10'h2d1 == _T_40[9:0] ? 4'h3 : _GEN_891; // @[Filter.scala 230:62]
  wire [3:0] _GEN_893 = 10'h2d2 == _T_40[9:0] ? 4'h8 : _GEN_892; // @[Filter.scala 230:62]
  wire [3:0] _GEN_894 = 10'h2d3 == _T_40[9:0] ? 4'h6 : _GEN_893; // @[Filter.scala 230:62]
  wire [3:0] _GEN_895 = 10'h2d4 == _T_40[9:0] ? 4'h6 : _GEN_894; // @[Filter.scala 230:62]
  wire [3:0] _GEN_896 = 10'h2d5 == _T_40[9:0] ? 4'h7 : _GEN_895; // @[Filter.scala 230:62]
  wire [3:0] _GEN_897 = 10'h2d6 == _T_40[9:0] ? 4'h7 : _GEN_896; // @[Filter.scala 230:62]
  wire [3:0] _GEN_898 = 10'h2d7 == _T_40[9:0] ? 4'h7 : _GEN_897; // @[Filter.scala 230:62]
  wire [3:0] _GEN_899 = 10'h2d8 == _T_40[9:0] ? 4'h6 : _GEN_898; // @[Filter.scala 230:62]
  wire [3:0] _GEN_900 = 10'h2d9 == _T_40[9:0] ? 4'h7 : _GEN_899; // @[Filter.scala 230:62]
  wire [3:0] _GEN_901 = 10'h2da == _T_40[9:0] ? 4'h5 : _GEN_900; // @[Filter.scala 230:62]
  wire [3:0] _GEN_902 = 10'h2db == _T_40[9:0] ? 4'h3 : _GEN_901; // @[Filter.scala 230:62]
  wire [3:0] _GEN_903 = 10'h2dc == _T_40[9:0] ? 4'h3 : _GEN_902; // @[Filter.scala 230:62]
  wire [3:0] _GEN_904 = 10'h2dd == _T_40[9:0] ? 4'h3 : _GEN_903; // @[Filter.scala 230:62]
  wire [3:0] _GEN_905 = 10'h2de == _T_40[9:0] ? 4'h3 : _GEN_904; // @[Filter.scala 230:62]
  wire [3:0] _GEN_906 = 10'h2df == _T_40[9:0] ? 4'h4 : _GEN_905; // @[Filter.scala 230:62]
  wire [3:0] _GEN_907 = 10'h2e0 == _T_40[9:0] ? 4'h3 : _GEN_906; // @[Filter.scala 230:62]
  wire [3:0] _GEN_908 = 10'h2e1 == _T_40[9:0] ? 4'h3 : _GEN_907; // @[Filter.scala 230:62]
  wire [3:0] _GEN_909 = 10'h2e2 == _T_40[9:0] ? 4'h3 : _GEN_908; // @[Filter.scala 230:62]
  wire [3:0] _GEN_910 = 10'h2e3 == _T_40[9:0] ? 4'h3 : _GEN_909; // @[Filter.scala 230:62]
  wire [3:0] _GEN_911 = 10'h2e4 == _T_40[9:0] ? 4'h3 : _GEN_910; // @[Filter.scala 230:62]
  wire [3:0] _GEN_912 = 10'h2e5 == _T_40[9:0] ? 4'h3 : _GEN_911; // @[Filter.scala 230:62]
  wire [3:0] _GEN_913 = 10'h2e6 == _T_40[9:0] ? 4'h2 : _GEN_912; // @[Filter.scala 230:62]
  wire [3:0] _GEN_914 = 10'h2e7 == _T_40[9:0] ? 4'h2 : _GEN_913; // @[Filter.scala 230:62]
  wire [3:0] _GEN_915 = 10'h2e8 == _T_40[9:0] ? 4'h2 : _GEN_914; // @[Filter.scala 230:62]
  wire [3:0] _GEN_916 = 10'h2e9 == _T_40[9:0] ? 4'h2 : _GEN_915; // @[Filter.scala 230:62]
  wire [3:0] _GEN_917 = 10'h2ea == _T_40[9:0] ? 4'h2 : _GEN_916; // @[Filter.scala 230:62]
  wire [3:0] _GEN_918 = 10'h2eb == _T_40[9:0] ? 4'h2 : _GEN_917; // @[Filter.scala 230:62]
  wire [3:0] _GEN_919 = 10'h2ec == _T_40[9:0] ? 4'h3 : _GEN_918; // @[Filter.scala 230:62]
  wire [3:0] _GEN_920 = 10'h2ed == _T_40[9:0] ? 4'h4 : _GEN_919; // @[Filter.scala 230:62]
  wire [3:0] _GEN_921 = 10'h2ee == _T_40[9:0] ? 4'h3 : _GEN_920; // @[Filter.scala 230:62]
  wire [3:0] _GEN_922 = 10'h2ef == _T_40[9:0] ? 4'h3 : _GEN_921; // @[Filter.scala 230:62]
  wire [3:0] _GEN_923 = 10'h2f0 == _T_40[9:0] ? 4'h6 : _GEN_922; // @[Filter.scala 230:62]
  wire [3:0] _GEN_924 = 10'h2f1 == _T_40[9:0] ? 4'h3 : _GEN_923; // @[Filter.scala 230:62]
  wire [3:0] _GEN_925 = 10'h2f2 == _T_40[9:0] ? 4'h3 : _GEN_924; // @[Filter.scala 230:62]
  wire [3:0] _GEN_926 = 10'h2f3 == _T_40[9:0] ? 4'h3 : _GEN_925; // @[Filter.scala 230:62]
  wire [3:0] _GEN_927 = 10'h2f4 == _T_40[9:0] ? 4'h3 : _GEN_926; // @[Filter.scala 230:62]
  wire [3:0] _GEN_928 = 10'h2f5 == _T_40[9:0] ? 4'h3 : _GEN_927; // @[Filter.scala 230:62]
  wire [3:0] _GEN_929 = 10'h2f6 == _T_40[9:0] ? 4'h3 : _GEN_928; // @[Filter.scala 230:62]
  wire [3:0] _GEN_930 = 10'h2f7 == _T_40[9:0] ? 4'h3 : _GEN_929; // @[Filter.scala 230:62]
  wire [3:0] _GEN_931 = 10'h2f8 == _T_40[9:0] ? 4'h8 : _GEN_930; // @[Filter.scala 230:62]
  wire [3:0] _GEN_932 = 10'h2f9 == _T_40[9:0] ? 4'h6 : _GEN_931; // @[Filter.scala 230:62]
  wire [3:0] _GEN_933 = 10'h2fa == _T_40[9:0] ? 4'h7 : _GEN_932; // @[Filter.scala 230:62]
  wire [3:0] _GEN_934 = 10'h2fb == _T_40[9:0] ? 4'h7 : _GEN_933; // @[Filter.scala 230:62]
  wire [3:0] _GEN_935 = 10'h2fc == _T_40[9:0] ? 4'h6 : _GEN_934; // @[Filter.scala 230:62]
  wire [3:0] _GEN_936 = 10'h2fd == _T_40[9:0] ? 4'h6 : _GEN_935; // @[Filter.scala 230:62]
  wire [3:0] _GEN_937 = 10'h2fe == _T_40[9:0] ? 4'h6 : _GEN_936; // @[Filter.scala 230:62]
  wire [3:0] _GEN_938 = 10'h2ff == _T_40[9:0] ? 4'h8 : _GEN_937; // @[Filter.scala 230:62]
  wire [3:0] _GEN_939 = 10'h300 == _T_40[9:0] ? 4'h9 : _GEN_938; // @[Filter.scala 230:62]
  wire [3:0] _GEN_940 = 10'h301 == _T_40[9:0] ? 4'h7 : _GEN_939; // @[Filter.scala 230:62]
  wire [3:0] _GEN_941 = 10'h302 == _T_40[9:0] ? 4'h4 : _GEN_940; // @[Filter.scala 230:62]
  wire [3:0] _GEN_942 = 10'h303 == _T_40[9:0] ? 4'h4 : _GEN_941; // @[Filter.scala 230:62]
  wire [3:0] _GEN_943 = 10'h304 == _T_40[9:0] ? 4'h3 : _GEN_942; // @[Filter.scala 230:62]
  wire [3:0] _GEN_944 = 10'h305 == _T_40[9:0] ? 4'h3 : _GEN_943; // @[Filter.scala 230:62]
  wire [3:0] _GEN_945 = 10'h306 == _T_40[9:0] ? 4'h3 : _GEN_944; // @[Filter.scala 230:62]
  wire [3:0] _GEN_946 = 10'h307 == _T_40[9:0] ? 4'h3 : _GEN_945; // @[Filter.scala 230:62]
  wire [3:0] _GEN_947 = 10'h308 == _T_40[9:0] ? 4'h3 : _GEN_946; // @[Filter.scala 230:62]
  wire [3:0] _GEN_948 = 10'h309 == _T_40[9:0] ? 4'h3 : _GEN_947; // @[Filter.scala 230:62]
  wire [3:0] _GEN_949 = 10'h30a == _T_40[9:0] ? 4'h3 : _GEN_948; // @[Filter.scala 230:62]
  wire [3:0] _GEN_950 = 10'h30b == _T_40[9:0] ? 4'h3 : _GEN_949; // @[Filter.scala 230:62]
  wire [3:0] _GEN_951 = 10'h30c == _T_40[9:0] ? 4'h2 : _GEN_950; // @[Filter.scala 230:62]
  wire [3:0] _GEN_952 = 10'h30d == _T_40[9:0] ? 4'h2 : _GEN_951; // @[Filter.scala 230:62]
  wire [3:0] _GEN_953 = 10'h30e == _T_40[9:0] ? 4'h2 : _GEN_952; // @[Filter.scala 230:62]
  wire [3:0] _GEN_954 = 10'h30f == _T_40[9:0] ? 4'h2 : _GEN_953; // @[Filter.scala 230:62]
  wire [3:0] _GEN_955 = 10'h310 == _T_40[9:0] ? 4'h2 : _GEN_954; // @[Filter.scala 230:62]
  wire [3:0] _GEN_956 = 10'h311 == _T_40[9:0] ? 4'h2 : _GEN_955; // @[Filter.scala 230:62]
  wire [3:0] _GEN_957 = 10'h312 == _T_40[9:0] ? 4'h3 : _GEN_956; // @[Filter.scala 230:62]
  wire [3:0] _GEN_958 = 10'h313 == _T_40[9:0] ? 4'h4 : _GEN_957; // @[Filter.scala 230:62]
  wire [3:0] _GEN_959 = 10'h314 == _T_40[9:0] ? 4'h3 : _GEN_958; // @[Filter.scala 230:62]
  wire [3:0] _GEN_960 = 10'h315 == _T_40[9:0] ? 4'h3 : _GEN_959; // @[Filter.scala 230:62]
  wire [3:0] _GEN_961 = 10'h316 == _T_40[9:0] ? 4'h5 : _GEN_960; // @[Filter.scala 230:62]
  wire [3:0] _GEN_962 = 10'h317 == _T_40[9:0] ? 4'h5 : _GEN_961; // @[Filter.scala 230:62]
  wire [3:0] _GEN_963 = 10'h318 == _T_40[9:0] ? 4'h3 : _GEN_962; // @[Filter.scala 230:62]
  wire [3:0] _GEN_964 = 10'h319 == _T_40[9:0] ? 4'h3 : _GEN_963; // @[Filter.scala 230:62]
  wire [3:0] _GEN_965 = 10'h31a == _T_40[9:0] ? 4'h3 : _GEN_964; // @[Filter.scala 230:62]
  wire [3:0] _GEN_966 = 10'h31b == _T_40[9:0] ? 4'h3 : _GEN_965; // @[Filter.scala 230:62]
  wire [3:0] _GEN_967 = 10'h31c == _T_40[9:0] ? 4'h3 : _GEN_966; // @[Filter.scala 230:62]
  wire [3:0] _GEN_968 = 10'h31d == _T_40[9:0] ? 4'h3 : _GEN_967; // @[Filter.scala 230:62]
  wire [4:0] _GEN_38954 = {{1'd0}, _GEN_968}; // @[Filter.scala 230:62]
  wire [8:0] _T_42 = _GEN_38954 * 5'h14; // @[Filter.scala 230:62]
  wire [3:0] _GEN_992 = 10'h17 == _T_40[9:0] ? 4'hb : 4'he; // @[Filter.scala 230:102]
  wire [3:0] _GEN_993 = 10'h18 == _T_40[9:0] ? 4'hc : _GEN_992; // @[Filter.scala 230:102]
  wire [3:0] _GEN_994 = 10'h19 == _T_40[9:0] ? 4'he : _GEN_993; // @[Filter.scala 230:102]
  wire [3:0] _GEN_995 = 10'h1a == _T_40[9:0] ? 4'he : _GEN_994; // @[Filter.scala 230:102]
  wire [3:0] _GEN_996 = 10'h1b == _T_40[9:0] ? 4'he : _GEN_995; // @[Filter.scala 230:102]
  wire [3:0] _GEN_997 = 10'h1c == _T_40[9:0] ? 4'he : _GEN_996; // @[Filter.scala 230:102]
  wire [3:0] _GEN_998 = 10'h1d == _T_40[9:0] ? 4'he : _GEN_997; // @[Filter.scala 230:102]
  wire [3:0] _GEN_999 = 10'h1e == _T_40[9:0] ? 4'he : _GEN_998; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1000 = 10'h1f == _T_40[9:0] ? 4'he : _GEN_999; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1001 = 10'h20 == _T_40[9:0] ? 4'he : _GEN_1000; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1002 = 10'h21 == _T_40[9:0] ? 4'he : _GEN_1001; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1003 = 10'h22 == _T_40[9:0] ? 4'he : _GEN_1002; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1004 = 10'h23 == _T_40[9:0] ? 4'he : _GEN_1003; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1005 = 10'h24 == _T_40[9:0] ? 4'he : _GEN_1004; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1006 = 10'h25 == _T_40[9:0] ? 4'he : _GEN_1005; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1007 = 10'h26 == _T_40[9:0] ? 4'he : _GEN_1006; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1008 = 10'h27 == _T_40[9:0] ? 4'he : _GEN_1007; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1009 = 10'h28 == _T_40[9:0] ? 4'he : _GEN_1008; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1010 = 10'h29 == _T_40[9:0] ? 4'he : _GEN_1009; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1011 = 10'h2a == _T_40[9:0] ? 4'he : _GEN_1010; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1012 = 10'h2b == _T_40[9:0] ? 4'he : _GEN_1011; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1013 = 10'h2c == _T_40[9:0] ? 4'he : _GEN_1012; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1014 = 10'h2d == _T_40[9:0] ? 4'he : _GEN_1013; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1015 = 10'h2e == _T_40[9:0] ? 4'he : _GEN_1014; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1016 = 10'h2f == _T_40[9:0] ? 4'he : _GEN_1015; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1017 = 10'h30 == _T_40[9:0] ? 4'he : _GEN_1016; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1018 = 10'h31 == _T_40[9:0] ? 4'he : _GEN_1017; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1019 = 10'h32 == _T_40[9:0] ? 4'he : _GEN_1018; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1020 = 10'h33 == _T_40[9:0] ? 4'he : _GEN_1019; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1021 = 10'h34 == _T_40[9:0] ? 4'he : _GEN_1020; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1022 = 10'h35 == _T_40[9:0] ? 4'he : _GEN_1021; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1023 = 10'h36 == _T_40[9:0] ? 4'he : _GEN_1022; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1024 = 10'h37 == _T_40[9:0] ? 4'he : _GEN_1023; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1025 = 10'h38 == _T_40[9:0] ? 4'he : _GEN_1024; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1026 = 10'h39 == _T_40[9:0] ? 4'he : _GEN_1025; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1027 = 10'h3a == _T_40[9:0] ? 4'he : _GEN_1026; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1028 = 10'h3b == _T_40[9:0] ? 4'he : _GEN_1027; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1029 = 10'h3c == _T_40[9:0] ? 4'ha : _GEN_1028; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1030 = 10'h3d == _T_40[9:0] ? 4'hc : _GEN_1029; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1031 = 10'h3e == _T_40[9:0] ? 4'hb : _GEN_1030; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1032 = 10'h3f == _T_40[9:0] ? 4'he : _GEN_1031; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1033 = 10'h40 == _T_40[9:0] ? 4'he : _GEN_1032; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1034 = 10'h41 == _T_40[9:0] ? 4'he : _GEN_1033; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1035 = 10'h42 == _T_40[9:0] ? 4'he : _GEN_1034; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1036 = 10'h43 == _T_40[9:0] ? 4'he : _GEN_1035; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1037 = 10'h44 == _T_40[9:0] ? 4'he : _GEN_1036; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1038 = 10'h45 == _T_40[9:0] ? 4'he : _GEN_1037; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1039 = 10'h46 == _T_40[9:0] ? 4'he : _GEN_1038; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1040 = 10'h47 == _T_40[9:0] ? 4'he : _GEN_1039; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1041 = 10'h48 == _T_40[9:0] ? 4'he : _GEN_1040; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1042 = 10'h49 == _T_40[9:0] ? 4'he : _GEN_1041; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1043 = 10'h4a == _T_40[9:0] ? 4'he : _GEN_1042; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1044 = 10'h4b == _T_40[9:0] ? 4'he : _GEN_1043; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1045 = 10'h4c == _T_40[9:0] ? 4'he : _GEN_1044; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1046 = 10'h4d == _T_40[9:0] ? 4'he : _GEN_1045; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1047 = 10'h4e == _T_40[9:0] ? 4'he : _GEN_1046; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1048 = 10'h4f == _T_40[9:0] ? 4'he : _GEN_1047; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1049 = 10'h50 == _T_40[9:0] ? 4'he : _GEN_1048; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1050 = 10'h51 == _T_40[9:0] ? 4'he : _GEN_1049; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1051 = 10'h52 == _T_40[9:0] ? 4'he : _GEN_1050; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1052 = 10'h53 == _T_40[9:0] ? 4'he : _GEN_1051; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1053 = 10'h54 == _T_40[9:0] ? 4'he : _GEN_1052; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1054 = 10'h55 == _T_40[9:0] ? 4'he : _GEN_1053; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1055 = 10'h56 == _T_40[9:0] ? 4'he : _GEN_1054; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1056 = 10'h57 == _T_40[9:0] ? 4'he : _GEN_1055; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1057 = 10'h58 == _T_40[9:0] ? 4'he : _GEN_1056; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1058 = 10'h59 == _T_40[9:0] ? 4'he : _GEN_1057; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1059 = 10'h5a == _T_40[9:0] ? 4'hc : _GEN_1058; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1060 = 10'h5b == _T_40[9:0] ? 4'hd : _GEN_1059; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1061 = 10'h5c == _T_40[9:0] ? 4'he : _GEN_1060; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1062 = 10'h5d == _T_40[9:0] ? 4'he : _GEN_1061; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1063 = 10'h5e == _T_40[9:0] ? 4'he : _GEN_1062; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1064 = 10'h5f == _T_40[9:0] ? 4'he : _GEN_1063; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1065 = 10'h60 == _T_40[9:0] ? 4'he : _GEN_1064; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1066 = 10'h61 == _T_40[9:0] ? 4'hd : _GEN_1065; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1067 = 10'h62 == _T_40[9:0] ? 4'hb : _GEN_1066; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1068 = 10'h63 == _T_40[9:0] ? 4'hc : _GEN_1067; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1069 = 10'h64 == _T_40[9:0] ? 4'ha : _GEN_1068; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1070 = 10'h65 == _T_40[9:0] ? 4'hd : _GEN_1069; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1071 = 10'h66 == _T_40[9:0] ? 4'he : _GEN_1070; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1072 = 10'h67 == _T_40[9:0] ? 4'he : _GEN_1071; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1073 = 10'h68 == _T_40[9:0] ? 4'he : _GEN_1072; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1074 = 10'h69 == _T_40[9:0] ? 4'he : _GEN_1073; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1075 = 10'h6a == _T_40[9:0] ? 4'he : _GEN_1074; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1076 = 10'h6b == _T_40[9:0] ? 4'hd : _GEN_1075; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1077 = 10'h6c == _T_40[9:0] ? 4'hc : _GEN_1076; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1078 = 10'h6d == _T_40[9:0] ? 4'hc : _GEN_1077; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1079 = 10'h6e == _T_40[9:0] ? 4'he : _GEN_1078; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1080 = 10'h6f == _T_40[9:0] ? 4'he : _GEN_1079; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1081 = 10'h70 == _T_40[9:0] ? 4'he : _GEN_1080; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1082 = 10'h71 == _T_40[9:0] ? 4'he : _GEN_1081; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1083 = 10'h72 == _T_40[9:0] ? 4'he : _GEN_1082; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1084 = 10'h73 == _T_40[9:0] ? 4'he : _GEN_1083; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1085 = 10'h74 == _T_40[9:0] ? 4'he : _GEN_1084; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1086 = 10'h75 == _T_40[9:0] ? 4'he : _GEN_1085; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1087 = 10'h76 == _T_40[9:0] ? 4'he : _GEN_1086; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1088 = 10'h77 == _T_40[9:0] ? 4'he : _GEN_1087; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1089 = 10'h78 == _T_40[9:0] ? 4'he : _GEN_1088; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1090 = 10'h79 == _T_40[9:0] ? 4'he : _GEN_1089; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1091 = 10'h7a == _T_40[9:0] ? 4'he : _GEN_1090; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1092 = 10'h7b == _T_40[9:0] ? 4'he : _GEN_1091; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1093 = 10'h7c == _T_40[9:0] ? 4'he : _GEN_1092; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1094 = 10'h7d == _T_40[9:0] ? 4'he : _GEN_1093; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1095 = 10'h7e == _T_40[9:0] ? 4'he : _GEN_1094; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1096 = 10'h7f == _T_40[9:0] ? 4'he : _GEN_1095; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1097 = 10'h80 == _T_40[9:0] ? 4'he : _GEN_1096; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1098 = 10'h81 == _T_40[9:0] ? 4'hb : _GEN_1097; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1099 = 10'h82 == _T_40[9:0] ? 4'hc : _GEN_1098; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1100 = 10'h83 == _T_40[9:0] ? 4'hc : _GEN_1099; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1101 = 10'h84 == _T_40[9:0] ? 4'he : _GEN_1100; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1102 = 10'h85 == _T_40[9:0] ? 4'he : _GEN_1101; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1103 = 10'h86 == _T_40[9:0] ? 4'he : _GEN_1102; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1104 = 10'h87 == _T_40[9:0] ? 4'ha : _GEN_1103; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1105 = 10'h88 == _T_40[9:0] ? 4'hd : _GEN_1104; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1106 = 10'h89 == _T_40[9:0] ? 4'hd : _GEN_1105; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1107 = 10'h8a == _T_40[9:0] ? 4'hc : _GEN_1106; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1108 = 10'h8b == _T_40[9:0] ? 4'he : _GEN_1107; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1109 = 10'h8c == _T_40[9:0] ? 4'he : _GEN_1108; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1110 = 10'h8d == _T_40[9:0] ? 4'he : _GEN_1109; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1111 = 10'h8e == _T_40[9:0] ? 4'he : _GEN_1110; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1112 = 10'h8f == _T_40[9:0] ? 4'hb : _GEN_1111; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1113 = 10'h90 == _T_40[9:0] ? 4'hc : _GEN_1112; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1114 = 10'h91 == _T_40[9:0] ? 4'hc : _GEN_1113; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1115 = 10'h92 == _T_40[9:0] ? 4'hd : _GEN_1114; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1116 = 10'h93 == _T_40[9:0] ? 4'he : _GEN_1115; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1117 = 10'h94 == _T_40[9:0] ? 4'he : _GEN_1116; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1118 = 10'h95 == _T_40[9:0] ? 4'he : _GEN_1117; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1119 = 10'h96 == _T_40[9:0] ? 4'he : _GEN_1118; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1120 = 10'h97 == _T_40[9:0] ? 4'he : _GEN_1119; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1121 = 10'h98 == _T_40[9:0] ? 4'he : _GEN_1120; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1122 = 10'h99 == _T_40[9:0] ? 4'he : _GEN_1121; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1123 = 10'h9a == _T_40[9:0] ? 4'he : _GEN_1122; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1124 = 10'h9b == _T_40[9:0] ? 4'he : _GEN_1123; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1125 = 10'h9c == _T_40[9:0] ? 4'he : _GEN_1124; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1126 = 10'h9d == _T_40[9:0] ? 4'he : _GEN_1125; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1127 = 10'h9e == _T_40[9:0] ? 4'he : _GEN_1126; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1128 = 10'h9f == _T_40[9:0] ? 4'he : _GEN_1127; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1129 = 10'ha0 == _T_40[9:0] ? 4'he : _GEN_1128; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1130 = 10'ha1 == _T_40[9:0] ? 4'he : _GEN_1129; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1131 = 10'ha2 == _T_40[9:0] ? 4'he : _GEN_1130; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1132 = 10'ha3 == _T_40[9:0] ? 4'he : _GEN_1131; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1133 = 10'ha4 == _T_40[9:0] ? 4'he : _GEN_1132; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1134 = 10'ha5 == _T_40[9:0] ? 4'he : _GEN_1133; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1135 = 10'ha6 == _T_40[9:0] ? 4'he : _GEN_1134; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1136 = 10'ha7 == _T_40[9:0] ? 4'he : _GEN_1135; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1137 = 10'ha8 == _T_40[9:0] ? 4'hb : _GEN_1136; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1138 = 10'ha9 == _T_40[9:0] ? 4'hc : _GEN_1137; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1139 = 10'haa == _T_40[9:0] ? 4'hb : _GEN_1138; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1140 = 10'hab == _T_40[9:0] ? 4'hc : _GEN_1139; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1141 = 10'hac == _T_40[9:0] ? 4'hd : _GEN_1140; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1142 = 10'had == _T_40[9:0] ? 4'ha : _GEN_1141; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1143 = 10'hae == _T_40[9:0] ? 4'hd : _GEN_1142; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1144 = 10'haf == _T_40[9:0] ? 4'hd : _GEN_1143; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1145 = 10'hb0 == _T_40[9:0] ? 4'hb : _GEN_1144; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1146 = 10'hb1 == _T_40[9:0] ? 4'hc : _GEN_1145; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1147 = 10'hb2 == _T_40[9:0] ? 4'he : _GEN_1146; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1148 = 10'hb3 == _T_40[9:0] ? 4'hb : _GEN_1147; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1149 = 10'hb4 == _T_40[9:0] ? 4'hc : _GEN_1148; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1150 = 10'hb5 == _T_40[9:0] ? 4'hd : _GEN_1149; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1151 = 10'hb6 == _T_40[9:0] ? 4'hd : _GEN_1150; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1152 = 10'hb7 == _T_40[9:0] ? 4'hc : _GEN_1151; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1153 = 10'hb8 == _T_40[9:0] ? 4'he : _GEN_1152; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1154 = 10'hb9 == _T_40[9:0] ? 4'he : _GEN_1153; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1155 = 10'hba == _T_40[9:0] ? 4'he : _GEN_1154; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1156 = 10'hbb == _T_40[9:0] ? 4'he : _GEN_1155; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1157 = 10'hbc == _T_40[9:0] ? 4'he : _GEN_1156; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1158 = 10'hbd == _T_40[9:0] ? 4'he : _GEN_1157; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1159 = 10'hbe == _T_40[9:0] ? 4'he : _GEN_1158; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1160 = 10'hbf == _T_40[9:0] ? 4'he : _GEN_1159; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1161 = 10'hc0 == _T_40[9:0] ? 4'he : _GEN_1160; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1162 = 10'hc1 == _T_40[9:0] ? 4'he : _GEN_1161; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1163 = 10'hc2 == _T_40[9:0] ? 4'he : _GEN_1162; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1164 = 10'hc3 == _T_40[9:0] ? 4'he : _GEN_1163; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1165 = 10'hc4 == _T_40[9:0] ? 4'he : _GEN_1164; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1166 = 10'hc5 == _T_40[9:0] ? 4'he : _GEN_1165; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1167 = 10'hc6 == _T_40[9:0] ? 4'he : _GEN_1166; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1168 = 10'hc7 == _T_40[9:0] ? 4'hd : _GEN_1167; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1169 = 10'hc8 == _T_40[9:0] ? 4'hb : _GEN_1168; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1170 = 10'hc9 == _T_40[9:0] ? 4'hc : _GEN_1169; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1171 = 10'hca == _T_40[9:0] ? 4'he : _GEN_1170; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1172 = 10'hcb == _T_40[9:0] ? 4'he : _GEN_1171; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1173 = 10'hcc == _T_40[9:0] ? 4'he : _GEN_1172; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1174 = 10'hcd == _T_40[9:0] ? 4'he : _GEN_1173; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1175 = 10'hce == _T_40[9:0] ? 4'hd : _GEN_1174; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1176 = 10'hcf == _T_40[9:0] ? 4'hb : _GEN_1175; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1177 = 10'hd0 == _T_40[9:0] ? 4'hc : _GEN_1176; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1178 = 10'hd1 == _T_40[9:0] ? 4'hc : _GEN_1177; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1179 = 10'hd2 == _T_40[9:0] ? 4'hb : _GEN_1178; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1180 = 10'hd3 == _T_40[9:0] ? 4'hd : _GEN_1179; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1181 = 10'hd4 == _T_40[9:0] ? 4'hd : _GEN_1180; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1182 = 10'hd5 == _T_40[9:0] ? 4'hd : _GEN_1181; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1183 = 10'hd6 == _T_40[9:0] ? 4'hd : _GEN_1182; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1184 = 10'hd7 == _T_40[9:0] ? 4'hc : _GEN_1183; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1185 = 10'hd8 == _T_40[9:0] ? 4'hc : _GEN_1184; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1186 = 10'hd9 == _T_40[9:0] ? 4'hc : _GEN_1185; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1187 = 10'hda == _T_40[9:0] ? 4'hd : _GEN_1186; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1188 = 10'hdb == _T_40[9:0] ? 4'hc : _GEN_1187; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1189 = 10'hdc == _T_40[9:0] ? 4'h9 : _GEN_1188; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1190 = 10'hdd == _T_40[9:0] ? 4'he : _GEN_1189; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1191 = 10'hde == _T_40[9:0] ? 4'he : _GEN_1190; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1192 = 10'hdf == _T_40[9:0] ? 4'he : _GEN_1191; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1193 = 10'he0 == _T_40[9:0] ? 4'he : _GEN_1192; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1194 = 10'he1 == _T_40[9:0] ? 4'he : _GEN_1193; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1195 = 10'he2 == _T_40[9:0] ? 4'he : _GEN_1194; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1196 = 10'he3 == _T_40[9:0] ? 4'h9 : _GEN_1195; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1197 = 10'he4 == _T_40[9:0] ? 4'he : _GEN_1196; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1198 = 10'he5 == _T_40[9:0] ? 4'he : _GEN_1197; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1199 = 10'he6 == _T_40[9:0] ? 4'he : _GEN_1198; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1200 = 10'he7 == _T_40[9:0] ? 4'he : _GEN_1199; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1201 = 10'he8 == _T_40[9:0] ? 4'he : _GEN_1200; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1202 = 10'he9 == _T_40[9:0] ? 4'he : _GEN_1201; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1203 = 10'hea == _T_40[9:0] ? 4'he : _GEN_1202; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1204 = 10'heb == _T_40[9:0] ? 4'hc : _GEN_1203; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1205 = 10'hec == _T_40[9:0] ? 4'h7 : _GEN_1204; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1206 = 10'hed == _T_40[9:0] ? 4'h1 : _GEN_1205; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1207 = 10'hee == _T_40[9:0] ? 4'h0 : _GEN_1206; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1208 = 10'hef == _T_40[9:0] ? 4'h0 : _GEN_1207; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1209 = 10'hf0 == _T_40[9:0] ? 4'h2 : _GEN_1208; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1210 = 10'hf1 == _T_40[9:0] ? 4'h9 : _GEN_1209; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1211 = 10'hf2 == _T_40[9:0] ? 4'he : _GEN_1210; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1212 = 10'hf3 == _T_40[9:0] ? 4'he : _GEN_1211; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1213 = 10'hf4 == _T_40[9:0] ? 4'he : _GEN_1212; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1214 = 10'hf5 == _T_40[9:0] ? 4'hc : _GEN_1213; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1215 = 10'hf6 == _T_40[9:0] ? 4'hc : _GEN_1214; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1216 = 10'hf7 == _T_40[9:0] ? 4'hd : _GEN_1215; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1217 = 10'hf8 == _T_40[9:0] ? 4'hd : _GEN_1216; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1218 = 10'hf9 == _T_40[9:0] ? 4'hd : _GEN_1217; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1219 = 10'hfa == _T_40[9:0] ? 4'hd : _GEN_1218; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1220 = 10'hfb == _T_40[9:0] ? 4'hd : _GEN_1219; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1221 = 10'hfc == _T_40[9:0] ? 4'hd : _GEN_1220; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1222 = 10'hfd == _T_40[9:0] ? 4'hd : _GEN_1221; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1223 = 10'hfe == _T_40[9:0] ? 4'hd : _GEN_1222; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1224 = 10'hff == _T_40[9:0] ? 4'hd : _GEN_1223; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1225 = 10'h100 == _T_40[9:0] ? 4'hd : _GEN_1224; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1226 = 10'h101 == _T_40[9:0] ? 4'h9 : _GEN_1225; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1227 = 10'h102 == _T_40[9:0] ? 4'h9 : _GEN_1226; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1228 = 10'h103 == _T_40[9:0] ? 4'he : _GEN_1227; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1229 = 10'h104 == _T_40[9:0] ? 4'he : _GEN_1228; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1230 = 10'h105 == _T_40[9:0] ? 4'he : _GEN_1229; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1231 = 10'h106 == _T_40[9:0] ? 4'he : _GEN_1230; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1232 = 10'h107 == _T_40[9:0] ? 4'he : _GEN_1231; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1233 = 10'h108 == _T_40[9:0] ? 4'he : _GEN_1232; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1234 = 10'h109 == _T_40[9:0] ? 4'h6 : _GEN_1233; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1235 = 10'h10a == _T_40[9:0] ? 4'he : _GEN_1234; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1236 = 10'h10b == _T_40[9:0] ? 4'he : _GEN_1235; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1237 = 10'h10c == _T_40[9:0] ? 4'he : _GEN_1236; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1238 = 10'h10d == _T_40[9:0] ? 4'he : _GEN_1237; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1239 = 10'h10e == _T_40[9:0] ? 4'he : _GEN_1238; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1240 = 10'h10f == _T_40[9:0] ? 4'ha : _GEN_1239; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1241 = 10'h110 == _T_40[9:0] ? 4'hd : _GEN_1240; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1242 = 10'h111 == _T_40[9:0] ? 4'h4 : _GEN_1241; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1243 = 10'h112 == _T_40[9:0] ? 4'h7 : _GEN_1242; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1244 = 10'h113 == _T_40[9:0] ? 4'h0 : _GEN_1243; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1245 = 10'h114 == _T_40[9:0] ? 4'h0 : _GEN_1244; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1246 = 10'h115 == _T_40[9:0] ? 4'h0 : _GEN_1245; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1247 = 10'h116 == _T_40[9:0] ? 4'h0 : _GEN_1246; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1248 = 10'h117 == _T_40[9:0] ? 4'h0 : _GEN_1247; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1249 = 10'h118 == _T_40[9:0] ? 4'ha : _GEN_1248; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1250 = 10'h119 == _T_40[9:0] ? 4'he : _GEN_1249; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1251 = 10'h11a == _T_40[9:0] ? 4'he : _GEN_1250; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1252 = 10'h11b == _T_40[9:0] ? 4'he : _GEN_1251; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1253 = 10'h11c == _T_40[9:0] ? 4'hb : _GEN_1252; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1254 = 10'h11d == _T_40[9:0] ? 4'hc : _GEN_1253; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1255 = 10'h11e == _T_40[9:0] ? 4'hd : _GEN_1254; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1256 = 10'h11f == _T_40[9:0] ? 4'hb : _GEN_1255; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1257 = 10'h120 == _T_40[9:0] ? 4'ha : _GEN_1256; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1258 = 10'h121 == _T_40[9:0] ? 4'hc : _GEN_1257; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1259 = 10'h122 == _T_40[9:0] ? 4'ha : _GEN_1258; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1260 = 10'h123 == _T_40[9:0] ? 4'ha : _GEN_1259; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1261 = 10'h124 == _T_40[9:0] ? 4'hd : _GEN_1260; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1262 = 10'h125 == _T_40[9:0] ? 4'hd : _GEN_1261; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1263 = 10'h126 == _T_40[9:0] ? 4'hb : _GEN_1262; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1264 = 10'h127 == _T_40[9:0] ? 4'h9 : _GEN_1263; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1265 = 10'h128 == _T_40[9:0] ? 4'h7 : _GEN_1264; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1266 = 10'h129 == _T_40[9:0] ? 4'hd : _GEN_1265; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1267 = 10'h12a == _T_40[9:0] ? 4'hc : _GEN_1266; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1268 = 10'h12b == _T_40[9:0] ? 4'hb : _GEN_1267; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1269 = 10'h12c == _T_40[9:0] ? 4'hc : _GEN_1268; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1270 = 10'h12d == _T_40[9:0] ? 4'hb : _GEN_1269; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1271 = 10'h12e == _T_40[9:0] ? 4'ha : _GEN_1270; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1272 = 10'h12f == _T_40[9:0] ? 4'h6 : _GEN_1271; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1273 = 10'h130 == _T_40[9:0] ? 4'he : _GEN_1272; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1274 = 10'h131 == _T_40[9:0] ? 4'hc : _GEN_1273; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1275 = 10'h132 == _T_40[9:0] ? 4'ha : _GEN_1274; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1276 = 10'h133 == _T_40[9:0] ? 4'h9 : _GEN_1275; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1277 = 10'h134 == _T_40[9:0] ? 4'hb : _GEN_1276; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1278 = 10'h135 == _T_40[9:0] ? 4'h8 : _GEN_1277; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1279 = 10'h136 == _T_40[9:0] ? 4'h8 : _GEN_1278; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1280 = 10'h137 == _T_40[9:0] ? 4'h4 : _GEN_1279; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1281 = 10'h138 == _T_40[9:0] ? 4'h7 : _GEN_1280; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1282 = 10'h139 == _T_40[9:0] ? 4'h0 : _GEN_1281; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1283 = 10'h13a == _T_40[9:0] ? 4'h0 : _GEN_1282; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1284 = 10'h13b == _T_40[9:0] ? 4'h0 : _GEN_1283; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1285 = 10'h13c == _T_40[9:0] ? 4'h0 : _GEN_1284; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1286 = 10'h13d == _T_40[9:0] ? 4'h0 : _GEN_1285; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1287 = 10'h13e == _T_40[9:0] ? 4'h4 : _GEN_1286; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1288 = 10'h13f == _T_40[9:0] ? 4'hc : _GEN_1287; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1289 = 10'h140 == _T_40[9:0] ? 4'he : _GEN_1288; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1290 = 10'h141 == _T_40[9:0] ? 4'he : _GEN_1289; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1291 = 10'h142 == _T_40[9:0] ? 4'he : _GEN_1290; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1292 = 10'h143 == _T_40[9:0] ? 4'hc : _GEN_1291; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1293 = 10'h144 == _T_40[9:0] ? 4'hd : _GEN_1292; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1294 = 10'h145 == _T_40[9:0] ? 4'hb : _GEN_1293; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1295 = 10'h146 == _T_40[9:0] ? 4'hb : _GEN_1294; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1296 = 10'h147 == _T_40[9:0] ? 4'ha : _GEN_1295; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1297 = 10'h148 == _T_40[9:0] ? 4'ha : _GEN_1296; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1298 = 10'h149 == _T_40[9:0] ? 4'hc : _GEN_1297; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1299 = 10'h14a == _T_40[9:0] ? 4'hd : _GEN_1298; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1300 = 10'h14b == _T_40[9:0] ? 4'hc : _GEN_1299; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1301 = 10'h14c == _T_40[9:0] ? 4'hd : _GEN_1300; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1302 = 10'h14d == _T_40[9:0] ? 4'h9 : _GEN_1301; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1303 = 10'h14e == _T_40[9:0] ? 4'h7 : _GEN_1302; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1304 = 10'h14f == _T_40[9:0] ? 4'ha : _GEN_1303; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1305 = 10'h150 == _T_40[9:0] ? 4'ha : _GEN_1304; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1306 = 10'h151 == _T_40[9:0] ? 4'hb : _GEN_1305; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1307 = 10'h152 == _T_40[9:0] ? 4'hb : _GEN_1306; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1308 = 10'h153 == _T_40[9:0] ? 4'hc : _GEN_1307; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1309 = 10'h154 == _T_40[9:0] ? 4'hb : _GEN_1308; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1310 = 10'h155 == _T_40[9:0] ? 4'h6 : _GEN_1309; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1311 = 10'h156 == _T_40[9:0] ? 4'hb : _GEN_1310; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1312 = 10'h157 == _T_40[9:0] ? 4'h7 : _GEN_1311; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1313 = 10'h158 == _T_40[9:0] ? 4'h7 : _GEN_1312; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1314 = 10'h159 == _T_40[9:0] ? 4'h7 : _GEN_1313; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1315 = 10'h15a == _T_40[9:0] ? 4'h7 : _GEN_1314; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1316 = 10'h15b == _T_40[9:0] ? 4'h7 : _GEN_1315; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1317 = 10'h15c == _T_40[9:0] ? 4'h7 : _GEN_1316; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1318 = 10'h15d == _T_40[9:0] ? 4'h6 : _GEN_1317; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1319 = 10'h15e == _T_40[9:0] ? 4'h7 : _GEN_1318; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1320 = 10'h15f == _T_40[9:0] ? 4'h0 : _GEN_1319; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1321 = 10'h160 == _T_40[9:0] ? 4'h0 : _GEN_1320; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1322 = 10'h161 == _T_40[9:0] ? 4'h0 : _GEN_1321; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1323 = 10'h162 == _T_40[9:0] ? 4'h0 : _GEN_1322; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1324 = 10'h163 == _T_40[9:0] ? 4'h2 : _GEN_1323; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1325 = 10'h164 == _T_40[9:0] ? 4'h4 : _GEN_1324; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1326 = 10'h165 == _T_40[9:0] ? 4'hb : _GEN_1325; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1327 = 10'h166 == _T_40[9:0] ? 4'hb : _GEN_1326; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1328 = 10'h167 == _T_40[9:0] ? 4'he : _GEN_1327; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1329 = 10'h168 == _T_40[9:0] ? 4'he : _GEN_1328; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1330 = 10'h169 == _T_40[9:0] ? 4'hc : _GEN_1329; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1331 = 10'h16a == _T_40[9:0] ? 4'hd : _GEN_1330; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1332 = 10'h16b == _T_40[9:0] ? 4'hd : _GEN_1331; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1333 = 10'h16c == _T_40[9:0] ? 4'ha : _GEN_1332; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1334 = 10'h16d == _T_40[9:0] ? 4'ha : _GEN_1333; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1335 = 10'h16e == _T_40[9:0] ? 4'ha : _GEN_1334; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1336 = 10'h16f == _T_40[9:0] ? 4'hd : _GEN_1335; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1337 = 10'h170 == _T_40[9:0] ? 4'hd : _GEN_1336; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1338 = 10'h171 == _T_40[9:0] ? 4'hd : _GEN_1337; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1339 = 10'h172 == _T_40[9:0] ? 4'he : _GEN_1338; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1340 = 10'h173 == _T_40[9:0] ? 4'h8 : _GEN_1339; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1341 = 10'h174 == _T_40[9:0] ? 4'h5 : _GEN_1340; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1342 = 10'h175 == _T_40[9:0] ? 4'h6 : _GEN_1341; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1343 = 10'h176 == _T_40[9:0] ? 4'h6 : _GEN_1342; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1344 = 10'h177 == _T_40[9:0] ? 4'h6 : _GEN_1343; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1345 = 10'h178 == _T_40[9:0] ? 4'h7 : _GEN_1344; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1346 = 10'h179 == _T_40[9:0] ? 4'h9 : _GEN_1345; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1347 = 10'h17a == _T_40[9:0] ? 4'h9 : _GEN_1346; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1348 = 10'h17b == _T_40[9:0] ? 4'h6 : _GEN_1347; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1349 = 10'h17c == _T_40[9:0] ? 4'h7 : _GEN_1348; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1350 = 10'h17d == _T_40[9:0] ? 4'h7 : _GEN_1349; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1351 = 10'h17e == _T_40[9:0] ? 4'h7 : _GEN_1350; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1352 = 10'h17f == _T_40[9:0] ? 4'h7 : _GEN_1351; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1353 = 10'h180 == _T_40[9:0] ? 4'h7 : _GEN_1352; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1354 = 10'h181 == _T_40[9:0] ? 4'h7 : _GEN_1353; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1355 = 10'h182 == _T_40[9:0] ? 4'h8 : _GEN_1354; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1356 = 10'h183 == _T_40[9:0] ? 4'h8 : _GEN_1355; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1357 = 10'h184 == _T_40[9:0] ? 4'h8 : _GEN_1356; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1358 = 10'h185 == _T_40[9:0] ? 4'h7 : _GEN_1357; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1359 = 10'h186 == _T_40[9:0] ? 4'h1 : _GEN_1358; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1360 = 10'h187 == _T_40[9:0] ? 4'h0 : _GEN_1359; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1361 = 10'h188 == _T_40[9:0] ? 4'h0 : _GEN_1360; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1362 = 10'h189 == _T_40[9:0] ? 4'h4 : _GEN_1361; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1363 = 10'h18a == _T_40[9:0] ? 4'h4 : _GEN_1362; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1364 = 10'h18b == _T_40[9:0] ? 4'hb : _GEN_1363; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1365 = 10'h18c == _T_40[9:0] ? 4'hb : _GEN_1364; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1366 = 10'h18d == _T_40[9:0] ? 4'hc : _GEN_1365; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1367 = 10'h18e == _T_40[9:0] ? 4'he : _GEN_1366; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1368 = 10'h18f == _T_40[9:0] ? 4'hb : _GEN_1367; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1369 = 10'h190 == _T_40[9:0] ? 4'hd : _GEN_1368; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1370 = 10'h191 == _T_40[9:0] ? 4'hc : _GEN_1369; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1371 = 10'h192 == _T_40[9:0] ? 4'h9 : _GEN_1370; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1372 = 10'h193 == _T_40[9:0] ? 4'ha : _GEN_1371; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1373 = 10'h194 == _T_40[9:0] ? 4'h9 : _GEN_1372; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1374 = 10'h195 == _T_40[9:0] ? 4'hd : _GEN_1373; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1375 = 10'h196 == _T_40[9:0] ? 4'hd : _GEN_1374; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1376 = 10'h197 == _T_40[9:0] ? 4'hb : _GEN_1375; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1377 = 10'h198 == _T_40[9:0] ? 4'he : _GEN_1376; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1378 = 10'h199 == _T_40[9:0] ? 4'h5 : _GEN_1377; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1379 = 10'h19a == _T_40[9:0] ? 4'h1 : _GEN_1378; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1380 = 10'h19b == _T_40[9:0] ? 4'h3 : _GEN_1379; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1381 = 10'h19c == _T_40[9:0] ? 4'h6 : _GEN_1380; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1382 = 10'h19d == _T_40[9:0] ? 4'h4 : _GEN_1381; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1383 = 10'h19e == _T_40[9:0] ? 4'h1 : _GEN_1382; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1384 = 10'h19f == _T_40[9:0] ? 4'h3 : _GEN_1383; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1385 = 10'h1a0 == _T_40[9:0] ? 4'h6 : _GEN_1384; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1386 = 10'h1a1 == _T_40[9:0] ? 4'h6 : _GEN_1385; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1387 = 10'h1a2 == _T_40[9:0] ? 4'h7 : _GEN_1386; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1388 = 10'h1a3 == _T_40[9:0] ? 4'h7 : _GEN_1387; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1389 = 10'h1a4 == _T_40[9:0] ? 4'h7 : _GEN_1388; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1390 = 10'h1a5 == _T_40[9:0] ? 4'h7 : _GEN_1389; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1391 = 10'h1a6 == _T_40[9:0] ? 4'h7 : _GEN_1390; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1392 = 10'h1a7 == _T_40[9:0] ? 4'h7 : _GEN_1391; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1393 = 10'h1a8 == _T_40[9:0] ? 4'h8 : _GEN_1392; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1394 = 10'h1a9 == _T_40[9:0] ? 4'h8 : _GEN_1393; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1395 = 10'h1aa == _T_40[9:0] ? 4'h7 : _GEN_1394; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1396 = 10'h1ab == _T_40[9:0] ? 4'h8 : _GEN_1395; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1397 = 10'h1ac == _T_40[9:0] ? 4'h8 : _GEN_1396; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1398 = 10'h1ad == _T_40[9:0] ? 4'h3 : _GEN_1397; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1399 = 10'h1ae == _T_40[9:0] ? 4'h2 : _GEN_1398; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1400 = 10'h1af == _T_40[9:0] ? 4'h8 : _GEN_1399; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1401 = 10'h1b0 == _T_40[9:0] ? 4'h6 : _GEN_1400; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1402 = 10'h1b1 == _T_40[9:0] ? 4'hb : _GEN_1401; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1403 = 10'h1b2 == _T_40[9:0] ? 4'hb : _GEN_1402; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1404 = 10'h1b3 == _T_40[9:0] ? 4'ha : _GEN_1403; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1405 = 10'h1b4 == _T_40[9:0] ? 4'he : _GEN_1404; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1406 = 10'h1b5 == _T_40[9:0] ? 4'hb : _GEN_1405; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1407 = 10'h1b6 == _T_40[9:0] ? 4'hc : _GEN_1406; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1408 = 10'h1b7 == _T_40[9:0] ? 4'ha : _GEN_1407; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1409 = 10'h1b8 == _T_40[9:0] ? 4'h9 : _GEN_1408; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1410 = 10'h1b9 == _T_40[9:0] ? 4'h9 : _GEN_1409; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1411 = 10'h1ba == _T_40[9:0] ? 4'h9 : _GEN_1410; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1412 = 10'h1bb == _T_40[9:0] ? 4'hb : _GEN_1411; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1413 = 10'h1bc == _T_40[9:0] ? 4'hd : _GEN_1412; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1414 = 10'h1bd == _T_40[9:0] ? 4'hd : _GEN_1413; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1415 = 10'h1be == _T_40[9:0] ? 4'he : _GEN_1414; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1416 = 10'h1bf == _T_40[9:0] ? 4'h7 : _GEN_1415; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1417 = 10'h1c0 == _T_40[9:0] ? 4'h6 : _GEN_1416; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1418 = 10'h1c1 == _T_40[9:0] ? 4'h6 : _GEN_1417; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1419 = 10'h1c2 == _T_40[9:0] ? 4'h5 : _GEN_1418; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1420 = 10'h1c3 == _T_40[9:0] ? 4'h5 : _GEN_1419; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1421 = 10'h1c4 == _T_40[9:0] ? 4'h4 : _GEN_1420; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1422 = 10'h1c5 == _T_40[9:0] ? 4'h5 : _GEN_1421; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1423 = 10'h1c6 == _T_40[9:0] ? 4'h6 : _GEN_1422; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1424 = 10'h1c7 == _T_40[9:0] ? 4'h6 : _GEN_1423; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1425 = 10'h1c8 == _T_40[9:0] ? 4'h7 : _GEN_1424; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1426 = 10'h1c9 == _T_40[9:0] ? 4'h7 : _GEN_1425; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1427 = 10'h1ca == _T_40[9:0] ? 4'h7 : _GEN_1426; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1428 = 10'h1cb == _T_40[9:0] ? 4'h7 : _GEN_1427; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1429 = 10'h1cc == _T_40[9:0] ? 4'h7 : _GEN_1428; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1430 = 10'h1cd == _T_40[9:0] ? 4'h8 : _GEN_1429; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1431 = 10'h1ce == _T_40[9:0] ? 4'h8 : _GEN_1430; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1432 = 10'h1cf == _T_40[9:0] ? 4'h8 : _GEN_1431; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1433 = 10'h1d0 == _T_40[9:0] ? 4'h5 : _GEN_1432; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1434 = 10'h1d1 == _T_40[9:0] ? 4'h8 : _GEN_1433; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1435 = 10'h1d2 == _T_40[9:0] ? 4'h8 : _GEN_1434; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1436 = 10'h1d3 == _T_40[9:0] ? 4'h8 : _GEN_1435; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1437 = 10'h1d4 == _T_40[9:0] ? 4'h8 : _GEN_1436; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1438 = 10'h1d5 == _T_40[9:0] ? 4'h7 : _GEN_1437; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1439 = 10'h1d6 == _T_40[9:0] ? 4'h9 : _GEN_1438; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1440 = 10'h1d7 == _T_40[9:0] ? 4'hb : _GEN_1439; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1441 = 10'h1d8 == _T_40[9:0] ? 4'hb : _GEN_1440; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1442 = 10'h1d9 == _T_40[9:0] ? 4'hb : _GEN_1441; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1443 = 10'h1da == _T_40[9:0] ? 4'ha : _GEN_1442; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1444 = 10'h1db == _T_40[9:0] ? 4'hc : _GEN_1443; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1445 = 10'h1dc == _T_40[9:0] ? 4'hb : _GEN_1444; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1446 = 10'h1dd == _T_40[9:0] ? 4'h5 : _GEN_1445; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1447 = 10'h1de == _T_40[9:0] ? 4'h9 : _GEN_1446; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1448 = 10'h1df == _T_40[9:0] ? 4'h9 : _GEN_1447; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1449 = 10'h1e0 == _T_40[9:0] ? 4'h9 : _GEN_1448; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1450 = 10'h1e1 == _T_40[9:0] ? 4'h7 : _GEN_1449; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1451 = 10'h1e2 == _T_40[9:0] ? 4'hc : _GEN_1450; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1452 = 10'h1e3 == _T_40[9:0] ? 4'hc : _GEN_1451; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1453 = 10'h1e4 == _T_40[9:0] ? 4'hd : _GEN_1452; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1454 = 10'h1e5 == _T_40[9:0] ? 4'h7 : _GEN_1453; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1455 = 10'h1e6 == _T_40[9:0] ? 4'h6 : _GEN_1454; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1456 = 10'h1e7 == _T_40[9:0] ? 4'h6 : _GEN_1455; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1457 = 10'h1e8 == _T_40[9:0] ? 4'h6 : _GEN_1456; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1458 = 10'h1e9 == _T_40[9:0] ? 4'h6 : _GEN_1457; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1459 = 10'h1ea == _T_40[9:0] ? 4'h6 : _GEN_1458; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1460 = 10'h1eb == _T_40[9:0] ? 4'h6 : _GEN_1459; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1461 = 10'h1ec == _T_40[9:0] ? 4'h6 : _GEN_1460; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1462 = 10'h1ed == _T_40[9:0] ? 4'h8 : _GEN_1461; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1463 = 10'h1ee == _T_40[9:0] ? 4'h7 : _GEN_1462; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1464 = 10'h1ef == _T_40[9:0] ? 4'h7 : _GEN_1463; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1465 = 10'h1f0 == _T_40[9:0] ? 4'h7 : _GEN_1464; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1466 = 10'h1f1 == _T_40[9:0] ? 4'h7 : _GEN_1465; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1467 = 10'h1f2 == _T_40[9:0] ? 4'h7 : _GEN_1466; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1468 = 10'h1f3 == _T_40[9:0] ? 4'h8 : _GEN_1467; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1469 = 10'h1f4 == _T_40[9:0] ? 4'h8 : _GEN_1468; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1470 = 10'h1f5 == _T_40[9:0] ? 4'h8 : _GEN_1469; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1471 = 10'h1f6 == _T_40[9:0] ? 4'ha : _GEN_1470; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1472 = 10'h1f7 == _T_40[9:0] ? 4'h8 : _GEN_1471; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1473 = 10'h1f8 == _T_40[9:0] ? 4'h8 : _GEN_1472; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1474 = 10'h1f9 == _T_40[9:0] ? 4'h9 : _GEN_1473; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1475 = 10'h1fa == _T_40[9:0] ? 4'h9 : _GEN_1474; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1476 = 10'h1fb == _T_40[9:0] ? 4'h8 : _GEN_1475; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1477 = 10'h1fc == _T_40[9:0] ? 4'hb : _GEN_1476; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1478 = 10'h1fd == _T_40[9:0] ? 4'hb : _GEN_1477; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1479 = 10'h1fe == _T_40[9:0] ? 4'hb : _GEN_1478; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1480 = 10'h1ff == _T_40[9:0] ? 4'ha : _GEN_1479; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1481 = 10'h200 == _T_40[9:0] ? 4'h3 : _GEN_1480; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1482 = 10'h201 == _T_40[9:0] ? 4'h9 : _GEN_1481; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1483 = 10'h202 == _T_40[9:0] ? 4'h5 : _GEN_1482; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1484 = 10'h203 == _T_40[9:0] ? 4'h3 : _GEN_1483; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1485 = 10'h204 == _T_40[9:0] ? 4'h4 : _GEN_1484; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1486 = 10'h205 == _T_40[9:0] ? 4'h4 : _GEN_1485; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1487 = 10'h206 == _T_40[9:0] ? 4'h4 : _GEN_1486; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1488 = 10'h207 == _T_40[9:0] ? 4'h4 : _GEN_1487; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1489 = 10'h208 == _T_40[9:0] ? 4'h8 : _GEN_1488; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1490 = 10'h209 == _T_40[9:0] ? 4'hc : _GEN_1489; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1491 = 10'h20a == _T_40[9:0] ? 4'hd : _GEN_1490; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1492 = 10'h20b == _T_40[9:0] ? 4'h7 : _GEN_1491; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1493 = 10'h20c == _T_40[9:0] ? 4'h6 : _GEN_1492; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1494 = 10'h20d == _T_40[9:0] ? 4'h6 : _GEN_1493; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1495 = 10'h20e == _T_40[9:0] ? 4'h6 : _GEN_1494; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1496 = 10'h20f == _T_40[9:0] ? 4'h5 : _GEN_1495; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1497 = 10'h210 == _T_40[9:0] ? 4'h6 : _GEN_1496; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1498 = 10'h211 == _T_40[9:0] ? 4'h6 : _GEN_1497; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1499 = 10'h212 == _T_40[9:0] ? 4'h7 : _GEN_1498; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1500 = 10'h213 == _T_40[9:0] ? 4'ha : _GEN_1499; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1501 = 10'h214 == _T_40[9:0] ? 4'h6 : _GEN_1500; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1502 = 10'h215 == _T_40[9:0] ? 4'h7 : _GEN_1501; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1503 = 10'h216 == _T_40[9:0] ? 4'h7 : _GEN_1502; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1504 = 10'h217 == _T_40[9:0] ? 4'h7 : _GEN_1503; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1505 = 10'h218 == _T_40[9:0] ? 4'h7 : _GEN_1504; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1506 = 10'h219 == _T_40[9:0] ? 4'h8 : _GEN_1505; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1507 = 10'h21a == _T_40[9:0] ? 4'h7 : _GEN_1506; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1508 = 10'h21b == _T_40[9:0] ? 4'h8 : _GEN_1507; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1509 = 10'h21c == _T_40[9:0] ? 4'hb : _GEN_1508; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1510 = 10'h21d == _T_40[9:0] ? 4'ha : _GEN_1509; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1511 = 10'h21e == _T_40[9:0] ? 4'h9 : _GEN_1510; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1512 = 10'h21f == _T_40[9:0] ? 4'h9 : _GEN_1511; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1513 = 10'h220 == _T_40[9:0] ? 4'h8 : _GEN_1512; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1514 = 10'h221 == _T_40[9:0] ? 4'h9 : _GEN_1513; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1515 = 10'h222 == _T_40[9:0] ? 4'hb : _GEN_1514; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1516 = 10'h223 == _T_40[9:0] ? 4'hb : _GEN_1515; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1517 = 10'h224 == _T_40[9:0] ? 4'hb : _GEN_1516; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1518 = 10'h225 == _T_40[9:0] ? 4'h8 : _GEN_1517; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1519 = 10'h226 == _T_40[9:0] ? 4'h1 : _GEN_1518; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1520 = 10'h227 == _T_40[9:0] ? 4'h3 : _GEN_1519; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1521 = 10'h228 == _T_40[9:0] ? 4'h3 : _GEN_1520; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1522 = 10'h229 == _T_40[9:0] ? 4'h3 : _GEN_1521; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1523 = 10'h22a == _T_40[9:0] ? 4'h3 : _GEN_1522; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1524 = 10'h22b == _T_40[9:0] ? 4'h3 : _GEN_1523; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1525 = 10'h22c == _T_40[9:0] ? 4'h3 : _GEN_1524; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1526 = 10'h22d == _T_40[9:0] ? 4'h3 : _GEN_1525; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1527 = 10'h22e == _T_40[9:0] ? 4'h3 : _GEN_1526; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1528 = 10'h22f == _T_40[9:0] ? 4'h9 : _GEN_1527; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1529 = 10'h230 == _T_40[9:0] ? 4'h6 : _GEN_1528; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1530 = 10'h231 == _T_40[9:0] ? 4'h7 : _GEN_1529; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1531 = 10'h232 == _T_40[9:0] ? 4'h6 : _GEN_1530; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1532 = 10'h233 == _T_40[9:0] ? 4'h7 : _GEN_1531; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1533 = 10'h234 == _T_40[9:0] ? 4'h7 : _GEN_1532; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1534 = 10'h235 == _T_40[9:0] ? 4'h6 : _GEN_1533; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1535 = 10'h236 == _T_40[9:0] ? 4'h6 : _GEN_1534; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1536 = 10'h237 == _T_40[9:0] ? 4'h6 : _GEN_1535; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1537 = 10'h238 == _T_40[9:0] ? 4'h6 : _GEN_1536; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1538 = 10'h239 == _T_40[9:0] ? 4'h8 : _GEN_1537; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1539 = 10'h23a == _T_40[9:0] ? 4'h6 : _GEN_1538; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1540 = 10'h23b == _T_40[9:0] ? 4'h7 : _GEN_1539; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1541 = 10'h23c == _T_40[9:0] ? 4'h7 : _GEN_1540; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1542 = 10'h23d == _T_40[9:0] ? 4'h7 : _GEN_1541; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1543 = 10'h23e == _T_40[9:0] ? 4'h7 : _GEN_1542; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1544 = 10'h23f == _T_40[9:0] ? 4'h7 : _GEN_1543; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1545 = 10'h240 == _T_40[9:0] ? 4'h7 : _GEN_1544; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1546 = 10'h241 == _T_40[9:0] ? 4'h8 : _GEN_1545; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1547 = 10'h242 == _T_40[9:0] ? 4'hb : _GEN_1546; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1548 = 10'h243 == _T_40[9:0] ? 4'hb : _GEN_1547; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1549 = 10'h244 == _T_40[9:0] ? 4'hb : _GEN_1548; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1550 = 10'h245 == _T_40[9:0] ? 4'ha : _GEN_1549; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1551 = 10'h246 == _T_40[9:0] ? 4'h9 : _GEN_1550; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1552 = 10'h247 == _T_40[9:0] ? 4'ha : _GEN_1551; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1553 = 10'h248 == _T_40[9:0] ? 4'hb : _GEN_1552; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1554 = 10'h249 == _T_40[9:0] ? 4'hb : _GEN_1553; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1555 = 10'h24a == _T_40[9:0] ? 4'ha : _GEN_1554; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1556 = 10'h24b == _T_40[9:0] ? 4'h2 : _GEN_1555; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1557 = 10'h24c == _T_40[9:0] ? 4'h0 : _GEN_1556; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1558 = 10'h24d == _T_40[9:0] ? 4'h2 : _GEN_1557; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1559 = 10'h24e == _T_40[9:0] ? 4'h3 : _GEN_1558; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1560 = 10'h24f == _T_40[9:0] ? 4'h3 : _GEN_1559; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1561 = 10'h250 == _T_40[9:0] ? 4'h3 : _GEN_1560; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1562 = 10'h251 == _T_40[9:0] ? 4'h3 : _GEN_1561; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1563 = 10'h252 == _T_40[9:0] ? 4'h3 : _GEN_1562; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1564 = 10'h253 == _T_40[9:0] ? 4'h3 : _GEN_1563; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1565 = 10'h254 == _T_40[9:0] ? 4'h3 : _GEN_1564; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1566 = 10'h255 == _T_40[9:0] ? 4'h5 : _GEN_1565; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1567 = 10'h256 == _T_40[9:0] ? 4'h6 : _GEN_1566; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1568 = 10'h257 == _T_40[9:0] ? 4'h8 : _GEN_1567; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1569 = 10'h258 == _T_40[9:0] ? 4'h5 : _GEN_1568; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1570 = 10'h259 == _T_40[9:0] ? 4'h6 : _GEN_1569; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1571 = 10'h25a == _T_40[9:0] ? 4'h6 : _GEN_1570; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1572 = 10'h25b == _T_40[9:0] ? 4'h5 : _GEN_1571; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1573 = 10'h25c == _T_40[9:0] ? 4'h6 : _GEN_1572; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1574 = 10'h25d == _T_40[9:0] ? 4'h6 : _GEN_1573; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1575 = 10'h25e == _T_40[9:0] ? 4'h9 : _GEN_1574; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1576 = 10'h25f == _T_40[9:0] ? 4'hc : _GEN_1575; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1577 = 10'h260 == _T_40[9:0] ? 4'h7 : _GEN_1576; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1578 = 10'h261 == _T_40[9:0] ? 4'h9 : _GEN_1577; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1579 = 10'h262 == _T_40[9:0] ? 4'ha : _GEN_1578; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1580 = 10'h263 == _T_40[9:0] ? 4'h8 : _GEN_1579; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1581 = 10'h264 == _T_40[9:0] ? 4'ha : _GEN_1580; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1582 = 10'h265 == _T_40[9:0] ? 4'h9 : _GEN_1581; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1583 = 10'h266 == _T_40[9:0] ? 4'h8 : _GEN_1582; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1584 = 10'h267 == _T_40[9:0] ? 4'h8 : _GEN_1583; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1585 = 10'h268 == _T_40[9:0] ? 4'ha : _GEN_1584; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1586 = 10'h269 == _T_40[9:0] ? 4'ha : _GEN_1585; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1587 = 10'h26a == _T_40[9:0] ? 4'hb : _GEN_1586; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1588 = 10'h26b == _T_40[9:0] ? 4'hb : _GEN_1587; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1589 = 10'h26c == _T_40[9:0] ? 4'hb : _GEN_1588; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1590 = 10'h26d == _T_40[9:0] ? 4'hb : _GEN_1589; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1591 = 10'h26e == _T_40[9:0] ? 4'hb : _GEN_1590; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1592 = 10'h26f == _T_40[9:0] ? 4'ha : _GEN_1591; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1593 = 10'h270 == _T_40[9:0] ? 4'h3 : _GEN_1592; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1594 = 10'h271 == _T_40[9:0] ? 4'h0 : _GEN_1593; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1595 = 10'h272 == _T_40[9:0] ? 4'h0 : _GEN_1594; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1596 = 10'h273 == _T_40[9:0] ? 4'h2 : _GEN_1595; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1597 = 10'h274 == _T_40[9:0] ? 4'h3 : _GEN_1596; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1598 = 10'h275 == _T_40[9:0] ? 4'h3 : _GEN_1597; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1599 = 10'h276 == _T_40[9:0] ? 4'h3 : _GEN_1598; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1600 = 10'h277 == _T_40[9:0] ? 4'h3 : _GEN_1599; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1601 = 10'h278 == _T_40[9:0] ? 4'h3 : _GEN_1600; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1602 = 10'h279 == _T_40[9:0] ? 4'h3 : _GEN_1601; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1603 = 10'h27a == _T_40[9:0] ? 4'h3 : _GEN_1602; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1604 = 10'h27b == _T_40[9:0] ? 4'h6 : _GEN_1603; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1605 = 10'h27c == _T_40[9:0] ? 4'h7 : _GEN_1604; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1606 = 10'h27d == _T_40[9:0] ? 4'h7 : _GEN_1605; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1607 = 10'h27e == _T_40[9:0] ? 4'h4 : _GEN_1606; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1608 = 10'h27f == _T_40[9:0] ? 4'h6 : _GEN_1607; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1609 = 10'h280 == _T_40[9:0] ? 4'h6 : _GEN_1608; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1610 = 10'h281 == _T_40[9:0] ? 4'h6 : _GEN_1609; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1611 = 10'h282 == _T_40[9:0] ? 4'h6 : _GEN_1610; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1612 = 10'h283 == _T_40[9:0] ? 4'ha : _GEN_1611; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1613 = 10'h284 == _T_40[9:0] ? 4'hc : _GEN_1612; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1614 = 10'h285 == _T_40[9:0] ? 4'hc : _GEN_1613; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1615 = 10'h286 == _T_40[9:0] ? 4'h8 : _GEN_1614; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1616 = 10'h287 == _T_40[9:0] ? 4'ha : _GEN_1615; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1617 = 10'h288 == _T_40[9:0] ? 4'ha : _GEN_1616; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1618 = 10'h289 == _T_40[9:0] ? 4'ha : _GEN_1617; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1619 = 10'h28a == _T_40[9:0] ? 4'hc : _GEN_1618; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1620 = 10'h28b == _T_40[9:0] ? 4'hb : _GEN_1619; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1621 = 10'h28c == _T_40[9:0] ? 4'ha : _GEN_1620; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1622 = 10'h28d == _T_40[9:0] ? 4'h7 : _GEN_1621; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1623 = 10'h28e == _T_40[9:0] ? 4'h2 : _GEN_1622; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1624 = 10'h28f == _T_40[9:0] ? 4'h5 : _GEN_1623; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1625 = 10'h290 == _T_40[9:0] ? 4'h8 : _GEN_1624; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1626 = 10'h291 == _T_40[9:0] ? 4'ha : _GEN_1625; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1627 = 10'h292 == _T_40[9:0] ? 4'ha : _GEN_1626; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1628 = 10'h293 == _T_40[9:0] ? 4'ha : _GEN_1627; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1629 = 10'h294 == _T_40[9:0] ? 4'h9 : _GEN_1628; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1630 = 10'h295 == _T_40[9:0] ? 4'h3 : _GEN_1629; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1631 = 10'h296 == _T_40[9:0] ? 4'h0 : _GEN_1630; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1632 = 10'h297 == _T_40[9:0] ? 4'h0 : _GEN_1631; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1633 = 10'h298 == _T_40[9:0] ? 4'h0 : _GEN_1632; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1634 = 10'h299 == _T_40[9:0] ? 4'h1 : _GEN_1633; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1635 = 10'h29a == _T_40[9:0] ? 4'h3 : _GEN_1634; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1636 = 10'h29b == _T_40[9:0] ? 4'h3 : _GEN_1635; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1637 = 10'h29c == _T_40[9:0] ? 4'h3 : _GEN_1636; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1638 = 10'h29d == _T_40[9:0] ? 4'h3 : _GEN_1637; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1639 = 10'h29e == _T_40[9:0] ? 4'h3 : _GEN_1638; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1640 = 10'h29f == _T_40[9:0] ? 4'h3 : _GEN_1639; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1641 = 10'h2a0 == _T_40[9:0] ? 4'h4 : _GEN_1640; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1642 = 10'h2a1 == _T_40[9:0] ? 4'h6 : _GEN_1641; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1643 = 10'h2a2 == _T_40[9:0] ? 4'h7 : _GEN_1642; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1644 = 10'h2a3 == _T_40[9:0] ? 4'h6 : _GEN_1643; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1645 = 10'h2a4 == _T_40[9:0] ? 4'h4 : _GEN_1644; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1646 = 10'h2a5 == _T_40[9:0] ? 4'h6 : _GEN_1645; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1647 = 10'h2a6 == _T_40[9:0] ? 4'h6 : _GEN_1646; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1648 = 10'h2a7 == _T_40[9:0] ? 4'h7 : _GEN_1647; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1649 = 10'h2a8 == _T_40[9:0] ? 4'ha : _GEN_1648; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1650 = 10'h2a9 == _T_40[9:0] ? 4'hb : _GEN_1649; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1651 = 10'h2aa == _T_40[9:0] ? 4'hb : _GEN_1650; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1652 = 10'h2ab == _T_40[9:0] ? 4'hb : _GEN_1651; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1653 = 10'h2ac == _T_40[9:0] ? 4'h8 : _GEN_1652; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1654 = 10'h2ad == _T_40[9:0] ? 4'hb : _GEN_1653; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1655 = 10'h2ae == _T_40[9:0] ? 4'ha : _GEN_1654; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1656 = 10'h2af == _T_40[9:0] ? 4'hb : _GEN_1655; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1657 = 10'h2b0 == _T_40[9:0] ? 4'hc : _GEN_1656; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1658 = 10'h2b1 == _T_40[9:0] ? 4'hb : _GEN_1657; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1659 = 10'h2b2 == _T_40[9:0] ? 4'ha : _GEN_1658; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1660 = 10'h2b3 == _T_40[9:0] ? 4'h6 : _GEN_1659; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1661 = 10'h2b4 == _T_40[9:0] ? 4'h0 : _GEN_1660; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1662 = 10'h2b5 == _T_40[9:0] ? 4'h0 : _GEN_1661; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1663 = 10'h2b6 == _T_40[9:0] ? 4'h0 : _GEN_1662; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1664 = 10'h2b7 == _T_40[9:0] ? 4'h1 : _GEN_1663; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1665 = 10'h2b8 == _T_40[9:0] ? 4'h5 : _GEN_1664; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1666 = 10'h2b9 == _T_40[9:0] ? 4'h9 : _GEN_1665; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1667 = 10'h2ba == _T_40[9:0] ? 4'h1 : _GEN_1666; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1668 = 10'h2bb == _T_40[9:0] ? 4'h0 : _GEN_1667; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1669 = 10'h2bc == _T_40[9:0] ? 4'h0 : _GEN_1668; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1670 = 10'h2bd == _T_40[9:0] ? 4'h0 : _GEN_1669; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1671 = 10'h2be == _T_40[9:0] ? 4'h0 : _GEN_1670; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1672 = 10'h2bf == _T_40[9:0] ? 4'h0 : _GEN_1671; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1673 = 10'h2c0 == _T_40[9:0] ? 4'h3 : _GEN_1672; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1674 = 10'h2c1 == _T_40[9:0] ? 4'h3 : _GEN_1673; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1675 = 10'h2c2 == _T_40[9:0] ? 4'h3 : _GEN_1674; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1676 = 10'h2c3 == _T_40[9:0] ? 4'h3 : _GEN_1675; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1677 = 10'h2c4 == _T_40[9:0] ? 4'h3 : _GEN_1676; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1678 = 10'h2c5 == _T_40[9:0] ? 4'h3 : _GEN_1677; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1679 = 10'h2c6 == _T_40[9:0] ? 4'h4 : _GEN_1678; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1680 = 10'h2c7 == _T_40[9:0] ? 4'h5 : _GEN_1679; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1681 = 10'h2c8 == _T_40[9:0] ? 4'h7 : _GEN_1680; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1682 = 10'h2c9 == _T_40[9:0] ? 4'h7 : _GEN_1681; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1683 = 10'h2ca == _T_40[9:0] ? 4'h4 : _GEN_1682; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1684 = 10'h2cb == _T_40[9:0] ? 4'h9 : _GEN_1683; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1685 = 10'h2cc == _T_40[9:0] ? 4'h9 : _GEN_1684; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1686 = 10'h2cd == _T_40[9:0] ? 4'hb : _GEN_1685; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1687 = 10'h2ce == _T_40[9:0] ? 4'hb : _GEN_1686; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1688 = 10'h2cf == _T_40[9:0] ? 4'hb : _GEN_1687; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1689 = 10'h2d0 == _T_40[9:0] ? 4'hb : _GEN_1688; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1690 = 10'h2d1 == _T_40[9:0] ? 4'hb : _GEN_1689; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1691 = 10'h2d2 == _T_40[9:0] ? 4'h8 : _GEN_1690; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1692 = 10'h2d3 == _T_40[9:0] ? 4'ha : _GEN_1691; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1693 = 10'h2d4 == _T_40[9:0] ? 4'hb : _GEN_1692; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1694 = 10'h2d5 == _T_40[9:0] ? 4'ha : _GEN_1693; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1695 = 10'h2d6 == _T_40[9:0] ? 4'ha : _GEN_1694; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1696 = 10'h2d7 == _T_40[9:0] ? 4'ha : _GEN_1695; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1697 = 10'h2d8 == _T_40[9:0] ? 4'ha : _GEN_1696; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1698 = 10'h2d9 == _T_40[9:0] ? 4'h7 : _GEN_1697; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1699 = 10'h2da == _T_40[9:0] ? 4'h2 : _GEN_1698; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1700 = 10'h2db == _T_40[9:0] ? 4'h0 : _GEN_1699; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1701 = 10'h2dc == _T_40[9:0] ? 4'h0 : _GEN_1700; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1702 = 10'h2dd == _T_40[9:0] ? 4'h0 : _GEN_1701; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1703 = 10'h2de == _T_40[9:0] ? 4'h0 : _GEN_1702; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1704 = 10'h2df == _T_40[9:0] ? 4'h2 : _GEN_1703; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1705 = 10'h2e0 == _T_40[9:0] ? 4'h0 : _GEN_1704; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1706 = 10'h2e1 == _T_40[9:0] ? 4'h0 : _GEN_1705; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1707 = 10'h2e2 == _T_40[9:0] ? 4'h0 : _GEN_1706; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1708 = 10'h2e3 == _T_40[9:0] ? 4'h0 : _GEN_1707; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1709 = 10'h2e4 == _T_40[9:0] ? 4'h0 : _GEN_1708; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1710 = 10'h2e5 == _T_40[9:0] ? 4'h0 : _GEN_1709; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1711 = 10'h2e6 == _T_40[9:0] ? 4'h2 : _GEN_1710; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1712 = 10'h2e7 == _T_40[9:0] ? 4'h3 : _GEN_1711; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1713 = 10'h2e8 == _T_40[9:0] ? 4'h3 : _GEN_1712; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1714 = 10'h2e9 == _T_40[9:0] ? 4'h3 : _GEN_1713; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1715 = 10'h2ea == _T_40[9:0] ? 4'h3 : _GEN_1714; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1716 = 10'h2eb == _T_40[9:0] ? 4'h3 : _GEN_1715; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1717 = 10'h2ec == _T_40[9:0] ? 4'h4 : _GEN_1716; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1718 = 10'h2ed == _T_40[9:0] ? 4'h5 : _GEN_1717; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1719 = 10'h2ee == _T_40[9:0] ? 4'h6 : _GEN_1718; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1720 = 10'h2ef == _T_40[9:0] ? 4'h8 : _GEN_1719; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1721 = 10'h2f0 == _T_40[9:0] ? 4'h4 : _GEN_1720; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1722 = 10'h2f1 == _T_40[9:0] ? 4'h9 : _GEN_1721; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1723 = 10'h2f2 == _T_40[9:0] ? 4'hb : _GEN_1722; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1724 = 10'h2f3 == _T_40[9:0] ? 4'hb : _GEN_1723; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1725 = 10'h2f4 == _T_40[9:0] ? 4'hb : _GEN_1724; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1726 = 10'h2f5 == _T_40[9:0] ? 4'hb : _GEN_1725; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1727 = 10'h2f6 == _T_40[9:0] ? 4'hb : _GEN_1726; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1728 = 10'h2f7 == _T_40[9:0] ? 4'hb : _GEN_1727; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1729 = 10'h2f8 == _T_40[9:0] ? 4'h8 : _GEN_1728; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1730 = 10'h2f9 == _T_40[9:0] ? 4'h9 : _GEN_1729; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1731 = 10'h2fa == _T_40[9:0] ? 4'hb : _GEN_1730; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1732 = 10'h2fb == _T_40[9:0] ? 4'hb : _GEN_1731; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1733 = 10'h2fc == _T_40[9:0] ? 4'ha : _GEN_1732; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1734 = 10'h2fd == _T_40[9:0] ? 4'ha : _GEN_1733; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1735 = 10'h2fe == _T_40[9:0] ? 4'h9 : _GEN_1734; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1736 = 10'h2ff == _T_40[9:0] ? 4'h8 : _GEN_1735; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1737 = 10'h300 == _T_40[9:0] ? 4'h8 : _GEN_1736; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1738 = 10'h301 == _T_40[9:0] ? 4'h6 : _GEN_1737; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1739 = 10'h302 == _T_40[9:0] ? 4'h1 : _GEN_1738; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1740 = 10'h303 == _T_40[9:0] ? 4'h0 : _GEN_1739; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1741 = 10'h304 == _T_40[9:0] ? 4'h0 : _GEN_1740; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1742 = 10'h305 == _T_40[9:0] ? 4'h0 : _GEN_1741; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1743 = 10'h306 == _T_40[9:0] ? 4'h0 : _GEN_1742; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1744 = 10'h307 == _T_40[9:0] ? 4'h0 : _GEN_1743; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1745 = 10'h308 == _T_40[9:0] ? 4'h0 : _GEN_1744; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1746 = 10'h309 == _T_40[9:0] ? 4'h0 : _GEN_1745; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1747 = 10'h30a == _T_40[9:0] ? 4'h0 : _GEN_1746; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1748 = 10'h30b == _T_40[9:0] ? 4'h0 : _GEN_1747; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1749 = 10'h30c == _T_40[9:0] ? 4'h2 : _GEN_1748; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1750 = 10'h30d == _T_40[9:0] ? 4'h3 : _GEN_1749; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1751 = 10'h30e == _T_40[9:0] ? 4'h3 : _GEN_1750; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1752 = 10'h30f == _T_40[9:0] ? 4'h3 : _GEN_1751; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1753 = 10'h310 == _T_40[9:0] ? 4'h3 : _GEN_1752; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1754 = 10'h311 == _T_40[9:0] ? 4'h3 : _GEN_1753; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1755 = 10'h312 == _T_40[9:0] ? 4'h4 : _GEN_1754; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1756 = 10'h313 == _T_40[9:0] ? 4'h5 : _GEN_1755; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1757 = 10'h314 == _T_40[9:0] ? 4'h5 : _GEN_1756; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1758 = 10'h315 == _T_40[9:0] ? 4'h8 : _GEN_1757; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1759 = 10'h316 == _T_40[9:0] ? 4'h4 : _GEN_1758; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1760 = 10'h317 == _T_40[9:0] ? 4'h6 : _GEN_1759; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1761 = 10'h318 == _T_40[9:0] ? 4'hb : _GEN_1760; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1762 = 10'h319 == _T_40[9:0] ? 4'hb : _GEN_1761; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1763 = 10'h31a == _T_40[9:0] ? 4'hb : _GEN_1762; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1764 = 10'h31b == _T_40[9:0] ? 4'hb : _GEN_1763; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1765 = 10'h31c == _T_40[9:0] ? 4'hb : _GEN_1764; // @[Filter.scala 230:102]
  wire [3:0] _GEN_1766 = 10'h31d == _T_40[9:0] ? 4'hb : _GEN_1765; // @[Filter.scala 230:102]
  wire [6:0] _GEN_38956 = {{3'd0}, _GEN_1766}; // @[Filter.scala 230:102]
  wire [10:0] _T_47 = _GEN_38956 * 7'h46; // @[Filter.scala 230:102]
  wire [10:0] _GEN_38957 = {{2'd0}, _T_42}; // @[Filter.scala 230:69]
  wire [10:0] _T_49 = _GEN_38957 + _T_47; // @[Filter.scala 230:69]
  wire [3:0] _GEN_1789 = 10'h16 == _T_40[9:0] ? 4'hb : 4'hc; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1790 = 10'h17 == _T_40[9:0] ? 4'h8 : _GEN_1789; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1791 = 10'h18 == _T_40[9:0] ? 4'ha : _GEN_1790; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1792 = 10'h19 == _T_40[9:0] ? 4'hc : _GEN_1791; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1793 = 10'h1a == _T_40[9:0] ? 4'hc : _GEN_1792; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1794 = 10'h1b == _T_40[9:0] ? 4'hc : _GEN_1793; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1795 = 10'h1c == _T_40[9:0] ? 4'hc : _GEN_1794; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1796 = 10'h1d == _T_40[9:0] ? 4'hc : _GEN_1795; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1797 = 10'h1e == _T_40[9:0] ? 4'hc : _GEN_1796; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1798 = 10'h1f == _T_40[9:0] ? 4'hc : _GEN_1797; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1799 = 10'h20 == _T_40[9:0] ? 4'hc : _GEN_1798; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1800 = 10'h21 == _T_40[9:0] ? 4'hc : _GEN_1799; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1801 = 10'h22 == _T_40[9:0] ? 4'hc : _GEN_1800; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1802 = 10'h23 == _T_40[9:0] ? 4'hc : _GEN_1801; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1803 = 10'h24 == _T_40[9:0] ? 4'hc : _GEN_1802; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1804 = 10'h25 == _T_40[9:0] ? 4'hc : _GEN_1803; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1805 = 10'h26 == _T_40[9:0] ? 4'hc : _GEN_1804; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1806 = 10'h27 == _T_40[9:0] ? 4'hc : _GEN_1805; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1807 = 10'h28 == _T_40[9:0] ? 4'hc : _GEN_1806; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1808 = 10'h29 == _T_40[9:0] ? 4'hc : _GEN_1807; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1809 = 10'h2a == _T_40[9:0] ? 4'hc : _GEN_1808; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1810 = 10'h2b == _T_40[9:0] ? 4'hc : _GEN_1809; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1811 = 10'h2c == _T_40[9:0] ? 4'hc : _GEN_1810; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1812 = 10'h2d == _T_40[9:0] ? 4'hc : _GEN_1811; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1813 = 10'h2e == _T_40[9:0] ? 4'hc : _GEN_1812; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1814 = 10'h2f == _T_40[9:0] ? 4'hc : _GEN_1813; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1815 = 10'h30 == _T_40[9:0] ? 4'hc : _GEN_1814; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1816 = 10'h31 == _T_40[9:0] ? 4'hc : _GEN_1815; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1817 = 10'h32 == _T_40[9:0] ? 4'hc : _GEN_1816; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1818 = 10'h33 == _T_40[9:0] ? 4'hc : _GEN_1817; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1819 = 10'h34 == _T_40[9:0] ? 4'hc : _GEN_1818; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1820 = 10'h35 == _T_40[9:0] ? 4'hc : _GEN_1819; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1821 = 10'h36 == _T_40[9:0] ? 4'hc : _GEN_1820; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1822 = 10'h37 == _T_40[9:0] ? 4'hc : _GEN_1821; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1823 = 10'h38 == _T_40[9:0] ? 4'hc : _GEN_1822; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1824 = 10'h39 == _T_40[9:0] ? 4'hc : _GEN_1823; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1825 = 10'h3a == _T_40[9:0] ? 4'hc : _GEN_1824; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1826 = 10'h3b == _T_40[9:0] ? 4'hc : _GEN_1825; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1827 = 10'h3c == _T_40[9:0] ? 4'h7 : _GEN_1826; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1828 = 10'h3d == _T_40[9:0] ? 4'h9 : _GEN_1827; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1829 = 10'h3e == _T_40[9:0] ? 4'h8 : _GEN_1828; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1830 = 10'h3f == _T_40[9:0] ? 4'hc : _GEN_1829; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1831 = 10'h40 == _T_40[9:0] ? 4'hc : _GEN_1830; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1832 = 10'h41 == _T_40[9:0] ? 4'hc : _GEN_1831; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1833 = 10'h42 == _T_40[9:0] ? 4'hc : _GEN_1832; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1834 = 10'h43 == _T_40[9:0] ? 4'hc : _GEN_1833; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1835 = 10'h44 == _T_40[9:0] ? 4'hc : _GEN_1834; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1836 = 10'h45 == _T_40[9:0] ? 4'hc : _GEN_1835; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1837 = 10'h46 == _T_40[9:0] ? 4'hc : _GEN_1836; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1838 = 10'h47 == _T_40[9:0] ? 4'hc : _GEN_1837; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1839 = 10'h48 == _T_40[9:0] ? 4'hc : _GEN_1838; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1840 = 10'h49 == _T_40[9:0] ? 4'hc : _GEN_1839; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1841 = 10'h4a == _T_40[9:0] ? 4'hc : _GEN_1840; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1842 = 10'h4b == _T_40[9:0] ? 4'hc : _GEN_1841; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1843 = 10'h4c == _T_40[9:0] ? 4'hc : _GEN_1842; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1844 = 10'h4d == _T_40[9:0] ? 4'hc : _GEN_1843; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1845 = 10'h4e == _T_40[9:0] ? 4'hc : _GEN_1844; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1846 = 10'h4f == _T_40[9:0] ? 4'hc : _GEN_1845; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1847 = 10'h50 == _T_40[9:0] ? 4'hc : _GEN_1846; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1848 = 10'h51 == _T_40[9:0] ? 4'hc : _GEN_1847; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1849 = 10'h52 == _T_40[9:0] ? 4'hc : _GEN_1848; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1850 = 10'h53 == _T_40[9:0] ? 4'hc : _GEN_1849; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1851 = 10'h54 == _T_40[9:0] ? 4'hc : _GEN_1850; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1852 = 10'h55 == _T_40[9:0] ? 4'hc : _GEN_1851; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1853 = 10'h56 == _T_40[9:0] ? 4'hc : _GEN_1852; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1854 = 10'h57 == _T_40[9:0] ? 4'hc : _GEN_1853; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1855 = 10'h58 == _T_40[9:0] ? 4'hc : _GEN_1854; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1856 = 10'h59 == _T_40[9:0] ? 4'hc : _GEN_1855; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1857 = 10'h5a == _T_40[9:0] ? 4'h9 : _GEN_1856; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1858 = 10'h5b == _T_40[9:0] ? 4'ha : _GEN_1857; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1859 = 10'h5c == _T_40[9:0] ? 4'hc : _GEN_1858; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1860 = 10'h5d == _T_40[9:0] ? 4'hc : _GEN_1859; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1861 = 10'h5e == _T_40[9:0] ? 4'hc : _GEN_1860; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1862 = 10'h5f == _T_40[9:0] ? 4'hc : _GEN_1861; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1863 = 10'h60 == _T_40[9:0] ? 4'hc : _GEN_1862; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1864 = 10'h61 == _T_40[9:0] ? 4'hb : _GEN_1863; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1865 = 10'h62 == _T_40[9:0] ? 4'h8 : _GEN_1864; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1866 = 10'h63 == _T_40[9:0] ? 4'h9 : _GEN_1865; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1867 = 10'h64 == _T_40[9:0] ? 4'h7 : _GEN_1866; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1868 = 10'h65 == _T_40[9:0] ? 4'hb : _GEN_1867; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1869 = 10'h66 == _T_40[9:0] ? 4'hc : _GEN_1868; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1870 = 10'h67 == _T_40[9:0] ? 4'hc : _GEN_1869; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1871 = 10'h68 == _T_40[9:0] ? 4'hc : _GEN_1870; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1872 = 10'h69 == _T_40[9:0] ? 4'hc : _GEN_1871; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1873 = 10'h6a == _T_40[9:0] ? 4'hc : _GEN_1872; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1874 = 10'h6b == _T_40[9:0] ? 4'hb : _GEN_1873; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1875 = 10'h6c == _T_40[9:0] ? 4'h9 : _GEN_1874; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1876 = 10'h6d == _T_40[9:0] ? 4'ha : _GEN_1875; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1877 = 10'h6e == _T_40[9:0] ? 4'hc : _GEN_1876; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1878 = 10'h6f == _T_40[9:0] ? 4'hc : _GEN_1877; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1879 = 10'h70 == _T_40[9:0] ? 4'hc : _GEN_1878; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1880 = 10'h71 == _T_40[9:0] ? 4'hc : _GEN_1879; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1881 = 10'h72 == _T_40[9:0] ? 4'hc : _GEN_1880; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1882 = 10'h73 == _T_40[9:0] ? 4'hc : _GEN_1881; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1883 = 10'h74 == _T_40[9:0] ? 4'hc : _GEN_1882; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1884 = 10'h75 == _T_40[9:0] ? 4'hc : _GEN_1883; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1885 = 10'h76 == _T_40[9:0] ? 4'hc : _GEN_1884; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1886 = 10'h77 == _T_40[9:0] ? 4'hc : _GEN_1885; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1887 = 10'h78 == _T_40[9:0] ? 4'hc : _GEN_1886; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1888 = 10'h79 == _T_40[9:0] ? 4'hc : _GEN_1887; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1889 = 10'h7a == _T_40[9:0] ? 4'hc : _GEN_1888; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1890 = 10'h7b == _T_40[9:0] ? 4'hc : _GEN_1889; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1891 = 10'h7c == _T_40[9:0] ? 4'hc : _GEN_1890; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1892 = 10'h7d == _T_40[9:0] ? 4'hc : _GEN_1891; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1893 = 10'h7e == _T_40[9:0] ? 4'hc : _GEN_1892; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1894 = 10'h7f == _T_40[9:0] ? 4'hc : _GEN_1893; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1895 = 10'h80 == _T_40[9:0] ? 4'hc : _GEN_1894; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1896 = 10'h81 == _T_40[9:0] ? 4'h9 : _GEN_1895; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1897 = 10'h82 == _T_40[9:0] ? 4'h9 : _GEN_1896; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1898 = 10'h83 == _T_40[9:0] ? 4'h9 : _GEN_1897; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1899 = 10'h84 == _T_40[9:0] ? 4'hc : _GEN_1898; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1900 = 10'h85 == _T_40[9:0] ? 4'hc : _GEN_1899; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1901 = 10'h86 == _T_40[9:0] ? 4'hc : _GEN_1900; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1902 = 10'h87 == _T_40[9:0] ? 4'h8 : _GEN_1901; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1903 = 10'h88 == _T_40[9:0] ? 4'h9 : _GEN_1902; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1904 = 10'h89 == _T_40[9:0] ? 4'h9 : _GEN_1903; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1905 = 10'h8a == _T_40[9:0] ? 4'h9 : _GEN_1904; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1906 = 10'h8b == _T_40[9:0] ? 4'hc : _GEN_1905; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1907 = 10'h8c == _T_40[9:0] ? 4'hc : _GEN_1906; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1908 = 10'h8d == _T_40[9:0] ? 4'hc : _GEN_1907; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1909 = 10'h8e == _T_40[9:0] ? 4'hc : _GEN_1908; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1910 = 10'h8f == _T_40[9:0] ? 4'h9 : _GEN_1909; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1911 = 10'h90 == _T_40[9:0] ? 4'h9 : _GEN_1910; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1912 = 10'h91 == _T_40[9:0] ? 4'h9 : _GEN_1911; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1913 = 10'h92 == _T_40[9:0] ? 4'ha : _GEN_1912; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1914 = 10'h93 == _T_40[9:0] ? 4'hc : _GEN_1913; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1915 = 10'h94 == _T_40[9:0] ? 4'hc : _GEN_1914; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1916 = 10'h95 == _T_40[9:0] ? 4'hc : _GEN_1915; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1917 = 10'h96 == _T_40[9:0] ? 4'hc : _GEN_1916; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1918 = 10'h97 == _T_40[9:0] ? 4'hc : _GEN_1917; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1919 = 10'h98 == _T_40[9:0] ? 4'hc : _GEN_1918; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1920 = 10'h99 == _T_40[9:0] ? 4'hc : _GEN_1919; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1921 = 10'h9a == _T_40[9:0] ? 4'hc : _GEN_1920; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1922 = 10'h9b == _T_40[9:0] ? 4'hc : _GEN_1921; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1923 = 10'h9c == _T_40[9:0] ? 4'hc : _GEN_1922; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1924 = 10'h9d == _T_40[9:0] ? 4'hc : _GEN_1923; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1925 = 10'h9e == _T_40[9:0] ? 4'hc : _GEN_1924; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1926 = 10'h9f == _T_40[9:0] ? 4'hc : _GEN_1925; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1927 = 10'ha0 == _T_40[9:0] ? 4'hc : _GEN_1926; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1928 = 10'ha1 == _T_40[9:0] ? 4'hc : _GEN_1927; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1929 = 10'ha2 == _T_40[9:0] ? 4'hc : _GEN_1928; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1930 = 10'ha3 == _T_40[9:0] ? 4'hc : _GEN_1929; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1931 = 10'ha4 == _T_40[9:0] ? 4'hc : _GEN_1930; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1932 = 10'ha5 == _T_40[9:0] ? 4'hc : _GEN_1931; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1933 = 10'ha6 == _T_40[9:0] ? 4'hc : _GEN_1932; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1934 = 10'ha7 == _T_40[9:0] ? 4'hc : _GEN_1933; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1935 = 10'ha8 == _T_40[9:0] ? 4'h9 : _GEN_1934; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1936 = 10'ha9 == _T_40[9:0] ? 4'h8 : _GEN_1935; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1937 = 10'haa == _T_40[9:0] ? 4'h8 : _GEN_1936; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1938 = 10'hab == _T_40[9:0] ? 4'ha : _GEN_1937; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1939 = 10'hac == _T_40[9:0] ? 4'hb : _GEN_1938; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1940 = 10'had == _T_40[9:0] ? 4'h7 : _GEN_1939; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1941 = 10'hae == _T_40[9:0] ? 4'h9 : _GEN_1940; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1942 = 10'haf == _T_40[9:0] ? 4'h9 : _GEN_1941; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1943 = 10'hb0 == _T_40[9:0] ? 4'h8 : _GEN_1942; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1944 = 10'hb1 == _T_40[9:0] ? 4'h9 : _GEN_1943; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1945 = 10'hb2 == _T_40[9:0] ? 4'hc : _GEN_1944; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1946 = 10'hb3 == _T_40[9:0] ? 4'h9 : _GEN_1945; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1947 = 10'hb4 == _T_40[9:0] ? 4'h9 : _GEN_1946; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1948 = 10'hb5 == _T_40[9:0] ? 4'h9 : _GEN_1947; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1949 = 10'hb6 == _T_40[9:0] ? 4'h9 : _GEN_1948; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1950 = 10'hb7 == _T_40[9:0] ? 4'ha : _GEN_1949; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1951 = 10'hb8 == _T_40[9:0] ? 4'hc : _GEN_1950; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1952 = 10'hb9 == _T_40[9:0] ? 4'hc : _GEN_1951; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1953 = 10'hba == _T_40[9:0] ? 4'hc : _GEN_1952; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1954 = 10'hbb == _T_40[9:0] ? 4'hc : _GEN_1953; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1955 = 10'hbc == _T_40[9:0] ? 4'hc : _GEN_1954; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1956 = 10'hbd == _T_40[9:0] ? 4'hb : _GEN_1955; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1957 = 10'hbe == _T_40[9:0] ? 4'hc : _GEN_1956; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1958 = 10'hbf == _T_40[9:0] ? 4'hc : _GEN_1957; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1959 = 10'hc0 == _T_40[9:0] ? 4'hc : _GEN_1958; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1960 = 10'hc1 == _T_40[9:0] ? 4'hc : _GEN_1959; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1961 = 10'hc2 == _T_40[9:0] ? 4'hc : _GEN_1960; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1962 = 10'hc3 == _T_40[9:0] ? 4'hc : _GEN_1961; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1963 = 10'hc4 == _T_40[9:0] ? 4'hc : _GEN_1962; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1964 = 10'hc5 == _T_40[9:0] ? 4'hc : _GEN_1963; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1965 = 10'hc6 == _T_40[9:0] ? 4'hb : _GEN_1964; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1966 = 10'hc7 == _T_40[9:0] ? 4'hb : _GEN_1965; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1967 = 10'hc8 == _T_40[9:0] ? 4'ha : _GEN_1966; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1968 = 10'hc9 == _T_40[9:0] ? 4'ha : _GEN_1967; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1969 = 10'hca == _T_40[9:0] ? 4'hb : _GEN_1968; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1970 = 10'hcb == _T_40[9:0] ? 4'hc : _GEN_1969; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1971 = 10'hcc == _T_40[9:0] ? 4'hc : _GEN_1970; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1972 = 10'hcd == _T_40[9:0] ? 4'hc : _GEN_1971; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1973 = 10'hce == _T_40[9:0] ? 4'ha : _GEN_1972; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1974 = 10'hcf == _T_40[9:0] ? 4'h8 : _GEN_1973; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1975 = 10'hd0 == _T_40[9:0] ? 4'h9 : _GEN_1974; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1976 = 10'hd1 == _T_40[9:0] ? 4'h8 : _GEN_1975; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1977 = 10'hd2 == _T_40[9:0] ? 4'h9 : _GEN_1976; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1978 = 10'hd3 == _T_40[9:0] ? 4'h9 : _GEN_1977; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1979 = 10'hd4 == _T_40[9:0] ? 4'h9 : _GEN_1978; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1980 = 10'hd5 == _T_40[9:0] ? 4'h9 : _GEN_1979; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1981 = 10'hd6 == _T_40[9:0] ? 4'ha : _GEN_1980; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1982 = 10'hd7 == _T_40[9:0] ? 4'h9 : _GEN_1981; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1983 = 10'hd8 == _T_40[9:0] ? 4'h9 : _GEN_1982; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1984 = 10'hd9 == _T_40[9:0] ? 4'h9 : _GEN_1983; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1985 = 10'hda == _T_40[9:0] ? 4'ha : _GEN_1984; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1986 = 10'hdb == _T_40[9:0] ? 4'h9 : _GEN_1985; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1987 = 10'hdc == _T_40[9:0] ? 4'h7 : _GEN_1986; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1988 = 10'hdd == _T_40[9:0] ? 4'hc : _GEN_1987; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1989 = 10'hde == _T_40[9:0] ? 4'hc : _GEN_1988; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1990 = 10'hdf == _T_40[9:0] ? 4'hc : _GEN_1989; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1991 = 10'he0 == _T_40[9:0] ? 4'hc : _GEN_1990; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1992 = 10'he1 == _T_40[9:0] ? 4'hc : _GEN_1991; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1993 = 10'he2 == _T_40[9:0] ? 4'hc : _GEN_1992; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1994 = 10'he3 == _T_40[9:0] ? 4'h8 : _GEN_1993; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1995 = 10'he4 == _T_40[9:0] ? 4'hc : _GEN_1994; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1996 = 10'he5 == _T_40[9:0] ? 4'hc : _GEN_1995; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1997 = 10'he6 == _T_40[9:0] ? 4'hc : _GEN_1996; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1998 = 10'he7 == _T_40[9:0] ? 4'hc : _GEN_1997; // @[Filter.scala 230:142]
  wire [3:0] _GEN_1999 = 10'he8 == _T_40[9:0] ? 4'hc : _GEN_1998; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2000 = 10'he9 == _T_40[9:0] ? 4'hc : _GEN_1999; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2001 = 10'hea == _T_40[9:0] ? 4'hc : _GEN_2000; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2002 = 10'heb == _T_40[9:0] ? 4'ha : _GEN_2001; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2003 = 10'hec == _T_40[9:0] ? 4'h7 : _GEN_2002; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2004 = 10'hed == _T_40[9:0] ? 4'h3 : _GEN_2003; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2005 = 10'hee == _T_40[9:0] ? 4'h3 : _GEN_2004; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2006 = 10'hef == _T_40[9:0] ? 4'h3 : _GEN_2005; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2007 = 10'hf0 == _T_40[9:0] ? 4'h3 : _GEN_2006; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2008 = 10'hf1 == _T_40[9:0] ? 4'h8 : _GEN_2007; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2009 = 10'hf2 == _T_40[9:0] ? 4'hc : _GEN_2008; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2010 = 10'hf3 == _T_40[9:0] ? 4'hc : _GEN_2009; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2011 = 10'hf4 == _T_40[9:0] ? 4'hc : _GEN_2010; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2012 = 10'hf5 == _T_40[9:0] ? 4'h9 : _GEN_2011; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2013 = 10'hf6 == _T_40[9:0] ? 4'h9 : _GEN_2012; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2014 = 10'hf7 == _T_40[9:0] ? 4'h9 : _GEN_2013; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2015 = 10'hf8 == _T_40[9:0] ? 4'h9 : _GEN_2014; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2016 = 10'hf9 == _T_40[9:0] ? 4'ha : _GEN_2015; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2017 = 10'hfa == _T_40[9:0] ? 4'h9 : _GEN_2016; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2018 = 10'hfb == _T_40[9:0] ? 4'h9 : _GEN_2017; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2019 = 10'hfc == _T_40[9:0] ? 4'h9 : _GEN_2018; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2020 = 10'hfd == _T_40[9:0] ? 4'h9 : _GEN_2019; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2021 = 10'hfe == _T_40[9:0] ? 4'h9 : _GEN_2020; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2022 = 10'hff == _T_40[9:0] ? 4'ha : _GEN_2021; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2023 = 10'h100 == _T_40[9:0] ? 4'ha : _GEN_2022; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2024 = 10'h101 == _T_40[9:0] ? 4'h7 : _GEN_2023; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2025 = 10'h102 == _T_40[9:0] ? 4'h9 : _GEN_2024; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2026 = 10'h103 == _T_40[9:0] ? 4'hc : _GEN_2025; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2027 = 10'h104 == _T_40[9:0] ? 4'hc : _GEN_2026; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2028 = 10'h105 == _T_40[9:0] ? 4'hb : _GEN_2027; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2029 = 10'h106 == _T_40[9:0] ? 4'hb : _GEN_2028; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2030 = 10'h107 == _T_40[9:0] ? 4'hb : _GEN_2029; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2031 = 10'h108 == _T_40[9:0] ? 4'hb : _GEN_2030; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2032 = 10'h109 == _T_40[9:0] ? 4'h7 : _GEN_2031; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2033 = 10'h10a == _T_40[9:0] ? 4'hc : _GEN_2032; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2034 = 10'h10b == _T_40[9:0] ? 4'hc : _GEN_2033; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2035 = 10'h10c == _T_40[9:0] ? 4'hc : _GEN_2034; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2036 = 10'h10d == _T_40[9:0] ? 4'hc : _GEN_2035; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2037 = 10'h10e == _T_40[9:0] ? 4'hc : _GEN_2036; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2038 = 10'h10f == _T_40[9:0] ? 4'h9 : _GEN_2037; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2039 = 10'h110 == _T_40[9:0] ? 4'hb : _GEN_2038; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2040 = 10'h111 == _T_40[9:0] ? 4'h4 : _GEN_2039; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2041 = 10'h112 == _T_40[9:0] ? 4'h7 : _GEN_2040; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2042 = 10'h113 == _T_40[9:0] ? 4'h3 : _GEN_2041; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2043 = 10'h114 == _T_40[9:0] ? 4'h3 : _GEN_2042; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2044 = 10'h115 == _T_40[9:0] ? 4'h3 : _GEN_2043; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2045 = 10'h116 == _T_40[9:0] ? 4'h3 : _GEN_2044; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2046 = 10'h117 == _T_40[9:0] ? 4'h2 : _GEN_2045; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2047 = 10'h118 == _T_40[9:0] ? 4'h9 : _GEN_2046; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2048 = 10'h119 == _T_40[9:0] ? 4'hc : _GEN_2047; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2049 = 10'h11a == _T_40[9:0] ? 4'hc : _GEN_2048; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2050 = 10'h11b == _T_40[9:0] ? 4'hc : _GEN_2049; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2051 = 10'h11c == _T_40[9:0] ? 4'h9 : _GEN_2050; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2052 = 10'h11d == _T_40[9:0] ? 4'h9 : _GEN_2051; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2053 = 10'h11e == _T_40[9:0] ? 4'h9 : _GEN_2052; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2054 = 10'h11f == _T_40[9:0] ? 4'h8 : _GEN_2053; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2055 = 10'h120 == _T_40[9:0] ? 4'h7 : _GEN_2054; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2056 = 10'h121 == _T_40[9:0] ? 4'h9 : _GEN_2055; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2057 = 10'h122 == _T_40[9:0] ? 4'h7 : _GEN_2056; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2058 = 10'h123 == _T_40[9:0] ? 4'h7 : _GEN_2057; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2059 = 10'h124 == _T_40[9:0] ? 4'h9 : _GEN_2058; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2060 = 10'h125 == _T_40[9:0] ? 4'h9 : _GEN_2059; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2061 = 10'h126 == _T_40[9:0] ? 4'h8 : _GEN_2060; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2062 = 10'h127 == _T_40[9:0] ? 4'h9 : _GEN_2061; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2063 = 10'h128 == _T_40[9:0] ? 4'h8 : _GEN_2062; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2064 = 10'h129 == _T_40[9:0] ? 4'ha : _GEN_2063; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2065 = 10'h12a == _T_40[9:0] ? 4'h5 : _GEN_2064; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2066 = 10'h12b == _T_40[9:0] ? 4'h3 : _GEN_2065; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2067 = 10'h12c == _T_40[9:0] ? 4'h3 : _GEN_2066; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2068 = 10'h12d == _T_40[9:0] ? 4'h3 : _GEN_2067; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2069 = 10'h12e == _T_40[9:0] ? 4'h5 : _GEN_2068; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2070 = 10'h12f == _T_40[9:0] ? 4'h8 : _GEN_2069; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2071 = 10'h130 == _T_40[9:0] ? 4'hc : _GEN_2070; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2072 = 10'h131 == _T_40[9:0] ? 4'hb : _GEN_2071; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2073 = 10'h132 == _T_40[9:0] ? 4'h9 : _GEN_2072; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2074 = 10'h133 == _T_40[9:0] ? 4'h8 : _GEN_2073; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2075 = 10'h134 == _T_40[9:0] ? 4'h9 : _GEN_2074; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2076 = 10'h135 == _T_40[9:0] ? 4'h7 : _GEN_2075; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2077 = 10'h136 == _T_40[9:0] ? 4'h7 : _GEN_2076; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2078 = 10'h137 == _T_40[9:0] ? 4'h5 : _GEN_2077; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2079 = 10'h138 == _T_40[9:0] ? 4'h7 : _GEN_2078; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2080 = 10'h139 == _T_40[9:0] ? 4'h3 : _GEN_2079; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2081 = 10'h13a == _T_40[9:0] ? 4'h3 : _GEN_2080; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2082 = 10'h13b == _T_40[9:0] ? 4'h3 : _GEN_2081; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2083 = 10'h13c == _T_40[9:0] ? 4'h3 : _GEN_2082; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2084 = 10'h13d == _T_40[9:0] ? 4'h3 : _GEN_2083; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2085 = 10'h13e == _T_40[9:0] ? 4'h5 : _GEN_2084; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2086 = 10'h13f == _T_40[9:0] ? 4'ha : _GEN_2085; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2087 = 10'h140 == _T_40[9:0] ? 4'hc : _GEN_2086; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2088 = 10'h141 == _T_40[9:0] ? 4'hc : _GEN_2087; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2089 = 10'h142 == _T_40[9:0] ? 4'hc : _GEN_2088; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2090 = 10'h143 == _T_40[9:0] ? 4'h9 : _GEN_2089; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2091 = 10'h144 == _T_40[9:0] ? 4'h9 : _GEN_2090; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2092 = 10'h145 == _T_40[9:0] ? 4'h8 : _GEN_2091; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2093 = 10'h146 == _T_40[9:0] ? 4'h8 : _GEN_2092; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2094 = 10'h147 == _T_40[9:0] ? 4'h7 : _GEN_2093; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2095 = 10'h148 == _T_40[9:0] ? 4'h8 : _GEN_2094; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2096 = 10'h149 == _T_40[9:0] ? 4'h9 : _GEN_2095; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2097 = 10'h14a == _T_40[9:0] ? 4'ha : _GEN_2096; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2098 = 10'h14b == _T_40[9:0] ? 4'h9 : _GEN_2097; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2099 = 10'h14c == _T_40[9:0] ? 4'ha : _GEN_2098; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2100 = 10'h14d == _T_40[9:0] ? 4'h9 : _GEN_2099; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2101 = 10'h14e == _T_40[9:0] ? 4'h7 : _GEN_2100; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2102 = 10'h14f == _T_40[9:0] ? 4'h3 : _GEN_2101; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2103 = 10'h150 == _T_40[9:0] ? 4'h3 : _GEN_2102; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2104 = 10'h151 == _T_40[9:0] ? 4'h3 : _GEN_2103; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2105 = 10'h152 == _T_40[9:0] ? 4'h3 : _GEN_2104; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2106 = 10'h153 == _T_40[9:0] ? 4'h3 : _GEN_2105; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2107 = 10'h154 == _T_40[9:0] ? 4'h3 : _GEN_2106; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2108 = 10'h155 == _T_40[9:0] ? 4'h8 : _GEN_2107; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2109 = 10'h156 == _T_40[9:0] ? 4'ha : _GEN_2108; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2110 = 10'h157 == _T_40[9:0] ? 4'h7 : _GEN_2109; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2111 = 10'h158 == _T_40[9:0] ? 4'h7 : _GEN_2110; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2112 = 10'h159 == _T_40[9:0] ? 4'h7 : _GEN_2111; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2113 = 10'h15a == _T_40[9:0] ? 4'h7 : _GEN_2112; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2114 = 10'h15b == _T_40[9:0] ? 4'h7 : _GEN_2113; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2115 = 10'h15c == _T_40[9:0] ? 4'h7 : _GEN_2114; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2116 = 10'h15d == _T_40[9:0] ? 4'h7 : _GEN_2115; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2117 = 10'h15e == _T_40[9:0] ? 4'h7 : _GEN_2116; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2118 = 10'h15f == _T_40[9:0] ? 4'h3 : _GEN_2117; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2119 = 10'h160 == _T_40[9:0] ? 4'h3 : _GEN_2118; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2120 = 10'h161 == _T_40[9:0] ? 4'h3 : _GEN_2119; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2121 = 10'h162 == _T_40[9:0] ? 4'h3 : _GEN_2120; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2122 = 10'h163 == _T_40[9:0] ? 4'h3 : _GEN_2121; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2123 = 10'h164 == _T_40[9:0] ? 4'h4 : _GEN_2122; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2124 = 10'h165 == _T_40[9:0] ? 4'ha : _GEN_2123; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2125 = 10'h166 == _T_40[9:0] ? 4'ha : _GEN_2124; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2126 = 10'h167 == _T_40[9:0] ? 4'hc : _GEN_2125; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2127 = 10'h168 == _T_40[9:0] ? 4'hc : _GEN_2126; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2128 = 10'h169 == _T_40[9:0] ? 4'h9 : _GEN_2127; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2129 = 10'h16a == _T_40[9:0] ? 4'h9 : _GEN_2128; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2130 = 10'h16b == _T_40[9:0] ? 4'ha : _GEN_2129; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2131 = 10'h16c == _T_40[9:0] ? 4'h7 : _GEN_2130; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2132 = 10'h16d == _T_40[9:0] ? 4'h7 : _GEN_2131; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2133 = 10'h16e == _T_40[9:0] ? 4'h7 : _GEN_2132; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2134 = 10'h16f == _T_40[9:0] ? 4'ha : _GEN_2133; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2135 = 10'h170 == _T_40[9:0] ? 4'ha : _GEN_2134; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2136 = 10'h171 == _T_40[9:0] ? 4'ha : _GEN_2135; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2137 = 10'h172 == _T_40[9:0] ? 4'hc : _GEN_2136; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2138 = 10'h173 == _T_40[9:0] ? 4'h8 : _GEN_2137; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2139 = 10'h174 == _T_40[9:0] ? 4'h5 : _GEN_2138; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2140 = 10'h175 == _T_40[9:0] ? 4'h8 : _GEN_2139; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2141 = 10'h176 == _T_40[9:0] ? 4'h7 : _GEN_2140; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2142 = 10'h177 == _T_40[9:0] ? 4'h8 : _GEN_2141; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2143 = 10'h178 == _T_40[9:0] ? 4'h7 : _GEN_2142; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2144 = 10'h179 == _T_40[9:0] ? 4'h5 : _GEN_2143; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2145 = 10'h17a == _T_40[9:0] ? 4'h5 : _GEN_2144; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2146 = 10'h17b == _T_40[9:0] ? 4'h7 : _GEN_2145; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2147 = 10'h17c == _T_40[9:0] ? 4'h7 : _GEN_2146; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2148 = 10'h17d == _T_40[9:0] ? 4'h7 : _GEN_2147; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2149 = 10'h17e == _T_40[9:0] ? 4'h7 : _GEN_2148; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2150 = 10'h17f == _T_40[9:0] ? 4'h7 : _GEN_2149; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2151 = 10'h180 == _T_40[9:0] ? 4'h7 : _GEN_2150; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2152 = 10'h181 == _T_40[9:0] ? 4'h7 : _GEN_2151; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2153 = 10'h182 == _T_40[9:0] ? 4'h7 : _GEN_2152; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2154 = 10'h183 == _T_40[9:0] ? 4'h7 : _GEN_2153; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2155 = 10'h184 == _T_40[9:0] ? 4'h7 : _GEN_2154; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2156 = 10'h185 == _T_40[9:0] ? 4'h5 : _GEN_2155; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2157 = 10'h186 == _T_40[9:0] ? 4'h3 : _GEN_2156; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2158 = 10'h187 == _T_40[9:0] ? 4'h3 : _GEN_2157; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2159 = 10'h188 == _T_40[9:0] ? 4'h3 : _GEN_2158; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2160 = 10'h189 == _T_40[9:0] ? 4'h4 : _GEN_2159; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2161 = 10'h18a == _T_40[9:0] ? 4'h5 : _GEN_2160; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2162 = 10'h18b == _T_40[9:0] ? 4'ha : _GEN_2161; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2163 = 10'h18c == _T_40[9:0] ? 4'ha : _GEN_2162; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2164 = 10'h18d == _T_40[9:0] ? 4'ha : _GEN_2163; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2165 = 10'h18e == _T_40[9:0] ? 4'hc : _GEN_2164; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2166 = 10'h18f == _T_40[9:0] ? 4'h8 : _GEN_2165; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2167 = 10'h190 == _T_40[9:0] ? 4'h9 : _GEN_2166; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2168 = 10'h191 == _T_40[9:0] ? 4'h8 : _GEN_2167; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2169 = 10'h192 == _T_40[9:0] ? 4'h7 : _GEN_2168; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2170 = 10'h193 == _T_40[9:0] ? 4'h7 : _GEN_2169; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2171 = 10'h194 == _T_40[9:0] ? 4'h7 : _GEN_2170; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2172 = 10'h195 == _T_40[9:0] ? 4'h9 : _GEN_2171; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2173 = 10'h196 == _T_40[9:0] ? 4'ha : _GEN_2172; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2174 = 10'h197 == _T_40[9:0] ? 4'h8 : _GEN_2173; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2175 = 10'h198 == _T_40[9:0] ? 4'hc : _GEN_2174; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2176 = 10'h199 == _T_40[9:0] ? 4'h5 : _GEN_2175; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2177 = 10'h19a == _T_40[9:0] ? 4'h1 : _GEN_2176; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2178 = 10'h19b == _T_40[9:0] ? 4'h4 : _GEN_2177; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2179 = 10'h19c == _T_40[9:0] ? 4'h7 : _GEN_2178; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2180 = 10'h19d == _T_40[9:0] ? 4'h5 : _GEN_2179; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2181 = 10'h19e == _T_40[9:0] ? 4'h2 : _GEN_2180; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2182 = 10'h19f == _T_40[9:0] ? 4'h3 : _GEN_2181; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2183 = 10'h1a0 == _T_40[9:0] ? 4'h7 : _GEN_2182; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2184 = 10'h1a1 == _T_40[9:0] ? 4'h7 : _GEN_2183; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2185 = 10'h1a2 == _T_40[9:0] ? 4'h7 : _GEN_2184; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2186 = 10'h1a3 == _T_40[9:0] ? 4'h7 : _GEN_2185; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2187 = 10'h1a4 == _T_40[9:0] ? 4'h7 : _GEN_2186; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2188 = 10'h1a5 == _T_40[9:0] ? 4'h7 : _GEN_2187; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2189 = 10'h1a6 == _T_40[9:0] ? 4'h7 : _GEN_2188; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2190 = 10'h1a7 == _T_40[9:0] ? 4'h7 : _GEN_2189; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2191 = 10'h1a8 == _T_40[9:0] ? 4'h8 : _GEN_2190; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2192 = 10'h1a9 == _T_40[9:0] ? 4'h8 : _GEN_2191; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2193 = 10'h1aa == _T_40[9:0] ? 4'h6 : _GEN_2192; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2194 = 10'h1ab == _T_40[9:0] ? 4'h6 : _GEN_2193; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2195 = 10'h1ac == _T_40[9:0] ? 4'h5 : _GEN_2194; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2196 = 10'h1ad == _T_40[9:0] ? 4'h4 : _GEN_2195; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2197 = 10'h1ae == _T_40[9:0] ? 4'h3 : _GEN_2196; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2198 = 10'h1af == _T_40[9:0] ? 4'h6 : _GEN_2197; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2199 = 10'h1b0 == _T_40[9:0] ? 4'h6 : _GEN_2198; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2200 = 10'h1b1 == _T_40[9:0] ? 4'ha : _GEN_2199; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2201 = 10'h1b2 == _T_40[9:0] ? 4'ha : _GEN_2200; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2202 = 10'h1b3 == _T_40[9:0] ? 4'h9 : _GEN_2201; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2203 = 10'h1b4 == _T_40[9:0] ? 4'hb : _GEN_2202; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2204 = 10'h1b5 == _T_40[9:0] ? 4'h8 : _GEN_2203; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2205 = 10'h1b6 == _T_40[9:0] ? 4'h8 : _GEN_2204; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2206 = 10'h1b7 == _T_40[9:0] ? 4'h7 : _GEN_2205; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2207 = 10'h1b8 == _T_40[9:0] ? 4'h6 : _GEN_2206; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2208 = 10'h1b9 == _T_40[9:0] ? 4'h7 : _GEN_2207; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2209 = 10'h1ba == _T_40[9:0] ? 4'h6 : _GEN_2208; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2210 = 10'h1bb == _T_40[9:0] ? 4'h8 : _GEN_2209; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2211 = 10'h1bc == _T_40[9:0] ? 4'ha : _GEN_2210; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2212 = 10'h1bd == _T_40[9:0] ? 4'h9 : _GEN_2211; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2213 = 10'h1be == _T_40[9:0] ? 4'hc : _GEN_2212; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2214 = 10'h1bf == _T_40[9:0] ? 4'h7 : _GEN_2213; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2215 = 10'h1c0 == _T_40[9:0] ? 4'h6 : _GEN_2214; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2216 = 10'h1c1 == _T_40[9:0] ? 4'h7 : _GEN_2215; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2217 = 10'h1c2 == _T_40[9:0] ? 4'h7 : _GEN_2216; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2218 = 10'h1c3 == _T_40[9:0] ? 4'h6 : _GEN_2217; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2219 = 10'h1c4 == _T_40[9:0] ? 4'h5 : _GEN_2218; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2220 = 10'h1c5 == _T_40[9:0] ? 4'h6 : _GEN_2219; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2221 = 10'h1c6 == _T_40[9:0] ? 4'h8 : _GEN_2220; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2222 = 10'h1c7 == _T_40[9:0] ? 4'h7 : _GEN_2221; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2223 = 10'h1c8 == _T_40[9:0] ? 4'h7 : _GEN_2222; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2224 = 10'h1c9 == _T_40[9:0] ? 4'h7 : _GEN_2223; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2225 = 10'h1ca == _T_40[9:0] ? 4'h7 : _GEN_2224; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2226 = 10'h1cb == _T_40[9:0] ? 4'h7 : _GEN_2225; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2227 = 10'h1cc == _T_40[9:0] ? 4'h7 : _GEN_2226; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2228 = 10'h1cd == _T_40[9:0] ? 4'h8 : _GEN_2227; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2229 = 10'h1ce == _T_40[9:0] ? 4'h8 : _GEN_2228; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2230 = 10'h1cf == _T_40[9:0] ? 4'h8 : _GEN_2229; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2231 = 10'h1d0 == _T_40[9:0] ? 4'h5 : _GEN_2230; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2232 = 10'h1d1 == _T_40[9:0] ? 4'h6 : _GEN_2231; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2233 = 10'h1d2 == _T_40[9:0] ? 4'h7 : _GEN_2232; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2234 = 10'h1d3 == _T_40[9:0] ? 4'h7 : _GEN_2233; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2235 = 10'h1d4 == _T_40[9:0] ? 4'h7 : _GEN_2234; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2236 = 10'h1d5 == _T_40[9:0] ? 4'h6 : _GEN_2235; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2237 = 10'h1d6 == _T_40[9:0] ? 4'h8 : _GEN_2236; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2238 = 10'h1d7 == _T_40[9:0] ? 4'ha : _GEN_2237; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2239 = 10'h1d8 == _T_40[9:0] ? 4'ha : _GEN_2238; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2240 = 10'h1d9 == _T_40[9:0] ? 4'ha : _GEN_2239; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2241 = 10'h1da == _T_40[9:0] ? 4'h8 : _GEN_2240; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2242 = 10'h1db == _T_40[9:0] ? 4'h9 : _GEN_2241; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2243 = 10'h1dc == _T_40[9:0] ? 4'h9 : _GEN_2242; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2244 = 10'h1dd == _T_40[9:0] ? 4'h5 : _GEN_2243; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2245 = 10'h1de == _T_40[9:0] ? 4'h7 : _GEN_2244; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2246 = 10'h1df == _T_40[9:0] ? 4'h7 : _GEN_2245; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2247 = 10'h1e0 == _T_40[9:0] ? 4'h7 : _GEN_2246; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2248 = 10'h1e1 == _T_40[9:0] ? 4'h6 : _GEN_2247; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2249 = 10'h1e2 == _T_40[9:0] ? 4'h9 : _GEN_2248; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2250 = 10'h1e3 == _T_40[9:0] ? 4'h9 : _GEN_2249; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2251 = 10'h1e4 == _T_40[9:0] ? 4'hb : _GEN_2250; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2252 = 10'h1e5 == _T_40[9:0] ? 4'h8 : _GEN_2251; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2253 = 10'h1e6 == _T_40[9:0] ? 4'h7 : _GEN_2252; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2254 = 10'h1e7 == _T_40[9:0] ? 4'h8 : _GEN_2253; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2255 = 10'h1e8 == _T_40[9:0] ? 4'h8 : _GEN_2254; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2256 = 10'h1e9 == _T_40[9:0] ? 4'h8 : _GEN_2255; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2257 = 10'h1ea == _T_40[9:0] ? 4'h8 : _GEN_2256; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2258 = 10'h1eb == _T_40[9:0] ? 4'h8 : _GEN_2257; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2259 = 10'h1ec == _T_40[9:0] ? 4'h8 : _GEN_2258; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2260 = 10'h1ed == _T_40[9:0] ? 4'h6 : _GEN_2259; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2261 = 10'h1ee == _T_40[9:0] ? 4'h7 : _GEN_2260; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2262 = 10'h1ef == _T_40[9:0] ? 4'h7 : _GEN_2261; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2263 = 10'h1f0 == _T_40[9:0] ? 4'h7 : _GEN_2262; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2264 = 10'h1f1 == _T_40[9:0] ? 4'h7 : _GEN_2263; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2265 = 10'h1f2 == _T_40[9:0] ? 4'h7 : _GEN_2264; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2266 = 10'h1f3 == _T_40[9:0] ? 4'h8 : _GEN_2265; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2267 = 10'h1f4 == _T_40[9:0] ? 4'h8 : _GEN_2266; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2268 = 10'h1f5 == _T_40[9:0] ? 4'h8 : _GEN_2267; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2269 = 10'h1f6 == _T_40[9:0] ? 4'ha : _GEN_2268; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2270 = 10'h1f7 == _T_40[9:0] ? 4'h6 : _GEN_2269; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2271 = 10'h1f8 == _T_40[9:0] ? 4'h6 : _GEN_2270; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2272 = 10'h1f9 == _T_40[9:0] ? 4'h8 : _GEN_2271; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2273 = 10'h1fa == _T_40[9:0] ? 4'h8 : _GEN_2272; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2274 = 10'h1fb == _T_40[9:0] ? 4'h6 : _GEN_2273; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2275 = 10'h1fc == _T_40[9:0] ? 4'ha : _GEN_2274; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2276 = 10'h1fd == _T_40[9:0] ? 4'hb : _GEN_2275; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2277 = 10'h1fe == _T_40[9:0] ? 4'ha : _GEN_2276; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2278 = 10'h1ff == _T_40[9:0] ? 4'ha : _GEN_2277; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2279 = 10'h200 == _T_40[9:0] ? 4'h4 : _GEN_2278; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2280 = 10'h201 == _T_40[9:0] ? 4'h7 : _GEN_2279; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2281 = 10'h202 == _T_40[9:0] ? 4'h6 : _GEN_2280; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2282 = 10'h203 == _T_40[9:0] ? 4'h6 : _GEN_2281; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2283 = 10'h204 == _T_40[9:0] ? 4'h5 : _GEN_2282; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2284 = 10'h205 == _T_40[9:0] ? 4'h6 : _GEN_2283; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2285 = 10'h206 == _T_40[9:0] ? 4'h6 : _GEN_2284; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2286 = 10'h207 == _T_40[9:0] ? 4'h5 : _GEN_2285; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2287 = 10'h208 == _T_40[9:0] ? 4'h7 : _GEN_2286; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2288 = 10'h209 == _T_40[9:0] ? 4'h9 : _GEN_2287; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2289 = 10'h20a == _T_40[9:0] ? 4'hb : _GEN_2288; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2290 = 10'h20b == _T_40[9:0] ? 4'h7 : _GEN_2289; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2291 = 10'h20c == _T_40[9:0] ? 4'h7 : _GEN_2290; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2292 = 10'h20d == _T_40[9:0] ? 4'h7 : _GEN_2291; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2293 = 10'h20e == _T_40[9:0] ? 4'h7 : _GEN_2292; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2294 = 10'h20f == _T_40[9:0] ? 4'h7 : _GEN_2293; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2295 = 10'h210 == _T_40[9:0] ? 4'h7 : _GEN_2294; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2296 = 10'h211 == _T_40[9:0] ? 4'h8 : _GEN_2295; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2297 = 10'h212 == _T_40[9:0] ? 4'h8 : _GEN_2296; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2298 = 10'h213 == _T_40[9:0] ? 4'h9 : _GEN_2297; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2299 = 10'h214 == _T_40[9:0] ? 4'h6 : _GEN_2298; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2300 = 10'h215 == _T_40[9:0] ? 4'h7 : _GEN_2299; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2301 = 10'h216 == _T_40[9:0] ? 4'h7 : _GEN_2300; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2302 = 10'h217 == _T_40[9:0] ? 4'h7 : _GEN_2301; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2303 = 10'h218 == _T_40[9:0] ? 4'h7 : _GEN_2302; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2304 = 10'h219 == _T_40[9:0] ? 4'h8 : _GEN_2303; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2305 = 10'h21a == _T_40[9:0] ? 4'h7 : _GEN_2304; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2306 = 10'h21b == _T_40[9:0] ? 4'h8 : _GEN_2305; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2307 = 10'h21c == _T_40[9:0] ? 4'ha : _GEN_2306; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2308 = 10'h21d == _T_40[9:0] ? 4'ha : _GEN_2307; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2309 = 10'h21e == _T_40[9:0] ? 4'h7 : _GEN_2308; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2310 = 10'h21f == _T_40[9:0] ? 4'h6 : _GEN_2309; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2311 = 10'h220 == _T_40[9:0] ? 4'h6 : _GEN_2310; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2312 = 10'h221 == _T_40[9:0] ? 4'h7 : _GEN_2311; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2313 = 10'h222 == _T_40[9:0] ? 4'ha : _GEN_2312; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2314 = 10'h223 == _T_40[9:0] ? 4'ha : _GEN_2313; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2315 = 10'h224 == _T_40[9:0] ? 4'ha : _GEN_2314; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2316 = 10'h225 == _T_40[9:0] ? 4'h8 : _GEN_2315; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2317 = 10'h226 == _T_40[9:0] ? 4'h3 : _GEN_2316; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2318 = 10'h227 == _T_40[9:0] ? 4'h4 : _GEN_2317; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2319 = 10'h228 == _T_40[9:0] ? 4'h6 : _GEN_2318; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2320 = 10'h229 == _T_40[9:0] ? 4'h6 : _GEN_2319; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2321 = 10'h22a == _T_40[9:0] ? 4'h6 : _GEN_2320; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2322 = 10'h22b == _T_40[9:0] ? 4'h6 : _GEN_2321; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2323 = 10'h22c == _T_40[9:0] ? 4'h5 : _GEN_2322; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2324 = 10'h22d == _T_40[9:0] ? 4'h6 : _GEN_2323; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2325 = 10'h22e == _T_40[9:0] ? 4'h6 : _GEN_2324; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2326 = 10'h22f == _T_40[9:0] ? 4'h8 : _GEN_2325; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2327 = 10'h230 == _T_40[9:0] ? 4'h7 : _GEN_2326; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2328 = 10'h231 == _T_40[9:0] ? 4'h5 : _GEN_2327; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2329 = 10'h232 == _T_40[9:0] ? 4'h6 : _GEN_2328; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2330 = 10'h233 == _T_40[9:0] ? 4'h8 : _GEN_2329; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2331 = 10'h234 == _T_40[9:0] ? 4'h8 : _GEN_2330; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2332 = 10'h235 == _T_40[9:0] ? 4'h8 : _GEN_2331; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2333 = 10'h236 == _T_40[9:0] ? 4'h8 : _GEN_2332; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2334 = 10'h237 == _T_40[9:0] ? 4'h8 : _GEN_2333; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2335 = 10'h238 == _T_40[9:0] ? 4'h8 : _GEN_2334; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2336 = 10'h239 == _T_40[9:0] ? 4'h6 : _GEN_2335; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2337 = 10'h23a == _T_40[9:0] ? 4'h6 : _GEN_2336; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2338 = 10'h23b == _T_40[9:0] ? 4'h7 : _GEN_2337; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2339 = 10'h23c == _T_40[9:0] ? 4'h6 : _GEN_2338; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2340 = 10'h23d == _T_40[9:0] ? 4'h7 : _GEN_2339; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2341 = 10'h23e == _T_40[9:0] ? 4'h7 : _GEN_2340; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2342 = 10'h23f == _T_40[9:0] ? 4'h6 : _GEN_2341; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2343 = 10'h240 == _T_40[9:0] ? 4'h6 : _GEN_2342; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2344 = 10'h241 == _T_40[9:0] ? 4'h8 : _GEN_2343; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2345 = 10'h242 == _T_40[9:0] ? 4'ha : _GEN_2344; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2346 = 10'h243 == _T_40[9:0] ? 4'ha : _GEN_2345; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2347 = 10'h244 == _T_40[9:0] ? 4'ha : _GEN_2346; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2348 = 10'h245 == _T_40[9:0] ? 4'h8 : _GEN_2347; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2349 = 10'h246 == _T_40[9:0] ? 4'h8 : _GEN_2348; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2350 = 10'h247 == _T_40[9:0] ? 4'h9 : _GEN_2349; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2351 = 10'h248 == _T_40[9:0] ? 4'ha : _GEN_2350; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2352 = 10'h249 == _T_40[9:0] ? 4'ha : _GEN_2351; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2353 = 10'h24a == _T_40[9:0] ? 4'ha : _GEN_2352; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2354 = 10'h24b == _T_40[9:0] ? 4'h4 : _GEN_2353; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2355 = 10'h24c == _T_40[9:0] ? 4'h3 : _GEN_2354; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2356 = 10'h24d == _T_40[9:0] ? 4'h4 : _GEN_2355; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2357 = 10'h24e == _T_40[9:0] ? 4'h5 : _GEN_2356; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2358 = 10'h24f == _T_40[9:0] ? 4'h5 : _GEN_2357; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2359 = 10'h250 == _T_40[9:0] ? 4'h5 : _GEN_2358; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2360 = 10'h251 == _T_40[9:0] ? 4'h5 : _GEN_2359; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2361 = 10'h252 == _T_40[9:0] ? 4'h5 : _GEN_2360; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2362 = 10'h253 == _T_40[9:0] ? 4'h5 : _GEN_2361; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2363 = 10'h254 == _T_40[9:0] ? 4'h5 : _GEN_2362; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2364 = 10'h255 == _T_40[9:0] ? 4'h6 : _GEN_2363; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2365 = 10'h256 == _T_40[9:0] ? 4'h7 : _GEN_2364; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2366 = 10'h257 == _T_40[9:0] ? 4'h3 : _GEN_2365; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2367 = 10'h258 == _T_40[9:0] ? 4'h6 : _GEN_2366; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2368 = 10'h259 == _T_40[9:0] ? 4'h7 : _GEN_2367; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2369 = 10'h25a == _T_40[9:0] ? 4'h7 : _GEN_2368; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2370 = 10'h25b == _T_40[9:0] ? 4'h7 : _GEN_2369; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2371 = 10'h25c == _T_40[9:0] ? 4'h8 : _GEN_2370; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2372 = 10'h25d == _T_40[9:0] ? 4'h8 : _GEN_2371; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2373 = 10'h25e == _T_40[9:0] ? 4'h4 : _GEN_2372; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2374 = 10'h25f == _T_40[9:0] ? 4'h3 : _GEN_2373; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2375 = 10'h260 == _T_40[9:0] ? 4'h7 : _GEN_2374; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2376 = 10'h261 == _T_40[9:0] ? 4'h7 : _GEN_2375; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2377 = 10'h262 == _T_40[9:0] ? 4'h7 : _GEN_2376; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2378 = 10'h263 == _T_40[9:0] ? 4'h6 : _GEN_2377; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2379 = 10'h264 == _T_40[9:0] ? 4'h7 : _GEN_2378; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2380 = 10'h265 == _T_40[9:0] ? 4'h6 : _GEN_2379; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2381 = 10'h266 == _T_40[9:0] ? 4'h5 : _GEN_2380; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2382 = 10'h267 == _T_40[9:0] ? 4'h7 : _GEN_2381; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2383 = 10'h268 == _T_40[9:0] ? 4'ha : _GEN_2382; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2384 = 10'h269 == _T_40[9:0] ? 4'ha : _GEN_2383; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2385 = 10'h26a == _T_40[9:0] ? 4'ha : _GEN_2384; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2386 = 10'h26b == _T_40[9:0] ? 4'ha : _GEN_2385; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2387 = 10'h26c == _T_40[9:0] ? 4'ha : _GEN_2386; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2388 = 10'h26d == _T_40[9:0] ? 4'ha : _GEN_2387; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2389 = 10'h26e == _T_40[9:0] ? 4'ha : _GEN_2388; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2390 = 10'h26f == _T_40[9:0] ? 4'ha : _GEN_2389; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2391 = 10'h270 == _T_40[9:0] ? 4'h5 : _GEN_2390; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2392 = 10'h271 == _T_40[9:0] ? 4'h3 : _GEN_2391; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2393 = 10'h272 == _T_40[9:0] ? 4'h3 : _GEN_2392; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2394 = 10'h273 == _T_40[9:0] ? 4'h4 : _GEN_2393; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2395 = 10'h274 == _T_40[9:0] ? 4'h6 : _GEN_2394; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2396 = 10'h275 == _T_40[9:0] ? 4'h5 : _GEN_2395; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2397 = 10'h276 == _T_40[9:0] ? 4'h6 : _GEN_2396; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2398 = 10'h277 == _T_40[9:0] ? 4'h5 : _GEN_2397; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2399 = 10'h278 == _T_40[9:0] ? 4'h6 : _GEN_2398; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2400 = 10'h279 == _T_40[9:0] ? 4'h6 : _GEN_2399; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2401 = 10'h27a == _T_40[9:0] ? 4'h6 : _GEN_2400; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2402 = 10'h27b == _T_40[9:0] ? 4'h8 : _GEN_2401; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2403 = 10'h27c == _T_40[9:0] ? 4'h6 : _GEN_2402; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2404 = 10'h27d == _T_40[9:0] ? 4'h2 : _GEN_2403; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2405 = 10'h27e == _T_40[9:0] ? 4'h5 : _GEN_2404; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2406 = 10'h27f == _T_40[9:0] ? 4'h7 : _GEN_2405; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2407 = 10'h280 == _T_40[9:0] ? 4'h7 : _GEN_2406; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2408 = 10'h281 == _T_40[9:0] ? 4'h8 : _GEN_2407; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2409 = 10'h282 == _T_40[9:0] ? 4'h7 : _GEN_2408; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2410 = 10'h283 == _T_40[9:0] ? 4'h3 : _GEN_2409; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2411 = 10'h284 == _T_40[9:0] ? 4'h3 : _GEN_2410; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2412 = 10'h285 == _T_40[9:0] ? 4'h3 : _GEN_2411; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2413 = 10'h286 == _T_40[9:0] ? 4'h7 : _GEN_2412; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2414 = 10'h287 == _T_40[9:0] ? 4'h7 : _GEN_2413; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2415 = 10'h288 == _T_40[9:0] ? 4'h7 : _GEN_2414; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2416 = 10'h289 == _T_40[9:0] ? 4'h7 : _GEN_2415; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2417 = 10'h28a == _T_40[9:0] ? 4'h8 : _GEN_2416; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2418 = 10'h28b == _T_40[9:0] ? 4'h8 : _GEN_2417; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2419 = 10'h28c == _T_40[9:0] ? 4'h7 : _GEN_2418; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2420 = 10'h28d == _T_40[9:0] ? 4'h6 : _GEN_2419; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2421 = 10'h28e == _T_40[9:0] ? 4'h3 : _GEN_2420; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2422 = 10'h28f == _T_40[9:0] ? 4'h6 : _GEN_2421; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2423 = 10'h290 == _T_40[9:0] ? 4'h8 : _GEN_2422; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2424 = 10'h291 == _T_40[9:0] ? 4'ha : _GEN_2423; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2425 = 10'h292 == _T_40[9:0] ? 4'ha : _GEN_2424; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2426 = 10'h293 == _T_40[9:0] ? 4'ha : _GEN_2425; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2427 = 10'h294 == _T_40[9:0] ? 4'h9 : _GEN_2426; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2428 = 10'h295 == _T_40[9:0] ? 4'h4 : _GEN_2427; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2429 = 10'h296 == _T_40[9:0] ? 4'h3 : _GEN_2428; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2430 = 10'h297 == _T_40[9:0] ? 4'h3 : _GEN_2429; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2431 = 10'h298 == _T_40[9:0] ? 4'h3 : _GEN_2430; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2432 = 10'h299 == _T_40[9:0] ? 4'h4 : _GEN_2431; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2433 = 10'h29a == _T_40[9:0] ? 4'h5 : _GEN_2432; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2434 = 10'h29b == _T_40[9:0] ? 4'h5 : _GEN_2433; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2435 = 10'h29c == _T_40[9:0] ? 4'h5 : _GEN_2434; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2436 = 10'h29d == _T_40[9:0] ? 4'h5 : _GEN_2435; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2437 = 10'h29e == _T_40[9:0] ? 4'h5 : _GEN_2436; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2438 = 10'h29f == _T_40[9:0] ? 4'h5 : _GEN_2437; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2439 = 10'h2a0 == _T_40[9:0] ? 4'h6 : _GEN_2438; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2440 = 10'h2a1 == _T_40[9:0] ? 4'h7 : _GEN_2439; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2441 = 10'h2a2 == _T_40[9:0] ? 4'h5 : _GEN_2440; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2442 = 10'h2a3 == _T_40[9:0] ? 4'h2 : _GEN_2441; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2443 = 10'h2a4 == _T_40[9:0] ? 4'h3 : _GEN_2442; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2444 = 10'h2a5 == _T_40[9:0] ? 4'h7 : _GEN_2443; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2445 = 10'h2a6 == _T_40[9:0] ? 4'h8 : _GEN_2444; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2446 = 10'h2a7 == _T_40[9:0] ? 4'h7 : _GEN_2445; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2447 = 10'h2a8 == _T_40[9:0] ? 4'h3 : _GEN_2446; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2448 = 10'h2a9 == _T_40[9:0] ? 4'h2 : _GEN_2447; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2449 = 10'h2aa == _T_40[9:0] ? 4'h3 : _GEN_2448; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2450 = 10'h2ab == _T_40[9:0] ? 4'h3 : _GEN_2449; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2451 = 10'h2ac == _T_40[9:0] ? 4'h7 : _GEN_2450; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2452 = 10'h2ad == _T_40[9:0] ? 4'h8 : _GEN_2451; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2453 = 10'h2ae == _T_40[9:0] ? 4'h7 : _GEN_2452; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2454 = 10'h2af == _T_40[9:0] ? 4'h8 : _GEN_2453; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2455 = 10'h2b0 == _T_40[9:0] ? 4'h8 : _GEN_2454; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2456 = 10'h2b1 == _T_40[9:0] ? 4'h8 : _GEN_2455; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2457 = 10'h2b2 == _T_40[9:0] ? 4'h7 : _GEN_2456; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2458 = 10'h2b3 == _T_40[9:0] ? 4'h6 : _GEN_2457; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2459 = 10'h2b4 == _T_40[9:0] ? 4'h2 : _GEN_2458; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2460 = 10'h2b5 == _T_40[9:0] ? 4'h2 : _GEN_2459; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2461 = 10'h2b6 == _T_40[9:0] ? 4'h3 : _GEN_2460; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2462 = 10'h2b7 == _T_40[9:0] ? 4'h3 : _GEN_2461; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2463 = 10'h2b8 == _T_40[9:0] ? 4'h6 : _GEN_2462; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2464 = 10'h2b9 == _T_40[9:0] ? 4'h9 : _GEN_2463; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2465 = 10'h2ba == _T_40[9:0] ? 4'h3 : _GEN_2464; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2466 = 10'h2bb == _T_40[9:0] ? 4'h3 : _GEN_2465; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2467 = 10'h2bc == _T_40[9:0] ? 4'h3 : _GEN_2466; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2468 = 10'h2bd == _T_40[9:0] ? 4'h2 : _GEN_2467; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2469 = 10'h2be == _T_40[9:0] ? 4'h3 : _GEN_2468; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2470 = 10'h2bf == _T_40[9:0] ? 4'h3 : _GEN_2469; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2471 = 10'h2c0 == _T_40[9:0] ? 4'h5 : _GEN_2470; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2472 = 10'h2c1 == _T_40[9:0] ? 4'h5 : _GEN_2471; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2473 = 10'h2c2 == _T_40[9:0] ? 4'h5 : _GEN_2472; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2474 = 10'h2c3 == _T_40[9:0] ? 4'h5 : _GEN_2473; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2475 = 10'h2c4 == _T_40[9:0] ? 4'h5 : _GEN_2474; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2476 = 10'h2c5 == _T_40[9:0] ? 4'h5 : _GEN_2475; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2477 = 10'h2c6 == _T_40[9:0] ? 4'h6 : _GEN_2476; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2478 = 10'h2c7 == _T_40[9:0] ? 4'h7 : _GEN_2477; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2479 = 10'h2c8 == _T_40[9:0] ? 4'h5 : _GEN_2478; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2480 = 10'h2c9 == _T_40[9:0] ? 4'h2 : _GEN_2479; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2481 = 10'h2ca == _T_40[9:0] ? 4'h2 : _GEN_2480; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2482 = 10'h2cb == _T_40[9:0] ? 4'h3 : _GEN_2481; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2483 = 10'h2cc == _T_40[9:0] ? 4'h3 : _GEN_2482; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2484 = 10'h2cd == _T_40[9:0] ? 4'h2 : _GEN_2483; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2485 = 10'h2ce == _T_40[9:0] ? 4'h2 : _GEN_2484; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2486 = 10'h2cf == _T_40[9:0] ? 4'h2 : _GEN_2485; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2487 = 10'h2d0 == _T_40[9:0] ? 4'h2 : _GEN_2486; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2488 = 10'h2d1 == _T_40[9:0] ? 4'h2 : _GEN_2487; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2489 = 10'h2d2 == _T_40[9:0] ? 4'h7 : _GEN_2488; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2490 = 10'h2d3 == _T_40[9:0] ? 4'h7 : _GEN_2489; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2491 = 10'h2d4 == _T_40[9:0] ? 4'h8 : _GEN_2490; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2492 = 10'h2d5 == _T_40[9:0] ? 4'h8 : _GEN_2491; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2493 = 10'h2d6 == _T_40[9:0] ? 4'h8 : _GEN_2492; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2494 = 10'h2d7 == _T_40[9:0] ? 4'h8 : _GEN_2493; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2495 = 10'h2d8 == _T_40[9:0] ? 4'h7 : _GEN_2494; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2496 = 10'h2d9 == _T_40[9:0] ? 4'h6 : _GEN_2495; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2497 = 10'h2da == _T_40[9:0] ? 4'h4 : _GEN_2496; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2498 = 10'h2db == _T_40[9:0] ? 4'h2 : _GEN_2497; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2499 = 10'h2dc == _T_40[9:0] ? 4'h2 : _GEN_2498; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2500 = 10'h2dd == _T_40[9:0] ? 4'h3 : _GEN_2499; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2501 = 10'h2de == _T_40[9:0] ? 4'h3 : _GEN_2500; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2502 = 10'h2df == _T_40[9:0] ? 4'h3 : _GEN_2501; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2503 = 10'h2e0 == _T_40[9:0] ? 4'h3 : _GEN_2502; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2504 = 10'h2e1 == _T_40[9:0] ? 4'h3 : _GEN_2503; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2505 = 10'h2e2 == _T_40[9:0] ? 4'h3 : _GEN_2504; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2506 = 10'h2e3 == _T_40[9:0] ? 4'h2 : _GEN_2505; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2507 = 10'h2e4 == _T_40[9:0] ? 4'h3 : _GEN_2506; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2508 = 10'h2e5 == _T_40[9:0] ? 4'h2 : _GEN_2507; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2509 = 10'h2e6 == _T_40[9:0] ? 4'h5 : _GEN_2508; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2510 = 10'h2e7 == _T_40[9:0] ? 4'h5 : _GEN_2509; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2511 = 10'h2e8 == _T_40[9:0] ? 4'h5 : _GEN_2510; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2512 = 10'h2e9 == _T_40[9:0] ? 4'h5 : _GEN_2511; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2513 = 10'h2ea == _T_40[9:0] ? 4'h5 : _GEN_2512; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2514 = 10'h2eb == _T_40[9:0] ? 4'h5 : _GEN_2513; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2515 = 10'h2ec == _T_40[9:0] ? 4'h6 : _GEN_2514; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2516 = 10'h2ed == _T_40[9:0] ? 4'h7 : _GEN_2515; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2517 = 10'h2ee == _T_40[9:0] ? 4'h6 : _GEN_2516; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2518 = 10'h2ef == _T_40[9:0] ? 4'h2 : _GEN_2517; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2519 = 10'h2f0 == _T_40[9:0] ? 4'h2 : _GEN_2518; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2520 = 10'h2f1 == _T_40[9:0] ? 4'h2 : _GEN_2519; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2521 = 10'h2f2 == _T_40[9:0] ? 4'h2 : _GEN_2520; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2522 = 10'h2f3 == _T_40[9:0] ? 4'h2 : _GEN_2521; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2523 = 10'h2f4 == _T_40[9:0] ? 4'h2 : _GEN_2522; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2524 = 10'h2f5 == _T_40[9:0] ? 4'h2 : _GEN_2523; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2525 = 10'h2f6 == _T_40[9:0] ? 4'h2 : _GEN_2524; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2526 = 10'h2f7 == _T_40[9:0] ? 4'h2 : _GEN_2525; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2527 = 10'h2f8 == _T_40[9:0] ? 4'h7 : _GEN_2526; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2528 = 10'h2f9 == _T_40[9:0] ? 4'h7 : _GEN_2527; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2529 = 10'h2fa == _T_40[9:0] ? 4'h8 : _GEN_2528; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2530 = 10'h2fb == _T_40[9:0] ? 4'h8 : _GEN_2529; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2531 = 10'h2fc == _T_40[9:0] ? 4'h7 : _GEN_2530; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2532 = 10'h2fd == _T_40[9:0] ? 4'h7 : _GEN_2531; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2533 = 10'h2fe == _T_40[9:0] ? 4'h7 : _GEN_2532; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2534 = 10'h2ff == _T_40[9:0] ? 4'h7 : _GEN_2533; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2535 = 10'h300 == _T_40[9:0] ? 4'h8 : _GEN_2534; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2536 = 10'h301 == _T_40[9:0] ? 4'h7 : _GEN_2535; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2537 = 10'h302 == _T_40[9:0] ? 4'h3 : _GEN_2536; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2538 = 10'h303 == _T_40[9:0] ? 4'h3 : _GEN_2537; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2539 = 10'h304 == _T_40[9:0] ? 4'h2 : _GEN_2538; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2540 = 10'h305 == _T_40[9:0] ? 4'h2 : _GEN_2539; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2541 = 10'h306 == _T_40[9:0] ? 4'h2 : _GEN_2540; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2542 = 10'h307 == _T_40[9:0] ? 4'h2 : _GEN_2541; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2543 = 10'h308 == _T_40[9:0] ? 4'h2 : _GEN_2542; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2544 = 10'h309 == _T_40[9:0] ? 4'h2 : _GEN_2543; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2545 = 10'h30a == _T_40[9:0] ? 4'h2 : _GEN_2544; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2546 = 10'h30b == _T_40[9:0] ? 4'h3 : _GEN_2545; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2547 = 10'h30c == _T_40[9:0] ? 4'h4 : _GEN_2546; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2548 = 10'h30d == _T_40[9:0] ? 4'h5 : _GEN_2547; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2549 = 10'h30e == _T_40[9:0] ? 4'h5 : _GEN_2548; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2550 = 10'h30f == _T_40[9:0] ? 4'h5 : _GEN_2549; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2551 = 10'h310 == _T_40[9:0] ? 4'h5 : _GEN_2550; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2552 = 10'h311 == _T_40[9:0] ? 4'h5 : _GEN_2551; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2553 = 10'h312 == _T_40[9:0] ? 4'h6 : _GEN_2552; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2554 = 10'h313 == _T_40[9:0] ? 4'h7 : _GEN_2553; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2555 = 10'h314 == _T_40[9:0] ? 4'h7 : _GEN_2554; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2556 = 10'h315 == _T_40[9:0] ? 4'h3 : _GEN_2555; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2557 = 10'h316 == _T_40[9:0] ? 4'h2 : _GEN_2556; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2558 = 10'h317 == _T_40[9:0] ? 4'h2 : _GEN_2557; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2559 = 10'h318 == _T_40[9:0] ? 4'h2 : _GEN_2558; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2560 = 10'h319 == _T_40[9:0] ? 4'h2 : _GEN_2559; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2561 = 10'h31a == _T_40[9:0] ? 4'h2 : _GEN_2560; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2562 = 10'h31b == _T_40[9:0] ? 4'h2 : _GEN_2561; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2563 = 10'h31c == _T_40[9:0] ? 4'h2 : _GEN_2562; // @[Filter.scala 230:142]
  wire [3:0] _GEN_2564 = 10'h31d == _T_40[9:0] ? 4'h2 : _GEN_2563; // @[Filter.scala 230:142]
  wire [7:0] _T_54 = _GEN_2564 * 4'ha; // @[Filter.scala 230:142]
  wire [10:0] _GEN_38959 = {{3'd0}, _T_54}; // @[Filter.scala 230:109]
  wire [10:0] _T_56 = _T_49 + _GEN_38959; // @[Filter.scala 230:109]
  wire [10:0] _T_57 = _T_56 / 11'h64; // @[Filter.scala 230:150]
  wire  _T_59 = _T_30 >= 6'h20; // @[Filter.scala 233:31]
  wire  _T_63 = _T_37 >= 32'h12; // @[Filter.scala 233:63]
  wire  _T_64 = _T_59 | _T_63; // @[Filter.scala 233:58]
  wire [10:0] _GEN_3363 = io_SPI_distort ? _T_57 : {{7'd0}, _GEN_968}; // @[Filter.scala 235:35]
  wire [10:0] _GEN_3364 = _T_64 ? 11'h0 : _GEN_3363; // @[Filter.scala 233:80]
  wire [10:0] _GEN_4163 = io_SPI_distort ? _T_57 : {{7'd0}, _GEN_1766}; // @[Filter.scala 235:35]
  wire [10:0] _GEN_4164 = _T_64 ? 11'h0 : _GEN_4163; // @[Filter.scala 233:80]
  wire [10:0] _GEN_4963 = io_SPI_distort ? _T_57 : {{7'd0}, _GEN_2564}; // @[Filter.scala 235:35]
  wire [10:0] _GEN_4964 = _T_64 ? 11'h0 : _GEN_4963; // @[Filter.scala 233:80]
  wire [31:0] _T_92 = pixelIndex + 32'h1; // @[Filter.scala 228:31]
  wire [31:0] _GEN_1 = _T_92 % 32'h20; // @[Filter.scala 228:38]
  wire [5:0] _T_93 = _GEN_1[5:0]; // @[Filter.scala 228:38]
  wire [5:0] _T_95 = _T_93 + _GEN_38951; // @[Filter.scala 228:53]
  wire [5:0] _T_97 = _T_95 - 6'h1; // @[Filter.scala 228:69]
  wire [31:0] _T_100 = _T_92 / 32'h20; // @[Filter.scala 229:38]
  wire [31:0] _T_102 = _T_100 + _GEN_38952; // @[Filter.scala 229:53]
  wire [31:0] _T_104 = _T_102 - 32'h1; // @[Filter.scala 229:69]
  wire [37:0] _T_105 = _T_104 * 32'h20; // @[Filter.scala 230:42]
  wire [37:0] _GEN_38965 = {{32'd0}, _T_97}; // @[Filter.scala 230:57]
  wire [37:0] _T_107 = _T_105 + _GEN_38965; // @[Filter.scala 230:57]
  wire [3:0] _GEN_4987 = 10'h16 == _T_107[9:0] ? 4'h9 : 4'ha; // @[Filter.scala 230:62]
  wire [3:0] _GEN_4988 = 10'h17 == _T_107[9:0] ? 4'h3 : _GEN_4987; // @[Filter.scala 230:62]
  wire [3:0] _GEN_4989 = 10'h18 == _T_107[9:0] ? 4'h6 : _GEN_4988; // @[Filter.scala 230:62]
  wire [3:0] _GEN_4990 = 10'h19 == _T_107[9:0] ? 4'ha : _GEN_4989; // @[Filter.scala 230:62]
  wire [3:0] _GEN_4991 = 10'h1a == _T_107[9:0] ? 4'ha : _GEN_4990; // @[Filter.scala 230:62]
  wire [3:0] _GEN_4992 = 10'h1b == _T_107[9:0] ? 4'ha : _GEN_4991; // @[Filter.scala 230:62]
  wire [3:0] _GEN_4993 = 10'h1c == _T_107[9:0] ? 4'ha : _GEN_4992; // @[Filter.scala 230:62]
  wire [3:0] _GEN_4994 = 10'h1d == _T_107[9:0] ? 4'ha : _GEN_4993; // @[Filter.scala 230:62]
  wire [3:0] _GEN_4995 = 10'h1e == _T_107[9:0] ? 4'ha : _GEN_4994; // @[Filter.scala 230:62]
  wire [3:0] _GEN_4996 = 10'h1f == _T_107[9:0] ? 4'ha : _GEN_4995; // @[Filter.scala 230:62]
  wire [3:0] _GEN_4997 = 10'h20 == _T_107[9:0] ? 4'ha : _GEN_4996; // @[Filter.scala 230:62]
  wire [3:0] _GEN_4998 = 10'h21 == _T_107[9:0] ? 4'ha : _GEN_4997; // @[Filter.scala 230:62]
  wire [3:0] _GEN_4999 = 10'h22 == _T_107[9:0] ? 4'ha : _GEN_4998; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5000 = 10'h23 == _T_107[9:0] ? 4'ha : _GEN_4999; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5001 = 10'h24 == _T_107[9:0] ? 4'ha : _GEN_5000; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5002 = 10'h25 == _T_107[9:0] ? 4'ha : _GEN_5001; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5003 = 10'h26 == _T_107[9:0] ? 4'ha : _GEN_5002; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5004 = 10'h27 == _T_107[9:0] ? 4'ha : _GEN_5003; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5005 = 10'h28 == _T_107[9:0] ? 4'ha : _GEN_5004; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5006 = 10'h29 == _T_107[9:0] ? 4'ha : _GEN_5005; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5007 = 10'h2a == _T_107[9:0] ? 4'ha : _GEN_5006; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5008 = 10'h2b == _T_107[9:0] ? 4'ha : _GEN_5007; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5009 = 10'h2c == _T_107[9:0] ? 4'ha : _GEN_5008; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5010 = 10'h2d == _T_107[9:0] ? 4'ha : _GEN_5009; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5011 = 10'h2e == _T_107[9:0] ? 4'ha : _GEN_5010; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5012 = 10'h2f == _T_107[9:0] ? 4'ha : _GEN_5011; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5013 = 10'h30 == _T_107[9:0] ? 4'ha : _GEN_5012; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5014 = 10'h31 == _T_107[9:0] ? 4'ha : _GEN_5013; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5015 = 10'h32 == _T_107[9:0] ? 4'ha : _GEN_5014; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5016 = 10'h33 == _T_107[9:0] ? 4'ha : _GEN_5015; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5017 = 10'h34 == _T_107[9:0] ? 4'ha : _GEN_5016; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5018 = 10'h35 == _T_107[9:0] ? 4'ha : _GEN_5017; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5019 = 10'h36 == _T_107[9:0] ? 4'ha : _GEN_5018; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5020 = 10'h37 == _T_107[9:0] ? 4'ha : _GEN_5019; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5021 = 10'h38 == _T_107[9:0] ? 4'ha : _GEN_5020; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5022 = 10'h39 == _T_107[9:0] ? 4'ha : _GEN_5021; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5023 = 10'h3a == _T_107[9:0] ? 4'ha : _GEN_5022; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5024 = 10'h3b == _T_107[9:0] ? 4'h9 : _GEN_5023; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5025 = 10'h3c == _T_107[9:0] ? 4'h4 : _GEN_5024; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5026 = 10'h3d == _T_107[9:0] ? 4'h3 : _GEN_5025; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5027 = 10'h3e == _T_107[9:0] ? 4'h4 : _GEN_5026; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5028 = 10'h3f == _T_107[9:0] ? 4'ha : _GEN_5027; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5029 = 10'h40 == _T_107[9:0] ? 4'ha : _GEN_5028; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5030 = 10'h41 == _T_107[9:0] ? 4'ha : _GEN_5029; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5031 = 10'h42 == _T_107[9:0] ? 4'ha : _GEN_5030; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5032 = 10'h43 == _T_107[9:0] ? 4'ha : _GEN_5031; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5033 = 10'h44 == _T_107[9:0] ? 4'ha : _GEN_5032; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5034 = 10'h45 == _T_107[9:0] ? 4'ha : _GEN_5033; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5035 = 10'h46 == _T_107[9:0] ? 4'ha : _GEN_5034; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5036 = 10'h47 == _T_107[9:0] ? 4'ha : _GEN_5035; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5037 = 10'h48 == _T_107[9:0] ? 4'ha : _GEN_5036; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5038 = 10'h49 == _T_107[9:0] ? 4'ha : _GEN_5037; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5039 = 10'h4a == _T_107[9:0] ? 4'ha : _GEN_5038; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5040 = 10'h4b == _T_107[9:0] ? 4'ha : _GEN_5039; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5041 = 10'h4c == _T_107[9:0] ? 4'ha : _GEN_5040; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5042 = 10'h4d == _T_107[9:0] ? 4'ha : _GEN_5041; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5043 = 10'h4e == _T_107[9:0] ? 4'ha : _GEN_5042; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5044 = 10'h4f == _T_107[9:0] ? 4'ha : _GEN_5043; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5045 = 10'h50 == _T_107[9:0] ? 4'ha : _GEN_5044; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5046 = 10'h51 == _T_107[9:0] ? 4'ha : _GEN_5045; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5047 = 10'h52 == _T_107[9:0] ? 4'ha : _GEN_5046; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5048 = 10'h53 == _T_107[9:0] ? 4'ha : _GEN_5047; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5049 = 10'h54 == _T_107[9:0] ? 4'ha : _GEN_5048; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5050 = 10'h55 == _T_107[9:0] ? 4'ha : _GEN_5049; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5051 = 10'h56 == _T_107[9:0] ? 4'ha : _GEN_5050; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5052 = 10'h57 == _T_107[9:0] ? 4'ha : _GEN_5051; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5053 = 10'h58 == _T_107[9:0] ? 4'ha : _GEN_5052; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5054 = 10'h59 == _T_107[9:0] ? 4'ha : _GEN_5053; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5055 = 10'h5a == _T_107[9:0] ? 4'h7 : _GEN_5054; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5056 = 10'h5b == _T_107[9:0] ? 4'h7 : _GEN_5055; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5057 = 10'h5c == _T_107[9:0] ? 4'ha : _GEN_5056; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5058 = 10'h5d == _T_107[9:0] ? 4'ha : _GEN_5057; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5059 = 10'h5e == _T_107[9:0] ? 4'ha : _GEN_5058; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5060 = 10'h5f == _T_107[9:0] ? 4'ha : _GEN_5059; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5061 = 10'h60 == _T_107[9:0] ? 4'ha : _GEN_5060; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5062 = 10'h61 == _T_107[9:0] ? 4'h8 : _GEN_5061; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5063 = 10'h62 == _T_107[9:0] ? 4'h3 : _GEN_5062; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5064 = 10'h63 == _T_107[9:0] ? 4'h3 : _GEN_5063; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5065 = 10'h64 == _T_107[9:0] ? 4'h3 : _GEN_5064; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5066 = 10'h65 == _T_107[9:0] ? 4'h9 : _GEN_5065; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5067 = 10'h66 == _T_107[9:0] ? 4'ha : _GEN_5066; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5068 = 10'h67 == _T_107[9:0] ? 4'ha : _GEN_5067; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5069 = 10'h68 == _T_107[9:0] ? 4'ha : _GEN_5068; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5070 = 10'h69 == _T_107[9:0] ? 4'ha : _GEN_5069; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5071 = 10'h6a == _T_107[9:0] ? 4'ha : _GEN_5070; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5072 = 10'h6b == _T_107[9:0] ? 4'h8 : _GEN_5071; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5073 = 10'h6c == _T_107[9:0] ? 4'h5 : _GEN_5072; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5074 = 10'h6d == _T_107[9:0] ? 4'h8 : _GEN_5073; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5075 = 10'h6e == _T_107[9:0] ? 4'ha : _GEN_5074; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5076 = 10'h6f == _T_107[9:0] ? 4'ha : _GEN_5075; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5077 = 10'h70 == _T_107[9:0] ? 4'ha : _GEN_5076; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5078 = 10'h71 == _T_107[9:0] ? 4'ha : _GEN_5077; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5079 = 10'h72 == _T_107[9:0] ? 4'ha : _GEN_5078; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5080 = 10'h73 == _T_107[9:0] ? 4'ha : _GEN_5079; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5081 = 10'h74 == _T_107[9:0] ? 4'ha : _GEN_5080; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5082 = 10'h75 == _T_107[9:0] ? 4'ha : _GEN_5081; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5083 = 10'h76 == _T_107[9:0] ? 4'ha : _GEN_5082; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5084 = 10'h77 == _T_107[9:0] ? 4'ha : _GEN_5083; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5085 = 10'h78 == _T_107[9:0] ? 4'ha : _GEN_5084; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5086 = 10'h79 == _T_107[9:0] ? 4'ha : _GEN_5085; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5087 = 10'h7a == _T_107[9:0] ? 4'ha : _GEN_5086; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5088 = 10'h7b == _T_107[9:0] ? 4'ha : _GEN_5087; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5089 = 10'h7c == _T_107[9:0] ? 4'ha : _GEN_5088; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5090 = 10'h7d == _T_107[9:0] ? 4'ha : _GEN_5089; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5091 = 10'h7e == _T_107[9:0] ? 4'ha : _GEN_5090; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5092 = 10'h7f == _T_107[9:0] ? 4'ha : _GEN_5091; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5093 = 10'h80 == _T_107[9:0] ? 4'ha : _GEN_5092; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5094 = 10'h81 == _T_107[9:0] ? 4'h5 : _GEN_5093; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5095 = 10'h82 == _T_107[9:0] ? 4'h5 : _GEN_5094; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5096 = 10'h83 == _T_107[9:0] ? 4'h7 : _GEN_5095; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5097 = 10'h84 == _T_107[9:0] ? 4'ha : _GEN_5096; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5098 = 10'h85 == _T_107[9:0] ? 4'ha : _GEN_5097; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5099 = 10'h86 == _T_107[9:0] ? 4'ha : _GEN_5098; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5100 = 10'h87 == _T_107[9:0] ? 4'h5 : _GEN_5099; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5101 = 10'h88 == _T_107[9:0] ? 4'h3 : _GEN_5100; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5102 = 10'h89 == _T_107[9:0] ? 4'h3 : _GEN_5101; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5103 = 10'h8a == _T_107[9:0] ? 4'h4 : _GEN_5102; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5104 = 10'h8b == _T_107[9:0] ? 4'h9 : _GEN_5103; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5105 = 10'h8c == _T_107[9:0] ? 4'ha : _GEN_5104; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5106 = 10'h8d == _T_107[9:0] ? 4'ha : _GEN_5105; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5107 = 10'h8e == _T_107[9:0] ? 4'ha : _GEN_5106; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5108 = 10'h8f == _T_107[9:0] ? 4'h6 : _GEN_5107; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5109 = 10'h90 == _T_107[9:0] ? 4'h4 : _GEN_5108; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5110 = 10'h91 == _T_107[9:0] ? 4'h3 : _GEN_5109; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5111 = 10'h92 == _T_107[9:0] ? 4'h7 : _GEN_5110; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5112 = 10'h93 == _T_107[9:0] ? 4'ha : _GEN_5111; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5113 = 10'h94 == _T_107[9:0] ? 4'ha : _GEN_5112; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5114 = 10'h95 == _T_107[9:0] ? 4'ha : _GEN_5113; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5115 = 10'h96 == _T_107[9:0] ? 4'ha : _GEN_5114; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5116 = 10'h97 == _T_107[9:0] ? 4'ha : _GEN_5115; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5117 = 10'h98 == _T_107[9:0] ? 4'ha : _GEN_5116; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5118 = 10'h99 == _T_107[9:0] ? 4'ha : _GEN_5117; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5119 = 10'h9a == _T_107[9:0] ? 4'ha : _GEN_5118; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5120 = 10'h9b == _T_107[9:0] ? 4'ha : _GEN_5119; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5121 = 10'h9c == _T_107[9:0] ? 4'ha : _GEN_5120; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5122 = 10'h9d == _T_107[9:0] ? 4'ha : _GEN_5121; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5123 = 10'h9e == _T_107[9:0] ? 4'ha : _GEN_5122; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5124 = 10'h9f == _T_107[9:0] ? 4'ha : _GEN_5123; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5125 = 10'ha0 == _T_107[9:0] ? 4'ha : _GEN_5124; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5126 = 10'ha1 == _T_107[9:0] ? 4'ha : _GEN_5125; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5127 = 10'ha2 == _T_107[9:0] ? 4'ha : _GEN_5126; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5128 = 10'ha3 == _T_107[9:0] ? 4'ha : _GEN_5127; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5129 = 10'ha4 == _T_107[9:0] ? 4'ha : _GEN_5128; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5130 = 10'ha5 == _T_107[9:0] ? 4'ha : _GEN_5129; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5131 = 10'ha6 == _T_107[9:0] ? 4'ha : _GEN_5130; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5132 = 10'ha7 == _T_107[9:0] ? 4'h9 : _GEN_5131; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5133 = 10'ha8 == _T_107[9:0] ? 4'h4 : _GEN_5132; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5134 = 10'ha9 == _T_107[9:0] ? 4'h3 : _GEN_5133; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5135 = 10'haa == _T_107[9:0] ? 4'h4 : _GEN_5134; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5136 = 10'hab == _T_107[9:0] ? 4'h7 : _GEN_5135; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5137 = 10'hac == _T_107[9:0] ? 4'h8 : _GEN_5136; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5138 = 10'had == _T_107[9:0] ? 4'h3 : _GEN_5137; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5139 = 10'hae == _T_107[9:0] ? 4'h3 : _GEN_5138; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5140 = 10'haf == _T_107[9:0] ? 4'h3 : _GEN_5139; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5141 = 10'hb0 == _T_107[9:0] ? 4'h3 : _GEN_5140; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5142 = 10'hb1 == _T_107[9:0] ? 4'h7 : _GEN_5141; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5143 = 10'hb2 == _T_107[9:0] ? 4'h9 : _GEN_5142; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5144 = 10'hb3 == _T_107[9:0] ? 4'h6 : _GEN_5143; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5145 = 10'hb4 == _T_107[9:0] ? 4'h4 : _GEN_5144; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5146 = 10'hb5 == _T_107[9:0] ? 4'h3 : _GEN_5145; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5147 = 10'hb6 == _T_107[9:0] ? 4'h3 : _GEN_5146; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5148 = 10'hb7 == _T_107[9:0] ? 4'h6 : _GEN_5147; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5149 = 10'hb8 == _T_107[9:0] ? 4'ha : _GEN_5148; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5150 = 10'hb9 == _T_107[9:0] ? 4'ha : _GEN_5149; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5151 = 10'hba == _T_107[9:0] ? 4'ha : _GEN_5150; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5152 = 10'hbb == _T_107[9:0] ? 4'ha : _GEN_5151; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5153 = 10'hbc == _T_107[9:0] ? 4'ha : _GEN_5152; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5154 = 10'hbd == _T_107[9:0] ? 4'h9 : _GEN_5153; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5155 = 10'hbe == _T_107[9:0] ? 4'ha : _GEN_5154; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5156 = 10'hbf == _T_107[9:0] ? 4'ha : _GEN_5155; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5157 = 10'hc0 == _T_107[9:0] ? 4'ha : _GEN_5156; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5158 = 10'hc1 == _T_107[9:0] ? 4'ha : _GEN_5157; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5159 = 10'hc2 == _T_107[9:0] ? 4'ha : _GEN_5158; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5160 = 10'hc3 == _T_107[9:0] ? 4'ha : _GEN_5159; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5161 = 10'hc4 == _T_107[9:0] ? 4'ha : _GEN_5160; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5162 = 10'hc5 == _T_107[9:0] ? 4'ha : _GEN_5161; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5163 = 10'hc6 == _T_107[9:0] ? 4'ha : _GEN_5162; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5164 = 10'hc7 == _T_107[9:0] ? 4'h9 : _GEN_5163; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5165 = 10'hc8 == _T_107[9:0] ? 4'h8 : _GEN_5164; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5166 = 10'hc9 == _T_107[9:0] ? 4'h8 : _GEN_5165; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5167 = 10'hca == _T_107[9:0] ? 4'h9 : _GEN_5166; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5168 = 10'hcb == _T_107[9:0] ? 4'ha : _GEN_5167; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5169 = 10'hcc == _T_107[9:0] ? 4'ha : _GEN_5168; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5170 = 10'hcd == _T_107[9:0] ? 4'ha : _GEN_5169; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5171 = 10'hce == _T_107[9:0] ? 4'h8 : _GEN_5170; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5172 = 10'hcf == _T_107[9:0] ? 4'h3 : _GEN_5171; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5173 = 10'hd0 == _T_107[9:0] ? 4'h3 : _GEN_5172; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5174 = 10'hd1 == _T_107[9:0] ? 4'h3 : _GEN_5173; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5175 = 10'hd2 == _T_107[9:0] ? 4'h4 : _GEN_5174; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5176 = 10'hd3 == _T_107[9:0] ? 4'h3 : _GEN_5175; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5177 = 10'hd4 == _T_107[9:0] ? 4'h3 : _GEN_5176; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5178 = 10'hd5 == _T_107[9:0] ? 4'h3 : _GEN_5177; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5179 = 10'hd6 == _T_107[9:0] ? 4'h3 : _GEN_5178; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5180 = 10'hd7 == _T_107[9:0] ? 4'h5 : _GEN_5179; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5181 = 10'hd8 == _T_107[9:0] ? 4'h4 : _GEN_5180; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5182 = 10'hd9 == _T_107[9:0] ? 4'h3 : _GEN_5181; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5183 = 10'hda == _T_107[9:0] ? 4'h3 : _GEN_5182; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5184 = 10'hdb == _T_107[9:0] ? 4'h3 : _GEN_5183; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5185 = 10'hdc == _T_107[9:0] ? 4'h4 : _GEN_5184; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5186 = 10'hdd == _T_107[9:0] ? 4'ha : _GEN_5185; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5187 = 10'hde == _T_107[9:0] ? 4'ha : _GEN_5186; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5188 = 10'hdf == _T_107[9:0] ? 4'ha : _GEN_5187; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5189 = 10'he0 == _T_107[9:0] ? 4'ha : _GEN_5188; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5190 = 10'he1 == _T_107[9:0] ? 4'ha : _GEN_5189; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5191 = 10'he2 == _T_107[9:0] ? 4'ha : _GEN_5190; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5192 = 10'he3 == _T_107[9:0] ? 4'h5 : _GEN_5191; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5193 = 10'he4 == _T_107[9:0] ? 4'ha : _GEN_5192; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5194 = 10'he5 == _T_107[9:0] ? 4'ha : _GEN_5193; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5195 = 10'he6 == _T_107[9:0] ? 4'ha : _GEN_5194; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5196 = 10'he7 == _T_107[9:0] ? 4'ha : _GEN_5195; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5197 = 10'he8 == _T_107[9:0] ? 4'ha : _GEN_5196; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5198 = 10'he9 == _T_107[9:0] ? 4'ha : _GEN_5197; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5199 = 10'hea == _T_107[9:0] ? 4'ha : _GEN_5198; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5200 = 10'heb == _T_107[9:0] ? 4'h9 : _GEN_5199; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5201 = 10'hec == _T_107[9:0] ? 4'h7 : _GEN_5200; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5202 = 10'hed == _T_107[9:0] ? 4'h3 : _GEN_5201; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5203 = 10'hee == _T_107[9:0] ? 4'h3 : _GEN_5202; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5204 = 10'hef == _T_107[9:0] ? 4'h3 : _GEN_5203; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5205 = 10'hf0 == _T_107[9:0] ? 4'h4 : _GEN_5204; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5206 = 10'hf1 == _T_107[9:0] ? 4'h7 : _GEN_5205; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5207 = 10'hf2 == _T_107[9:0] ? 4'ha : _GEN_5206; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5208 = 10'hf3 == _T_107[9:0] ? 4'ha : _GEN_5207; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5209 = 10'hf4 == _T_107[9:0] ? 4'ha : _GEN_5208; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5210 = 10'hf5 == _T_107[9:0] ? 4'h7 : _GEN_5209; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5211 = 10'hf6 == _T_107[9:0] ? 4'h3 : _GEN_5210; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5212 = 10'hf7 == _T_107[9:0] ? 4'h3 : _GEN_5211; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5213 = 10'hf8 == _T_107[9:0] ? 4'h3 : _GEN_5212; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5214 = 10'hf9 == _T_107[9:0] ? 4'h3 : _GEN_5213; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5215 = 10'hfa == _T_107[9:0] ? 4'h3 : _GEN_5214; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5216 = 10'hfb == _T_107[9:0] ? 4'h3 : _GEN_5215; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5217 = 10'hfc == _T_107[9:0] ? 4'h3 : _GEN_5216; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5218 = 10'hfd == _T_107[9:0] ? 4'h3 : _GEN_5217; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5219 = 10'hfe == _T_107[9:0] ? 4'h3 : _GEN_5218; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5220 = 10'hff == _T_107[9:0] ? 4'h3 : _GEN_5219; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5221 = 10'h100 == _T_107[9:0] ? 4'h3 : _GEN_5220; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5222 = 10'h101 == _T_107[9:0] ? 4'h4 : _GEN_5221; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5223 = 10'h102 == _T_107[9:0] ? 4'h6 : _GEN_5222; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5224 = 10'h103 == _T_107[9:0] ? 4'ha : _GEN_5223; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5225 = 10'h104 == _T_107[9:0] ? 4'ha : _GEN_5224; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5226 = 10'h105 == _T_107[9:0] ? 4'h9 : _GEN_5225; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5227 = 10'h106 == _T_107[9:0] ? 4'h9 : _GEN_5226; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5228 = 10'h107 == _T_107[9:0] ? 4'h9 : _GEN_5227; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5229 = 10'h108 == _T_107[9:0] ? 4'h9 : _GEN_5228; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5230 = 10'h109 == _T_107[9:0] ? 4'h3 : _GEN_5229; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5231 = 10'h10a == _T_107[9:0] ? 4'ha : _GEN_5230; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5232 = 10'h10b == _T_107[9:0] ? 4'ha : _GEN_5231; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5233 = 10'h10c == _T_107[9:0] ? 4'ha : _GEN_5232; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5234 = 10'h10d == _T_107[9:0] ? 4'ha : _GEN_5233; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5235 = 10'h10e == _T_107[9:0] ? 4'ha : _GEN_5234; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5236 = 10'h10f == _T_107[9:0] ? 4'h9 : _GEN_5235; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5237 = 10'h110 == _T_107[9:0] ? 4'h9 : _GEN_5236; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5238 = 10'h111 == _T_107[9:0] ? 4'h4 : _GEN_5237; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5239 = 10'h112 == _T_107[9:0] ? 4'h8 : _GEN_5238; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5240 = 10'h113 == _T_107[9:0] ? 4'h3 : _GEN_5239; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5241 = 10'h114 == _T_107[9:0] ? 4'h3 : _GEN_5240; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5242 = 10'h115 == _T_107[9:0] ? 4'h4 : _GEN_5241; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5243 = 10'h116 == _T_107[9:0] ? 4'h4 : _GEN_5242; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5244 = 10'h117 == _T_107[9:0] ? 4'h3 : _GEN_5243; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5245 = 10'h118 == _T_107[9:0] ? 4'h8 : _GEN_5244; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5246 = 10'h119 == _T_107[9:0] ? 4'ha : _GEN_5245; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5247 = 10'h11a == _T_107[9:0] ? 4'ha : _GEN_5246; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5248 = 10'h11b == _T_107[9:0] ? 4'ha : _GEN_5247; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5249 = 10'h11c == _T_107[9:0] ? 4'h6 : _GEN_5248; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5250 = 10'h11d == _T_107[9:0] ? 4'h3 : _GEN_5249; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5251 = 10'h11e == _T_107[9:0] ? 4'h3 : _GEN_5250; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5252 = 10'h11f == _T_107[9:0] ? 4'h3 : _GEN_5251; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5253 = 10'h120 == _T_107[9:0] ? 4'h3 : _GEN_5252; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5254 = 10'h121 == _T_107[9:0] ? 4'h3 : _GEN_5253; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5255 = 10'h122 == _T_107[9:0] ? 4'h3 : _GEN_5254; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5256 = 10'h123 == _T_107[9:0] ? 4'h3 : _GEN_5255; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5257 = 10'h124 == _T_107[9:0] ? 4'h3 : _GEN_5256; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5258 = 10'h125 == _T_107[9:0] ? 4'h3 : _GEN_5257; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5259 = 10'h126 == _T_107[9:0] ? 4'h4 : _GEN_5258; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5260 = 10'h127 == _T_107[9:0] ? 4'h6 : _GEN_5259; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5261 = 10'h128 == _T_107[9:0] ? 4'h5 : _GEN_5260; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5262 = 10'h129 == _T_107[9:0] ? 4'h8 : _GEN_5261; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5263 = 10'h12a == _T_107[9:0] ? 4'h5 : _GEN_5262; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5264 = 10'h12b == _T_107[9:0] ? 4'h3 : _GEN_5263; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5265 = 10'h12c == _T_107[9:0] ? 4'h3 : _GEN_5264; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5266 = 10'h12d == _T_107[9:0] ? 4'h3 : _GEN_5265; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5267 = 10'h12e == _T_107[9:0] ? 4'h4 : _GEN_5266; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5268 = 10'h12f == _T_107[9:0] ? 4'h4 : _GEN_5267; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5269 = 10'h130 == _T_107[9:0] ? 4'ha : _GEN_5268; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5270 = 10'h131 == _T_107[9:0] ? 4'h9 : _GEN_5269; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5271 = 10'h132 == _T_107[9:0] ? 4'h9 : _GEN_5270; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5272 = 10'h133 == _T_107[9:0] ? 4'h8 : _GEN_5271; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5273 = 10'h134 == _T_107[9:0] ? 4'h9 : _GEN_5272; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5274 = 10'h135 == _T_107[9:0] ? 4'h8 : _GEN_5273; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5275 = 10'h136 == _T_107[9:0] ? 4'h7 : _GEN_5274; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5276 = 10'h137 == _T_107[9:0] ? 4'h6 : _GEN_5275; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5277 = 10'h138 == _T_107[9:0] ? 4'h8 : _GEN_5276; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5278 = 10'h139 == _T_107[9:0] ? 4'h3 : _GEN_5277; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5279 = 10'h13a == _T_107[9:0] ? 4'h3 : _GEN_5278; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5280 = 10'h13b == _T_107[9:0] ? 4'h4 : _GEN_5279; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5281 = 10'h13c == _T_107[9:0] ? 4'h4 : _GEN_5280; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5282 = 10'h13d == _T_107[9:0] ? 4'h3 : _GEN_5281; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5283 = 10'h13e == _T_107[9:0] ? 4'h5 : _GEN_5282; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5284 = 10'h13f == _T_107[9:0] ? 4'h9 : _GEN_5283; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5285 = 10'h140 == _T_107[9:0] ? 4'ha : _GEN_5284; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5286 = 10'h141 == _T_107[9:0] ? 4'ha : _GEN_5285; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5287 = 10'h142 == _T_107[9:0] ? 4'ha : _GEN_5286; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5288 = 10'h143 == _T_107[9:0] ? 4'h5 : _GEN_5287; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5289 = 10'h144 == _T_107[9:0] ? 4'h3 : _GEN_5288; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5290 = 10'h145 == _T_107[9:0] ? 4'h3 : _GEN_5289; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5291 = 10'h146 == _T_107[9:0] ? 4'h3 : _GEN_5290; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5292 = 10'h147 == _T_107[9:0] ? 4'h4 : _GEN_5291; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5293 = 10'h148 == _T_107[9:0] ? 4'h3 : _GEN_5292; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5294 = 10'h149 == _T_107[9:0] ? 4'h3 : _GEN_5293; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5295 = 10'h14a == _T_107[9:0] ? 4'h3 : _GEN_5294; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5296 = 10'h14b == _T_107[9:0] ? 4'h6 : _GEN_5295; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5297 = 10'h14c == _T_107[9:0] ? 4'h8 : _GEN_5296; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5298 = 10'h14d == _T_107[9:0] ? 4'h5 : _GEN_5297; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5299 = 10'h14e == _T_107[9:0] ? 4'h4 : _GEN_5298; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5300 = 10'h14f == _T_107[9:0] ? 4'h3 : _GEN_5299; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5301 = 10'h150 == _T_107[9:0] ? 4'h3 : _GEN_5300; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5302 = 10'h151 == _T_107[9:0] ? 4'h3 : _GEN_5301; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5303 = 10'h152 == _T_107[9:0] ? 4'h3 : _GEN_5302; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5304 = 10'h153 == _T_107[9:0] ? 4'h3 : _GEN_5303; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5305 = 10'h154 == _T_107[9:0] ? 4'h3 : _GEN_5304; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5306 = 10'h155 == _T_107[9:0] ? 4'h4 : _GEN_5305; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5307 = 10'h156 == _T_107[9:0] ? 4'h9 : _GEN_5306; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5308 = 10'h157 == _T_107[9:0] ? 4'h8 : _GEN_5307; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5309 = 10'h158 == _T_107[9:0] ? 4'h8 : _GEN_5308; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5310 = 10'h159 == _T_107[9:0] ? 4'h8 : _GEN_5309; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5311 = 10'h15a == _T_107[9:0] ? 4'h8 : _GEN_5310; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5312 = 10'h15b == _T_107[9:0] ? 4'h8 : _GEN_5311; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5313 = 10'h15c == _T_107[9:0] ? 4'h7 : _GEN_5312; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5314 = 10'h15d == _T_107[9:0] ? 4'h7 : _GEN_5313; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5315 = 10'h15e == _T_107[9:0] ? 4'h8 : _GEN_5314; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5316 = 10'h15f == _T_107[9:0] ? 4'h3 : _GEN_5315; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5317 = 10'h160 == _T_107[9:0] ? 4'h4 : _GEN_5316; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5318 = 10'h161 == _T_107[9:0] ? 4'h4 : _GEN_5317; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5319 = 10'h162 == _T_107[9:0] ? 4'h4 : _GEN_5318; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5320 = 10'h163 == _T_107[9:0] ? 4'h4 : _GEN_5319; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5321 = 10'h164 == _T_107[9:0] ? 4'h5 : _GEN_5320; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5322 = 10'h165 == _T_107[9:0] ? 4'ha : _GEN_5321; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5323 = 10'h166 == _T_107[9:0] ? 4'h9 : _GEN_5322; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5324 = 10'h167 == _T_107[9:0] ? 4'ha : _GEN_5323; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5325 = 10'h168 == _T_107[9:0] ? 4'ha : _GEN_5324; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5326 = 10'h169 == _T_107[9:0] ? 4'h6 : _GEN_5325; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5327 = 10'h16a == _T_107[9:0] ? 4'h3 : _GEN_5326; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5328 = 10'h16b == _T_107[9:0] ? 4'h3 : _GEN_5327; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5329 = 10'h16c == _T_107[9:0] ? 4'h3 : _GEN_5328; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5330 = 10'h16d == _T_107[9:0] ? 4'h4 : _GEN_5329; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5331 = 10'h16e == _T_107[9:0] ? 4'h3 : _GEN_5330; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5332 = 10'h16f == _T_107[9:0] ? 4'h3 : _GEN_5331; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5333 = 10'h170 == _T_107[9:0] ? 4'h3 : _GEN_5332; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5334 = 10'h171 == _T_107[9:0] ? 4'h7 : _GEN_5333; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5335 = 10'h172 == _T_107[9:0] ? 4'ha : _GEN_5334; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5336 = 10'h173 == _T_107[9:0] ? 4'h5 : _GEN_5335; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5337 = 10'h174 == _T_107[9:0] ? 4'h3 : _GEN_5336; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5338 = 10'h175 == _T_107[9:0] ? 4'h4 : _GEN_5337; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5339 = 10'h176 == _T_107[9:0] ? 4'h4 : _GEN_5338; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5340 = 10'h177 == _T_107[9:0] ? 4'h4 : _GEN_5339; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5341 = 10'h178 == _T_107[9:0] ? 4'h4 : _GEN_5340; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5342 = 10'h179 == _T_107[9:0] ? 4'h3 : _GEN_5341; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5343 = 10'h17a == _T_107[9:0] ? 4'h3 : _GEN_5342; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5344 = 10'h17b == _T_107[9:0] ? 4'h3 : _GEN_5343; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5345 = 10'h17c == _T_107[9:0] ? 4'h8 : _GEN_5344; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5346 = 10'h17d == _T_107[9:0] ? 4'h8 : _GEN_5345; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5347 = 10'h17e == _T_107[9:0] ? 4'h8 : _GEN_5346; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5348 = 10'h17f == _T_107[9:0] ? 4'h8 : _GEN_5347; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5349 = 10'h180 == _T_107[9:0] ? 4'h8 : _GEN_5348; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5350 = 10'h181 == _T_107[9:0] ? 4'h8 : _GEN_5349; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5351 = 10'h182 == _T_107[9:0] ? 4'h8 : _GEN_5350; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5352 = 10'h183 == _T_107[9:0] ? 4'h8 : _GEN_5351; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5353 = 10'h184 == _T_107[9:0] ? 4'h8 : _GEN_5352; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5354 = 10'h185 == _T_107[9:0] ? 4'h5 : _GEN_5353; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5355 = 10'h186 == _T_107[9:0] ? 4'h3 : _GEN_5354; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5356 = 10'h187 == _T_107[9:0] ? 4'h4 : _GEN_5355; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5357 = 10'h188 == _T_107[9:0] ? 4'h4 : _GEN_5356; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5358 = 10'h189 == _T_107[9:0] ? 4'h4 : _GEN_5357; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5359 = 10'h18a == _T_107[9:0] ? 4'h5 : _GEN_5358; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5360 = 10'h18b == _T_107[9:0] ? 4'ha : _GEN_5359; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5361 = 10'h18c == _T_107[9:0] ? 4'ha : _GEN_5360; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5362 = 10'h18d == _T_107[9:0] ? 4'h9 : _GEN_5361; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5363 = 10'h18e == _T_107[9:0] ? 4'ha : _GEN_5362; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5364 = 10'h18f == _T_107[9:0] ? 4'h4 : _GEN_5363; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5365 = 10'h190 == _T_107[9:0] ? 4'h3 : _GEN_5364; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5366 = 10'h191 == _T_107[9:0] ? 4'h3 : _GEN_5365; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5367 = 10'h192 == _T_107[9:0] ? 4'h5 : _GEN_5366; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5368 = 10'h193 == _T_107[9:0] ? 4'h6 : _GEN_5367; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5369 = 10'h194 == _T_107[9:0] ? 4'h5 : _GEN_5368; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5370 = 10'h195 == _T_107[9:0] ? 4'h3 : _GEN_5369; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5371 = 10'h196 == _T_107[9:0] ? 4'h3 : _GEN_5370; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5372 = 10'h197 == _T_107[9:0] ? 4'h5 : _GEN_5371; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5373 = 10'h198 == _T_107[9:0] ? 4'ha : _GEN_5372; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5374 = 10'h199 == _T_107[9:0] ? 4'h3 : _GEN_5373; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5375 = 10'h19a == _T_107[9:0] ? 4'h1 : _GEN_5374; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5376 = 10'h19b == _T_107[9:0] ? 4'h2 : _GEN_5375; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5377 = 10'h19c == _T_107[9:0] ? 4'h4 : _GEN_5376; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5378 = 10'h19d == _T_107[9:0] ? 4'h3 : _GEN_5377; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5379 = 10'h19e == _T_107[9:0] ? 4'h1 : _GEN_5378; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5380 = 10'h19f == _T_107[9:0] ? 4'h2 : _GEN_5379; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5381 = 10'h1a0 == _T_107[9:0] ? 4'h3 : _GEN_5380; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5382 = 10'h1a1 == _T_107[9:0] ? 4'h4 : _GEN_5381; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5383 = 10'h1a2 == _T_107[9:0] ? 4'h8 : _GEN_5382; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5384 = 10'h1a3 == _T_107[9:0] ? 4'h8 : _GEN_5383; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5385 = 10'h1a4 == _T_107[9:0] ? 4'h8 : _GEN_5384; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5386 = 10'h1a5 == _T_107[9:0] ? 4'h8 : _GEN_5385; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5387 = 10'h1a6 == _T_107[9:0] ? 4'h7 : _GEN_5386; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5388 = 10'h1a7 == _T_107[9:0] ? 4'h8 : _GEN_5387; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5389 = 10'h1a8 == _T_107[9:0] ? 4'h8 : _GEN_5388; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5390 = 10'h1a9 == _T_107[9:0] ? 4'h8 : _GEN_5389; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5391 = 10'h1aa == _T_107[9:0] ? 4'h7 : _GEN_5390; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5392 = 10'h1ab == _T_107[9:0] ? 4'h4 : _GEN_5391; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5393 = 10'h1ac == _T_107[9:0] ? 4'h4 : _GEN_5392; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5394 = 10'h1ad == _T_107[9:0] ? 4'h3 : _GEN_5393; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5395 = 10'h1ae == _T_107[9:0] ? 4'h3 : _GEN_5394; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5396 = 10'h1af == _T_107[9:0] ? 4'h4 : _GEN_5395; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5397 = 10'h1b0 == _T_107[9:0] ? 4'h6 : _GEN_5396; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5398 = 10'h1b1 == _T_107[9:0] ? 4'ha : _GEN_5397; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5399 = 10'h1b2 == _T_107[9:0] ? 4'ha : _GEN_5398; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5400 = 10'h1b3 == _T_107[9:0] ? 4'h9 : _GEN_5399; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5401 = 10'h1b4 == _T_107[9:0] ? 4'h9 : _GEN_5400; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5402 = 10'h1b5 == _T_107[9:0] ? 4'h3 : _GEN_5401; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5403 = 10'h1b6 == _T_107[9:0] ? 4'h3 : _GEN_5402; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5404 = 10'h1b7 == _T_107[9:0] ? 4'h4 : _GEN_5403; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5405 = 10'h1b8 == _T_107[9:0] ? 4'h5 : _GEN_5404; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5406 = 10'h1b9 == _T_107[9:0] ? 4'h6 : _GEN_5405; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5407 = 10'h1ba == _T_107[9:0] ? 4'h4 : _GEN_5406; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5408 = 10'h1bb == _T_107[9:0] ? 4'h3 : _GEN_5407; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5409 = 10'h1bc == _T_107[9:0] ? 4'h3 : _GEN_5408; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5410 = 10'h1bd == _T_107[9:0] ? 4'h4 : _GEN_5409; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5411 = 10'h1be == _T_107[9:0] ? 4'ha : _GEN_5410; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5412 = 10'h1bf == _T_107[9:0] ? 4'h4 : _GEN_5411; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5413 = 10'h1c0 == _T_107[9:0] ? 4'h5 : _GEN_5412; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5414 = 10'h1c1 == _T_107[9:0] ? 4'h5 : _GEN_5413; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5415 = 10'h1c2 == _T_107[9:0] ? 4'h4 : _GEN_5414; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5416 = 10'h1c3 == _T_107[9:0] ? 4'h5 : _GEN_5415; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5417 = 10'h1c4 == _T_107[9:0] ? 4'h4 : _GEN_5416; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5418 = 10'h1c5 == _T_107[9:0] ? 4'h3 : _GEN_5417; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5419 = 10'h1c6 == _T_107[9:0] ? 4'h4 : _GEN_5418; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5420 = 10'h1c7 == _T_107[9:0] ? 4'h3 : _GEN_5419; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5421 = 10'h1c8 == _T_107[9:0] ? 4'h8 : _GEN_5420; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5422 = 10'h1c9 == _T_107[9:0] ? 4'h8 : _GEN_5421; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5423 = 10'h1ca == _T_107[9:0] ? 4'h8 : _GEN_5422; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5424 = 10'h1cb == _T_107[9:0] ? 4'h8 : _GEN_5423; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5425 = 10'h1cc == _T_107[9:0] ? 4'h8 : _GEN_5424; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5426 = 10'h1cd == _T_107[9:0] ? 4'h8 : _GEN_5425; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5427 = 10'h1ce == _T_107[9:0] ? 4'h8 : _GEN_5426; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5428 = 10'h1cf == _T_107[9:0] ? 4'h8 : _GEN_5427; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5429 = 10'h1d0 == _T_107[9:0] ? 4'h5 : _GEN_5428; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5430 = 10'h1d1 == _T_107[9:0] ? 4'h4 : _GEN_5429; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5431 = 10'h1d2 == _T_107[9:0] ? 4'h6 : _GEN_5430; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5432 = 10'h1d3 == _T_107[9:0] ? 4'h6 : _GEN_5431; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5433 = 10'h1d4 == _T_107[9:0] ? 4'h6 : _GEN_5432; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5434 = 10'h1d5 == _T_107[9:0] ? 4'h5 : _GEN_5433; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5435 = 10'h1d6 == _T_107[9:0] ? 4'h8 : _GEN_5434; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5436 = 10'h1d7 == _T_107[9:0] ? 4'ha : _GEN_5435; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5437 = 10'h1d8 == _T_107[9:0] ? 4'ha : _GEN_5436; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5438 = 10'h1d9 == _T_107[9:0] ? 4'ha : _GEN_5437; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5439 = 10'h1da == _T_107[9:0] ? 4'h6 : _GEN_5438; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5440 = 10'h1db == _T_107[9:0] ? 4'h3 : _GEN_5439; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5441 = 10'h1dc == _T_107[9:0] ? 4'h5 : _GEN_5440; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5442 = 10'h1dd == _T_107[9:0] ? 4'h2 : _GEN_5441; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5443 = 10'h1de == _T_107[9:0] ? 4'h5 : _GEN_5442; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5444 = 10'h1df == _T_107[9:0] ? 4'h5 : _GEN_5443; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5445 = 10'h1e0 == _T_107[9:0] ? 4'h5 : _GEN_5444; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5446 = 10'h1e1 == _T_107[9:0] ? 4'h3 : _GEN_5445; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5447 = 10'h1e2 == _T_107[9:0] ? 4'h3 : _GEN_5446; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5448 = 10'h1e3 == _T_107[9:0] ? 4'h3 : _GEN_5447; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5449 = 10'h1e4 == _T_107[9:0] ? 4'h9 : _GEN_5448; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5450 = 10'h1e5 == _T_107[9:0] ? 4'h4 : _GEN_5449; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5451 = 10'h1e6 == _T_107[9:0] ? 4'h4 : _GEN_5450; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5452 = 10'h1e7 == _T_107[9:0] ? 4'h4 : _GEN_5451; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5453 = 10'h1e8 == _T_107[9:0] ? 4'h4 : _GEN_5452; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5454 = 10'h1e9 == _T_107[9:0] ? 4'h4 : _GEN_5453; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5455 = 10'h1ea == _T_107[9:0] ? 4'h4 : _GEN_5454; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5456 = 10'h1eb == _T_107[9:0] ? 4'h4 : _GEN_5455; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5457 = 10'h1ec == _T_107[9:0] ? 4'h4 : _GEN_5456; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5458 = 10'h1ed == _T_107[9:0] ? 4'h4 : _GEN_5457; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5459 = 10'h1ee == _T_107[9:0] ? 4'h8 : _GEN_5458; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5460 = 10'h1ef == _T_107[9:0] ? 4'h8 : _GEN_5459; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5461 = 10'h1f0 == _T_107[9:0] ? 4'h8 : _GEN_5460; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5462 = 10'h1f1 == _T_107[9:0] ? 4'h8 : _GEN_5461; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5463 = 10'h1f2 == _T_107[9:0] ? 4'h8 : _GEN_5462; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5464 = 10'h1f3 == _T_107[9:0] ? 4'h8 : _GEN_5463; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5465 = 10'h1f4 == _T_107[9:0] ? 4'h9 : _GEN_5464; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5466 = 10'h1f5 == _T_107[9:0] ? 4'h9 : _GEN_5465; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5467 = 10'h1f6 == _T_107[9:0] ? 4'ha : _GEN_5466; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5468 = 10'h1f7 == _T_107[9:0] ? 4'h5 : _GEN_5467; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5469 = 10'h1f8 == _T_107[9:0] ? 4'h5 : _GEN_5468; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5470 = 10'h1f9 == _T_107[9:0] ? 4'h7 : _GEN_5469; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5471 = 10'h1fa == _T_107[9:0] ? 4'h7 : _GEN_5470; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5472 = 10'h1fb == _T_107[9:0] ? 4'h5 : _GEN_5471; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5473 = 10'h1fc == _T_107[9:0] ? 4'ha : _GEN_5472; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5474 = 10'h1fd == _T_107[9:0] ? 4'hb : _GEN_5473; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5475 = 10'h1fe == _T_107[9:0] ? 4'hb : _GEN_5474; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5476 = 10'h1ff == _T_107[9:0] ? 4'ha : _GEN_5475; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5477 = 10'h200 == _T_107[9:0] ? 4'h4 : _GEN_5476; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5478 = 10'h201 == _T_107[9:0] ? 4'h3 : _GEN_5477; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5479 = 10'h202 == _T_107[9:0] ? 4'h2 : _GEN_5478; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5480 = 10'h203 == _T_107[9:0] ? 4'h2 : _GEN_5479; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5481 = 10'h204 == _T_107[9:0] ? 4'h2 : _GEN_5480; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5482 = 10'h205 == _T_107[9:0] ? 4'h2 : _GEN_5481; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5483 = 10'h206 == _T_107[9:0] ? 4'h2 : _GEN_5482; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5484 = 10'h207 == _T_107[9:0] ? 4'h2 : _GEN_5483; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5485 = 10'h208 == _T_107[9:0] ? 4'h3 : _GEN_5484; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5486 = 10'h209 == _T_107[9:0] ? 4'h3 : _GEN_5485; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5487 = 10'h20a == _T_107[9:0] ? 4'h8 : _GEN_5486; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5488 = 10'h20b == _T_107[9:0] ? 4'h4 : _GEN_5487; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5489 = 10'h20c == _T_107[9:0] ? 4'h4 : _GEN_5488; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5490 = 10'h20d == _T_107[9:0] ? 4'h4 : _GEN_5489; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5491 = 10'h20e == _T_107[9:0] ? 4'h4 : _GEN_5490; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5492 = 10'h20f == _T_107[9:0] ? 4'h4 : _GEN_5491; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5493 = 10'h210 == _T_107[9:0] ? 4'h4 : _GEN_5492; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5494 = 10'h211 == _T_107[9:0] ? 4'h4 : _GEN_5493; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5495 = 10'h212 == _T_107[9:0] ? 4'h4 : _GEN_5494; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5496 = 10'h213 == _T_107[9:0] ? 4'h6 : _GEN_5495; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5497 = 10'h214 == _T_107[9:0] ? 4'h7 : _GEN_5496; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5498 = 10'h215 == _T_107[9:0] ? 4'h8 : _GEN_5497; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5499 = 10'h216 == _T_107[9:0] ? 4'h8 : _GEN_5498; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5500 = 10'h217 == _T_107[9:0] ? 4'h8 : _GEN_5499; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5501 = 10'h218 == _T_107[9:0] ? 4'h8 : _GEN_5500; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5502 = 10'h219 == _T_107[9:0] ? 4'h8 : _GEN_5501; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5503 = 10'h21a == _T_107[9:0] ? 4'h8 : _GEN_5502; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5504 = 10'h21b == _T_107[9:0] ? 4'h8 : _GEN_5503; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5505 = 10'h21c == _T_107[9:0] ? 4'ha : _GEN_5504; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5506 = 10'h21d == _T_107[9:0] ? 4'h9 : _GEN_5505; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5507 = 10'h21e == _T_107[9:0] ? 4'h6 : _GEN_5506; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5508 = 10'h21f == _T_107[9:0] ? 4'h4 : _GEN_5507; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5509 = 10'h220 == _T_107[9:0] ? 4'h4 : _GEN_5508; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5510 = 10'h221 == _T_107[9:0] ? 4'h5 : _GEN_5509; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5511 = 10'h222 == _T_107[9:0] ? 4'ha : _GEN_5510; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5512 = 10'h223 == _T_107[9:0] ? 4'ha : _GEN_5511; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5513 = 10'h224 == _T_107[9:0] ? 4'ha : _GEN_5512; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5514 = 10'h225 == _T_107[9:0] ? 4'h8 : _GEN_5513; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5515 = 10'h226 == _T_107[9:0] ? 4'h4 : _GEN_5514; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5516 = 10'h227 == _T_107[9:0] ? 4'h2 : _GEN_5515; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5517 = 10'h228 == _T_107[9:0] ? 4'h2 : _GEN_5516; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5518 = 10'h229 == _T_107[9:0] ? 4'h2 : _GEN_5517; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5519 = 10'h22a == _T_107[9:0] ? 4'h2 : _GEN_5518; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5520 = 10'h22b == _T_107[9:0] ? 4'h2 : _GEN_5519; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5521 = 10'h22c == _T_107[9:0] ? 4'h2 : _GEN_5520; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5522 = 10'h22d == _T_107[9:0] ? 4'h2 : _GEN_5521; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5523 = 10'h22e == _T_107[9:0] ? 4'h2 : _GEN_5522; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5524 = 10'h22f == _T_107[9:0] ? 4'h3 : _GEN_5523; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5525 = 10'h230 == _T_107[9:0] ? 4'h3 : _GEN_5524; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5526 = 10'h231 == _T_107[9:0] ? 4'h3 : _GEN_5525; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5527 = 10'h232 == _T_107[9:0] ? 4'h4 : _GEN_5526; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5528 = 10'h233 == _T_107[9:0] ? 4'h6 : _GEN_5527; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5529 = 10'h234 == _T_107[9:0] ? 4'h6 : _GEN_5528; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5530 = 10'h235 == _T_107[9:0] ? 4'h4 : _GEN_5529; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5531 = 10'h236 == _T_107[9:0] ? 4'h4 : _GEN_5530; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5532 = 10'h237 == _T_107[9:0] ? 4'h4 : _GEN_5531; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5533 = 10'h238 == _T_107[9:0] ? 4'h4 : _GEN_5532; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5534 = 10'h239 == _T_107[9:0] ? 4'h3 : _GEN_5533; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5535 = 10'h23a == _T_107[9:0] ? 4'h7 : _GEN_5534; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5536 = 10'h23b == _T_107[9:0] ? 4'h7 : _GEN_5535; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5537 = 10'h23c == _T_107[9:0] ? 4'h7 : _GEN_5536; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5538 = 10'h23d == _T_107[9:0] ? 4'h7 : _GEN_5537; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5539 = 10'h23e == _T_107[9:0] ? 4'h7 : _GEN_5538; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5540 = 10'h23f == _T_107[9:0] ? 4'h7 : _GEN_5539; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5541 = 10'h240 == _T_107[9:0] ? 4'h7 : _GEN_5540; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5542 = 10'h241 == _T_107[9:0] ? 4'h8 : _GEN_5541; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5543 = 10'h242 == _T_107[9:0] ? 4'ha : _GEN_5542; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5544 = 10'h243 == _T_107[9:0] ? 4'ha : _GEN_5543; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5545 = 10'h244 == _T_107[9:0] ? 4'ha : _GEN_5544; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5546 = 10'h245 == _T_107[9:0] ? 4'h8 : _GEN_5545; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5547 = 10'h246 == _T_107[9:0] ? 4'h7 : _GEN_5546; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5548 = 10'h247 == _T_107[9:0] ? 4'h8 : _GEN_5547; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5549 = 10'h248 == _T_107[9:0] ? 4'ha : _GEN_5548; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5550 = 10'h249 == _T_107[9:0] ? 4'ha : _GEN_5549; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5551 = 10'h24a == _T_107[9:0] ? 4'ha : _GEN_5550; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5552 = 10'h24b == _T_107[9:0] ? 4'h4 : _GEN_5551; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5553 = 10'h24c == _T_107[9:0] ? 4'h4 : _GEN_5552; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5554 = 10'h24d == _T_107[9:0] ? 4'h2 : _GEN_5553; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5555 = 10'h24e == _T_107[9:0] ? 4'h2 : _GEN_5554; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5556 = 10'h24f == _T_107[9:0] ? 4'h2 : _GEN_5555; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5557 = 10'h250 == _T_107[9:0] ? 4'h2 : _GEN_5556; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5558 = 10'h251 == _T_107[9:0] ? 4'h2 : _GEN_5557; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5559 = 10'h252 == _T_107[9:0] ? 4'h2 : _GEN_5558; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5560 = 10'h253 == _T_107[9:0] ? 4'h2 : _GEN_5559; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5561 = 10'h254 == _T_107[9:0] ? 4'h2 : _GEN_5560; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5562 = 10'h255 == _T_107[9:0] ? 4'h3 : _GEN_5561; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5563 = 10'h256 == _T_107[9:0] ? 4'h4 : _GEN_5562; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5564 = 10'h257 == _T_107[9:0] ? 4'h3 : _GEN_5563; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5565 = 10'h258 == _T_107[9:0] ? 4'h4 : _GEN_5564; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5566 = 10'h259 == _T_107[9:0] ? 4'h4 : _GEN_5565; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5567 = 10'h25a == _T_107[9:0] ? 4'h4 : _GEN_5566; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5568 = 10'h25b == _T_107[9:0] ? 4'h3 : _GEN_5567; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5569 = 10'h25c == _T_107[9:0] ? 4'h4 : _GEN_5568; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5570 = 10'h25d == _T_107[9:0] ? 4'h4 : _GEN_5569; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5571 = 10'h25e == _T_107[9:0] ? 4'h3 : _GEN_5570; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5572 = 10'h25f == _T_107[9:0] ? 4'h3 : _GEN_5571; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5573 = 10'h260 == _T_107[9:0] ? 4'h8 : _GEN_5572; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5574 = 10'h261 == _T_107[9:0] ? 4'h7 : _GEN_5573; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5575 = 10'h262 == _T_107[9:0] ? 4'h6 : _GEN_5574; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5576 = 10'h263 == _T_107[9:0] ? 4'h5 : _GEN_5575; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5577 = 10'h264 == _T_107[9:0] ? 4'h6 : _GEN_5576; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5578 = 10'h265 == _T_107[9:0] ? 4'h5 : _GEN_5577; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5579 = 10'h266 == _T_107[9:0] ? 4'h5 : _GEN_5578; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5580 = 10'h267 == _T_107[9:0] ? 4'h7 : _GEN_5579; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5581 = 10'h268 == _T_107[9:0] ? 4'ha : _GEN_5580; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5582 = 10'h269 == _T_107[9:0] ? 4'ha : _GEN_5581; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5583 = 10'h26a == _T_107[9:0] ? 4'ha : _GEN_5582; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5584 = 10'h26b == _T_107[9:0] ? 4'ha : _GEN_5583; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5585 = 10'h26c == _T_107[9:0] ? 4'ha : _GEN_5584; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5586 = 10'h26d == _T_107[9:0] ? 4'ha : _GEN_5585; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5587 = 10'h26e == _T_107[9:0] ? 4'ha : _GEN_5586; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5588 = 10'h26f == _T_107[9:0] ? 4'ha : _GEN_5587; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5589 = 10'h270 == _T_107[9:0] ? 4'h5 : _GEN_5588; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5590 = 10'h271 == _T_107[9:0] ? 4'h4 : _GEN_5589; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5591 = 10'h272 == _T_107[9:0] ? 4'h3 : _GEN_5590; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5592 = 10'h273 == _T_107[9:0] ? 4'h2 : _GEN_5591; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5593 = 10'h274 == _T_107[9:0] ? 4'h2 : _GEN_5592; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5594 = 10'h275 == _T_107[9:0] ? 4'h2 : _GEN_5593; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5595 = 10'h276 == _T_107[9:0] ? 4'h2 : _GEN_5594; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5596 = 10'h277 == _T_107[9:0] ? 4'h2 : _GEN_5595; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5597 = 10'h278 == _T_107[9:0] ? 4'h2 : _GEN_5596; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5598 = 10'h279 == _T_107[9:0] ? 4'h2 : _GEN_5597; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5599 = 10'h27a == _T_107[9:0] ? 4'h2 : _GEN_5598; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5600 = 10'h27b == _T_107[9:0] ? 4'h4 : _GEN_5599; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5601 = 10'h27c == _T_107[9:0] ? 4'h3 : _GEN_5600; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5602 = 10'h27d == _T_107[9:0] ? 4'h4 : _GEN_5601; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5603 = 10'h27e == _T_107[9:0] ? 4'h5 : _GEN_5602; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5604 = 10'h27f == _T_107[9:0] ? 4'h4 : _GEN_5603; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5605 = 10'h280 == _T_107[9:0] ? 4'h4 : _GEN_5604; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5606 = 10'h281 == _T_107[9:0] ? 4'h4 : _GEN_5605; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5607 = 10'h282 == _T_107[9:0] ? 4'h4 : _GEN_5606; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5608 = 10'h283 == _T_107[9:0] ? 4'h3 : _GEN_5607; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5609 = 10'h284 == _T_107[9:0] ? 4'h3 : _GEN_5608; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5610 = 10'h285 == _T_107[9:0] ? 4'h3 : _GEN_5609; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5611 = 10'h286 == _T_107[9:0] ? 4'h8 : _GEN_5610; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5612 = 10'h287 == _T_107[9:0] ? 4'h6 : _GEN_5611; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5613 = 10'h288 == _T_107[9:0] ? 4'h6 : _GEN_5612; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5614 = 10'h289 == _T_107[9:0] ? 4'h6 : _GEN_5613; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5615 = 10'h28a == _T_107[9:0] ? 4'h7 : _GEN_5614; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5616 = 10'h28b == _T_107[9:0] ? 4'h7 : _GEN_5615; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5617 = 10'h28c == _T_107[9:0] ? 4'h6 : _GEN_5616; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5618 = 10'h28d == _T_107[9:0] ? 4'h6 : _GEN_5617; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5619 = 10'h28e == _T_107[9:0] ? 4'h4 : _GEN_5618; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5620 = 10'h28f == _T_107[9:0] ? 4'h7 : _GEN_5619; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5621 = 10'h290 == _T_107[9:0] ? 4'h9 : _GEN_5620; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5622 = 10'h291 == _T_107[9:0] ? 4'ha : _GEN_5621; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5623 = 10'h292 == _T_107[9:0] ? 4'ha : _GEN_5622; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5624 = 10'h293 == _T_107[9:0] ? 4'ha : _GEN_5623; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5625 = 10'h294 == _T_107[9:0] ? 4'h9 : _GEN_5624; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5626 = 10'h295 == _T_107[9:0] ? 4'h5 : _GEN_5625; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5627 = 10'h296 == _T_107[9:0] ? 4'h4 : _GEN_5626; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5628 = 10'h297 == _T_107[9:0] ? 4'h4 : _GEN_5627; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5629 = 10'h298 == _T_107[9:0] ? 4'h3 : _GEN_5628; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5630 = 10'h299 == _T_107[9:0] ? 4'h3 : _GEN_5629; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5631 = 10'h29a == _T_107[9:0] ? 4'h2 : _GEN_5630; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5632 = 10'h29b == _T_107[9:0] ? 4'h2 : _GEN_5631; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5633 = 10'h29c == _T_107[9:0] ? 4'h2 : _GEN_5632; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5634 = 10'h29d == _T_107[9:0] ? 4'h2 : _GEN_5633; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5635 = 10'h29e == _T_107[9:0] ? 4'h2 : _GEN_5634; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5636 = 10'h29f == _T_107[9:0] ? 4'h2 : _GEN_5635; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5637 = 10'h2a0 == _T_107[9:0] ? 4'h2 : _GEN_5636; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5638 = 10'h2a1 == _T_107[9:0] ? 4'h4 : _GEN_5637; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5639 = 10'h2a2 == _T_107[9:0] ? 4'h3 : _GEN_5638; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5640 = 10'h2a3 == _T_107[9:0] ? 4'h4 : _GEN_5639; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5641 = 10'h2a4 == _T_107[9:0] ? 4'h5 : _GEN_5640; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5642 = 10'h2a5 == _T_107[9:0] ? 4'h4 : _GEN_5641; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5643 = 10'h2a6 == _T_107[9:0] ? 4'h4 : _GEN_5642; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5644 = 10'h2a7 == _T_107[9:0] ? 4'h4 : _GEN_5643; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5645 = 10'h2a8 == _T_107[9:0] ? 4'h3 : _GEN_5644; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5646 = 10'h2a9 == _T_107[9:0] ? 4'h3 : _GEN_5645; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5647 = 10'h2aa == _T_107[9:0] ? 4'h3 : _GEN_5646; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5648 = 10'h2ab == _T_107[9:0] ? 4'h3 : _GEN_5647; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5649 = 10'h2ac == _T_107[9:0] ? 4'h8 : _GEN_5648; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5650 = 10'h2ad == _T_107[9:0] ? 4'h7 : _GEN_5649; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5651 = 10'h2ae == _T_107[9:0] ? 4'h5 : _GEN_5650; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5652 = 10'h2af == _T_107[9:0] ? 4'h6 : _GEN_5651; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5653 = 10'h2b0 == _T_107[9:0] ? 4'h7 : _GEN_5652; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5654 = 10'h2b1 == _T_107[9:0] ? 4'h6 : _GEN_5653; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5655 = 10'h2b2 == _T_107[9:0] ? 4'h6 : _GEN_5654; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5656 = 10'h2b3 == _T_107[9:0] ? 4'h6 : _GEN_5655; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5657 = 10'h2b4 == _T_107[9:0] ? 4'h3 : _GEN_5656; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5658 = 10'h2b5 == _T_107[9:0] ? 4'h3 : _GEN_5657; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5659 = 10'h2b6 == _T_107[9:0] ? 4'h3 : _GEN_5658; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5660 = 10'h2b7 == _T_107[9:0] ? 4'h4 : _GEN_5659; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5661 = 10'h2b8 == _T_107[9:0] ? 4'h6 : _GEN_5660; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5662 = 10'h2b9 == _T_107[9:0] ? 4'h9 : _GEN_5661; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5663 = 10'h2ba == _T_107[9:0] ? 4'h4 : _GEN_5662; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5664 = 10'h2bb == _T_107[9:0] ? 4'h3 : _GEN_5663; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5665 = 10'h2bc == _T_107[9:0] ? 4'h4 : _GEN_5664; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5666 = 10'h2bd == _T_107[9:0] ? 4'h3 : _GEN_5665; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5667 = 10'h2be == _T_107[9:0] ? 4'h3 : _GEN_5666; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5668 = 10'h2bf == _T_107[9:0] ? 4'h3 : _GEN_5667; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5669 = 10'h2c0 == _T_107[9:0] ? 4'h2 : _GEN_5668; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5670 = 10'h2c1 == _T_107[9:0] ? 4'h2 : _GEN_5669; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5671 = 10'h2c2 == _T_107[9:0] ? 4'h2 : _GEN_5670; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5672 = 10'h2c3 == _T_107[9:0] ? 4'h2 : _GEN_5671; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5673 = 10'h2c4 == _T_107[9:0] ? 4'h2 : _GEN_5672; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5674 = 10'h2c5 == _T_107[9:0] ? 4'h2 : _GEN_5673; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5675 = 10'h2c6 == _T_107[9:0] ? 4'h2 : _GEN_5674; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5676 = 10'h2c7 == _T_107[9:0] ? 4'h4 : _GEN_5675; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5677 = 10'h2c8 == _T_107[9:0] ? 4'h3 : _GEN_5676; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5678 = 10'h2c9 == _T_107[9:0] ? 4'h4 : _GEN_5677; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5679 = 10'h2ca == _T_107[9:0] ? 4'h5 : _GEN_5678; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5680 = 10'h2cb == _T_107[9:0] ? 4'h3 : _GEN_5679; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5681 = 10'h2cc == _T_107[9:0] ? 4'h3 : _GEN_5680; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5682 = 10'h2cd == _T_107[9:0] ? 4'h3 : _GEN_5681; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5683 = 10'h2ce == _T_107[9:0] ? 4'h3 : _GEN_5682; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5684 = 10'h2cf == _T_107[9:0] ? 4'h3 : _GEN_5683; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5685 = 10'h2d0 == _T_107[9:0] ? 4'h3 : _GEN_5684; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5686 = 10'h2d1 == _T_107[9:0] ? 4'h3 : _GEN_5685; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5687 = 10'h2d2 == _T_107[9:0] ? 4'h8 : _GEN_5686; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5688 = 10'h2d3 == _T_107[9:0] ? 4'h6 : _GEN_5687; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5689 = 10'h2d4 == _T_107[9:0] ? 4'h6 : _GEN_5688; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5690 = 10'h2d5 == _T_107[9:0] ? 4'h7 : _GEN_5689; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5691 = 10'h2d6 == _T_107[9:0] ? 4'h7 : _GEN_5690; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5692 = 10'h2d7 == _T_107[9:0] ? 4'h7 : _GEN_5691; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5693 = 10'h2d8 == _T_107[9:0] ? 4'h6 : _GEN_5692; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5694 = 10'h2d9 == _T_107[9:0] ? 4'h7 : _GEN_5693; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5695 = 10'h2da == _T_107[9:0] ? 4'h5 : _GEN_5694; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5696 = 10'h2db == _T_107[9:0] ? 4'h3 : _GEN_5695; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5697 = 10'h2dc == _T_107[9:0] ? 4'h3 : _GEN_5696; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5698 = 10'h2dd == _T_107[9:0] ? 4'h3 : _GEN_5697; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5699 = 10'h2de == _T_107[9:0] ? 4'h3 : _GEN_5698; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5700 = 10'h2df == _T_107[9:0] ? 4'h4 : _GEN_5699; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5701 = 10'h2e0 == _T_107[9:0] ? 4'h3 : _GEN_5700; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5702 = 10'h2e1 == _T_107[9:0] ? 4'h3 : _GEN_5701; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5703 = 10'h2e2 == _T_107[9:0] ? 4'h3 : _GEN_5702; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5704 = 10'h2e3 == _T_107[9:0] ? 4'h3 : _GEN_5703; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5705 = 10'h2e4 == _T_107[9:0] ? 4'h3 : _GEN_5704; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5706 = 10'h2e5 == _T_107[9:0] ? 4'h3 : _GEN_5705; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5707 = 10'h2e6 == _T_107[9:0] ? 4'h2 : _GEN_5706; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5708 = 10'h2e7 == _T_107[9:0] ? 4'h2 : _GEN_5707; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5709 = 10'h2e8 == _T_107[9:0] ? 4'h2 : _GEN_5708; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5710 = 10'h2e9 == _T_107[9:0] ? 4'h2 : _GEN_5709; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5711 = 10'h2ea == _T_107[9:0] ? 4'h2 : _GEN_5710; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5712 = 10'h2eb == _T_107[9:0] ? 4'h2 : _GEN_5711; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5713 = 10'h2ec == _T_107[9:0] ? 4'h3 : _GEN_5712; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5714 = 10'h2ed == _T_107[9:0] ? 4'h4 : _GEN_5713; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5715 = 10'h2ee == _T_107[9:0] ? 4'h3 : _GEN_5714; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5716 = 10'h2ef == _T_107[9:0] ? 4'h3 : _GEN_5715; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5717 = 10'h2f0 == _T_107[9:0] ? 4'h6 : _GEN_5716; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5718 = 10'h2f1 == _T_107[9:0] ? 4'h3 : _GEN_5717; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5719 = 10'h2f2 == _T_107[9:0] ? 4'h3 : _GEN_5718; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5720 = 10'h2f3 == _T_107[9:0] ? 4'h3 : _GEN_5719; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5721 = 10'h2f4 == _T_107[9:0] ? 4'h3 : _GEN_5720; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5722 = 10'h2f5 == _T_107[9:0] ? 4'h3 : _GEN_5721; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5723 = 10'h2f6 == _T_107[9:0] ? 4'h3 : _GEN_5722; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5724 = 10'h2f7 == _T_107[9:0] ? 4'h3 : _GEN_5723; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5725 = 10'h2f8 == _T_107[9:0] ? 4'h8 : _GEN_5724; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5726 = 10'h2f9 == _T_107[9:0] ? 4'h6 : _GEN_5725; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5727 = 10'h2fa == _T_107[9:0] ? 4'h7 : _GEN_5726; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5728 = 10'h2fb == _T_107[9:0] ? 4'h7 : _GEN_5727; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5729 = 10'h2fc == _T_107[9:0] ? 4'h6 : _GEN_5728; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5730 = 10'h2fd == _T_107[9:0] ? 4'h6 : _GEN_5729; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5731 = 10'h2fe == _T_107[9:0] ? 4'h6 : _GEN_5730; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5732 = 10'h2ff == _T_107[9:0] ? 4'h8 : _GEN_5731; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5733 = 10'h300 == _T_107[9:0] ? 4'h9 : _GEN_5732; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5734 = 10'h301 == _T_107[9:0] ? 4'h7 : _GEN_5733; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5735 = 10'h302 == _T_107[9:0] ? 4'h4 : _GEN_5734; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5736 = 10'h303 == _T_107[9:0] ? 4'h4 : _GEN_5735; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5737 = 10'h304 == _T_107[9:0] ? 4'h3 : _GEN_5736; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5738 = 10'h305 == _T_107[9:0] ? 4'h3 : _GEN_5737; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5739 = 10'h306 == _T_107[9:0] ? 4'h3 : _GEN_5738; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5740 = 10'h307 == _T_107[9:0] ? 4'h3 : _GEN_5739; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5741 = 10'h308 == _T_107[9:0] ? 4'h3 : _GEN_5740; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5742 = 10'h309 == _T_107[9:0] ? 4'h3 : _GEN_5741; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5743 = 10'h30a == _T_107[9:0] ? 4'h3 : _GEN_5742; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5744 = 10'h30b == _T_107[9:0] ? 4'h3 : _GEN_5743; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5745 = 10'h30c == _T_107[9:0] ? 4'h2 : _GEN_5744; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5746 = 10'h30d == _T_107[9:0] ? 4'h2 : _GEN_5745; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5747 = 10'h30e == _T_107[9:0] ? 4'h2 : _GEN_5746; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5748 = 10'h30f == _T_107[9:0] ? 4'h2 : _GEN_5747; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5749 = 10'h310 == _T_107[9:0] ? 4'h2 : _GEN_5748; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5750 = 10'h311 == _T_107[9:0] ? 4'h2 : _GEN_5749; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5751 = 10'h312 == _T_107[9:0] ? 4'h3 : _GEN_5750; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5752 = 10'h313 == _T_107[9:0] ? 4'h4 : _GEN_5751; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5753 = 10'h314 == _T_107[9:0] ? 4'h3 : _GEN_5752; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5754 = 10'h315 == _T_107[9:0] ? 4'h3 : _GEN_5753; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5755 = 10'h316 == _T_107[9:0] ? 4'h5 : _GEN_5754; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5756 = 10'h317 == _T_107[9:0] ? 4'h5 : _GEN_5755; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5757 = 10'h318 == _T_107[9:0] ? 4'h3 : _GEN_5756; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5758 = 10'h319 == _T_107[9:0] ? 4'h3 : _GEN_5757; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5759 = 10'h31a == _T_107[9:0] ? 4'h3 : _GEN_5758; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5760 = 10'h31b == _T_107[9:0] ? 4'h3 : _GEN_5759; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5761 = 10'h31c == _T_107[9:0] ? 4'h3 : _GEN_5760; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5762 = 10'h31d == _T_107[9:0] ? 4'h3 : _GEN_5761; // @[Filter.scala 230:62]
  wire [4:0] _GEN_38966 = {{1'd0}, _GEN_5762}; // @[Filter.scala 230:62]
  wire [8:0] _T_109 = _GEN_38966 * 5'h14; // @[Filter.scala 230:62]
  wire [3:0] _GEN_5786 = 10'h17 == _T_107[9:0] ? 4'hb : 4'he; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5787 = 10'h18 == _T_107[9:0] ? 4'hc : _GEN_5786; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5788 = 10'h19 == _T_107[9:0] ? 4'he : _GEN_5787; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5789 = 10'h1a == _T_107[9:0] ? 4'he : _GEN_5788; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5790 = 10'h1b == _T_107[9:0] ? 4'he : _GEN_5789; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5791 = 10'h1c == _T_107[9:0] ? 4'he : _GEN_5790; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5792 = 10'h1d == _T_107[9:0] ? 4'he : _GEN_5791; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5793 = 10'h1e == _T_107[9:0] ? 4'he : _GEN_5792; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5794 = 10'h1f == _T_107[9:0] ? 4'he : _GEN_5793; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5795 = 10'h20 == _T_107[9:0] ? 4'he : _GEN_5794; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5796 = 10'h21 == _T_107[9:0] ? 4'he : _GEN_5795; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5797 = 10'h22 == _T_107[9:0] ? 4'he : _GEN_5796; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5798 = 10'h23 == _T_107[9:0] ? 4'he : _GEN_5797; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5799 = 10'h24 == _T_107[9:0] ? 4'he : _GEN_5798; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5800 = 10'h25 == _T_107[9:0] ? 4'he : _GEN_5799; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5801 = 10'h26 == _T_107[9:0] ? 4'he : _GEN_5800; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5802 = 10'h27 == _T_107[9:0] ? 4'he : _GEN_5801; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5803 = 10'h28 == _T_107[9:0] ? 4'he : _GEN_5802; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5804 = 10'h29 == _T_107[9:0] ? 4'he : _GEN_5803; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5805 = 10'h2a == _T_107[9:0] ? 4'he : _GEN_5804; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5806 = 10'h2b == _T_107[9:0] ? 4'he : _GEN_5805; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5807 = 10'h2c == _T_107[9:0] ? 4'he : _GEN_5806; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5808 = 10'h2d == _T_107[9:0] ? 4'he : _GEN_5807; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5809 = 10'h2e == _T_107[9:0] ? 4'he : _GEN_5808; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5810 = 10'h2f == _T_107[9:0] ? 4'he : _GEN_5809; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5811 = 10'h30 == _T_107[9:0] ? 4'he : _GEN_5810; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5812 = 10'h31 == _T_107[9:0] ? 4'he : _GEN_5811; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5813 = 10'h32 == _T_107[9:0] ? 4'he : _GEN_5812; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5814 = 10'h33 == _T_107[9:0] ? 4'he : _GEN_5813; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5815 = 10'h34 == _T_107[9:0] ? 4'he : _GEN_5814; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5816 = 10'h35 == _T_107[9:0] ? 4'he : _GEN_5815; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5817 = 10'h36 == _T_107[9:0] ? 4'he : _GEN_5816; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5818 = 10'h37 == _T_107[9:0] ? 4'he : _GEN_5817; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5819 = 10'h38 == _T_107[9:0] ? 4'he : _GEN_5818; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5820 = 10'h39 == _T_107[9:0] ? 4'he : _GEN_5819; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5821 = 10'h3a == _T_107[9:0] ? 4'he : _GEN_5820; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5822 = 10'h3b == _T_107[9:0] ? 4'he : _GEN_5821; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5823 = 10'h3c == _T_107[9:0] ? 4'ha : _GEN_5822; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5824 = 10'h3d == _T_107[9:0] ? 4'hc : _GEN_5823; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5825 = 10'h3e == _T_107[9:0] ? 4'hb : _GEN_5824; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5826 = 10'h3f == _T_107[9:0] ? 4'he : _GEN_5825; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5827 = 10'h40 == _T_107[9:0] ? 4'he : _GEN_5826; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5828 = 10'h41 == _T_107[9:0] ? 4'he : _GEN_5827; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5829 = 10'h42 == _T_107[9:0] ? 4'he : _GEN_5828; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5830 = 10'h43 == _T_107[9:0] ? 4'he : _GEN_5829; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5831 = 10'h44 == _T_107[9:0] ? 4'he : _GEN_5830; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5832 = 10'h45 == _T_107[9:0] ? 4'he : _GEN_5831; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5833 = 10'h46 == _T_107[9:0] ? 4'he : _GEN_5832; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5834 = 10'h47 == _T_107[9:0] ? 4'he : _GEN_5833; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5835 = 10'h48 == _T_107[9:0] ? 4'he : _GEN_5834; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5836 = 10'h49 == _T_107[9:0] ? 4'he : _GEN_5835; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5837 = 10'h4a == _T_107[9:0] ? 4'he : _GEN_5836; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5838 = 10'h4b == _T_107[9:0] ? 4'he : _GEN_5837; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5839 = 10'h4c == _T_107[9:0] ? 4'he : _GEN_5838; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5840 = 10'h4d == _T_107[9:0] ? 4'he : _GEN_5839; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5841 = 10'h4e == _T_107[9:0] ? 4'he : _GEN_5840; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5842 = 10'h4f == _T_107[9:0] ? 4'he : _GEN_5841; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5843 = 10'h50 == _T_107[9:0] ? 4'he : _GEN_5842; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5844 = 10'h51 == _T_107[9:0] ? 4'he : _GEN_5843; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5845 = 10'h52 == _T_107[9:0] ? 4'he : _GEN_5844; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5846 = 10'h53 == _T_107[9:0] ? 4'he : _GEN_5845; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5847 = 10'h54 == _T_107[9:0] ? 4'he : _GEN_5846; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5848 = 10'h55 == _T_107[9:0] ? 4'he : _GEN_5847; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5849 = 10'h56 == _T_107[9:0] ? 4'he : _GEN_5848; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5850 = 10'h57 == _T_107[9:0] ? 4'he : _GEN_5849; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5851 = 10'h58 == _T_107[9:0] ? 4'he : _GEN_5850; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5852 = 10'h59 == _T_107[9:0] ? 4'he : _GEN_5851; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5853 = 10'h5a == _T_107[9:0] ? 4'hc : _GEN_5852; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5854 = 10'h5b == _T_107[9:0] ? 4'hd : _GEN_5853; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5855 = 10'h5c == _T_107[9:0] ? 4'he : _GEN_5854; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5856 = 10'h5d == _T_107[9:0] ? 4'he : _GEN_5855; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5857 = 10'h5e == _T_107[9:0] ? 4'he : _GEN_5856; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5858 = 10'h5f == _T_107[9:0] ? 4'he : _GEN_5857; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5859 = 10'h60 == _T_107[9:0] ? 4'he : _GEN_5858; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5860 = 10'h61 == _T_107[9:0] ? 4'hd : _GEN_5859; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5861 = 10'h62 == _T_107[9:0] ? 4'hb : _GEN_5860; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5862 = 10'h63 == _T_107[9:0] ? 4'hc : _GEN_5861; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5863 = 10'h64 == _T_107[9:0] ? 4'ha : _GEN_5862; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5864 = 10'h65 == _T_107[9:0] ? 4'hd : _GEN_5863; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5865 = 10'h66 == _T_107[9:0] ? 4'he : _GEN_5864; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5866 = 10'h67 == _T_107[9:0] ? 4'he : _GEN_5865; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5867 = 10'h68 == _T_107[9:0] ? 4'he : _GEN_5866; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5868 = 10'h69 == _T_107[9:0] ? 4'he : _GEN_5867; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5869 = 10'h6a == _T_107[9:0] ? 4'he : _GEN_5868; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5870 = 10'h6b == _T_107[9:0] ? 4'hd : _GEN_5869; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5871 = 10'h6c == _T_107[9:0] ? 4'hc : _GEN_5870; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5872 = 10'h6d == _T_107[9:0] ? 4'hc : _GEN_5871; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5873 = 10'h6e == _T_107[9:0] ? 4'he : _GEN_5872; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5874 = 10'h6f == _T_107[9:0] ? 4'he : _GEN_5873; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5875 = 10'h70 == _T_107[9:0] ? 4'he : _GEN_5874; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5876 = 10'h71 == _T_107[9:0] ? 4'he : _GEN_5875; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5877 = 10'h72 == _T_107[9:0] ? 4'he : _GEN_5876; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5878 = 10'h73 == _T_107[9:0] ? 4'he : _GEN_5877; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5879 = 10'h74 == _T_107[9:0] ? 4'he : _GEN_5878; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5880 = 10'h75 == _T_107[9:0] ? 4'he : _GEN_5879; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5881 = 10'h76 == _T_107[9:0] ? 4'he : _GEN_5880; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5882 = 10'h77 == _T_107[9:0] ? 4'he : _GEN_5881; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5883 = 10'h78 == _T_107[9:0] ? 4'he : _GEN_5882; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5884 = 10'h79 == _T_107[9:0] ? 4'he : _GEN_5883; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5885 = 10'h7a == _T_107[9:0] ? 4'he : _GEN_5884; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5886 = 10'h7b == _T_107[9:0] ? 4'he : _GEN_5885; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5887 = 10'h7c == _T_107[9:0] ? 4'he : _GEN_5886; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5888 = 10'h7d == _T_107[9:0] ? 4'he : _GEN_5887; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5889 = 10'h7e == _T_107[9:0] ? 4'he : _GEN_5888; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5890 = 10'h7f == _T_107[9:0] ? 4'he : _GEN_5889; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5891 = 10'h80 == _T_107[9:0] ? 4'he : _GEN_5890; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5892 = 10'h81 == _T_107[9:0] ? 4'hb : _GEN_5891; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5893 = 10'h82 == _T_107[9:0] ? 4'hc : _GEN_5892; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5894 = 10'h83 == _T_107[9:0] ? 4'hc : _GEN_5893; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5895 = 10'h84 == _T_107[9:0] ? 4'he : _GEN_5894; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5896 = 10'h85 == _T_107[9:0] ? 4'he : _GEN_5895; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5897 = 10'h86 == _T_107[9:0] ? 4'he : _GEN_5896; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5898 = 10'h87 == _T_107[9:0] ? 4'ha : _GEN_5897; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5899 = 10'h88 == _T_107[9:0] ? 4'hd : _GEN_5898; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5900 = 10'h89 == _T_107[9:0] ? 4'hd : _GEN_5899; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5901 = 10'h8a == _T_107[9:0] ? 4'hc : _GEN_5900; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5902 = 10'h8b == _T_107[9:0] ? 4'he : _GEN_5901; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5903 = 10'h8c == _T_107[9:0] ? 4'he : _GEN_5902; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5904 = 10'h8d == _T_107[9:0] ? 4'he : _GEN_5903; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5905 = 10'h8e == _T_107[9:0] ? 4'he : _GEN_5904; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5906 = 10'h8f == _T_107[9:0] ? 4'hb : _GEN_5905; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5907 = 10'h90 == _T_107[9:0] ? 4'hc : _GEN_5906; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5908 = 10'h91 == _T_107[9:0] ? 4'hc : _GEN_5907; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5909 = 10'h92 == _T_107[9:0] ? 4'hd : _GEN_5908; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5910 = 10'h93 == _T_107[9:0] ? 4'he : _GEN_5909; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5911 = 10'h94 == _T_107[9:0] ? 4'he : _GEN_5910; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5912 = 10'h95 == _T_107[9:0] ? 4'he : _GEN_5911; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5913 = 10'h96 == _T_107[9:0] ? 4'he : _GEN_5912; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5914 = 10'h97 == _T_107[9:0] ? 4'he : _GEN_5913; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5915 = 10'h98 == _T_107[9:0] ? 4'he : _GEN_5914; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5916 = 10'h99 == _T_107[9:0] ? 4'he : _GEN_5915; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5917 = 10'h9a == _T_107[9:0] ? 4'he : _GEN_5916; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5918 = 10'h9b == _T_107[9:0] ? 4'he : _GEN_5917; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5919 = 10'h9c == _T_107[9:0] ? 4'he : _GEN_5918; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5920 = 10'h9d == _T_107[9:0] ? 4'he : _GEN_5919; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5921 = 10'h9e == _T_107[9:0] ? 4'he : _GEN_5920; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5922 = 10'h9f == _T_107[9:0] ? 4'he : _GEN_5921; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5923 = 10'ha0 == _T_107[9:0] ? 4'he : _GEN_5922; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5924 = 10'ha1 == _T_107[9:0] ? 4'he : _GEN_5923; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5925 = 10'ha2 == _T_107[9:0] ? 4'he : _GEN_5924; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5926 = 10'ha3 == _T_107[9:0] ? 4'he : _GEN_5925; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5927 = 10'ha4 == _T_107[9:0] ? 4'he : _GEN_5926; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5928 = 10'ha5 == _T_107[9:0] ? 4'he : _GEN_5927; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5929 = 10'ha6 == _T_107[9:0] ? 4'he : _GEN_5928; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5930 = 10'ha7 == _T_107[9:0] ? 4'he : _GEN_5929; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5931 = 10'ha8 == _T_107[9:0] ? 4'hb : _GEN_5930; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5932 = 10'ha9 == _T_107[9:0] ? 4'hc : _GEN_5931; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5933 = 10'haa == _T_107[9:0] ? 4'hb : _GEN_5932; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5934 = 10'hab == _T_107[9:0] ? 4'hc : _GEN_5933; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5935 = 10'hac == _T_107[9:0] ? 4'hd : _GEN_5934; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5936 = 10'had == _T_107[9:0] ? 4'ha : _GEN_5935; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5937 = 10'hae == _T_107[9:0] ? 4'hd : _GEN_5936; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5938 = 10'haf == _T_107[9:0] ? 4'hd : _GEN_5937; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5939 = 10'hb0 == _T_107[9:0] ? 4'hb : _GEN_5938; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5940 = 10'hb1 == _T_107[9:0] ? 4'hc : _GEN_5939; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5941 = 10'hb2 == _T_107[9:0] ? 4'he : _GEN_5940; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5942 = 10'hb3 == _T_107[9:0] ? 4'hb : _GEN_5941; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5943 = 10'hb4 == _T_107[9:0] ? 4'hc : _GEN_5942; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5944 = 10'hb5 == _T_107[9:0] ? 4'hd : _GEN_5943; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5945 = 10'hb6 == _T_107[9:0] ? 4'hd : _GEN_5944; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5946 = 10'hb7 == _T_107[9:0] ? 4'hc : _GEN_5945; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5947 = 10'hb8 == _T_107[9:0] ? 4'he : _GEN_5946; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5948 = 10'hb9 == _T_107[9:0] ? 4'he : _GEN_5947; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5949 = 10'hba == _T_107[9:0] ? 4'he : _GEN_5948; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5950 = 10'hbb == _T_107[9:0] ? 4'he : _GEN_5949; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5951 = 10'hbc == _T_107[9:0] ? 4'he : _GEN_5950; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5952 = 10'hbd == _T_107[9:0] ? 4'he : _GEN_5951; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5953 = 10'hbe == _T_107[9:0] ? 4'he : _GEN_5952; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5954 = 10'hbf == _T_107[9:0] ? 4'he : _GEN_5953; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5955 = 10'hc0 == _T_107[9:0] ? 4'he : _GEN_5954; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5956 = 10'hc1 == _T_107[9:0] ? 4'he : _GEN_5955; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5957 = 10'hc2 == _T_107[9:0] ? 4'he : _GEN_5956; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5958 = 10'hc3 == _T_107[9:0] ? 4'he : _GEN_5957; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5959 = 10'hc4 == _T_107[9:0] ? 4'he : _GEN_5958; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5960 = 10'hc5 == _T_107[9:0] ? 4'he : _GEN_5959; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5961 = 10'hc6 == _T_107[9:0] ? 4'he : _GEN_5960; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5962 = 10'hc7 == _T_107[9:0] ? 4'hd : _GEN_5961; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5963 = 10'hc8 == _T_107[9:0] ? 4'hb : _GEN_5962; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5964 = 10'hc9 == _T_107[9:0] ? 4'hc : _GEN_5963; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5965 = 10'hca == _T_107[9:0] ? 4'he : _GEN_5964; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5966 = 10'hcb == _T_107[9:0] ? 4'he : _GEN_5965; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5967 = 10'hcc == _T_107[9:0] ? 4'he : _GEN_5966; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5968 = 10'hcd == _T_107[9:0] ? 4'he : _GEN_5967; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5969 = 10'hce == _T_107[9:0] ? 4'hd : _GEN_5968; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5970 = 10'hcf == _T_107[9:0] ? 4'hb : _GEN_5969; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5971 = 10'hd0 == _T_107[9:0] ? 4'hc : _GEN_5970; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5972 = 10'hd1 == _T_107[9:0] ? 4'hc : _GEN_5971; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5973 = 10'hd2 == _T_107[9:0] ? 4'hb : _GEN_5972; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5974 = 10'hd3 == _T_107[9:0] ? 4'hd : _GEN_5973; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5975 = 10'hd4 == _T_107[9:0] ? 4'hd : _GEN_5974; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5976 = 10'hd5 == _T_107[9:0] ? 4'hd : _GEN_5975; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5977 = 10'hd6 == _T_107[9:0] ? 4'hd : _GEN_5976; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5978 = 10'hd7 == _T_107[9:0] ? 4'hc : _GEN_5977; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5979 = 10'hd8 == _T_107[9:0] ? 4'hc : _GEN_5978; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5980 = 10'hd9 == _T_107[9:0] ? 4'hc : _GEN_5979; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5981 = 10'hda == _T_107[9:0] ? 4'hd : _GEN_5980; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5982 = 10'hdb == _T_107[9:0] ? 4'hc : _GEN_5981; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5983 = 10'hdc == _T_107[9:0] ? 4'h9 : _GEN_5982; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5984 = 10'hdd == _T_107[9:0] ? 4'he : _GEN_5983; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5985 = 10'hde == _T_107[9:0] ? 4'he : _GEN_5984; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5986 = 10'hdf == _T_107[9:0] ? 4'he : _GEN_5985; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5987 = 10'he0 == _T_107[9:0] ? 4'he : _GEN_5986; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5988 = 10'he1 == _T_107[9:0] ? 4'he : _GEN_5987; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5989 = 10'he2 == _T_107[9:0] ? 4'he : _GEN_5988; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5990 = 10'he3 == _T_107[9:0] ? 4'h9 : _GEN_5989; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5991 = 10'he4 == _T_107[9:0] ? 4'he : _GEN_5990; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5992 = 10'he5 == _T_107[9:0] ? 4'he : _GEN_5991; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5993 = 10'he6 == _T_107[9:0] ? 4'he : _GEN_5992; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5994 = 10'he7 == _T_107[9:0] ? 4'he : _GEN_5993; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5995 = 10'he8 == _T_107[9:0] ? 4'he : _GEN_5994; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5996 = 10'he9 == _T_107[9:0] ? 4'he : _GEN_5995; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5997 = 10'hea == _T_107[9:0] ? 4'he : _GEN_5996; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5998 = 10'heb == _T_107[9:0] ? 4'hc : _GEN_5997; // @[Filter.scala 230:102]
  wire [3:0] _GEN_5999 = 10'hec == _T_107[9:0] ? 4'h7 : _GEN_5998; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6000 = 10'hed == _T_107[9:0] ? 4'h1 : _GEN_5999; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6001 = 10'hee == _T_107[9:0] ? 4'h0 : _GEN_6000; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6002 = 10'hef == _T_107[9:0] ? 4'h0 : _GEN_6001; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6003 = 10'hf0 == _T_107[9:0] ? 4'h2 : _GEN_6002; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6004 = 10'hf1 == _T_107[9:0] ? 4'h9 : _GEN_6003; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6005 = 10'hf2 == _T_107[9:0] ? 4'he : _GEN_6004; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6006 = 10'hf3 == _T_107[9:0] ? 4'he : _GEN_6005; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6007 = 10'hf4 == _T_107[9:0] ? 4'he : _GEN_6006; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6008 = 10'hf5 == _T_107[9:0] ? 4'hc : _GEN_6007; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6009 = 10'hf6 == _T_107[9:0] ? 4'hc : _GEN_6008; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6010 = 10'hf7 == _T_107[9:0] ? 4'hd : _GEN_6009; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6011 = 10'hf8 == _T_107[9:0] ? 4'hd : _GEN_6010; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6012 = 10'hf9 == _T_107[9:0] ? 4'hd : _GEN_6011; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6013 = 10'hfa == _T_107[9:0] ? 4'hd : _GEN_6012; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6014 = 10'hfb == _T_107[9:0] ? 4'hd : _GEN_6013; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6015 = 10'hfc == _T_107[9:0] ? 4'hd : _GEN_6014; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6016 = 10'hfd == _T_107[9:0] ? 4'hd : _GEN_6015; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6017 = 10'hfe == _T_107[9:0] ? 4'hd : _GEN_6016; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6018 = 10'hff == _T_107[9:0] ? 4'hd : _GEN_6017; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6019 = 10'h100 == _T_107[9:0] ? 4'hd : _GEN_6018; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6020 = 10'h101 == _T_107[9:0] ? 4'h9 : _GEN_6019; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6021 = 10'h102 == _T_107[9:0] ? 4'h9 : _GEN_6020; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6022 = 10'h103 == _T_107[9:0] ? 4'he : _GEN_6021; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6023 = 10'h104 == _T_107[9:0] ? 4'he : _GEN_6022; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6024 = 10'h105 == _T_107[9:0] ? 4'he : _GEN_6023; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6025 = 10'h106 == _T_107[9:0] ? 4'he : _GEN_6024; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6026 = 10'h107 == _T_107[9:0] ? 4'he : _GEN_6025; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6027 = 10'h108 == _T_107[9:0] ? 4'he : _GEN_6026; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6028 = 10'h109 == _T_107[9:0] ? 4'h6 : _GEN_6027; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6029 = 10'h10a == _T_107[9:0] ? 4'he : _GEN_6028; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6030 = 10'h10b == _T_107[9:0] ? 4'he : _GEN_6029; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6031 = 10'h10c == _T_107[9:0] ? 4'he : _GEN_6030; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6032 = 10'h10d == _T_107[9:0] ? 4'he : _GEN_6031; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6033 = 10'h10e == _T_107[9:0] ? 4'he : _GEN_6032; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6034 = 10'h10f == _T_107[9:0] ? 4'ha : _GEN_6033; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6035 = 10'h110 == _T_107[9:0] ? 4'hd : _GEN_6034; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6036 = 10'h111 == _T_107[9:0] ? 4'h4 : _GEN_6035; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6037 = 10'h112 == _T_107[9:0] ? 4'h7 : _GEN_6036; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6038 = 10'h113 == _T_107[9:0] ? 4'h0 : _GEN_6037; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6039 = 10'h114 == _T_107[9:0] ? 4'h0 : _GEN_6038; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6040 = 10'h115 == _T_107[9:0] ? 4'h0 : _GEN_6039; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6041 = 10'h116 == _T_107[9:0] ? 4'h0 : _GEN_6040; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6042 = 10'h117 == _T_107[9:0] ? 4'h0 : _GEN_6041; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6043 = 10'h118 == _T_107[9:0] ? 4'ha : _GEN_6042; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6044 = 10'h119 == _T_107[9:0] ? 4'he : _GEN_6043; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6045 = 10'h11a == _T_107[9:0] ? 4'he : _GEN_6044; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6046 = 10'h11b == _T_107[9:0] ? 4'he : _GEN_6045; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6047 = 10'h11c == _T_107[9:0] ? 4'hb : _GEN_6046; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6048 = 10'h11d == _T_107[9:0] ? 4'hc : _GEN_6047; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6049 = 10'h11e == _T_107[9:0] ? 4'hd : _GEN_6048; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6050 = 10'h11f == _T_107[9:0] ? 4'hb : _GEN_6049; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6051 = 10'h120 == _T_107[9:0] ? 4'ha : _GEN_6050; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6052 = 10'h121 == _T_107[9:0] ? 4'hc : _GEN_6051; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6053 = 10'h122 == _T_107[9:0] ? 4'ha : _GEN_6052; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6054 = 10'h123 == _T_107[9:0] ? 4'ha : _GEN_6053; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6055 = 10'h124 == _T_107[9:0] ? 4'hd : _GEN_6054; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6056 = 10'h125 == _T_107[9:0] ? 4'hd : _GEN_6055; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6057 = 10'h126 == _T_107[9:0] ? 4'hb : _GEN_6056; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6058 = 10'h127 == _T_107[9:0] ? 4'h9 : _GEN_6057; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6059 = 10'h128 == _T_107[9:0] ? 4'h7 : _GEN_6058; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6060 = 10'h129 == _T_107[9:0] ? 4'hd : _GEN_6059; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6061 = 10'h12a == _T_107[9:0] ? 4'hc : _GEN_6060; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6062 = 10'h12b == _T_107[9:0] ? 4'hb : _GEN_6061; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6063 = 10'h12c == _T_107[9:0] ? 4'hc : _GEN_6062; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6064 = 10'h12d == _T_107[9:0] ? 4'hb : _GEN_6063; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6065 = 10'h12e == _T_107[9:0] ? 4'ha : _GEN_6064; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6066 = 10'h12f == _T_107[9:0] ? 4'h6 : _GEN_6065; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6067 = 10'h130 == _T_107[9:0] ? 4'he : _GEN_6066; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6068 = 10'h131 == _T_107[9:0] ? 4'hc : _GEN_6067; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6069 = 10'h132 == _T_107[9:0] ? 4'ha : _GEN_6068; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6070 = 10'h133 == _T_107[9:0] ? 4'h9 : _GEN_6069; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6071 = 10'h134 == _T_107[9:0] ? 4'hb : _GEN_6070; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6072 = 10'h135 == _T_107[9:0] ? 4'h8 : _GEN_6071; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6073 = 10'h136 == _T_107[9:0] ? 4'h8 : _GEN_6072; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6074 = 10'h137 == _T_107[9:0] ? 4'h4 : _GEN_6073; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6075 = 10'h138 == _T_107[9:0] ? 4'h7 : _GEN_6074; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6076 = 10'h139 == _T_107[9:0] ? 4'h0 : _GEN_6075; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6077 = 10'h13a == _T_107[9:0] ? 4'h0 : _GEN_6076; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6078 = 10'h13b == _T_107[9:0] ? 4'h0 : _GEN_6077; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6079 = 10'h13c == _T_107[9:0] ? 4'h0 : _GEN_6078; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6080 = 10'h13d == _T_107[9:0] ? 4'h0 : _GEN_6079; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6081 = 10'h13e == _T_107[9:0] ? 4'h4 : _GEN_6080; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6082 = 10'h13f == _T_107[9:0] ? 4'hc : _GEN_6081; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6083 = 10'h140 == _T_107[9:0] ? 4'he : _GEN_6082; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6084 = 10'h141 == _T_107[9:0] ? 4'he : _GEN_6083; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6085 = 10'h142 == _T_107[9:0] ? 4'he : _GEN_6084; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6086 = 10'h143 == _T_107[9:0] ? 4'hc : _GEN_6085; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6087 = 10'h144 == _T_107[9:0] ? 4'hd : _GEN_6086; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6088 = 10'h145 == _T_107[9:0] ? 4'hb : _GEN_6087; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6089 = 10'h146 == _T_107[9:0] ? 4'hb : _GEN_6088; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6090 = 10'h147 == _T_107[9:0] ? 4'ha : _GEN_6089; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6091 = 10'h148 == _T_107[9:0] ? 4'ha : _GEN_6090; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6092 = 10'h149 == _T_107[9:0] ? 4'hc : _GEN_6091; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6093 = 10'h14a == _T_107[9:0] ? 4'hd : _GEN_6092; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6094 = 10'h14b == _T_107[9:0] ? 4'hc : _GEN_6093; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6095 = 10'h14c == _T_107[9:0] ? 4'hd : _GEN_6094; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6096 = 10'h14d == _T_107[9:0] ? 4'h9 : _GEN_6095; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6097 = 10'h14e == _T_107[9:0] ? 4'h7 : _GEN_6096; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6098 = 10'h14f == _T_107[9:0] ? 4'ha : _GEN_6097; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6099 = 10'h150 == _T_107[9:0] ? 4'ha : _GEN_6098; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6100 = 10'h151 == _T_107[9:0] ? 4'hb : _GEN_6099; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6101 = 10'h152 == _T_107[9:0] ? 4'hb : _GEN_6100; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6102 = 10'h153 == _T_107[9:0] ? 4'hc : _GEN_6101; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6103 = 10'h154 == _T_107[9:0] ? 4'hb : _GEN_6102; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6104 = 10'h155 == _T_107[9:0] ? 4'h6 : _GEN_6103; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6105 = 10'h156 == _T_107[9:0] ? 4'hb : _GEN_6104; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6106 = 10'h157 == _T_107[9:0] ? 4'h7 : _GEN_6105; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6107 = 10'h158 == _T_107[9:0] ? 4'h7 : _GEN_6106; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6108 = 10'h159 == _T_107[9:0] ? 4'h7 : _GEN_6107; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6109 = 10'h15a == _T_107[9:0] ? 4'h7 : _GEN_6108; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6110 = 10'h15b == _T_107[9:0] ? 4'h7 : _GEN_6109; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6111 = 10'h15c == _T_107[9:0] ? 4'h7 : _GEN_6110; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6112 = 10'h15d == _T_107[9:0] ? 4'h6 : _GEN_6111; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6113 = 10'h15e == _T_107[9:0] ? 4'h7 : _GEN_6112; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6114 = 10'h15f == _T_107[9:0] ? 4'h0 : _GEN_6113; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6115 = 10'h160 == _T_107[9:0] ? 4'h0 : _GEN_6114; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6116 = 10'h161 == _T_107[9:0] ? 4'h0 : _GEN_6115; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6117 = 10'h162 == _T_107[9:0] ? 4'h0 : _GEN_6116; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6118 = 10'h163 == _T_107[9:0] ? 4'h2 : _GEN_6117; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6119 = 10'h164 == _T_107[9:0] ? 4'h4 : _GEN_6118; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6120 = 10'h165 == _T_107[9:0] ? 4'hb : _GEN_6119; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6121 = 10'h166 == _T_107[9:0] ? 4'hb : _GEN_6120; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6122 = 10'h167 == _T_107[9:0] ? 4'he : _GEN_6121; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6123 = 10'h168 == _T_107[9:0] ? 4'he : _GEN_6122; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6124 = 10'h169 == _T_107[9:0] ? 4'hc : _GEN_6123; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6125 = 10'h16a == _T_107[9:0] ? 4'hd : _GEN_6124; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6126 = 10'h16b == _T_107[9:0] ? 4'hd : _GEN_6125; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6127 = 10'h16c == _T_107[9:0] ? 4'ha : _GEN_6126; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6128 = 10'h16d == _T_107[9:0] ? 4'ha : _GEN_6127; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6129 = 10'h16e == _T_107[9:0] ? 4'ha : _GEN_6128; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6130 = 10'h16f == _T_107[9:0] ? 4'hd : _GEN_6129; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6131 = 10'h170 == _T_107[9:0] ? 4'hd : _GEN_6130; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6132 = 10'h171 == _T_107[9:0] ? 4'hd : _GEN_6131; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6133 = 10'h172 == _T_107[9:0] ? 4'he : _GEN_6132; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6134 = 10'h173 == _T_107[9:0] ? 4'h8 : _GEN_6133; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6135 = 10'h174 == _T_107[9:0] ? 4'h5 : _GEN_6134; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6136 = 10'h175 == _T_107[9:0] ? 4'h6 : _GEN_6135; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6137 = 10'h176 == _T_107[9:0] ? 4'h6 : _GEN_6136; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6138 = 10'h177 == _T_107[9:0] ? 4'h6 : _GEN_6137; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6139 = 10'h178 == _T_107[9:0] ? 4'h7 : _GEN_6138; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6140 = 10'h179 == _T_107[9:0] ? 4'h9 : _GEN_6139; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6141 = 10'h17a == _T_107[9:0] ? 4'h9 : _GEN_6140; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6142 = 10'h17b == _T_107[9:0] ? 4'h6 : _GEN_6141; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6143 = 10'h17c == _T_107[9:0] ? 4'h7 : _GEN_6142; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6144 = 10'h17d == _T_107[9:0] ? 4'h7 : _GEN_6143; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6145 = 10'h17e == _T_107[9:0] ? 4'h7 : _GEN_6144; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6146 = 10'h17f == _T_107[9:0] ? 4'h7 : _GEN_6145; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6147 = 10'h180 == _T_107[9:0] ? 4'h7 : _GEN_6146; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6148 = 10'h181 == _T_107[9:0] ? 4'h7 : _GEN_6147; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6149 = 10'h182 == _T_107[9:0] ? 4'h8 : _GEN_6148; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6150 = 10'h183 == _T_107[9:0] ? 4'h8 : _GEN_6149; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6151 = 10'h184 == _T_107[9:0] ? 4'h8 : _GEN_6150; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6152 = 10'h185 == _T_107[9:0] ? 4'h7 : _GEN_6151; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6153 = 10'h186 == _T_107[9:0] ? 4'h1 : _GEN_6152; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6154 = 10'h187 == _T_107[9:0] ? 4'h0 : _GEN_6153; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6155 = 10'h188 == _T_107[9:0] ? 4'h0 : _GEN_6154; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6156 = 10'h189 == _T_107[9:0] ? 4'h4 : _GEN_6155; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6157 = 10'h18a == _T_107[9:0] ? 4'h4 : _GEN_6156; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6158 = 10'h18b == _T_107[9:0] ? 4'hb : _GEN_6157; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6159 = 10'h18c == _T_107[9:0] ? 4'hb : _GEN_6158; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6160 = 10'h18d == _T_107[9:0] ? 4'hc : _GEN_6159; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6161 = 10'h18e == _T_107[9:0] ? 4'he : _GEN_6160; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6162 = 10'h18f == _T_107[9:0] ? 4'hb : _GEN_6161; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6163 = 10'h190 == _T_107[9:0] ? 4'hd : _GEN_6162; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6164 = 10'h191 == _T_107[9:0] ? 4'hc : _GEN_6163; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6165 = 10'h192 == _T_107[9:0] ? 4'h9 : _GEN_6164; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6166 = 10'h193 == _T_107[9:0] ? 4'ha : _GEN_6165; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6167 = 10'h194 == _T_107[9:0] ? 4'h9 : _GEN_6166; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6168 = 10'h195 == _T_107[9:0] ? 4'hd : _GEN_6167; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6169 = 10'h196 == _T_107[9:0] ? 4'hd : _GEN_6168; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6170 = 10'h197 == _T_107[9:0] ? 4'hb : _GEN_6169; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6171 = 10'h198 == _T_107[9:0] ? 4'he : _GEN_6170; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6172 = 10'h199 == _T_107[9:0] ? 4'h5 : _GEN_6171; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6173 = 10'h19a == _T_107[9:0] ? 4'h1 : _GEN_6172; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6174 = 10'h19b == _T_107[9:0] ? 4'h3 : _GEN_6173; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6175 = 10'h19c == _T_107[9:0] ? 4'h6 : _GEN_6174; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6176 = 10'h19d == _T_107[9:0] ? 4'h4 : _GEN_6175; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6177 = 10'h19e == _T_107[9:0] ? 4'h1 : _GEN_6176; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6178 = 10'h19f == _T_107[9:0] ? 4'h3 : _GEN_6177; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6179 = 10'h1a0 == _T_107[9:0] ? 4'h6 : _GEN_6178; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6180 = 10'h1a1 == _T_107[9:0] ? 4'h6 : _GEN_6179; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6181 = 10'h1a2 == _T_107[9:0] ? 4'h7 : _GEN_6180; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6182 = 10'h1a3 == _T_107[9:0] ? 4'h7 : _GEN_6181; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6183 = 10'h1a4 == _T_107[9:0] ? 4'h7 : _GEN_6182; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6184 = 10'h1a5 == _T_107[9:0] ? 4'h7 : _GEN_6183; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6185 = 10'h1a6 == _T_107[9:0] ? 4'h7 : _GEN_6184; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6186 = 10'h1a7 == _T_107[9:0] ? 4'h7 : _GEN_6185; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6187 = 10'h1a8 == _T_107[9:0] ? 4'h8 : _GEN_6186; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6188 = 10'h1a9 == _T_107[9:0] ? 4'h8 : _GEN_6187; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6189 = 10'h1aa == _T_107[9:0] ? 4'h7 : _GEN_6188; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6190 = 10'h1ab == _T_107[9:0] ? 4'h8 : _GEN_6189; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6191 = 10'h1ac == _T_107[9:0] ? 4'h8 : _GEN_6190; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6192 = 10'h1ad == _T_107[9:0] ? 4'h3 : _GEN_6191; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6193 = 10'h1ae == _T_107[9:0] ? 4'h2 : _GEN_6192; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6194 = 10'h1af == _T_107[9:0] ? 4'h8 : _GEN_6193; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6195 = 10'h1b0 == _T_107[9:0] ? 4'h6 : _GEN_6194; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6196 = 10'h1b1 == _T_107[9:0] ? 4'hb : _GEN_6195; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6197 = 10'h1b2 == _T_107[9:0] ? 4'hb : _GEN_6196; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6198 = 10'h1b3 == _T_107[9:0] ? 4'ha : _GEN_6197; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6199 = 10'h1b4 == _T_107[9:0] ? 4'he : _GEN_6198; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6200 = 10'h1b5 == _T_107[9:0] ? 4'hb : _GEN_6199; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6201 = 10'h1b6 == _T_107[9:0] ? 4'hc : _GEN_6200; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6202 = 10'h1b7 == _T_107[9:0] ? 4'ha : _GEN_6201; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6203 = 10'h1b8 == _T_107[9:0] ? 4'h9 : _GEN_6202; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6204 = 10'h1b9 == _T_107[9:0] ? 4'h9 : _GEN_6203; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6205 = 10'h1ba == _T_107[9:0] ? 4'h9 : _GEN_6204; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6206 = 10'h1bb == _T_107[9:0] ? 4'hb : _GEN_6205; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6207 = 10'h1bc == _T_107[9:0] ? 4'hd : _GEN_6206; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6208 = 10'h1bd == _T_107[9:0] ? 4'hd : _GEN_6207; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6209 = 10'h1be == _T_107[9:0] ? 4'he : _GEN_6208; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6210 = 10'h1bf == _T_107[9:0] ? 4'h7 : _GEN_6209; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6211 = 10'h1c0 == _T_107[9:0] ? 4'h6 : _GEN_6210; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6212 = 10'h1c1 == _T_107[9:0] ? 4'h6 : _GEN_6211; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6213 = 10'h1c2 == _T_107[9:0] ? 4'h5 : _GEN_6212; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6214 = 10'h1c3 == _T_107[9:0] ? 4'h5 : _GEN_6213; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6215 = 10'h1c4 == _T_107[9:0] ? 4'h4 : _GEN_6214; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6216 = 10'h1c5 == _T_107[9:0] ? 4'h5 : _GEN_6215; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6217 = 10'h1c6 == _T_107[9:0] ? 4'h6 : _GEN_6216; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6218 = 10'h1c7 == _T_107[9:0] ? 4'h6 : _GEN_6217; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6219 = 10'h1c8 == _T_107[9:0] ? 4'h7 : _GEN_6218; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6220 = 10'h1c9 == _T_107[9:0] ? 4'h7 : _GEN_6219; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6221 = 10'h1ca == _T_107[9:0] ? 4'h7 : _GEN_6220; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6222 = 10'h1cb == _T_107[9:0] ? 4'h7 : _GEN_6221; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6223 = 10'h1cc == _T_107[9:0] ? 4'h7 : _GEN_6222; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6224 = 10'h1cd == _T_107[9:0] ? 4'h8 : _GEN_6223; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6225 = 10'h1ce == _T_107[9:0] ? 4'h8 : _GEN_6224; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6226 = 10'h1cf == _T_107[9:0] ? 4'h8 : _GEN_6225; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6227 = 10'h1d0 == _T_107[9:0] ? 4'h5 : _GEN_6226; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6228 = 10'h1d1 == _T_107[9:0] ? 4'h8 : _GEN_6227; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6229 = 10'h1d2 == _T_107[9:0] ? 4'h8 : _GEN_6228; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6230 = 10'h1d3 == _T_107[9:0] ? 4'h8 : _GEN_6229; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6231 = 10'h1d4 == _T_107[9:0] ? 4'h8 : _GEN_6230; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6232 = 10'h1d5 == _T_107[9:0] ? 4'h7 : _GEN_6231; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6233 = 10'h1d6 == _T_107[9:0] ? 4'h9 : _GEN_6232; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6234 = 10'h1d7 == _T_107[9:0] ? 4'hb : _GEN_6233; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6235 = 10'h1d8 == _T_107[9:0] ? 4'hb : _GEN_6234; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6236 = 10'h1d9 == _T_107[9:0] ? 4'hb : _GEN_6235; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6237 = 10'h1da == _T_107[9:0] ? 4'ha : _GEN_6236; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6238 = 10'h1db == _T_107[9:0] ? 4'hc : _GEN_6237; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6239 = 10'h1dc == _T_107[9:0] ? 4'hb : _GEN_6238; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6240 = 10'h1dd == _T_107[9:0] ? 4'h5 : _GEN_6239; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6241 = 10'h1de == _T_107[9:0] ? 4'h9 : _GEN_6240; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6242 = 10'h1df == _T_107[9:0] ? 4'h9 : _GEN_6241; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6243 = 10'h1e0 == _T_107[9:0] ? 4'h9 : _GEN_6242; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6244 = 10'h1e1 == _T_107[9:0] ? 4'h7 : _GEN_6243; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6245 = 10'h1e2 == _T_107[9:0] ? 4'hc : _GEN_6244; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6246 = 10'h1e3 == _T_107[9:0] ? 4'hc : _GEN_6245; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6247 = 10'h1e4 == _T_107[9:0] ? 4'hd : _GEN_6246; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6248 = 10'h1e5 == _T_107[9:0] ? 4'h7 : _GEN_6247; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6249 = 10'h1e6 == _T_107[9:0] ? 4'h6 : _GEN_6248; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6250 = 10'h1e7 == _T_107[9:0] ? 4'h6 : _GEN_6249; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6251 = 10'h1e8 == _T_107[9:0] ? 4'h6 : _GEN_6250; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6252 = 10'h1e9 == _T_107[9:0] ? 4'h6 : _GEN_6251; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6253 = 10'h1ea == _T_107[9:0] ? 4'h6 : _GEN_6252; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6254 = 10'h1eb == _T_107[9:0] ? 4'h6 : _GEN_6253; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6255 = 10'h1ec == _T_107[9:0] ? 4'h6 : _GEN_6254; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6256 = 10'h1ed == _T_107[9:0] ? 4'h8 : _GEN_6255; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6257 = 10'h1ee == _T_107[9:0] ? 4'h7 : _GEN_6256; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6258 = 10'h1ef == _T_107[9:0] ? 4'h7 : _GEN_6257; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6259 = 10'h1f0 == _T_107[9:0] ? 4'h7 : _GEN_6258; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6260 = 10'h1f1 == _T_107[9:0] ? 4'h7 : _GEN_6259; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6261 = 10'h1f2 == _T_107[9:0] ? 4'h7 : _GEN_6260; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6262 = 10'h1f3 == _T_107[9:0] ? 4'h8 : _GEN_6261; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6263 = 10'h1f4 == _T_107[9:0] ? 4'h8 : _GEN_6262; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6264 = 10'h1f5 == _T_107[9:0] ? 4'h8 : _GEN_6263; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6265 = 10'h1f6 == _T_107[9:0] ? 4'ha : _GEN_6264; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6266 = 10'h1f7 == _T_107[9:0] ? 4'h8 : _GEN_6265; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6267 = 10'h1f8 == _T_107[9:0] ? 4'h8 : _GEN_6266; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6268 = 10'h1f9 == _T_107[9:0] ? 4'h9 : _GEN_6267; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6269 = 10'h1fa == _T_107[9:0] ? 4'h9 : _GEN_6268; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6270 = 10'h1fb == _T_107[9:0] ? 4'h8 : _GEN_6269; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6271 = 10'h1fc == _T_107[9:0] ? 4'hb : _GEN_6270; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6272 = 10'h1fd == _T_107[9:0] ? 4'hb : _GEN_6271; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6273 = 10'h1fe == _T_107[9:0] ? 4'hb : _GEN_6272; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6274 = 10'h1ff == _T_107[9:0] ? 4'ha : _GEN_6273; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6275 = 10'h200 == _T_107[9:0] ? 4'h3 : _GEN_6274; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6276 = 10'h201 == _T_107[9:0] ? 4'h9 : _GEN_6275; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6277 = 10'h202 == _T_107[9:0] ? 4'h5 : _GEN_6276; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6278 = 10'h203 == _T_107[9:0] ? 4'h3 : _GEN_6277; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6279 = 10'h204 == _T_107[9:0] ? 4'h4 : _GEN_6278; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6280 = 10'h205 == _T_107[9:0] ? 4'h4 : _GEN_6279; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6281 = 10'h206 == _T_107[9:0] ? 4'h4 : _GEN_6280; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6282 = 10'h207 == _T_107[9:0] ? 4'h4 : _GEN_6281; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6283 = 10'h208 == _T_107[9:0] ? 4'h8 : _GEN_6282; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6284 = 10'h209 == _T_107[9:0] ? 4'hc : _GEN_6283; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6285 = 10'h20a == _T_107[9:0] ? 4'hd : _GEN_6284; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6286 = 10'h20b == _T_107[9:0] ? 4'h7 : _GEN_6285; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6287 = 10'h20c == _T_107[9:0] ? 4'h6 : _GEN_6286; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6288 = 10'h20d == _T_107[9:0] ? 4'h6 : _GEN_6287; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6289 = 10'h20e == _T_107[9:0] ? 4'h6 : _GEN_6288; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6290 = 10'h20f == _T_107[9:0] ? 4'h5 : _GEN_6289; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6291 = 10'h210 == _T_107[9:0] ? 4'h6 : _GEN_6290; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6292 = 10'h211 == _T_107[9:0] ? 4'h6 : _GEN_6291; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6293 = 10'h212 == _T_107[9:0] ? 4'h7 : _GEN_6292; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6294 = 10'h213 == _T_107[9:0] ? 4'ha : _GEN_6293; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6295 = 10'h214 == _T_107[9:0] ? 4'h6 : _GEN_6294; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6296 = 10'h215 == _T_107[9:0] ? 4'h7 : _GEN_6295; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6297 = 10'h216 == _T_107[9:0] ? 4'h7 : _GEN_6296; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6298 = 10'h217 == _T_107[9:0] ? 4'h7 : _GEN_6297; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6299 = 10'h218 == _T_107[9:0] ? 4'h7 : _GEN_6298; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6300 = 10'h219 == _T_107[9:0] ? 4'h8 : _GEN_6299; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6301 = 10'h21a == _T_107[9:0] ? 4'h7 : _GEN_6300; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6302 = 10'h21b == _T_107[9:0] ? 4'h8 : _GEN_6301; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6303 = 10'h21c == _T_107[9:0] ? 4'hb : _GEN_6302; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6304 = 10'h21d == _T_107[9:0] ? 4'ha : _GEN_6303; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6305 = 10'h21e == _T_107[9:0] ? 4'h9 : _GEN_6304; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6306 = 10'h21f == _T_107[9:0] ? 4'h9 : _GEN_6305; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6307 = 10'h220 == _T_107[9:0] ? 4'h8 : _GEN_6306; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6308 = 10'h221 == _T_107[9:0] ? 4'h9 : _GEN_6307; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6309 = 10'h222 == _T_107[9:0] ? 4'hb : _GEN_6308; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6310 = 10'h223 == _T_107[9:0] ? 4'hb : _GEN_6309; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6311 = 10'h224 == _T_107[9:0] ? 4'hb : _GEN_6310; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6312 = 10'h225 == _T_107[9:0] ? 4'h8 : _GEN_6311; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6313 = 10'h226 == _T_107[9:0] ? 4'h1 : _GEN_6312; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6314 = 10'h227 == _T_107[9:0] ? 4'h3 : _GEN_6313; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6315 = 10'h228 == _T_107[9:0] ? 4'h3 : _GEN_6314; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6316 = 10'h229 == _T_107[9:0] ? 4'h3 : _GEN_6315; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6317 = 10'h22a == _T_107[9:0] ? 4'h3 : _GEN_6316; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6318 = 10'h22b == _T_107[9:0] ? 4'h3 : _GEN_6317; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6319 = 10'h22c == _T_107[9:0] ? 4'h3 : _GEN_6318; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6320 = 10'h22d == _T_107[9:0] ? 4'h3 : _GEN_6319; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6321 = 10'h22e == _T_107[9:0] ? 4'h3 : _GEN_6320; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6322 = 10'h22f == _T_107[9:0] ? 4'h9 : _GEN_6321; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6323 = 10'h230 == _T_107[9:0] ? 4'h6 : _GEN_6322; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6324 = 10'h231 == _T_107[9:0] ? 4'h7 : _GEN_6323; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6325 = 10'h232 == _T_107[9:0] ? 4'h6 : _GEN_6324; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6326 = 10'h233 == _T_107[9:0] ? 4'h7 : _GEN_6325; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6327 = 10'h234 == _T_107[9:0] ? 4'h7 : _GEN_6326; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6328 = 10'h235 == _T_107[9:0] ? 4'h6 : _GEN_6327; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6329 = 10'h236 == _T_107[9:0] ? 4'h6 : _GEN_6328; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6330 = 10'h237 == _T_107[9:0] ? 4'h6 : _GEN_6329; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6331 = 10'h238 == _T_107[9:0] ? 4'h6 : _GEN_6330; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6332 = 10'h239 == _T_107[9:0] ? 4'h8 : _GEN_6331; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6333 = 10'h23a == _T_107[9:0] ? 4'h6 : _GEN_6332; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6334 = 10'h23b == _T_107[9:0] ? 4'h7 : _GEN_6333; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6335 = 10'h23c == _T_107[9:0] ? 4'h7 : _GEN_6334; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6336 = 10'h23d == _T_107[9:0] ? 4'h7 : _GEN_6335; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6337 = 10'h23e == _T_107[9:0] ? 4'h7 : _GEN_6336; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6338 = 10'h23f == _T_107[9:0] ? 4'h7 : _GEN_6337; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6339 = 10'h240 == _T_107[9:0] ? 4'h7 : _GEN_6338; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6340 = 10'h241 == _T_107[9:0] ? 4'h8 : _GEN_6339; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6341 = 10'h242 == _T_107[9:0] ? 4'hb : _GEN_6340; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6342 = 10'h243 == _T_107[9:0] ? 4'hb : _GEN_6341; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6343 = 10'h244 == _T_107[9:0] ? 4'hb : _GEN_6342; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6344 = 10'h245 == _T_107[9:0] ? 4'ha : _GEN_6343; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6345 = 10'h246 == _T_107[9:0] ? 4'h9 : _GEN_6344; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6346 = 10'h247 == _T_107[9:0] ? 4'ha : _GEN_6345; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6347 = 10'h248 == _T_107[9:0] ? 4'hb : _GEN_6346; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6348 = 10'h249 == _T_107[9:0] ? 4'hb : _GEN_6347; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6349 = 10'h24a == _T_107[9:0] ? 4'ha : _GEN_6348; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6350 = 10'h24b == _T_107[9:0] ? 4'h2 : _GEN_6349; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6351 = 10'h24c == _T_107[9:0] ? 4'h0 : _GEN_6350; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6352 = 10'h24d == _T_107[9:0] ? 4'h2 : _GEN_6351; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6353 = 10'h24e == _T_107[9:0] ? 4'h3 : _GEN_6352; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6354 = 10'h24f == _T_107[9:0] ? 4'h3 : _GEN_6353; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6355 = 10'h250 == _T_107[9:0] ? 4'h3 : _GEN_6354; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6356 = 10'h251 == _T_107[9:0] ? 4'h3 : _GEN_6355; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6357 = 10'h252 == _T_107[9:0] ? 4'h3 : _GEN_6356; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6358 = 10'h253 == _T_107[9:0] ? 4'h3 : _GEN_6357; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6359 = 10'h254 == _T_107[9:0] ? 4'h3 : _GEN_6358; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6360 = 10'h255 == _T_107[9:0] ? 4'h5 : _GEN_6359; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6361 = 10'h256 == _T_107[9:0] ? 4'h6 : _GEN_6360; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6362 = 10'h257 == _T_107[9:0] ? 4'h8 : _GEN_6361; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6363 = 10'h258 == _T_107[9:0] ? 4'h5 : _GEN_6362; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6364 = 10'h259 == _T_107[9:0] ? 4'h6 : _GEN_6363; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6365 = 10'h25a == _T_107[9:0] ? 4'h6 : _GEN_6364; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6366 = 10'h25b == _T_107[9:0] ? 4'h5 : _GEN_6365; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6367 = 10'h25c == _T_107[9:0] ? 4'h6 : _GEN_6366; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6368 = 10'h25d == _T_107[9:0] ? 4'h6 : _GEN_6367; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6369 = 10'h25e == _T_107[9:0] ? 4'h9 : _GEN_6368; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6370 = 10'h25f == _T_107[9:0] ? 4'hc : _GEN_6369; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6371 = 10'h260 == _T_107[9:0] ? 4'h7 : _GEN_6370; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6372 = 10'h261 == _T_107[9:0] ? 4'h9 : _GEN_6371; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6373 = 10'h262 == _T_107[9:0] ? 4'ha : _GEN_6372; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6374 = 10'h263 == _T_107[9:0] ? 4'h8 : _GEN_6373; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6375 = 10'h264 == _T_107[9:0] ? 4'ha : _GEN_6374; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6376 = 10'h265 == _T_107[9:0] ? 4'h9 : _GEN_6375; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6377 = 10'h266 == _T_107[9:0] ? 4'h8 : _GEN_6376; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6378 = 10'h267 == _T_107[9:0] ? 4'h8 : _GEN_6377; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6379 = 10'h268 == _T_107[9:0] ? 4'ha : _GEN_6378; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6380 = 10'h269 == _T_107[9:0] ? 4'ha : _GEN_6379; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6381 = 10'h26a == _T_107[9:0] ? 4'hb : _GEN_6380; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6382 = 10'h26b == _T_107[9:0] ? 4'hb : _GEN_6381; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6383 = 10'h26c == _T_107[9:0] ? 4'hb : _GEN_6382; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6384 = 10'h26d == _T_107[9:0] ? 4'hb : _GEN_6383; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6385 = 10'h26e == _T_107[9:0] ? 4'hb : _GEN_6384; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6386 = 10'h26f == _T_107[9:0] ? 4'ha : _GEN_6385; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6387 = 10'h270 == _T_107[9:0] ? 4'h3 : _GEN_6386; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6388 = 10'h271 == _T_107[9:0] ? 4'h0 : _GEN_6387; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6389 = 10'h272 == _T_107[9:0] ? 4'h0 : _GEN_6388; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6390 = 10'h273 == _T_107[9:0] ? 4'h2 : _GEN_6389; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6391 = 10'h274 == _T_107[9:0] ? 4'h3 : _GEN_6390; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6392 = 10'h275 == _T_107[9:0] ? 4'h3 : _GEN_6391; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6393 = 10'h276 == _T_107[9:0] ? 4'h3 : _GEN_6392; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6394 = 10'h277 == _T_107[9:0] ? 4'h3 : _GEN_6393; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6395 = 10'h278 == _T_107[9:0] ? 4'h3 : _GEN_6394; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6396 = 10'h279 == _T_107[9:0] ? 4'h3 : _GEN_6395; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6397 = 10'h27a == _T_107[9:0] ? 4'h3 : _GEN_6396; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6398 = 10'h27b == _T_107[9:0] ? 4'h6 : _GEN_6397; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6399 = 10'h27c == _T_107[9:0] ? 4'h7 : _GEN_6398; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6400 = 10'h27d == _T_107[9:0] ? 4'h7 : _GEN_6399; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6401 = 10'h27e == _T_107[9:0] ? 4'h4 : _GEN_6400; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6402 = 10'h27f == _T_107[9:0] ? 4'h6 : _GEN_6401; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6403 = 10'h280 == _T_107[9:0] ? 4'h6 : _GEN_6402; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6404 = 10'h281 == _T_107[9:0] ? 4'h6 : _GEN_6403; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6405 = 10'h282 == _T_107[9:0] ? 4'h6 : _GEN_6404; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6406 = 10'h283 == _T_107[9:0] ? 4'ha : _GEN_6405; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6407 = 10'h284 == _T_107[9:0] ? 4'hc : _GEN_6406; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6408 = 10'h285 == _T_107[9:0] ? 4'hc : _GEN_6407; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6409 = 10'h286 == _T_107[9:0] ? 4'h8 : _GEN_6408; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6410 = 10'h287 == _T_107[9:0] ? 4'ha : _GEN_6409; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6411 = 10'h288 == _T_107[9:0] ? 4'ha : _GEN_6410; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6412 = 10'h289 == _T_107[9:0] ? 4'ha : _GEN_6411; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6413 = 10'h28a == _T_107[9:0] ? 4'hc : _GEN_6412; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6414 = 10'h28b == _T_107[9:0] ? 4'hb : _GEN_6413; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6415 = 10'h28c == _T_107[9:0] ? 4'ha : _GEN_6414; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6416 = 10'h28d == _T_107[9:0] ? 4'h7 : _GEN_6415; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6417 = 10'h28e == _T_107[9:0] ? 4'h2 : _GEN_6416; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6418 = 10'h28f == _T_107[9:0] ? 4'h5 : _GEN_6417; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6419 = 10'h290 == _T_107[9:0] ? 4'h8 : _GEN_6418; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6420 = 10'h291 == _T_107[9:0] ? 4'ha : _GEN_6419; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6421 = 10'h292 == _T_107[9:0] ? 4'ha : _GEN_6420; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6422 = 10'h293 == _T_107[9:0] ? 4'ha : _GEN_6421; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6423 = 10'h294 == _T_107[9:0] ? 4'h9 : _GEN_6422; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6424 = 10'h295 == _T_107[9:0] ? 4'h3 : _GEN_6423; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6425 = 10'h296 == _T_107[9:0] ? 4'h0 : _GEN_6424; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6426 = 10'h297 == _T_107[9:0] ? 4'h0 : _GEN_6425; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6427 = 10'h298 == _T_107[9:0] ? 4'h0 : _GEN_6426; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6428 = 10'h299 == _T_107[9:0] ? 4'h1 : _GEN_6427; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6429 = 10'h29a == _T_107[9:0] ? 4'h3 : _GEN_6428; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6430 = 10'h29b == _T_107[9:0] ? 4'h3 : _GEN_6429; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6431 = 10'h29c == _T_107[9:0] ? 4'h3 : _GEN_6430; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6432 = 10'h29d == _T_107[9:0] ? 4'h3 : _GEN_6431; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6433 = 10'h29e == _T_107[9:0] ? 4'h3 : _GEN_6432; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6434 = 10'h29f == _T_107[9:0] ? 4'h3 : _GEN_6433; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6435 = 10'h2a0 == _T_107[9:0] ? 4'h4 : _GEN_6434; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6436 = 10'h2a1 == _T_107[9:0] ? 4'h6 : _GEN_6435; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6437 = 10'h2a2 == _T_107[9:0] ? 4'h7 : _GEN_6436; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6438 = 10'h2a3 == _T_107[9:0] ? 4'h6 : _GEN_6437; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6439 = 10'h2a4 == _T_107[9:0] ? 4'h4 : _GEN_6438; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6440 = 10'h2a5 == _T_107[9:0] ? 4'h6 : _GEN_6439; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6441 = 10'h2a6 == _T_107[9:0] ? 4'h6 : _GEN_6440; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6442 = 10'h2a7 == _T_107[9:0] ? 4'h7 : _GEN_6441; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6443 = 10'h2a8 == _T_107[9:0] ? 4'ha : _GEN_6442; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6444 = 10'h2a9 == _T_107[9:0] ? 4'hb : _GEN_6443; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6445 = 10'h2aa == _T_107[9:0] ? 4'hb : _GEN_6444; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6446 = 10'h2ab == _T_107[9:0] ? 4'hb : _GEN_6445; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6447 = 10'h2ac == _T_107[9:0] ? 4'h8 : _GEN_6446; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6448 = 10'h2ad == _T_107[9:0] ? 4'hb : _GEN_6447; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6449 = 10'h2ae == _T_107[9:0] ? 4'ha : _GEN_6448; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6450 = 10'h2af == _T_107[9:0] ? 4'hb : _GEN_6449; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6451 = 10'h2b0 == _T_107[9:0] ? 4'hc : _GEN_6450; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6452 = 10'h2b1 == _T_107[9:0] ? 4'hb : _GEN_6451; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6453 = 10'h2b2 == _T_107[9:0] ? 4'ha : _GEN_6452; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6454 = 10'h2b3 == _T_107[9:0] ? 4'h6 : _GEN_6453; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6455 = 10'h2b4 == _T_107[9:0] ? 4'h0 : _GEN_6454; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6456 = 10'h2b5 == _T_107[9:0] ? 4'h0 : _GEN_6455; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6457 = 10'h2b6 == _T_107[9:0] ? 4'h0 : _GEN_6456; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6458 = 10'h2b7 == _T_107[9:0] ? 4'h1 : _GEN_6457; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6459 = 10'h2b8 == _T_107[9:0] ? 4'h5 : _GEN_6458; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6460 = 10'h2b9 == _T_107[9:0] ? 4'h9 : _GEN_6459; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6461 = 10'h2ba == _T_107[9:0] ? 4'h1 : _GEN_6460; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6462 = 10'h2bb == _T_107[9:0] ? 4'h0 : _GEN_6461; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6463 = 10'h2bc == _T_107[9:0] ? 4'h0 : _GEN_6462; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6464 = 10'h2bd == _T_107[9:0] ? 4'h0 : _GEN_6463; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6465 = 10'h2be == _T_107[9:0] ? 4'h0 : _GEN_6464; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6466 = 10'h2bf == _T_107[9:0] ? 4'h0 : _GEN_6465; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6467 = 10'h2c0 == _T_107[9:0] ? 4'h3 : _GEN_6466; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6468 = 10'h2c1 == _T_107[9:0] ? 4'h3 : _GEN_6467; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6469 = 10'h2c2 == _T_107[9:0] ? 4'h3 : _GEN_6468; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6470 = 10'h2c3 == _T_107[9:0] ? 4'h3 : _GEN_6469; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6471 = 10'h2c4 == _T_107[9:0] ? 4'h3 : _GEN_6470; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6472 = 10'h2c5 == _T_107[9:0] ? 4'h3 : _GEN_6471; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6473 = 10'h2c6 == _T_107[9:0] ? 4'h4 : _GEN_6472; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6474 = 10'h2c7 == _T_107[9:0] ? 4'h5 : _GEN_6473; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6475 = 10'h2c8 == _T_107[9:0] ? 4'h7 : _GEN_6474; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6476 = 10'h2c9 == _T_107[9:0] ? 4'h7 : _GEN_6475; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6477 = 10'h2ca == _T_107[9:0] ? 4'h4 : _GEN_6476; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6478 = 10'h2cb == _T_107[9:0] ? 4'h9 : _GEN_6477; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6479 = 10'h2cc == _T_107[9:0] ? 4'h9 : _GEN_6478; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6480 = 10'h2cd == _T_107[9:0] ? 4'hb : _GEN_6479; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6481 = 10'h2ce == _T_107[9:0] ? 4'hb : _GEN_6480; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6482 = 10'h2cf == _T_107[9:0] ? 4'hb : _GEN_6481; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6483 = 10'h2d0 == _T_107[9:0] ? 4'hb : _GEN_6482; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6484 = 10'h2d1 == _T_107[9:0] ? 4'hb : _GEN_6483; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6485 = 10'h2d2 == _T_107[9:0] ? 4'h8 : _GEN_6484; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6486 = 10'h2d3 == _T_107[9:0] ? 4'ha : _GEN_6485; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6487 = 10'h2d4 == _T_107[9:0] ? 4'hb : _GEN_6486; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6488 = 10'h2d5 == _T_107[9:0] ? 4'ha : _GEN_6487; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6489 = 10'h2d6 == _T_107[9:0] ? 4'ha : _GEN_6488; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6490 = 10'h2d7 == _T_107[9:0] ? 4'ha : _GEN_6489; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6491 = 10'h2d8 == _T_107[9:0] ? 4'ha : _GEN_6490; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6492 = 10'h2d9 == _T_107[9:0] ? 4'h7 : _GEN_6491; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6493 = 10'h2da == _T_107[9:0] ? 4'h2 : _GEN_6492; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6494 = 10'h2db == _T_107[9:0] ? 4'h0 : _GEN_6493; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6495 = 10'h2dc == _T_107[9:0] ? 4'h0 : _GEN_6494; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6496 = 10'h2dd == _T_107[9:0] ? 4'h0 : _GEN_6495; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6497 = 10'h2de == _T_107[9:0] ? 4'h0 : _GEN_6496; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6498 = 10'h2df == _T_107[9:0] ? 4'h2 : _GEN_6497; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6499 = 10'h2e0 == _T_107[9:0] ? 4'h0 : _GEN_6498; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6500 = 10'h2e1 == _T_107[9:0] ? 4'h0 : _GEN_6499; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6501 = 10'h2e2 == _T_107[9:0] ? 4'h0 : _GEN_6500; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6502 = 10'h2e3 == _T_107[9:0] ? 4'h0 : _GEN_6501; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6503 = 10'h2e4 == _T_107[9:0] ? 4'h0 : _GEN_6502; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6504 = 10'h2e5 == _T_107[9:0] ? 4'h0 : _GEN_6503; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6505 = 10'h2e6 == _T_107[9:0] ? 4'h2 : _GEN_6504; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6506 = 10'h2e7 == _T_107[9:0] ? 4'h3 : _GEN_6505; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6507 = 10'h2e8 == _T_107[9:0] ? 4'h3 : _GEN_6506; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6508 = 10'h2e9 == _T_107[9:0] ? 4'h3 : _GEN_6507; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6509 = 10'h2ea == _T_107[9:0] ? 4'h3 : _GEN_6508; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6510 = 10'h2eb == _T_107[9:0] ? 4'h3 : _GEN_6509; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6511 = 10'h2ec == _T_107[9:0] ? 4'h4 : _GEN_6510; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6512 = 10'h2ed == _T_107[9:0] ? 4'h5 : _GEN_6511; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6513 = 10'h2ee == _T_107[9:0] ? 4'h6 : _GEN_6512; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6514 = 10'h2ef == _T_107[9:0] ? 4'h8 : _GEN_6513; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6515 = 10'h2f0 == _T_107[9:0] ? 4'h4 : _GEN_6514; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6516 = 10'h2f1 == _T_107[9:0] ? 4'h9 : _GEN_6515; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6517 = 10'h2f2 == _T_107[9:0] ? 4'hb : _GEN_6516; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6518 = 10'h2f3 == _T_107[9:0] ? 4'hb : _GEN_6517; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6519 = 10'h2f4 == _T_107[9:0] ? 4'hb : _GEN_6518; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6520 = 10'h2f5 == _T_107[9:0] ? 4'hb : _GEN_6519; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6521 = 10'h2f6 == _T_107[9:0] ? 4'hb : _GEN_6520; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6522 = 10'h2f7 == _T_107[9:0] ? 4'hb : _GEN_6521; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6523 = 10'h2f8 == _T_107[9:0] ? 4'h8 : _GEN_6522; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6524 = 10'h2f9 == _T_107[9:0] ? 4'h9 : _GEN_6523; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6525 = 10'h2fa == _T_107[9:0] ? 4'hb : _GEN_6524; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6526 = 10'h2fb == _T_107[9:0] ? 4'hb : _GEN_6525; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6527 = 10'h2fc == _T_107[9:0] ? 4'ha : _GEN_6526; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6528 = 10'h2fd == _T_107[9:0] ? 4'ha : _GEN_6527; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6529 = 10'h2fe == _T_107[9:0] ? 4'h9 : _GEN_6528; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6530 = 10'h2ff == _T_107[9:0] ? 4'h8 : _GEN_6529; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6531 = 10'h300 == _T_107[9:0] ? 4'h8 : _GEN_6530; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6532 = 10'h301 == _T_107[9:0] ? 4'h6 : _GEN_6531; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6533 = 10'h302 == _T_107[9:0] ? 4'h1 : _GEN_6532; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6534 = 10'h303 == _T_107[9:0] ? 4'h0 : _GEN_6533; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6535 = 10'h304 == _T_107[9:0] ? 4'h0 : _GEN_6534; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6536 = 10'h305 == _T_107[9:0] ? 4'h0 : _GEN_6535; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6537 = 10'h306 == _T_107[9:0] ? 4'h0 : _GEN_6536; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6538 = 10'h307 == _T_107[9:0] ? 4'h0 : _GEN_6537; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6539 = 10'h308 == _T_107[9:0] ? 4'h0 : _GEN_6538; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6540 = 10'h309 == _T_107[9:0] ? 4'h0 : _GEN_6539; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6541 = 10'h30a == _T_107[9:0] ? 4'h0 : _GEN_6540; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6542 = 10'h30b == _T_107[9:0] ? 4'h0 : _GEN_6541; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6543 = 10'h30c == _T_107[9:0] ? 4'h2 : _GEN_6542; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6544 = 10'h30d == _T_107[9:0] ? 4'h3 : _GEN_6543; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6545 = 10'h30e == _T_107[9:0] ? 4'h3 : _GEN_6544; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6546 = 10'h30f == _T_107[9:0] ? 4'h3 : _GEN_6545; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6547 = 10'h310 == _T_107[9:0] ? 4'h3 : _GEN_6546; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6548 = 10'h311 == _T_107[9:0] ? 4'h3 : _GEN_6547; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6549 = 10'h312 == _T_107[9:0] ? 4'h4 : _GEN_6548; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6550 = 10'h313 == _T_107[9:0] ? 4'h5 : _GEN_6549; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6551 = 10'h314 == _T_107[9:0] ? 4'h5 : _GEN_6550; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6552 = 10'h315 == _T_107[9:0] ? 4'h8 : _GEN_6551; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6553 = 10'h316 == _T_107[9:0] ? 4'h4 : _GEN_6552; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6554 = 10'h317 == _T_107[9:0] ? 4'h6 : _GEN_6553; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6555 = 10'h318 == _T_107[9:0] ? 4'hb : _GEN_6554; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6556 = 10'h319 == _T_107[9:0] ? 4'hb : _GEN_6555; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6557 = 10'h31a == _T_107[9:0] ? 4'hb : _GEN_6556; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6558 = 10'h31b == _T_107[9:0] ? 4'hb : _GEN_6557; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6559 = 10'h31c == _T_107[9:0] ? 4'hb : _GEN_6558; // @[Filter.scala 230:102]
  wire [3:0] _GEN_6560 = 10'h31d == _T_107[9:0] ? 4'hb : _GEN_6559; // @[Filter.scala 230:102]
  wire [6:0] _GEN_38968 = {{3'd0}, _GEN_6560}; // @[Filter.scala 230:102]
  wire [10:0] _T_114 = _GEN_38968 * 7'h46; // @[Filter.scala 230:102]
  wire [10:0] _GEN_38969 = {{2'd0}, _T_109}; // @[Filter.scala 230:69]
  wire [10:0] _T_116 = _GEN_38969 + _T_114; // @[Filter.scala 230:69]
  wire [3:0] _GEN_6583 = 10'h16 == _T_107[9:0] ? 4'hb : 4'hc; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6584 = 10'h17 == _T_107[9:0] ? 4'h8 : _GEN_6583; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6585 = 10'h18 == _T_107[9:0] ? 4'ha : _GEN_6584; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6586 = 10'h19 == _T_107[9:0] ? 4'hc : _GEN_6585; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6587 = 10'h1a == _T_107[9:0] ? 4'hc : _GEN_6586; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6588 = 10'h1b == _T_107[9:0] ? 4'hc : _GEN_6587; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6589 = 10'h1c == _T_107[9:0] ? 4'hc : _GEN_6588; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6590 = 10'h1d == _T_107[9:0] ? 4'hc : _GEN_6589; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6591 = 10'h1e == _T_107[9:0] ? 4'hc : _GEN_6590; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6592 = 10'h1f == _T_107[9:0] ? 4'hc : _GEN_6591; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6593 = 10'h20 == _T_107[9:0] ? 4'hc : _GEN_6592; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6594 = 10'h21 == _T_107[9:0] ? 4'hc : _GEN_6593; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6595 = 10'h22 == _T_107[9:0] ? 4'hc : _GEN_6594; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6596 = 10'h23 == _T_107[9:0] ? 4'hc : _GEN_6595; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6597 = 10'h24 == _T_107[9:0] ? 4'hc : _GEN_6596; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6598 = 10'h25 == _T_107[9:0] ? 4'hc : _GEN_6597; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6599 = 10'h26 == _T_107[9:0] ? 4'hc : _GEN_6598; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6600 = 10'h27 == _T_107[9:0] ? 4'hc : _GEN_6599; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6601 = 10'h28 == _T_107[9:0] ? 4'hc : _GEN_6600; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6602 = 10'h29 == _T_107[9:0] ? 4'hc : _GEN_6601; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6603 = 10'h2a == _T_107[9:0] ? 4'hc : _GEN_6602; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6604 = 10'h2b == _T_107[9:0] ? 4'hc : _GEN_6603; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6605 = 10'h2c == _T_107[9:0] ? 4'hc : _GEN_6604; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6606 = 10'h2d == _T_107[9:0] ? 4'hc : _GEN_6605; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6607 = 10'h2e == _T_107[9:0] ? 4'hc : _GEN_6606; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6608 = 10'h2f == _T_107[9:0] ? 4'hc : _GEN_6607; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6609 = 10'h30 == _T_107[9:0] ? 4'hc : _GEN_6608; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6610 = 10'h31 == _T_107[9:0] ? 4'hc : _GEN_6609; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6611 = 10'h32 == _T_107[9:0] ? 4'hc : _GEN_6610; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6612 = 10'h33 == _T_107[9:0] ? 4'hc : _GEN_6611; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6613 = 10'h34 == _T_107[9:0] ? 4'hc : _GEN_6612; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6614 = 10'h35 == _T_107[9:0] ? 4'hc : _GEN_6613; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6615 = 10'h36 == _T_107[9:0] ? 4'hc : _GEN_6614; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6616 = 10'h37 == _T_107[9:0] ? 4'hc : _GEN_6615; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6617 = 10'h38 == _T_107[9:0] ? 4'hc : _GEN_6616; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6618 = 10'h39 == _T_107[9:0] ? 4'hc : _GEN_6617; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6619 = 10'h3a == _T_107[9:0] ? 4'hc : _GEN_6618; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6620 = 10'h3b == _T_107[9:0] ? 4'hc : _GEN_6619; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6621 = 10'h3c == _T_107[9:0] ? 4'h7 : _GEN_6620; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6622 = 10'h3d == _T_107[9:0] ? 4'h9 : _GEN_6621; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6623 = 10'h3e == _T_107[9:0] ? 4'h8 : _GEN_6622; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6624 = 10'h3f == _T_107[9:0] ? 4'hc : _GEN_6623; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6625 = 10'h40 == _T_107[9:0] ? 4'hc : _GEN_6624; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6626 = 10'h41 == _T_107[9:0] ? 4'hc : _GEN_6625; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6627 = 10'h42 == _T_107[9:0] ? 4'hc : _GEN_6626; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6628 = 10'h43 == _T_107[9:0] ? 4'hc : _GEN_6627; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6629 = 10'h44 == _T_107[9:0] ? 4'hc : _GEN_6628; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6630 = 10'h45 == _T_107[9:0] ? 4'hc : _GEN_6629; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6631 = 10'h46 == _T_107[9:0] ? 4'hc : _GEN_6630; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6632 = 10'h47 == _T_107[9:0] ? 4'hc : _GEN_6631; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6633 = 10'h48 == _T_107[9:0] ? 4'hc : _GEN_6632; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6634 = 10'h49 == _T_107[9:0] ? 4'hc : _GEN_6633; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6635 = 10'h4a == _T_107[9:0] ? 4'hc : _GEN_6634; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6636 = 10'h4b == _T_107[9:0] ? 4'hc : _GEN_6635; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6637 = 10'h4c == _T_107[9:0] ? 4'hc : _GEN_6636; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6638 = 10'h4d == _T_107[9:0] ? 4'hc : _GEN_6637; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6639 = 10'h4e == _T_107[9:0] ? 4'hc : _GEN_6638; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6640 = 10'h4f == _T_107[9:0] ? 4'hc : _GEN_6639; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6641 = 10'h50 == _T_107[9:0] ? 4'hc : _GEN_6640; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6642 = 10'h51 == _T_107[9:0] ? 4'hc : _GEN_6641; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6643 = 10'h52 == _T_107[9:0] ? 4'hc : _GEN_6642; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6644 = 10'h53 == _T_107[9:0] ? 4'hc : _GEN_6643; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6645 = 10'h54 == _T_107[9:0] ? 4'hc : _GEN_6644; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6646 = 10'h55 == _T_107[9:0] ? 4'hc : _GEN_6645; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6647 = 10'h56 == _T_107[9:0] ? 4'hc : _GEN_6646; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6648 = 10'h57 == _T_107[9:0] ? 4'hc : _GEN_6647; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6649 = 10'h58 == _T_107[9:0] ? 4'hc : _GEN_6648; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6650 = 10'h59 == _T_107[9:0] ? 4'hc : _GEN_6649; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6651 = 10'h5a == _T_107[9:0] ? 4'h9 : _GEN_6650; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6652 = 10'h5b == _T_107[9:0] ? 4'ha : _GEN_6651; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6653 = 10'h5c == _T_107[9:0] ? 4'hc : _GEN_6652; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6654 = 10'h5d == _T_107[9:0] ? 4'hc : _GEN_6653; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6655 = 10'h5e == _T_107[9:0] ? 4'hc : _GEN_6654; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6656 = 10'h5f == _T_107[9:0] ? 4'hc : _GEN_6655; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6657 = 10'h60 == _T_107[9:0] ? 4'hc : _GEN_6656; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6658 = 10'h61 == _T_107[9:0] ? 4'hb : _GEN_6657; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6659 = 10'h62 == _T_107[9:0] ? 4'h8 : _GEN_6658; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6660 = 10'h63 == _T_107[9:0] ? 4'h9 : _GEN_6659; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6661 = 10'h64 == _T_107[9:0] ? 4'h7 : _GEN_6660; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6662 = 10'h65 == _T_107[9:0] ? 4'hb : _GEN_6661; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6663 = 10'h66 == _T_107[9:0] ? 4'hc : _GEN_6662; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6664 = 10'h67 == _T_107[9:0] ? 4'hc : _GEN_6663; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6665 = 10'h68 == _T_107[9:0] ? 4'hc : _GEN_6664; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6666 = 10'h69 == _T_107[9:0] ? 4'hc : _GEN_6665; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6667 = 10'h6a == _T_107[9:0] ? 4'hc : _GEN_6666; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6668 = 10'h6b == _T_107[9:0] ? 4'hb : _GEN_6667; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6669 = 10'h6c == _T_107[9:0] ? 4'h9 : _GEN_6668; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6670 = 10'h6d == _T_107[9:0] ? 4'ha : _GEN_6669; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6671 = 10'h6e == _T_107[9:0] ? 4'hc : _GEN_6670; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6672 = 10'h6f == _T_107[9:0] ? 4'hc : _GEN_6671; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6673 = 10'h70 == _T_107[9:0] ? 4'hc : _GEN_6672; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6674 = 10'h71 == _T_107[9:0] ? 4'hc : _GEN_6673; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6675 = 10'h72 == _T_107[9:0] ? 4'hc : _GEN_6674; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6676 = 10'h73 == _T_107[9:0] ? 4'hc : _GEN_6675; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6677 = 10'h74 == _T_107[9:0] ? 4'hc : _GEN_6676; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6678 = 10'h75 == _T_107[9:0] ? 4'hc : _GEN_6677; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6679 = 10'h76 == _T_107[9:0] ? 4'hc : _GEN_6678; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6680 = 10'h77 == _T_107[9:0] ? 4'hc : _GEN_6679; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6681 = 10'h78 == _T_107[9:0] ? 4'hc : _GEN_6680; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6682 = 10'h79 == _T_107[9:0] ? 4'hc : _GEN_6681; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6683 = 10'h7a == _T_107[9:0] ? 4'hc : _GEN_6682; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6684 = 10'h7b == _T_107[9:0] ? 4'hc : _GEN_6683; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6685 = 10'h7c == _T_107[9:0] ? 4'hc : _GEN_6684; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6686 = 10'h7d == _T_107[9:0] ? 4'hc : _GEN_6685; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6687 = 10'h7e == _T_107[9:0] ? 4'hc : _GEN_6686; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6688 = 10'h7f == _T_107[9:0] ? 4'hc : _GEN_6687; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6689 = 10'h80 == _T_107[9:0] ? 4'hc : _GEN_6688; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6690 = 10'h81 == _T_107[9:0] ? 4'h9 : _GEN_6689; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6691 = 10'h82 == _T_107[9:0] ? 4'h9 : _GEN_6690; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6692 = 10'h83 == _T_107[9:0] ? 4'h9 : _GEN_6691; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6693 = 10'h84 == _T_107[9:0] ? 4'hc : _GEN_6692; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6694 = 10'h85 == _T_107[9:0] ? 4'hc : _GEN_6693; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6695 = 10'h86 == _T_107[9:0] ? 4'hc : _GEN_6694; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6696 = 10'h87 == _T_107[9:0] ? 4'h8 : _GEN_6695; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6697 = 10'h88 == _T_107[9:0] ? 4'h9 : _GEN_6696; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6698 = 10'h89 == _T_107[9:0] ? 4'h9 : _GEN_6697; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6699 = 10'h8a == _T_107[9:0] ? 4'h9 : _GEN_6698; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6700 = 10'h8b == _T_107[9:0] ? 4'hc : _GEN_6699; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6701 = 10'h8c == _T_107[9:0] ? 4'hc : _GEN_6700; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6702 = 10'h8d == _T_107[9:0] ? 4'hc : _GEN_6701; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6703 = 10'h8e == _T_107[9:0] ? 4'hc : _GEN_6702; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6704 = 10'h8f == _T_107[9:0] ? 4'h9 : _GEN_6703; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6705 = 10'h90 == _T_107[9:0] ? 4'h9 : _GEN_6704; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6706 = 10'h91 == _T_107[9:0] ? 4'h9 : _GEN_6705; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6707 = 10'h92 == _T_107[9:0] ? 4'ha : _GEN_6706; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6708 = 10'h93 == _T_107[9:0] ? 4'hc : _GEN_6707; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6709 = 10'h94 == _T_107[9:0] ? 4'hc : _GEN_6708; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6710 = 10'h95 == _T_107[9:0] ? 4'hc : _GEN_6709; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6711 = 10'h96 == _T_107[9:0] ? 4'hc : _GEN_6710; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6712 = 10'h97 == _T_107[9:0] ? 4'hc : _GEN_6711; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6713 = 10'h98 == _T_107[9:0] ? 4'hc : _GEN_6712; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6714 = 10'h99 == _T_107[9:0] ? 4'hc : _GEN_6713; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6715 = 10'h9a == _T_107[9:0] ? 4'hc : _GEN_6714; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6716 = 10'h9b == _T_107[9:0] ? 4'hc : _GEN_6715; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6717 = 10'h9c == _T_107[9:0] ? 4'hc : _GEN_6716; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6718 = 10'h9d == _T_107[9:0] ? 4'hc : _GEN_6717; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6719 = 10'h9e == _T_107[9:0] ? 4'hc : _GEN_6718; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6720 = 10'h9f == _T_107[9:0] ? 4'hc : _GEN_6719; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6721 = 10'ha0 == _T_107[9:0] ? 4'hc : _GEN_6720; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6722 = 10'ha1 == _T_107[9:0] ? 4'hc : _GEN_6721; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6723 = 10'ha2 == _T_107[9:0] ? 4'hc : _GEN_6722; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6724 = 10'ha3 == _T_107[9:0] ? 4'hc : _GEN_6723; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6725 = 10'ha4 == _T_107[9:0] ? 4'hc : _GEN_6724; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6726 = 10'ha5 == _T_107[9:0] ? 4'hc : _GEN_6725; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6727 = 10'ha6 == _T_107[9:0] ? 4'hc : _GEN_6726; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6728 = 10'ha7 == _T_107[9:0] ? 4'hc : _GEN_6727; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6729 = 10'ha8 == _T_107[9:0] ? 4'h9 : _GEN_6728; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6730 = 10'ha9 == _T_107[9:0] ? 4'h8 : _GEN_6729; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6731 = 10'haa == _T_107[9:0] ? 4'h8 : _GEN_6730; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6732 = 10'hab == _T_107[9:0] ? 4'ha : _GEN_6731; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6733 = 10'hac == _T_107[9:0] ? 4'hb : _GEN_6732; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6734 = 10'had == _T_107[9:0] ? 4'h7 : _GEN_6733; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6735 = 10'hae == _T_107[9:0] ? 4'h9 : _GEN_6734; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6736 = 10'haf == _T_107[9:0] ? 4'h9 : _GEN_6735; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6737 = 10'hb0 == _T_107[9:0] ? 4'h8 : _GEN_6736; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6738 = 10'hb1 == _T_107[9:0] ? 4'h9 : _GEN_6737; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6739 = 10'hb2 == _T_107[9:0] ? 4'hc : _GEN_6738; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6740 = 10'hb3 == _T_107[9:0] ? 4'h9 : _GEN_6739; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6741 = 10'hb4 == _T_107[9:0] ? 4'h9 : _GEN_6740; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6742 = 10'hb5 == _T_107[9:0] ? 4'h9 : _GEN_6741; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6743 = 10'hb6 == _T_107[9:0] ? 4'h9 : _GEN_6742; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6744 = 10'hb7 == _T_107[9:0] ? 4'ha : _GEN_6743; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6745 = 10'hb8 == _T_107[9:0] ? 4'hc : _GEN_6744; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6746 = 10'hb9 == _T_107[9:0] ? 4'hc : _GEN_6745; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6747 = 10'hba == _T_107[9:0] ? 4'hc : _GEN_6746; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6748 = 10'hbb == _T_107[9:0] ? 4'hc : _GEN_6747; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6749 = 10'hbc == _T_107[9:0] ? 4'hc : _GEN_6748; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6750 = 10'hbd == _T_107[9:0] ? 4'hb : _GEN_6749; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6751 = 10'hbe == _T_107[9:0] ? 4'hc : _GEN_6750; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6752 = 10'hbf == _T_107[9:0] ? 4'hc : _GEN_6751; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6753 = 10'hc0 == _T_107[9:0] ? 4'hc : _GEN_6752; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6754 = 10'hc1 == _T_107[9:0] ? 4'hc : _GEN_6753; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6755 = 10'hc2 == _T_107[9:0] ? 4'hc : _GEN_6754; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6756 = 10'hc3 == _T_107[9:0] ? 4'hc : _GEN_6755; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6757 = 10'hc4 == _T_107[9:0] ? 4'hc : _GEN_6756; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6758 = 10'hc5 == _T_107[9:0] ? 4'hc : _GEN_6757; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6759 = 10'hc6 == _T_107[9:0] ? 4'hb : _GEN_6758; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6760 = 10'hc7 == _T_107[9:0] ? 4'hb : _GEN_6759; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6761 = 10'hc8 == _T_107[9:0] ? 4'ha : _GEN_6760; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6762 = 10'hc9 == _T_107[9:0] ? 4'ha : _GEN_6761; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6763 = 10'hca == _T_107[9:0] ? 4'hb : _GEN_6762; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6764 = 10'hcb == _T_107[9:0] ? 4'hc : _GEN_6763; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6765 = 10'hcc == _T_107[9:0] ? 4'hc : _GEN_6764; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6766 = 10'hcd == _T_107[9:0] ? 4'hc : _GEN_6765; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6767 = 10'hce == _T_107[9:0] ? 4'ha : _GEN_6766; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6768 = 10'hcf == _T_107[9:0] ? 4'h8 : _GEN_6767; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6769 = 10'hd0 == _T_107[9:0] ? 4'h9 : _GEN_6768; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6770 = 10'hd1 == _T_107[9:0] ? 4'h8 : _GEN_6769; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6771 = 10'hd2 == _T_107[9:0] ? 4'h9 : _GEN_6770; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6772 = 10'hd3 == _T_107[9:0] ? 4'h9 : _GEN_6771; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6773 = 10'hd4 == _T_107[9:0] ? 4'h9 : _GEN_6772; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6774 = 10'hd5 == _T_107[9:0] ? 4'h9 : _GEN_6773; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6775 = 10'hd6 == _T_107[9:0] ? 4'ha : _GEN_6774; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6776 = 10'hd7 == _T_107[9:0] ? 4'h9 : _GEN_6775; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6777 = 10'hd8 == _T_107[9:0] ? 4'h9 : _GEN_6776; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6778 = 10'hd9 == _T_107[9:0] ? 4'h9 : _GEN_6777; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6779 = 10'hda == _T_107[9:0] ? 4'ha : _GEN_6778; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6780 = 10'hdb == _T_107[9:0] ? 4'h9 : _GEN_6779; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6781 = 10'hdc == _T_107[9:0] ? 4'h7 : _GEN_6780; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6782 = 10'hdd == _T_107[9:0] ? 4'hc : _GEN_6781; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6783 = 10'hde == _T_107[9:0] ? 4'hc : _GEN_6782; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6784 = 10'hdf == _T_107[9:0] ? 4'hc : _GEN_6783; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6785 = 10'he0 == _T_107[9:0] ? 4'hc : _GEN_6784; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6786 = 10'he1 == _T_107[9:0] ? 4'hc : _GEN_6785; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6787 = 10'he2 == _T_107[9:0] ? 4'hc : _GEN_6786; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6788 = 10'he3 == _T_107[9:0] ? 4'h8 : _GEN_6787; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6789 = 10'he4 == _T_107[9:0] ? 4'hc : _GEN_6788; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6790 = 10'he5 == _T_107[9:0] ? 4'hc : _GEN_6789; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6791 = 10'he6 == _T_107[9:0] ? 4'hc : _GEN_6790; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6792 = 10'he7 == _T_107[9:0] ? 4'hc : _GEN_6791; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6793 = 10'he8 == _T_107[9:0] ? 4'hc : _GEN_6792; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6794 = 10'he9 == _T_107[9:0] ? 4'hc : _GEN_6793; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6795 = 10'hea == _T_107[9:0] ? 4'hc : _GEN_6794; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6796 = 10'heb == _T_107[9:0] ? 4'ha : _GEN_6795; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6797 = 10'hec == _T_107[9:0] ? 4'h7 : _GEN_6796; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6798 = 10'hed == _T_107[9:0] ? 4'h3 : _GEN_6797; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6799 = 10'hee == _T_107[9:0] ? 4'h3 : _GEN_6798; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6800 = 10'hef == _T_107[9:0] ? 4'h3 : _GEN_6799; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6801 = 10'hf0 == _T_107[9:0] ? 4'h3 : _GEN_6800; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6802 = 10'hf1 == _T_107[9:0] ? 4'h8 : _GEN_6801; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6803 = 10'hf2 == _T_107[9:0] ? 4'hc : _GEN_6802; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6804 = 10'hf3 == _T_107[9:0] ? 4'hc : _GEN_6803; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6805 = 10'hf4 == _T_107[9:0] ? 4'hc : _GEN_6804; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6806 = 10'hf5 == _T_107[9:0] ? 4'h9 : _GEN_6805; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6807 = 10'hf6 == _T_107[9:0] ? 4'h9 : _GEN_6806; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6808 = 10'hf7 == _T_107[9:0] ? 4'h9 : _GEN_6807; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6809 = 10'hf8 == _T_107[9:0] ? 4'h9 : _GEN_6808; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6810 = 10'hf9 == _T_107[9:0] ? 4'ha : _GEN_6809; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6811 = 10'hfa == _T_107[9:0] ? 4'h9 : _GEN_6810; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6812 = 10'hfb == _T_107[9:0] ? 4'h9 : _GEN_6811; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6813 = 10'hfc == _T_107[9:0] ? 4'h9 : _GEN_6812; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6814 = 10'hfd == _T_107[9:0] ? 4'h9 : _GEN_6813; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6815 = 10'hfe == _T_107[9:0] ? 4'h9 : _GEN_6814; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6816 = 10'hff == _T_107[9:0] ? 4'ha : _GEN_6815; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6817 = 10'h100 == _T_107[9:0] ? 4'ha : _GEN_6816; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6818 = 10'h101 == _T_107[9:0] ? 4'h7 : _GEN_6817; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6819 = 10'h102 == _T_107[9:0] ? 4'h9 : _GEN_6818; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6820 = 10'h103 == _T_107[9:0] ? 4'hc : _GEN_6819; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6821 = 10'h104 == _T_107[9:0] ? 4'hc : _GEN_6820; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6822 = 10'h105 == _T_107[9:0] ? 4'hb : _GEN_6821; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6823 = 10'h106 == _T_107[9:0] ? 4'hb : _GEN_6822; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6824 = 10'h107 == _T_107[9:0] ? 4'hb : _GEN_6823; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6825 = 10'h108 == _T_107[9:0] ? 4'hb : _GEN_6824; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6826 = 10'h109 == _T_107[9:0] ? 4'h7 : _GEN_6825; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6827 = 10'h10a == _T_107[9:0] ? 4'hc : _GEN_6826; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6828 = 10'h10b == _T_107[9:0] ? 4'hc : _GEN_6827; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6829 = 10'h10c == _T_107[9:0] ? 4'hc : _GEN_6828; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6830 = 10'h10d == _T_107[9:0] ? 4'hc : _GEN_6829; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6831 = 10'h10e == _T_107[9:0] ? 4'hc : _GEN_6830; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6832 = 10'h10f == _T_107[9:0] ? 4'h9 : _GEN_6831; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6833 = 10'h110 == _T_107[9:0] ? 4'hb : _GEN_6832; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6834 = 10'h111 == _T_107[9:0] ? 4'h4 : _GEN_6833; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6835 = 10'h112 == _T_107[9:0] ? 4'h7 : _GEN_6834; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6836 = 10'h113 == _T_107[9:0] ? 4'h3 : _GEN_6835; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6837 = 10'h114 == _T_107[9:0] ? 4'h3 : _GEN_6836; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6838 = 10'h115 == _T_107[9:0] ? 4'h3 : _GEN_6837; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6839 = 10'h116 == _T_107[9:0] ? 4'h3 : _GEN_6838; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6840 = 10'h117 == _T_107[9:0] ? 4'h2 : _GEN_6839; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6841 = 10'h118 == _T_107[9:0] ? 4'h9 : _GEN_6840; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6842 = 10'h119 == _T_107[9:0] ? 4'hc : _GEN_6841; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6843 = 10'h11a == _T_107[9:0] ? 4'hc : _GEN_6842; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6844 = 10'h11b == _T_107[9:0] ? 4'hc : _GEN_6843; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6845 = 10'h11c == _T_107[9:0] ? 4'h9 : _GEN_6844; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6846 = 10'h11d == _T_107[9:0] ? 4'h9 : _GEN_6845; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6847 = 10'h11e == _T_107[9:0] ? 4'h9 : _GEN_6846; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6848 = 10'h11f == _T_107[9:0] ? 4'h8 : _GEN_6847; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6849 = 10'h120 == _T_107[9:0] ? 4'h7 : _GEN_6848; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6850 = 10'h121 == _T_107[9:0] ? 4'h9 : _GEN_6849; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6851 = 10'h122 == _T_107[9:0] ? 4'h7 : _GEN_6850; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6852 = 10'h123 == _T_107[9:0] ? 4'h7 : _GEN_6851; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6853 = 10'h124 == _T_107[9:0] ? 4'h9 : _GEN_6852; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6854 = 10'h125 == _T_107[9:0] ? 4'h9 : _GEN_6853; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6855 = 10'h126 == _T_107[9:0] ? 4'h8 : _GEN_6854; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6856 = 10'h127 == _T_107[9:0] ? 4'h9 : _GEN_6855; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6857 = 10'h128 == _T_107[9:0] ? 4'h8 : _GEN_6856; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6858 = 10'h129 == _T_107[9:0] ? 4'ha : _GEN_6857; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6859 = 10'h12a == _T_107[9:0] ? 4'h5 : _GEN_6858; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6860 = 10'h12b == _T_107[9:0] ? 4'h3 : _GEN_6859; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6861 = 10'h12c == _T_107[9:0] ? 4'h3 : _GEN_6860; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6862 = 10'h12d == _T_107[9:0] ? 4'h3 : _GEN_6861; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6863 = 10'h12e == _T_107[9:0] ? 4'h5 : _GEN_6862; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6864 = 10'h12f == _T_107[9:0] ? 4'h8 : _GEN_6863; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6865 = 10'h130 == _T_107[9:0] ? 4'hc : _GEN_6864; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6866 = 10'h131 == _T_107[9:0] ? 4'hb : _GEN_6865; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6867 = 10'h132 == _T_107[9:0] ? 4'h9 : _GEN_6866; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6868 = 10'h133 == _T_107[9:0] ? 4'h8 : _GEN_6867; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6869 = 10'h134 == _T_107[9:0] ? 4'h9 : _GEN_6868; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6870 = 10'h135 == _T_107[9:0] ? 4'h7 : _GEN_6869; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6871 = 10'h136 == _T_107[9:0] ? 4'h7 : _GEN_6870; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6872 = 10'h137 == _T_107[9:0] ? 4'h5 : _GEN_6871; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6873 = 10'h138 == _T_107[9:0] ? 4'h7 : _GEN_6872; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6874 = 10'h139 == _T_107[9:0] ? 4'h3 : _GEN_6873; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6875 = 10'h13a == _T_107[9:0] ? 4'h3 : _GEN_6874; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6876 = 10'h13b == _T_107[9:0] ? 4'h3 : _GEN_6875; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6877 = 10'h13c == _T_107[9:0] ? 4'h3 : _GEN_6876; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6878 = 10'h13d == _T_107[9:0] ? 4'h3 : _GEN_6877; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6879 = 10'h13e == _T_107[9:0] ? 4'h5 : _GEN_6878; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6880 = 10'h13f == _T_107[9:0] ? 4'ha : _GEN_6879; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6881 = 10'h140 == _T_107[9:0] ? 4'hc : _GEN_6880; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6882 = 10'h141 == _T_107[9:0] ? 4'hc : _GEN_6881; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6883 = 10'h142 == _T_107[9:0] ? 4'hc : _GEN_6882; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6884 = 10'h143 == _T_107[9:0] ? 4'h9 : _GEN_6883; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6885 = 10'h144 == _T_107[9:0] ? 4'h9 : _GEN_6884; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6886 = 10'h145 == _T_107[9:0] ? 4'h8 : _GEN_6885; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6887 = 10'h146 == _T_107[9:0] ? 4'h8 : _GEN_6886; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6888 = 10'h147 == _T_107[9:0] ? 4'h7 : _GEN_6887; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6889 = 10'h148 == _T_107[9:0] ? 4'h8 : _GEN_6888; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6890 = 10'h149 == _T_107[9:0] ? 4'h9 : _GEN_6889; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6891 = 10'h14a == _T_107[9:0] ? 4'ha : _GEN_6890; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6892 = 10'h14b == _T_107[9:0] ? 4'h9 : _GEN_6891; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6893 = 10'h14c == _T_107[9:0] ? 4'ha : _GEN_6892; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6894 = 10'h14d == _T_107[9:0] ? 4'h9 : _GEN_6893; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6895 = 10'h14e == _T_107[9:0] ? 4'h7 : _GEN_6894; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6896 = 10'h14f == _T_107[9:0] ? 4'h3 : _GEN_6895; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6897 = 10'h150 == _T_107[9:0] ? 4'h3 : _GEN_6896; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6898 = 10'h151 == _T_107[9:0] ? 4'h3 : _GEN_6897; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6899 = 10'h152 == _T_107[9:0] ? 4'h3 : _GEN_6898; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6900 = 10'h153 == _T_107[9:0] ? 4'h3 : _GEN_6899; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6901 = 10'h154 == _T_107[9:0] ? 4'h3 : _GEN_6900; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6902 = 10'h155 == _T_107[9:0] ? 4'h8 : _GEN_6901; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6903 = 10'h156 == _T_107[9:0] ? 4'ha : _GEN_6902; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6904 = 10'h157 == _T_107[9:0] ? 4'h7 : _GEN_6903; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6905 = 10'h158 == _T_107[9:0] ? 4'h7 : _GEN_6904; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6906 = 10'h159 == _T_107[9:0] ? 4'h7 : _GEN_6905; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6907 = 10'h15a == _T_107[9:0] ? 4'h7 : _GEN_6906; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6908 = 10'h15b == _T_107[9:0] ? 4'h7 : _GEN_6907; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6909 = 10'h15c == _T_107[9:0] ? 4'h7 : _GEN_6908; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6910 = 10'h15d == _T_107[9:0] ? 4'h7 : _GEN_6909; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6911 = 10'h15e == _T_107[9:0] ? 4'h7 : _GEN_6910; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6912 = 10'h15f == _T_107[9:0] ? 4'h3 : _GEN_6911; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6913 = 10'h160 == _T_107[9:0] ? 4'h3 : _GEN_6912; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6914 = 10'h161 == _T_107[9:0] ? 4'h3 : _GEN_6913; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6915 = 10'h162 == _T_107[9:0] ? 4'h3 : _GEN_6914; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6916 = 10'h163 == _T_107[9:0] ? 4'h3 : _GEN_6915; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6917 = 10'h164 == _T_107[9:0] ? 4'h4 : _GEN_6916; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6918 = 10'h165 == _T_107[9:0] ? 4'ha : _GEN_6917; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6919 = 10'h166 == _T_107[9:0] ? 4'ha : _GEN_6918; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6920 = 10'h167 == _T_107[9:0] ? 4'hc : _GEN_6919; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6921 = 10'h168 == _T_107[9:0] ? 4'hc : _GEN_6920; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6922 = 10'h169 == _T_107[9:0] ? 4'h9 : _GEN_6921; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6923 = 10'h16a == _T_107[9:0] ? 4'h9 : _GEN_6922; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6924 = 10'h16b == _T_107[9:0] ? 4'ha : _GEN_6923; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6925 = 10'h16c == _T_107[9:0] ? 4'h7 : _GEN_6924; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6926 = 10'h16d == _T_107[9:0] ? 4'h7 : _GEN_6925; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6927 = 10'h16e == _T_107[9:0] ? 4'h7 : _GEN_6926; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6928 = 10'h16f == _T_107[9:0] ? 4'ha : _GEN_6927; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6929 = 10'h170 == _T_107[9:0] ? 4'ha : _GEN_6928; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6930 = 10'h171 == _T_107[9:0] ? 4'ha : _GEN_6929; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6931 = 10'h172 == _T_107[9:0] ? 4'hc : _GEN_6930; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6932 = 10'h173 == _T_107[9:0] ? 4'h8 : _GEN_6931; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6933 = 10'h174 == _T_107[9:0] ? 4'h5 : _GEN_6932; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6934 = 10'h175 == _T_107[9:0] ? 4'h8 : _GEN_6933; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6935 = 10'h176 == _T_107[9:0] ? 4'h7 : _GEN_6934; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6936 = 10'h177 == _T_107[9:0] ? 4'h8 : _GEN_6935; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6937 = 10'h178 == _T_107[9:0] ? 4'h7 : _GEN_6936; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6938 = 10'h179 == _T_107[9:0] ? 4'h5 : _GEN_6937; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6939 = 10'h17a == _T_107[9:0] ? 4'h5 : _GEN_6938; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6940 = 10'h17b == _T_107[9:0] ? 4'h7 : _GEN_6939; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6941 = 10'h17c == _T_107[9:0] ? 4'h7 : _GEN_6940; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6942 = 10'h17d == _T_107[9:0] ? 4'h7 : _GEN_6941; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6943 = 10'h17e == _T_107[9:0] ? 4'h7 : _GEN_6942; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6944 = 10'h17f == _T_107[9:0] ? 4'h7 : _GEN_6943; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6945 = 10'h180 == _T_107[9:0] ? 4'h7 : _GEN_6944; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6946 = 10'h181 == _T_107[9:0] ? 4'h7 : _GEN_6945; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6947 = 10'h182 == _T_107[9:0] ? 4'h7 : _GEN_6946; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6948 = 10'h183 == _T_107[9:0] ? 4'h7 : _GEN_6947; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6949 = 10'h184 == _T_107[9:0] ? 4'h7 : _GEN_6948; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6950 = 10'h185 == _T_107[9:0] ? 4'h5 : _GEN_6949; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6951 = 10'h186 == _T_107[9:0] ? 4'h3 : _GEN_6950; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6952 = 10'h187 == _T_107[9:0] ? 4'h3 : _GEN_6951; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6953 = 10'h188 == _T_107[9:0] ? 4'h3 : _GEN_6952; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6954 = 10'h189 == _T_107[9:0] ? 4'h4 : _GEN_6953; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6955 = 10'h18a == _T_107[9:0] ? 4'h5 : _GEN_6954; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6956 = 10'h18b == _T_107[9:0] ? 4'ha : _GEN_6955; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6957 = 10'h18c == _T_107[9:0] ? 4'ha : _GEN_6956; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6958 = 10'h18d == _T_107[9:0] ? 4'ha : _GEN_6957; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6959 = 10'h18e == _T_107[9:0] ? 4'hc : _GEN_6958; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6960 = 10'h18f == _T_107[9:0] ? 4'h8 : _GEN_6959; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6961 = 10'h190 == _T_107[9:0] ? 4'h9 : _GEN_6960; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6962 = 10'h191 == _T_107[9:0] ? 4'h8 : _GEN_6961; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6963 = 10'h192 == _T_107[9:0] ? 4'h7 : _GEN_6962; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6964 = 10'h193 == _T_107[9:0] ? 4'h7 : _GEN_6963; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6965 = 10'h194 == _T_107[9:0] ? 4'h7 : _GEN_6964; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6966 = 10'h195 == _T_107[9:0] ? 4'h9 : _GEN_6965; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6967 = 10'h196 == _T_107[9:0] ? 4'ha : _GEN_6966; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6968 = 10'h197 == _T_107[9:0] ? 4'h8 : _GEN_6967; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6969 = 10'h198 == _T_107[9:0] ? 4'hc : _GEN_6968; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6970 = 10'h199 == _T_107[9:0] ? 4'h5 : _GEN_6969; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6971 = 10'h19a == _T_107[9:0] ? 4'h1 : _GEN_6970; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6972 = 10'h19b == _T_107[9:0] ? 4'h4 : _GEN_6971; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6973 = 10'h19c == _T_107[9:0] ? 4'h7 : _GEN_6972; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6974 = 10'h19d == _T_107[9:0] ? 4'h5 : _GEN_6973; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6975 = 10'h19e == _T_107[9:0] ? 4'h2 : _GEN_6974; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6976 = 10'h19f == _T_107[9:0] ? 4'h3 : _GEN_6975; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6977 = 10'h1a0 == _T_107[9:0] ? 4'h7 : _GEN_6976; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6978 = 10'h1a1 == _T_107[9:0] ? 4'h7 : _GEN_6977; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6979 = 10'h1a2 == _T_107[9:0] ? 4'h7 : _GEN_6978; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6980 = 10'h1a3 == _T_107[9:0] ? 4'h7 : _GEN_6979; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6981 = 10'h1a4 == _T_107[9:0] ? 4'h7 : _GEN_6980; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6982 = 10'h1a5 == _T_107[9:0] ? 4'h7 : _GEN_6981; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6983 = 10'h1a6 == _T_107[9:0] ? 4'h7 : _GEN_6982; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6984 = 10'h1a7 == _T_107[9:0] ? 4'h7 : _GEN_6983; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6985 = 10'h1a8 == _T_107[9:0] ? 4'h8 : _GEN_6984; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6986 = 10'h1a9 == _T_107[9:0] ? 4'h8 : _GEN_6985; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6987 = 10'h1aa == _T_107[9:0] ? 4'h6 : _GEN_6986; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6988 = 10'h1ab == _T_107[9:0] ? 4'h6 : _GEN_6987; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6989 = 10'h1ac == _T_107[9:0] ? 4'h5 : _GEN_6988; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6990 = 10'h1ad == _T_107[9:0] ? 4'h4 : _GEN_6989; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6991 = 10'h1ae == _T_107[9:0] ? 4'h3 : _GEN_6990; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6992 = 10'h1af == _T_107[9:0] ? 4'h6 : _GEN_6991; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6993 = 10'h1b0 == _T_107[9:0] ? 4'h6 : _GEN_6992; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6994 = 10'h1b1 == _T_107[9:0] ? 4'ha : _GEN_6993; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6995 = 10'h1b2 == _T_107[9:0] ? 4'ha : _GEN_6994; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6996 = 10'h1b3 == _T_107[9:0] ? 4'h9 : _GEN_6995; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6997 = 10'h1b4 == _T_107[9:0] ? 4'hb : _GEN_6996; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6998 = 10'h1b5 == _T_107[9:0] ? 4'h8 : _GEN_6997; // @[Filter.scala 230:142]
  wire [3:0] _GEN_6999 = 10'h1b6 == _T_107[9:0] ? 4'h8 : _GEN_6998; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7000 = 10'h1b7 == _T_107[9:0] ? 4'h7 : _GEN_6999; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7001 = 10'h1b8 == _T_107[9:0] ? 4'h6 : _GEN_7000; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7002 = 10'h1b9 == _T_107[9:0] ? 4'h7 : _GEN_7001; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7003 = 10'h1ba == _T_107[9:0] ? 4'h6 : _GEN_7002; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7004 = 10'h1bb == _T_107[9:0] ? 4'h8 : _GEN_7003; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7005 = 10'h1bc == _T_107[9:0] ? 4'ha : _GEN_7004; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7006 = 10'h1bd == _T_107[9:0] ? 4'h9 : _GEN_7005; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7007 = 10'h1be == _T_107[9:0] ? 4'hc : _GEN_7006; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7008 = 10'h1bf == _T_107[9:0] ? 4'h7 : _GEN_7007; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7009 = 10'h1c0 == _T_107[9:0] ? 4'h6 : _GEN_7008; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7010 = 10'h1c1 == _T_107[9:0] ? 4'h7 : _GEN_7009; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7011 = 10'h1c2 == _T_107[9:0] ? 4'h7 : _GEN_7010; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7012 = 10'h1c3 == _T_107[9:0] ? 4'h6 : _GEN_7011; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7013 = 10'h1c4 == _T_107[9:0] ? 4'h5 : _GEN_7012; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7014 = 10'h1c5 == _T_107[9:0] ? 4'h6 : _GEN_7013; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7015 = 10'h1c6 == _T_107[9:0] ? 4'h8 : _GEN_7014; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7016 = 10'h1c7 == _T_107[9:0] ? 4'h7 : _GEN_7015; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7017 = 10'h1c8 == _T_107[9:0] ? 4'h7 : _GEN_7016; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7018 = 10'h1c9 == _T_107[9:0] ? 4'h7 : _GEN_7017; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7019 = 10'h1ca == _T_107[9:0] ? 4'h7 : _GEN_7018; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7020 = 10'h1cb == _T_107[9:0] ? 4'h7 : _GEN_7019; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7021 = 10'h1cc == _T_107[9:0] ? 4'h7 : _GEN_7020; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7022 = 10'h1cd == _T_107[9:0] ? 4'h8 : _GEN_7021; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7023 = 10'h1ce == _T_107[9:0] ? 4'h8 : _GEN_7022; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7024 = 10'h1cf == _T_107[9:0] ? 4'h8 : _GEN_7023; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7025 = 10'h1d0 == _T_107[9:0] ? 4'h5 : _GEN_7024; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7026 = 10'h1d1 == _T_107[9:0] ? 4'h6 : _GEN_7025; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7027 = 10'h1d2 == _T_107[9:0] ? 4'h7 : _GEN_7026; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7028 = 10'h1d3 == _T_107[9:0] ? 4'h7 : _GEN_7027; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7029 = 10'h1d4 == _T_107[9:0] ? 4'h7 : _GEN_7028; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7030 = 10'h1d5 == _T_107[9:0] ? 4'h6 : _GEN_7029; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7031 = 10'h1d6 == _T_107[9:0] ? 4'h8 : _GEN_7030; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7032 = 10'h1d7 == _T_107[9:0] ? 4'ha : _GEN_7031; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7033 = 10'h1d8 == _T_107[9:0] ? 4'ha : _GEN_7032; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7034 = 10'h1d9 == _T_107[9:0] ? 4'ha : _GEN_7033; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7035 = 10'h1da == _T_107[9:0] ? 4'h8 : _GEN_7034; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7036 = 10'h1db == _T_107[9:0] ? 4'h9 : _GEN_7035; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7037 = 10'h1dc == _T_107[9:0] ? 4'h9 : _GEN_7036; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7038 = 10'h1dd == _T_107[9:0] ? 4'h5 : _GEN_7037; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7039 = 10'h1de == _T_107[9:0] ? 4'h7 : _GEN_7038; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7040 = 10'h1df == _T_107[9:0] ? 4'h7 : _GEN_7039; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7041 = 10'h1e0 == _T_107[9:0] ? 4'h7 : _GEN_7040; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7042 = 10'h1e1 == _T_107[9:0] ? 4'h6 : _GEN_7041; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7043 = 10'h1e2 == _T_107[9:0] ? 4'h9 : _GEN_7042; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7044 = 10'h1e3 == _T_107[9:0] ? 4'h9 : _GEN_7043; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7045 = 10'h1e4 == _T_107[9:0] ? 4'hb : _GEN_7044; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7046 = 10'h1e5 == _T_107[9:0] ? 4'h8 : _GEN_7045; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7047 = 10'h1e6 == _T_107[9:0] ? 4'h7 : _GEN_7046; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7048 = 10'h1e7 == _T_107[9:0] ? 4'h8 : _GEN_7047; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7049 = 10'h1e8 == _T_107[9:0] ? 4'h8 : _GEN_7048; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7050 = 10'h1e9 == _T_107[9:0] ? 4'h8 : _GEN_7049; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7051 = 10'h1ea == _T_107[9:0] ? 4'h8 : _GEN_7050; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7052 = 10'h1eb == _T_107[9:0] ? 4'h8 : _GEN_7051; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7053 = 10'h1ec == _T_107[9:0] ? 4'h8 : _GEN_7052; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7054 = 10'h1ed == _T_107[9:0] ? 4'h6 : _GEN_7053; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7055 = 10'h1ee == _T_107[9:0] ? 4'h7 : _GEN_7054; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7056 = 10'h1ef == _T_107[9:0] ? 4'h7 : _GEN_7055; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7057 = 10'h1f0 == _T_107[9:0] ? 4'h7 : _GEN_7056; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7058 = 10'h1f1 == _T_107[9:0] ? 4'h7 : _GEN_7057; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7059 = 10'h1f2 == _T_107[9:0] ? 4'h7 : _GEN_7058; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7060 = 10'h1f3 == _T_107[9:0] ? 4'h8 : _GEN_7059; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7061 = 10'h1f4 == _T_107[9:0] ? 4'h8 : _GEN_7060; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7062 = 10'h1f5 == _T_107[9:0] ? 4'h8 : _GEN_7061; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7063 = 10'h1f6 == _T_107[9:0] ? 4'ha : _GEN_7062; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7064 = 10'h1f7 == _T_107[9:0] ? 4'h6 : _GEN_7063; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7065 = 10'h1f8 == _T_107[9:0] ? 4'h6 : _GEN_7064; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7066 = 10'h1f9 == _T_107[9:0] ? 4'h8 : _GEN_7065; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7067 = 10'h1fa == _T_107[9:0] ? 4'h8 : _GEN_7066; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7068 = 10'h1fb == _T_107[9:0] ? 4'h6 : _GEN_7067; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7069 = 10'h1fc == _T_107[9:0] ? 4'ha : _GEN_7068; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7070 = 10'h1fd == _T_107[9:0] ? 4'hb : _GEN_7069; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7071 = 10'h1fe == _T_107[9:0] ? 4'ha : _GEN_7070; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7072 = 10'h1ff == _T_107[9:0] ? 4'ha : _GEN_7071; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7073 = 10'h200 == _T_107[9:0] ? 4'h4 : _GEN_7072; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7074 = 10'h201 == _T_107[9:0] ? 4'h7 : _GEN_7073; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7075 = 10'h202 == _T_107[9:0] ? 4'h6 : _GEN_7074; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7076 = 10'h203 == _T_107[9:0] ? 4'h6 : _GEN_7075; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7077 = 10'h204 == _T_107[9:0] ? 4'h5 : _GEN_7076; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7078 = 10'h205 == _T_107[9:0] ? 4'h6 : _GEN_7077; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7079 = 10'h206 == _T_107[9:0] ? 4'h6 : _GEN_7078; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7080 = 10'h207 == _T_107[9:0] ? 4'h5 : _GEN_7079; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7081 = 10'h208 == _T_107[9:0] ? 4'h7 : _GEN_7080; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7082 = 10'h209 == _T_107[9:0] ? 4'h9 : _GEN_7081; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7083 = 10'h20a == _T_107[9:0] ? 4'hb : _GEN_7082; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7084 = 10'h20b == _T_107[9:0] ? 4'h7 : _GEN_7083; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7085 = 10'h20c == _T_107[9:0] ? 4'h7 : _GEN_7084; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7086 = 10'h20d == _T_107[9:0] ? 4'h7 : _GEN_7085; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7087 = 10'h20e == _T_107[9:0] ? 4'h7 : _GEN_7086; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7088 = 10'h20f == _T_107[9:0] ? 4'h7 : _GEN_7087; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7089 = 10'h210 == _T_107[9:0] ? 4'h7 : _GEN_7088; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7090 = 10'h211 == _T_107[9:0] ? 4'h8 : _GEN_7089; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7091 = 10'h212 == _T_107[9:0] ? 4'h8 : _GEN_7090; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7092 = 10'h213 == _T_107[9:0] ? 4'h9 : _GEN_7091; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7093 = 10'h214 == _T_107[9:0] ? 4'h6 : _GEN_7092; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7094 = 10'h215 == _T_107[9:0] ? 4'h7 : _GEN_7093; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7095 = 10'h216 == _T_107[9:0] ? 4'h7 : _GEN_7094; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7096 = 10'h217 == _T_107[9:0] ? 4'h7 : _GEN_7095; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7097 = 10'h218 == _T_107[9:0] ? 4'h7 : _GEN_7096; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7098 = 10'h219 == _T_107[9:0] ? 4'h8 : _GEN_7097; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7099 = 10'h21a == _T_107[9:0] ? 4'h7 : _GEN_7098; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7100 = 10'h21b == _T_107[9:0] ? 4'h8 : _GEN_7099; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7101 = 10'h21c == _T_107[9:0] ? 4'ha : _GEN_7100; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7102 = 10'h21d == _T_107[9:0] ? 4'ha : _GEN_7101; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7103 = 10'h21e == _T_107[9:0] ? 4'h7 : _GEN_7102; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7104 = 10'h21f == _T_107[9:0] ? 4'h6 : _GEN_7103; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7105 = 10'h220 == _T_107[9:0] ? 4'h6 : _GEN_7104; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7106 = 10'h221 == _T_107[9:0] ? 4'h7 : _GEN_7105; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7107 = 10'h222 == _T_107[9:0] ? 4'ha : _GEN_7106; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7108 = 10'h223 == _T_107[9:0] ? 4'ha : _GEN_7107; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7109 = 10'h224 == _T_107[9:0] ? 4'ha : _GEN_7108; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7110 = 10'h225 == _T_107[9:0] ? 4'h8 : _GEN_7109; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7111 = 10'h226 == _T_107[9:0] ? 4'h3 : _GEN_7110; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7112 = 10'h227 == _T_107[9:0] ? 4'h4 : _GEN_7111; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7113 = 10'h228 == _T_107[9:0] ? 4'h6 : _GEN_7112; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7114 = 10'h229 == _T_107[9:0] ? 4'h6 : _GEN_7113; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7115 = 10'h22a == _T_107[9:0] ? 4'h6 : _GEN_7114; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7116 = 10'h22b == _T_107[9:0] ? 4'h6 : _GEN_7115; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7117 = 10'h22c == _T_107[9:0] ? 4'h5 : _GEN_7116; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7118 = 10'h22d == _T_107[9:0] ? 4'h6 : _GEN_7117; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7119 = 10'h22e == _T_107[9:0] ? 4'h6 : _GEN_7118; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7120 = 10'h22f == _T_107[9:0] ? 4'h8 : _GEN_7119; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7121 = 10'h230 == _T_107[9:0] ? 4'h7 : _GEN_7120; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7122 = 10'h231 == _T_107[9:0] ? 4'h5 : _GEN_7121; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7123 = 10'h232 == _T_107[9:0] ? 4'h6 : _GEN_7122; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7124 = 10'h233 == _T_107[9:0] ? 4'h8 : _GEN_7123; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7125 = 10'h234 == _T_107[9:0] ? 4'h8 : _GEN_7124; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7126 = 10'h235 == _T_107[9:0] ? 4'h8 : _GEN_7125; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7127 = 10'h236 == _T_107[9:0] ? 4'h8 : _GEN_7126; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7128 = 10'h237 == _T_107[9:0] ? 4'h8 : _GEN_7127; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7129 = 10'h238 == _T_107[9:0] ? 4'h8 : _GEN_7128; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7130 = 10'h239 == _T_107[9:0] ? 4'h6 : _GEN_7129; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7131 = 10'h23a == _T_107[9:0] ? 4'h6 : _GEN_7130; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7132 = 10'h23b == _T_107[9:0] ? 4'h7 : _GEN_7131; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7133 = 10'h23c == _T_107[9:0] ? 4'h6 : _GEN_7132; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7134 = 10'h23d == _T_107[9:0] ? 4'h7 : _GEN_7133; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7135 = 10'h23e == _T_107[9:0] ? 4'h7 : _GEN_7134; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7136 = 10'h23f == _T_107[9:0] ? 4'h6 : _GEN_7135; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7137 = 10'h240 == _T_107[9:0] ? 4'h6 : _GEN_7136; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7138 = 10'h241 == _T_107[9:0] ? 4'h8 : _GEN_7137; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7139 = 10'h242 == _T_107[9:0] ? 4'ha : _GEN_7138; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7140 = 10'h243 == _T_107[9:0] ? 4'ha : _GEN_7139; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7141 = 10'h244 == _T_107[9:0] ? 4'ha : _GEN_7140; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7142 = 10'h245 == _T_107[9:0] ? 4'h8 : _GEN_7141; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7143 = 10'h246 == _T_107[9:0] ? 4'h8 : _GEN_7142; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7144 = 10'h247 == _T_107[9:0] ? 4'h9 : _GEN_7143; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7145 = 10'h248 == _T_107[9:0] ? 4'ha : _GEN_7144; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7146 = 10'h249 == _T_107[9:0] ? 4'ha : _GEN_7145; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7147 = 10'h24a == _T_107[9:0] ? 4'ha : _GEN_7146; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7148 = 10'h24b == _T_107[9:0] ? 4'h4 : _GEN_7147; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7149 = 10'h24c == _T_107[9:0] ? 4'h3 : _GEN_7148; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7150 = 10'h24d == _T_107[9:0] ? 4'h4 : _GEN_7149; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7151 = 10'h24e == _T_107[9:0] ? 4'h5 : _GEN_7150; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7152 = 10'h24f == _T_107[9:0] ? 4'h5 : _GEN_7151; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7153 = 10'h250 == _T_107[9:0] ? 4'h5 : _GEN_7152; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7154 = 10'h251 == _T_107[9:0] ? 4'h5 : _GEN_7153; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7155 = 10'h252 == _T_107[9:0] ? 4'h5 : _GEN_7154; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7156 = 10'h253 == _T_107[9:0] ? 4'h5 : _GEN_7155; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7157 = 10'h254 == _T_107[9:0] ? 4'h5 : _GEN_7156; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7158 = 10'h255 == _T_107[9:0] ? 4'h6 : _GEN_7157; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7159 = 10'h256 == _T_107[9:0] ? 4'h7 : _GEN_7158; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7160 = 10'h257 == _T_107[9:0] ? 4'h3 : _GEN_7159; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7161 = 10'h258 == _T_107[9:0] ? 4'h6 : _GEN_7160; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7162 = 10'h259 == _T_107[9:0] ? 4'h7 : _GEN_7161; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7163 = 10'h25a == _T_107[9:0] ? 4'h7 : _GEN_7162; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7164 = 10'h25b == _T_107[9:0] ? 4'h7 : _GEN_7163; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7165 = 10'h25c == _T_107[9:0] ? 4'h8 : _GEN_7164; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7166 = 10'h25d == _T_107[9:0] ? 4'h8 : _GEN_7165; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7167 = 10'h25e == _T_107[9:0] ? 4'h4 : _GEN_7166; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7168 = 10'h25f == _T_107[9:0] ? 4'h3 : _GEN_7167; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7169 = 10'h260 == _T_107[9:0] ? 4'h7 : _GEN_7168; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7170 = 10'h261 == _T_107[9:0] ? 4'h7 : _GEN_7169; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7171 = 10'h262 == _T_107[9:0] ? 4'h7 : _GEN_7170; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7172 = 10'h263 == _T_107[9:0] ? 4'h6 : _GEN_7171; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7173 = 10'h264 == _T_107[9:0] ? 4'h7 : _GEN_7172; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7174 = 10'h265 == _T_107[9:0] ? 4'h6 : _GEN_7173; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7175 = 10'h266 == _T_107[9:0] ? 4'h5 : _GEN_7174; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7176 = 10'h267 == _T_107[9:0] ? 4'h7 : _GEN_7175; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7177 = 10'h268 == _T_107[9:0] ? 4'ha : _GEN_7176; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7178 = 10'h269 == _T_107[9:0] ? 4'ha : _GEN_7177; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7179 = 10'h26a == _T_107[9:0] ? 4'ha : _GEN_7178; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7180 = 10'h26b == _T_107[9:0] ? 4'ha : _GEN_7179; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7181 = 10'h26c == _T_107[9:0] ? 4'ha : _GEN_7180; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7182 = 10'h26d == _T_107[9:0] ? 4'ha : _GEN_7181; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7183 = 10'h26e == _T_107[9:0] ? 4'ha : _GEN_7182; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7184 = 10'h26f == _T_107[9:0] ? 4'ha : _GEN_7183; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7185 = 10'h270 == _T_107[9:0] ? 4'h5 : _GEN_7184; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7186 = 10'h271 == _T_107[9:0] ? 4'h3 : _GEN_7185; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7187 = 10'h272 == _T_107[9:0] ? 4'h3 : _GEN_7186; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7188 = 10'h273 == _T_107[9:0] ? 4'h4 : _GEN_7187; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7189 = 10'h274 == _T_107[9:0] ? 4'h6 : _GEN_7188; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7190 = 10'h275 == _T_107[9:0] ? 4'h5 : _GEN_7189; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7191 = 10'h276 == _T_107[9:0] ? 4'h6 : _GEN_7190; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7192 = 10'h277 == _T_107[9:0] ? 4'h5 : _GEN_7191; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7193 = 10'h278 == _T_107[9:0] ? 4'h6 : _GEN_7192; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7194 = 10'h279 == _T_107[9:0] ? 4'h6 : _GEN_7193; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7195 = 10'h27a == _T_107[9:0] ? 4'h6 : _GEN_7194; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7196 = 10'h27b == _T_107[9:0] ? 4'h8 : _GEN_7195; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7197 = 10'h27c == _T_107[9:0] ? 4'h6 : _GEN_7196; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7198 = 10'h27d == _T_107[9:0] ? 4'h2 : _GEN_7197; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7199 = 10'h27e == _T_107[9:0] ? 4'h5 : _GEN_7198; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7200 = 10'h27f == _T_107[9:0] ? 4'h7 : _GEN_7199; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7201 = 10'h280 == _T_107[9:0] ? 4'h7 : _GEN_7200; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7202 = 10'h281 == _T_107[9:0] ? 4'h8 : _GEN_7201; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7203 = 10'h282 == _T_107[9:0] ? 4'h7 : _GEN_7202; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7204 = 10'h283 == _T_107[9:0] ? 4'h3 : _GEN_7203; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7205 = 10'h284 == _T_107[9:0] ? 4'h3 : _GEN_7204; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7206 = 10'h285 == _T_107[9:0] ? 4'h3 : _GEN_7205; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7207 = 10'h286 == _T_107[9:0] ? 4'h7 : _GEN_7206; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7208 = 10'h287 == _T_107[9:0] ? 4'h7 : _GEN_7207; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7209 = 10'h288 == _T_107[9:0] ? 4'h7 : _GEN_7208; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7210 = 10'h289 == _T_107[9:0] ? 4'h7 : _GEN_7209; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7211 = 10'h28a == _T_107[9:0] ? 4'h8 : _GEN_7210; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7212 = 10'h28b == _T_107[9:0] ? 4'h8 : _GEN_7211; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7213 = 10'h28c == _T_107[9:0] ? 4'h7 : _GEN_7212; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7214 = 10'h28d == _T_107[9:0] ? 4'h6 : _GEN_7213; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7215 = 10'h28e == _T_107[9:0] ? 4'h3 : _GEN_7214; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7216 = 10'h28f == _T_107[9:0] ? 4'h6 : _GEN_7215; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7217 = 10'h290 == _T_107[9:0] ? 4'h8 : _GEN_7216; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7218 = 10'h291 == _T_107[9:0] ? 4'ha : _GEN_7217; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7219 = 10'h292 == _T_107[9:0] ? 4'ha : _GEN_7218; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7220 = 10'h293 == _T_107[9:0] ? 4'ha : _GEN_7219; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7221 = 10'h294 == _T_107[9:0] ? 4'h9 : _GEN_7220; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7222 = 10'h295 == _T_107[9:0] ? 4'h4 : _GEN_7221; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7223 = 10'h296 == _T_107[9:0] ? 4'h3 : _GEN_7222; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7224 = 10'h297 == _T_107[9:0] ? 4'h3 : _GEN_7223; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7225 = 10'h298 == _T_107[9:0] ? 4'h3 : _GEN_7224; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7226 = 10'h299 == _T_107[9:0] ? 4'h4 : _GEN_7225; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7227 = 10'h29a == _T_107[9:0] ? 4'h5 : _GEN_7226; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7228 = 10'h29b == _T_107[9:0] ? 4'h5 : _GEN_7227; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7229 = 10'h29c == _T_107[9:0] ? 4'h5 : _GEN_7228; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7230 = 10'h29d == _T_107[9:0] ? 4'h5 : _GEN_7229; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7231 = 10'h29e == _T_107[9:0] ? 4'h5 : _GEN_7230; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7232 = 10'h29f == _T_107[9:0] ? 4'h5 : _GEN_7231; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7233 = 10'h2a0 == _T_107[9:0] ? 4'h6 : _GEN_7232; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7234 = 10'h2a1 == _T_107[9:0] ? 4'h7 : _GEN_7233; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7235 = 10'h2a2 == _T_107[9:0] ? 4'h5 : _GEN_7234; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7236 = 10'h2a3 == _T_107[9:0] ? 4'h2 : _GEN_7235; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7237 = 10'h2a4 == _T_107[9:0] ? 4'h3 : _GEN_7236; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7238 = 10'h2a5 == _T_107[9:0] ? 4'h7 : _GEN_7237; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7239 = 10'h2a6 == _T_107[9:0] ? 4'h8 : _GEN_7238; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7240 = 10'h2a7 == _T_107[9:0] ? 4'h7 : _GEN_7239; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7241 = 10'h2a8 == _T_107[9:0] ? 4'h3 : _GEN_7240; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7242 = 10'h2a9 == _T_107[9:0] ? 4'h2 : _GEN_7241; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7243 = 10'h2aa == _T_107[9:0] ? 4'h3 : _GEN_7242; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7244 = 10'h2ab == _T_107[9:0] ? 4'h3 : _GEN_7243; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7245 = 10'h2ac == _T_107[9:0] ? 4'h7 : _GEN_7244; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7246 = 10'h2ad == _T_107[9:0] ? 4'h8 : _GEN_7245; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7247 = 10'h2ae == _T_107[9:0] ? 4'h7 : _GEN_7246; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7248 = 10'h2af == _T_107[9:0] ? 4'h8 : _GEN_7247; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7249 = 10'h2b0 == _T_107[9:0] ? 4'h8 : _GEN_7248; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7250 = 10'h2b1 == _T_107[9:0] ? 4'h8 : _GEN_7249; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7251 = 10'h2b2 == _T_107[9:0] ? 4'h7 : _GEN_7250; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7252 = 10'h2b3 == _T_107[9:0] ? 4'h6 : _GEN_7251; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7253 = 10'h2b4 == _T_107[9:0] ? 4'h2 : _GEN_7252; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7254 = 10'h2b5 == _T_107[9:0] ? 4'h2 : _GEN_7253; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7255 = 10'h2b6 == _T_107[9:0] ? 4'h3 : _GEN_7254; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7256 = 10'h2b7 == _T_107[9:0] ? 4'h3 : _GEN_7255; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7257 = 10'h2b8 == _T_107[9:0] ? 4'h6 : _GEN_7256; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7258 = 10'h2b9 == _T_107[9:0] ? 4'h9 : _GEN_7257; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7259 = 10'h2ba == _T_107[9:0] ? 4'h3 : _GEN_7258; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7260 = 10'h2bb == _T_107[9:0] ? 4'h3 : _GEN_7259; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7261 = 10'h2bc == _T_107[9:0] ? 4'h3 : _GEN_7260; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7262 = 10'h2bd == _T_107[9:0] ? 4'h2 : _GEN_7261; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7263 = 10'h2be == _T_107[9:0] ? 4'h3 : _GEN_7262; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7264 = 10'h2bf == _T_107[9:0] ? 4'h3 : _GEN_7263; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7265 = 10'h2c0 == _T_107[9:0] ? 4'h5 : _GEN_7264; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7266 = 10'h2c1 == _T_107[9:0] ? 4'h5 : _GEN_7265; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7267 = 10'h2c2 == _T_107[9:0] ? 4'h5 : _GEN_7266; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7268 = 10'h2c3 == _T_107[9:0] ? 4'h5 : _GEN_7267; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7269 = 10'h2c4 == _T_107[9:0] ? 4'h5 : _GEN_7268; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7270 = 10'h2c5 == _T_107[9:0] ? 4'h5 : _GEN_7269; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7271 = 10'h2c6 == _T_107[9:0] ? 4'h6 : _GEN_7270; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7272 = 10'h2c7 == _T_107[9:0] ? 4'h7 : _GEN_7271; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7273 = 10'h2c8 == _T_107[9:0] ? 4'h5 : _GEN_7272; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7274 = 10'h2c9 == _T_107[9:0] ? 4'h2 : _GEN_7273; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7275 = 10'h2ca == _T_107[9:0] ? 4'h2 : _GEN_7274; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7276 = 10'h2cb == _T_107[9:0] ? 4'h3 : _GEN_7275; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7277 = 10'h2cc == _T_107[9:0] ? 4'h3 : _GEN_7276; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7278 = 10'h2cd == _T_107[9:0] ? 4'h2 : _GEN_7277; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7279 = 10'h2ce == _T_107[9:0] ? 4'h2 : _GEN_7278; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7280 = 10'h2cf == _T_107[9:0] ? 4'h2 : _GEN_7279; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7281 = 10'h2d0 == _T_107[9:0] ? 4'h2 : _GEN_7280; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7282 = 10'h2d1 == _T_107[9:0] ? 4'h2 : _GEN_7281; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7283 = 10'h2d2 == _T_107[9:0] ? 4'h7 : _GEN_7282; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7284 = 10'h2d3 == _T_107[9:0] ? 4'h7 : _GEN_7283; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7285 = 10'h2d4 == _T_107[9:0] ? 4'h8 : _GEN_7284; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7286 = 10'h2d5 == _T_107[9:0] ? 4'h8 : _GEN_7285; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7287 = 10'h2d6 == _T_107[9:0] ? 4'h8 : _GEN_7286; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7288 = 10'h2d7 == _T_107[9:0] ? 4'h8 : _GEN_7287; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7289 = 10'h2d8 == _T_107[9:0] ? 4'h7 : _GEN_7288; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7290 = 10'h2d9 == _T_107[9:0] ? 4'h6 : _GEN_7289; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7291 = 10'h2da == _T_107[9:0] ? 4'h4 : _GEN_7290; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7292 = 10'h2db == _T_107[9:0] ? 4'h2 : _GEN_7291; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7293 = 10'h2dc == _T_107[9:0] ? 4'h2 : _GEN_7292; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7294 = 10'h2dd == _T_107[9:0] ? 4'h3 : _GEN_7293; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7295 = 10'h2de == _T_107[9:0] ? 4'h3 : _GEN_7294; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7296 = 10'h2df == _T_107[9:0] ? 4'h3 : _GEN_7295; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7297 = 10'h2e0 == _T_107[9:0] ? 4'h3 : _GEN_7296; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7298 = 10'h2e1 == _T_107[9:0] ? 4'h3 : _GEN_7297; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7299 = 10'h2e2 == _T_107[9:0] ? 4'h3 : _GEN_7298; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7300 = 10'h2e3 == _T_107[9:0] ? 4'h2 : _GEN_7299; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7301 = 10'h2e4 == _T_107[9:0] ? 4'h3 : _GEN_7300; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7302 = 10'h2e5 == _T_107[9:0] ? 4'h2 : _GEN_7301; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7303 = 10'h2e6 == _T_107[9:0] ? 4'h5 : _GEN_7302; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7304 = 10'h2e7 == _T_107[9:0] ? 4'h5 : _GEN_7303; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7305 = 10'h2e8 == _T_107[9:0] ? 4'h5 : _GEN_7304; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7306 = 10'h2e9 == _T_107[9:0] ? 4'h5 : _GEN_7305; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7307 = 10'h2ea == _T_107[9:0] ? 4'h5 : _GEN_7306; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7308 = 10'h2eb == _T_107[9:0] ? 4'h5 : _GEN_7307; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7309 = 10'h2ec == _T_107[9:0] ? 4'h6 : _GEN_7308; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7310 = 10'h2ed == _T_107[9:0] ? 4'h7 : _GEN_7309; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7311 = 10'h2ee == _T_107[9:0] ? 4'h6 : _GEN_7310; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7312 = 10'h2ef == _T_107[9:0] ? 4'h2 : _GEN_7311; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7313 = 10'h2f0 == _T_107[9:0] ? 4'h2 : _GEN_7312; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7314 = 10'h2f1 == _T_107[9:0] ? 4'h2 : _GEN_7313; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7315 = 10'h2f2 == _T_107[9:0] ? 4'h2 : _GEN_7314; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7316 = 10'h2f3 == _T_107[9:0] ? 4'h2 : _GEN_7315; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7317 = 10'h2f4 == _T_107[9:0] ? 4'h2 : _GEN_7316; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7318 = 10'h2f5 == _T_107[9:0] ? 4'h2 : _GEN_7317; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7319 = 10'h2f6 == _T_107[9:0] ? 4'h2 : _GEN_7318; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7320 = 10'h2f7 == _T_107[9:0] ? 4'h2 : _GEN_7319; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7321 = 10'h2f8 == _T_107[9:0] ? 4'h7 : _GEN_7320; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7322 = 10'h2f9 == _T_107[9:0] ? 4'h7 : _GEN_7321; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7323 = 10'h2fa == _T_107[9:0] ? 4'h8 : _GEN_7322; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7324 = 10'h2fb == _T_107[9:0] ? 4'h8 : _GEN_7323; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7325 = 10'h2fc == _T_107[9:0] ? 4'h7 : _GEN_7324; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7326 = 10'h2fd == _T_107[9:0] ? 4'h7 : _GEN_7325; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7327 = 10'h2fe == _T_107[9:0] ? 4'h7 : _GEN_7326; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7328 = 10'h2ff == _T_107[9:0] ? 4'h7 : _GEN_7327; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7329 = 10'h300 == _T_107[9:0] ? 4'h8 : _GEN_7328; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7330 = 10'h301 == _T_107[9:0] ? 4'h7 : _GEN_7329; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7331 = 10'h302 == _T_107[9:0] ? 4'h3 : _GEN_7330; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7332 = 10'h303 == _T_107[9:0] ? 4'h3 : _GEN_7331; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7333 = 10'h304 == _T_107[9:0] ? 4'h2 : _GEN_7332; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7334 = 10'h305 == _T_107[9:0] ? 4'h2 : _GEN_7333; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7335 = 10'h306 == _T_107[9:0] ? 4'h2 : _GEN_7334; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7336 = 10'h307 == _T_107[9:0] ? 4'h2 : _GEN_7335; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7337 = 10'h308 == _T_107[9:0] ? 4'h2 : _GEN_7336; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7338 = 10'h309 == _T_107[9:0] ? 4'h2 : _GEN_7337; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7339 = 10'h30a == _T_107[9:0] ? 4'h2 : _GEN_7338; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7340 = 10'h30b == _T_107[9:0] ? 4'h3 : _GEN_7339; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7341 = 10'h30c == _T_107[9:0] ? 4'h4 : _GEN_7340; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7342 = 10'h30d == _T_107[9:0] ? 4'h5 : _GEN_7341; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7343 = 10'h30e == _T_107[9:0] ? 4'h5 : _GEN_7342; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7344 = 10'h30f == _T_107[9:0] ? 4'h5 : _GEN_7343; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7345 = 10'h310 == _T_107[9:0] ? 4'h5 : _GEN_7344; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7346 = 10'h311 == _T_107[9:0] ? 4'h5 : _GEN_7345; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7347 = 10'h312 == _T_107[9:0] ? 4'h6 : _GEN_7346; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7348 = 10'h313 == _T_107[9:0] ? 4'h7 : _GEN_7347; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7349 = 10'h314 == _T_107[9:0] ? 4'h7 : _GEN_7348; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7350 = 10'h315 == _T_107[9:0] ? 4'h3 : _GEN_7349; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7351 = 10'h316 == _T_107[9:0] ? 4'h2 : _GEN_7350; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7352 = 10'h317 == _T_107[9:0] ? 4'h2 : _GEN_7351; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7353 = 10'h318 == _T_107[9:0] ? 4'h2 : _GEN_7352; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7354 = 10'h319 == _T_107[9:0] ? 4'h2 : _GEN_7353; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7355 = 10'h31a == _T_107[9:0] ? 4'h2 : _GEN_7354; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7356 = 10'h31b == _T_107[9:0] ? 4'h2 : _GEN_7355; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7357 = 10'h31c == _T_107[9:0] ? 4'h2 : _GEN_7356; // @[Filter.scala 230:142]
  wire [3:0] _GEN_7358 = 10'h31d == _T_107[9:0] ? 4'h2 : _GEN_7357; // @[Filter.scala 230:142]
  wire [7:0] _T_121 = _GEN_7358 * 4'ha; // @[Filter.scala 230:142]
  wire [10:0] _GEN_38971 = {{3'd0}, _T_121}; // @[Filter.scala 230:109]
  wire [10:0] _T_123 = _T_116 + _GEN_38971; // @[Filter.scala 230:109]
  wire [10:0] _T_124 = _T_123 / 11'h64; // @[Filter.scala 230:150]
  wire  _T_126 = _T_97 >= 6'h20; // @[Filter.scala 233:31]
  wire  _T_130 = _T_104 >= 32'h12; // @[Filter.scala 233:63]
  wire  _T_131 = _T_126 | _T_130; // @[Filter.scala 233:58]
  wire [10:0] _GEN_8157 = io_SPI_distort ? _T_124 : {{7'd0}, _GEN_5762}; // @[Filter.scala 235:35]
  wire [10:0] _GEN_8158 = _T_131 ? 11'h0 : _GEN_8157; // @[Filter.scala 233:80]
  wire [10:0] _GEN_8957 = io_SPI_distort ? _T_124 : {{7'd0}, _GEN_6560}; // @[Filter.scala 235:35]
  wire [10:0] _GEN_8958 = _T_131 ? 11'h0 : _GEN_8957; // @[Filter.scala 233:80]
  wire [10:0] _GEN_9757 = io_SPI_distort ? _T_124 : {{7'd0}, _GEN_7358}; // @[Filter.scala 235:35]
  wire [10:0] _GEN_9758 = _T_131 ? 11'h0 : _GEN_9757; // @[Filter.scala 233:80]
  wire [31:0] _T_159 = pixelIndex + 32'h2; // @[Filter.scala 228:31]
  wire [31:0] _GEN_2 = _T_159 % 32'h20; // @[Filter.scala 228:38]
  wire [5:0] _T_160 = _GEN_2[5:0]; // @[Filter.scala 228:38]
  wire [5:0] _T_162 = _T_160 + _GEN_38951; // @[Filter.scala 228:53]
  wire [5:0] _T_164 = _T_162 - 6'h1; // @[Filter.scala 228:69]
  wire [31:0] _T_167 = _T_159 / 32'h20; // @[Filter.scala 229:38]
  wire [31:0] _T_169 = _T_167 + _GEN_38952; // @[Filter.scala 229:53]
  wire [31:0] _T_171 = _T_169 - 32'h1; // @[Filter.scala 229:69]
  wire [37:0] _T_172 = _T_171 * 32'h20; // @[Filter.scala 230:42]
  wire [37:0] _GEN_38977 = {{32'd0}, _T_164}; // @[Filter.scala 230:57]
  wire [37:0] _T_174 = _T_172 + _GEN_38977; // @[Filter.scala 230:57]
  wire [3:0] _GEN_9781 = 10'h16 == _T_174[9:0] ? 4'h9 : 4'ha; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9782 = 10'h17 == _T_174[9:0] ? 4'h3 : _GEN_9781; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9783 = 10'h18 == _T_174[9:0] ? 4'h6 : _GEN_9782; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9784 = 10'h19 == _T_174[9:0] ? 4'ha : _GEN_9783; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9785 = 10'h1a == _T_174[9:0] ? 4'ha : _GEN_9784; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9786 = 10'h1b == _T_174[9:0] ? 4'ha : _GEN_9785; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9787 = 10'h1c == _T_174[9:0] ? 4'ha : _GEN_9786; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9788 = 10'h1d == _T_174[9:0] ? 4'ha : _GEN_9787; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9789 = 10'h1e == _T_174[9:0] ? 4'ha : _GEN_9788; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9790 = 10'h1f == _T_174[9:0] ? 4'ha : _GEN_9789; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9791 = 10'h20 == _T_174[9:0] ? 4'ha : _GEN_9790; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9792 = 10'h21 == _T_174[9:0] ? 4'ha : _GEN_9791; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9793 = 10'h22 == _T_174[9:0] ? 4'ha : _GEN_9792; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9794 = 10'h23 == _T_174[9:0] ? 4'ha : _GEN_9793; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9795 = 10'h24 == _T_174[9:0] ? 4'ha : _GEN_9794; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9796 = 10'h25 == _T_174[9:0] ? 4'ha : _GEN_9795; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9797 = 10'h26 == _T_174[9:0] ? 4'ha : _GEN_9796; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9798 = 10'h27 == _T_174[9:0] ? 4'ha : _GEN_9797; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9799 = 10'h28 == _T_174[9:0] ? 4'ha : _GEN_9798; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9800 = 10'h29 == _T_174[9:0] ? 4'ha : _GEN_9799; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9801 = 10'h2a == _T_174[9:0] ? 4'ha : _GEN_9800; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9802 = 10'h2b == _T_174[9:0] ? 4'ha : _GEN_9801; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9803 = 10'h2c == _T_174[9:0] ? 4'ha : _GEN_9802; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9804 = 10'h2d == _T_174[9:0] ? 4'ha : _GEN_9803; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9805 = 10'h2e == _T_174[9:0] ? 4'ha : _GEN_9804; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9806 = 10'h2f == _T_174[9:0] ? 4'ha : _GEN_9805; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9807 = 10'h30 == _T_174[9:0] ? 4'ha : _GEN_9806; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9808 = 10'h31 == _T_174[9:0] ? 4'ha : _GEN_9807; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9809 = 10'h32 == _T_174[9:0] ? 4'ha : _GEN_9808; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9810 = 10'h33 == _T_174[9:0] ? 4'ha : _GEN_9809; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9811 = 10'h34 == _T_174[9:0] ? 4'ha : _GEN_9810; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9812 = 10'h35 == _T_174[9:0] ? 4'ha : _GEN_9811; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9813 = 10'h36 == _T_174[9:0] ? 4'ha : _GEN_9812; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9814 = 10'h37 == _T_174[9:0] ? 4'ha : _GEN_9813; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9815 = 10'h38 == _T_174[9:0] ? 4'ha : _GEN_9814; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9816 = 10'h39 == _T_174[9:0] ? 4'ha : _GEN_9815; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9817 = 10'h3a == _T_174[9:0] ? 4'ha : _GEN_9816; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9818 = 10'h3b == _T_174[9:0] ? 4'h9 : _GEN_9817; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9819 = 10'h3c == _T_174[9:0] ? 4'h4 : _GEN_9818; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9820 = 10'h3d == _T_174[9:0] ? 4'h3 : _GEN_9819; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9821 = 10'h3e == _T_174[9:0] ? 4'h4 : _GEN_9820; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9822 = 10'h3f == _T_174[9:0] ? 4'ha : _GEN_9821; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9823 = 10'h40 == _T_174[9:0] ? 4'ha : _GEN_9822; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9824 = 10'h41 == _T_174[9:0] ? 4'ha : _GEN_9823; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9825 = 10'h42 == _T_174[9:0] ? 4'ha : _GEN_9824; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9826 = 10'h43 == _T_174[9:0] ? 4'ha : _GEN_9825; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9827 = 10'h44 == _T_174[9:0] ? 4'ha : _GEN_9826; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9828 = 10'h45 == _T_174[9:0] ? 4'ha : _GEN_9827; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9829 = 10'h46 == _T_174[9:0] ? 4'ha : _GEN_9828; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9830 = 10'h47 == _T_174[9:0] ? 4'ha : _GEN_9829; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9831 = 10'h48 == _T_174[9:0] ? 4'ha : _GEN_9830; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9832 = 10'h49 == _T_174[9:0] ? 4'ha : _GEN_9831; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9833 = 10'h4a == _T_174[9:0] ? 4'ha : _GEN_9832; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9834 = 10'h4b == _T_174[9:0] ? 4'ha : _GEN_9833; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9835 = 10'h4c == _T_174[9:0] ? 4'ha : _GEN_9834; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9836 = 10'h4d == _T_174[9:0] ? 4'ha : _GEN_9835; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9837 = 10'h4e == _T_174[9:0] ? 4'ha : _GEN_9836; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9838 = 10'h4f == _T_174[9:0] ? 4'ha : _GEN_9837; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9839 = 10'h50 == _T_174[9:0] ? 4'ha : _GEN_9838; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9840 = 10'h51 == _T_174[9:0] ? 4'ha : _GEN_9839; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9841 = 10'h52 == _T_174[9:0] ? 4'ha : _GEN_9840; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9842 = 10'h53 == _T_174[9:0] ? 4'ha : _GEN_9841; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9843 = 10'h54 == _T_174[9:0] ? 4'ha : _GEN_9842; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9844 = 10'h55 == _T_174[9:0] ? 4'ha : _GEN_9843; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9845 = 10'h56 == _T_174[9:0] ? 4'ha : _GEN_9844; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9846 = 10'h57 == _T_174[9:0] ? 4'ha : _GEN_9845; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9847 = 10'h58 == _T_174[9:0] ? 4'ha : _GEN_9846; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9848 = 10'h59 == _T_174[9:0] ? 4'ha : _GEN_9847; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9849 = 10'h5a == _T_174[9:0] ? 4'h7 : _GEN_9848; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9850 = 10'h5b == _T_174[9:0] ? 4'h7 : _GEN_9849; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9851 = 10'h5c == _T_174[9:0] ? 4'ha : _GEN_9850; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9852 = 10'h5d == _T_174[9:0] ? 4'ha : _GEN_9851; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9853 = 10'h5e == _T_174[9:0] ? 4'ha : _GEN_9852; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9854 = 10'h5f == _T_174[9:0] ? 4'ha : _GEN_9853; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9855 = 10'h60 == _T_174[9:0] ? 4'ha : _GEN_9854; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9856 = 10'h61 == _T_174[9:0] ? 4'h8 : _GEN_9855; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9857 = 10'h62 == _T_174[9:0] ? 4'h3 : _GEN_9856; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9858 = 10'h63 == _T_174[9:0] ? 4'h3 : _GEN_9857; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9859 = 10'h64 == _T_174[9:0] ? 4'h3 : _GEN_9858; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9860 = 10'h65 == _T_174[9:0] ? 4'h9 : _GEN_9859; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9861 = 10'h66 == _T_174[9:0] ? 4'ha : _GEN_9860; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9862 = 10'h67 == _T_174[9:0] ? 4'ha : _GEN_9861; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9863 = 10'h68 == _T_174[9:0] ? 4'ha : _GEN_9862; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9864 = 10'h69 == _T_174[9:0] ? 4'ha : _GEN_9863; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9865 = 10'h6a == _T_174[9:0] ? 4'ha : _GEN_9864; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9866 = 10'h6b == _T_174[9:0] ? 4'h8 : _GEN_9865; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9867 = 10'h6c == _T_174[9:0] ? 4'h5 : _GEN_9866; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9868 = 10'h6d == _T_174[9:0] ? 4'h8 : _GEN_9867; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9869 = 10'h6e == _T_174[9:0] ? 4'ha : _GEN_9868; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9870 = 10'h6f == _T_174[9:0] ? 4'ha : _GEN_9869; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9871 = 10'h70 == _T_174[9:0] ? 4'ha : _GEN_9870; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9872 = 10'h71 == _T_174[9:0] ? 4'ha : _GEN_9871; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9873 = 10'h72 == _T_174[9:0] ? 4'ha : _GEN_9872; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9874 = 10'h73 == _T_174[9:0] ? 4'ha : _GEN_9873; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9875 = 10'h74 == _T_174[9:0] ? 4'ha : _GEN_9874; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9876 = 10'h75 == _T_174[9:0] ? 4'ha : _GEN_9875; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9877 = 10'h76 == _T_174[9:0] ? 4'ha : _GEN_9876; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9878 = 10'h77 == _T_174[9:0] ? 4'ha : _GEN_9877; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9879 = 10'h78 == _T_174[9:0] ? 4'ha : _GEN_9878; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9880 = 10'h79 == _T_174[9:0] ? 4'ha : _GEN_9879; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9881 = 10'h7a == _T_174[9:0] ? 4'ha : _GEN_9880; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9882 = 10'h7b == _T_174[9:0] ? 4'ha : _GEN_9881; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9883 = 10'h7c == _T_174[9:0] ? 4'ha : _GEN_9882; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9884 = 10'h7d == _T_174[9:0] ? 4'ha : _GEN_9883; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9885 = 10'h7e == _T_174[9:0] ? 4'ha : _GEN_9884; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9886 = 10'h7f == _T_174[9:0] ? 4'ha : _GEN_9885; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9887 = 10'h80 == _T_174[9:0] ? 4'ha : _GEN_9886; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9888 = 10'h81 == _T_174[9:0] ? 4'h5 : _GEN_9887; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9889 = 10'h82 == _T_174[9:0] ? 4'h5 : _GEN_9888; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9890 = 10'h83 == _T_174[9:0] ? 4'h7 : _GEN_9889; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9891 = 10'h84 == _T_174[9:0] ? 4'ha : _GEN_9890; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9892 = 10'h85 == _T_174[9:0] ? 4'ha : _GEN_9891; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9893 = 10'h86 == _T_174[9:0] ? 4'ha : _GEN_9892; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9894 = 10'h87 == _T_174[9:0] ? 4'h5 : _GEN_9893; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9895 = 10'h88 == _T_174[9:0] ? 4'h3 : _GEN_9894; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9896 = 10'h89 == _T_174[9:0] ? 4'h3 : _GEN_9895; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9897 = 10'h8a == _T_174[9:0] ? 4'h4 : _GEN_9896; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9898 = 10'h8b == _T_174[9:0] ? 4'h9 : _GEN_9897; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9899 = 10'h8c == _T_174[9:0] ? 4'ha : _GEN_9898; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9900 = 10'h8d == _T_174[9:0] ? 4'ha : _GEN_9899; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9901 = 10'h8e == _T_174[9:0] ? 4'ha : _GEN_9900; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9902 = 10'h8f == _T_174[9:0] ? 4'h6 : _GEN_9901; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9903 = 10'h90 == _T_174[9:0] ? 4'h4 : _GEN_9902; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9904 = 10'h91 == _T_174[9:0] ? 4'h3 : _GEN_9903; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9905 = 10'h92 == _T_174[9:0] ? 4'h7 : _GEN_9904; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9906 = 10'h93 == _T_174[9:0] ? 4'ha : _GEN_9905; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9907 = 10'h94 == _T_174[9:0] ? 4'ha : _GEN_9906; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9908 = 10'h95 == _T_174[9:0] ? 4'ha : _GEN_9907; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9909 = 10'h96 == _T_174[9:0] ? 4'ha : _GEN_9908; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9910 = 10'h97 == _T_174[9:0] ? 4'ha : _GEN_9909; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9911 = 10'h98 == _T_174[9:0] ? 4'ha : _GEN_9910; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9912 = 10'h99 == _T_174[9:0] ? 4'ha : _GEN_9911; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9913 = 10'h9a == _T_174[9:0] ? 4'ha : _GEN_9912; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9914 = 10'h9b == _T_174[9:0] ? 4'ha : _GEN_9913; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9915 = 10'h9c == _T_174[9:0] ? 4'ha : _GEN_9914; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9916 = 10'h9d == _T_174[9:0] ? 4'ha : _GEN_9915; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9917 = 10'h9e == _T_174[9:0] ? 4'ha : _GEN_9916; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9918 = 10'h9f == _T_174[9:0] ? 4'ha : _GEN_9917; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9919 = 10'ha0 == _T_174[9:0] ? 4'ha : _GEN_9918; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9920 = 10'ha1 == _T_174[9:0] ? 4'ha : _GEN_9919; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9921 = 10'ha2 == _T_174[9:0] ? 4'ha : _GEN_9920; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9922 = 10'ha3 == _T_174[9:0] ? 4'ha : _GEN_9921; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9923 = 10'ha4 == _T_174[9:0] ? 4'ha : _GEN_9922; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9924 = 10'ha5 == _T_174[9:0] ? 4'ha : _GEN_9923; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9925 = 10'ha6 == _T_174[9:0] ? 4'ha : _GEN_9924; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9926 = 10'ha7 == _T_174[9:0] ? 4'h9 : _GEN_9925; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9927 = 10'ha8 == _T_174[9:0] ? 4'h4 : _GEN_9926; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9928 = 10'ha9 == _T_174[9:0] ? 4'h3 : _GEN_9927; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9929 = 10'haa == _T_174[9:0] ? 4'h4 : _GEN_9928; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9930 = 10'hab == _T_174[9:0] ? 4'h7 : _GEN_9929; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9931 = 10'hac == _T_174[9:0] ? 4'h8 : _GEN_9930; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9932 = 10'had == _T_174[9:0] ? 4'h3 : _GEN_9931; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9933 = 10'hae == _T_174[9:0] ? 4'h3 : _GEN_9932; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9934 = 10'haf == _T_174[9:0] ? 4'h3 : _GEN_9933; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9935 = 10'hb0 == _T_174[9:0] ? 4'h3 : _GEN_9934; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9936 = 10'hb1 == _T_174[9:0] ? 4'h7 : _GEN_9935; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9937 = 10'hb2 == _T_174[9:0] ? 4'h9 : _GEN_9936; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9938 = 10'hb3 == _T_174[9:0] ? 4'h6 : _GEN_9937; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9939 = 10'hb4 == _T_174[9:0] ? 4'h4 : _GEN_9938; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9940 = 10'hb5 == _T_174[9:0] ? 4'h3 : _GEN_9939; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9941 = 10'hb6 == _T_174[9:0] ? 4'h3 : _GEN_9940; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9942 = 10'hb7 == _T_174[9:0] ? 4'h6 : _GEN_9941; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9943 = 10'hb8 == _T_174[9:0] ? 4'ha : _GEN_9942; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9944 = 10'hb9 == _T_174[9:0] ? 4'ha : _GEN_9943; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9945 = 10'hba == _T_174[9:0] ? 4'ha : _GEN_9944; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9946 = 10'hbb == _T_174[9:0] ? 4'ha : _GEN_9945; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9947 = 10'hbc == _T_174[9:0] ? 4'ha : _GEN_9946; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9948 = 10'hbd == _T_174[9:0] ? 4'h9 : _GEN_9947; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9949 = 10'hbe == _T_174[9:0] ? 4'ha : _GEN_9948; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9950 = 10'hbf == _T_174[9:0] ? 4'ha : _GEN_9949; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9951 = 10'hc0 == _T_174[9:0] ? 4'ha : _GEN_9950; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9952 = 10'hc1 == _T_174[9:0] ? 4'ha : _GEN_9951; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9953 = 10'hc2 == _T_174[9:0] ? 4'ha : _GEN_9952; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9954 = 10'hc3 == _T_174[9:0] ? 4'ha : _GEN_9953; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9955 = 10'hc4 == _T_174[9:0] ? 4'ha : _GEN_9954; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9956 = 10'hc5 == _T_174[9:0] ? 4'ha : _GEN_9955; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9957 = 10'hc6 == _T_174[9:0] ? 4'ha : _GEN_9956; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9958 = 10'hc7 == _T_174[9:0] ? 4'h9 : _GEN_9957; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9959 = 10'hc8 == _T_174[9:0] ? 4'h8 : _GEN_9958; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9960 = 10'hc9 == _T_174[9:0] ? 4'h8 : _GEN_9959; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9961 = 10'hca == _T_174[9:0] ? 4'h9 : _GEN_9960; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9962 = 10'hcb == _T_174[9:0] ? 4'ha : _GEN_9961; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9963 = 10'hcc == _T_174[9:0] ? 4'ha : _GEN_9962; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9964 = 10'hcd == _T_174[9:0] ? 4'ha : _GEN_9963; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9965 = 10'hce == _T_174[9:0] ? 4'h8 : _GEN_9964; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9966 = 10'hcf == _T_174[9:0] ? 4'h3 : _GEN_9965; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9967 = 10'hd0 == _T_174[9:0] ? 4'h3 : _GEN_9966; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9968 = 10'hd1 == _T_174[9:0] ? 4'h3 : _GEN_9967; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9969 = 10'hd2 == _T_174[9:0] ? 4'h4 : _GEN_9968; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9970 = 10'hd3 == _T_174[9:0] ? 4'h3 : _GEN_9969; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9971 = 10'hd4 == _T_174[9:0] ? 4'h3 : _GEN_9970; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9972 = 10'hd5 == _T_174[9:0] ? 4'h3 : _GEN_9971; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9973 = 10'hd6 == _T_174[9:0] ? 4'h3 : _GEN_9972; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9974 = 10'hd7 == _T_174[9:0] ? 4'h5 : _GEN_9973; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9975 = 10'hd8 == _T_174[9:0] ? 4'h4 : _GEN_9974; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9976 = 10'hd9 == _T_174[9:0] ? 4'h3 : _GEN_9975; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9977 = 10'hda == _T_174[9:0] ? 4'h3 : _GEN_9976; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9978 = 10'hdb == _T_174[9:0] ? 4'h3 : _GEN_9977; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9979 = 10'hdc == _T_174[9:0] ? 4'h4 : _GEN_9978; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9980 = 10'hdd == _T_174[9:0] ? 4'ha : _GEN_9979; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9981 = 10'hde == _T_174[9:0] ? 4'ha : _GEN_9980; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9982 = 10'hdf == _T_174[9:0] ? 4'ha : _GEN_9981; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9983 = 10'he0 == _T_174[9:0] ? 4'ha : _GEN_9982; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9984 = 10'he1 == _T_174[9:0] ? 4'ha : _GEN_9983; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9985 = 10'he2 == _T_174[9:0] ? 4'ha : _GEN_9984; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9986 = 10'he3 == _T_174[9:0] ? 4'h5 : _GEN_9985; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9987 = 10'he4 == _T_174[9:0] ? 4'ha : _GEN_9986; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9988 = 10'he5 == _T_174[9:0] ? 4'ha : _GEN_9987; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9989 = 10'he6 == _T_174[9:0] ? 4'ha : _GEN_9988; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9990 = 10'he7 == _T_174[9:0] ? 4'ha : _GEN_9989; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9991 = 10'he8 == _T_174[9:0] ? 4'ha : _GEN_9990; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9992 = 10'he9 == _T_174[9:0] ? 4'ha : _GEN_9991; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9993 = 10'hea == _T_174[9:0] ? 4'ha : _GEN_9992; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9994 = 10'heb == _T_174[9:0] ? 4'h9 : _GEN_9993; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9995 = 10'hec == _T_174[9:0] ? 4'h7 : _GEN_9994; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9996 = 10'hed == _T_174[9:0] ? 4'h3 : _GEN_9995; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9997 = 10'hee == _T_174[9:0] ? 4'h3 : _GEN_9996; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9998 = 10'hef == _T_174[9:0] ? 4'h3 : _GEN_9997; // @[Filter.scala 230:62]
  wire [3:0] _GEN_9999 = 10'hf0 == _T_174[9:0] ? 4'h4 : _GEN_9998; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10000 = 10'hf1 == _T_174[9:0] ? 4'h7 : _GEN_9999; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10001 = 10'hf2 == _T_174[9:0] ? 4'ha : _GEN_10000; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10002 = 10'hf3 == _T_174[9:0] ? 4'ha : _GEN_10001; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10003 = 10'hf4 == _T_174[9:0] ? 4'ha : _GEN_10002; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10004 = 10'hf5 == _T_174[9:0] ? 4'h7 : _GEN_10003; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10005 = 10'hf6 == _T_174[9:0] ? 4'h3 : _GEN_10004; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10006 = 10'hf7 == _T_174[9:0] ? 4'h3 : _GEN_10005; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10007 = 10'hf8 == _T_174[9:0] ? 4'h3 : _GEN_10006; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10008 = 10'hf9 == _T_174[9:0] ? 4'h3 : _GEN_10007; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10009 = 10'hfa == _T_174[9:0] ? 4'h3 : _GEN_10008; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10010 = 10'hfb == _T_174[9:0] ? 4'h3 : _GEN_10009; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10011 = 10'hfc == _T_174[9:0] ? 4'h3 : _GEN_10010; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10012 = 10'hfd == _T_174[9:0] ? 4'h3 : _GEN_10011; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10013 = 10'hfe == _T_174[9:0] ? 4'h3 : _GEN_10012; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10014 = 10'hff == _T_174[9:0] ? 4'h3 : _GEN_10013; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10015 = 10'h100 == _T_174[9:0] ? 4'h3 : _GEN_10014; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10016 = 10'h101 == _T_174[9:0] ? 4'h4 : _GEN_10015; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10017 = 10'h102 == _T_174[9:0] ? 4'h6 : _GEN_10016; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10018 = 10'h103 == _T_174[9:0] ? 4'ha : _GEN_10017; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10019 = 10'h104 == _T_174[9:0] ? 4'ha : _GEN_10018; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10020 = 10'h105 == _T_174[9:0] ? 4'h9 : _GEN_10019; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10021 = 10'h106 == _T_174[9:0] ? 4'h9 : _GEN_10020; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10022 = 10'h107 == _T_174[9:0] ? 4'h9 : _GEN_10021; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10023 = 10'h108 == _T_174[9:0] ? 4'h9 : _GEN_10022; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10024 = 10'h109 == _T_174[9:0] ? 4'h3 : _GEN_10023; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10025 = 10'h10a == _T_174[9:0] ? 4'ha : _GEN_10024; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10026 = 10'h10b == _T_174[9:0] ? 4'ha : _GEN_10025; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10027 = 10'h10c == _T_174[9:0] ? 4'ha : _GEN_10026; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10028 = 10'h10d == _T_174[9:0] ? 4'ha : _GEN_10027; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10029 = 10'h10e == _T_174[9:0] ? 4'ha : _GEN_10028; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10030 = 10'h10f == _T_174[9:0] ? 4'h9 : _GEN_10029; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10031 = 10'h110 == _T_174[9:0] ? 4'h9 : _GEN_10030; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10032 = 10'h111 == _T_174[9:0] ? 4'h4 : _GEN_10031; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10033 = 10'h112 == _T_174[9:0] ? 4'h8 : _GEN_10032; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10034 = 10'h113 == _T_174[9:0] ? 4'h3 : _GEN_10033; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10035 = 10'h114 == _T_174[9:0] ? 4'h3 : _GEN_10034; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10036 = 10'h115 == _T_174[9:0] ? 4'h4 : _GEN_10035; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10037 = 10'h116 == _T_174[9:0] ? 4'h4 : _GEN_10036; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10038 = 10'h117 == _T_174[9:0] ? 4'h3 : _GEN_10037; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10039 = 10'h118 == _T_174[9:0] ? 4'h8 : _GEN_10038; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10040 = 10'h119 == _T_174[9:0] ? 4'ha : _GEN_10039; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10041 = 10'h11a == _T_174[9:0] ? 4'ha : _GEN_10040; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10042 = 10'h11b == _T_174[9:0] ? 4'ha : _GEN_10041; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10043 = 10'h11c == _T_174[9:0] ? 4'h6 : _GEN_10042; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10044 = 10'h11d == _T_174[9:0] ? 4'h3 : _GEN_10043; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10045 = 10'h11e == _T_174[9:0] ? 4'h3 : _GEN_10044; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10046 = 10'h11f == _T_174[9:0] ? 4'h3 : _GEN_10045; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10047 = 10'h120 == _T_174[9:0] ? 4'h3 : _GEN_10046; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10048 = 10'h121 == _T_174[9:0] ? 4'h3 : _GEN_10047; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10049 = 10'h122 == _T_174[9:0] ? 4'h3 : _GEN_10048; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10050 = 10'h123 == _T_174[9:0] ? 4'h3 : _GEN_10049; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10051 = 10'h124 == _T_174[9:0] ? 4'h3 : _GEN_10050; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10052 = 10'h125 == _T_174[9:0] ? 4'h3 : _GEN_10051; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10053 = 10'h126 == _T_174[9:0] ? 4'h4 : _GEN_10052; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10054 = 10'h127 == _T_174[9:0] ? 4'h6 : _GEN_10053; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10055 = 10'h128 == _T_174[9:0] ? 4'h5 : _GEN_10054; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10056 = 10'h129 == _T_174[9:0] ? 4'h8 : _GEN_10055; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10057 = 10'h12a == _T_174[9:0] ? 4'h5 : _GEN_10056; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10058 = 10'h12b == _T_174[9:0] ? 4'h3 : _GEN_10057; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10059 = 10'h12c == _T_174[9:0] ? 4'h3 : _GEN_10058; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10060 = 10'h12d == _T_174[9:0] ? 4'h3 : _GEN_10059; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10061 = 10'h12e == _T_174[9:0] ? 4'h4 : _GEN_10060; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10062 = 10'h12f == _T_174[9:0] ? 4'h4 : _GEN_10061; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10063 = 10'h130 == _T_174[9:0] ? 4'ha : _GEN_10062; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10064 = 10'h131 == _T_174[9:0] ? 4'h9 : _GEN_10063; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10065 = 10'h132 == _T_174[9:0] ? 4'h9 : _GEN_10064; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10066 = 10'h133 == _T_174[9:0] ? 4'h8 : _GEN_10065; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10067 = 10'h134 == _T_174[9:0] ? 4'h9 : _GEN_10066; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10068 = 10'h135 == _T_174[9:0] ? 4'h8 : _GEN_10067; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10069 = 10'h136 == _T_174[9:0] ? 4'h7 : _GEN_10068; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10070 = 10'h137 == _T_174[9:0] ? 4'h6 : _GEN_10069; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10071 = 10'h138 == _T_174[9:0] ? 4'h8 : _GEN_10070; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10072 = 10'h139 == _T_174[9:0] ? 4'h3 : _GEN_10071; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10073 = 10'h13a == _T_174[9:0] ? 4'h3 : _GEN_10072; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10074 = 10'h13b == _T_174[9:0] ? 4'h4 : _GEN_10073; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10075 = 10'h13c == _T_174[9:0] ? 4'h4 : _GEN_10074; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10076 = 10'h13d == _T_174[9:0] ? 4'h3 : _GEN_10075; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10077 = 10'h13e == _T_174[9:0] ? 4'h5 : _GEN_10076; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10078 = 10'h13f == _T_174[9:0] ? 4'h9 : _GEN_10077; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10079 = 10'h140 == _T_174[9:0] ? 4'ha : _GEN_10078; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10080 = 10'h141 == _T_174[9:0] ? 4'ha : _GEN_10079; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10081 = 10'h142 == _T_174[9:0] ? 4'ha : _GEN_10080; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10082 = 10'h143 == _T_174[9:0] ? 4'h5 : _GEN_10081; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10083 = 10'h144 == _T_174[9:0] ? 4'h3 : _GEN_10082; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10084 = 10'h145 == _T_174[9:0] ? 4'h3 : _GEN_10083; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10085 = 10'h146 == _T_174[9:0] ? 4'h3 : _GEN_10084; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10086 = 10'h147 == _T_174[9:0] ? 4'h4 : _GEN_10085; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10087 = 10'h148 == _T_174[9:0] ? 4'h3 : _GEN_10086; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10088 = 10'h149 == _T_174[9:0] ? 4'h3 : _GEN_10087; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10089 = 10'h14a == _T_174[9:0] ? 4'h3 : _GEN_10088; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10090 = 10'h14b == _T_174[9:0] ? 4'h6 : _GEN_10089; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10091 = 10'h14c == _T_174[9:0] ? 4'h8 : _GEN_10090; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10092 = 10'h14d == _T_174[9:0] ? 4'h5 : _GEN_10091; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10093 = 10'h14e == _T_174[9:0] ? 4'h4 : _GEN_10092; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10094 = 10'h14f == _T_174[9:0] ? 4'h3 : _GEN_10093; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10095 = 10'h150 == _T_174[9:0] ? 4'h3 : _GEN_10094; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10096 = 10'h151 == _T_174[9:0] ? 4'h3 : _GEN_10095; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10097 = 10'h152 == _T_174[9:0] ? 4'h3 : _GEN_10096; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10098 = 10'h153 == _T_174[9:0] ? 4'h3 : _GEN_10097; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10099 = 10'h154 == _T_174[9:0] ? 4'h3 : _GEN_10098; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10100 = 10'h155 == _T_174[9:0] ? 4'h4 : _GEN_10099; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10101 = 10'h156 == _T_174[9:0] ? 4'h9 : _GEN_10100; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10102 = 10'h157 == _T_174[9:0] ? 4'h8 : _GEN_10101; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10103 = 10'h158 == _T_174[9:0] ? 4'h8 : _GEN_10102; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10104 = 10'h159 == _T_174[9:0] ? 4'h8 : _GEN_10103; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10105 = 10'h15a == _T_174[9:0] ? 4'h8 : _GEN_10104; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10106 = 10'h15b == _T_174[9:0] ? 4'h8 : _GEN_10105; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10107 = 10'h15c == _T_174[9:0] ? 4'h7 : _GEN_10106; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10108 = 10'h15d == _T_174[9:0] ? 4'h7 : _GEN_10107; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10109 = 10'h15e == _T_174[9:0] ? 4'h8 : _GEN_10108; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10110 = 10'h15f == _T_174[9:0] ? 4'h3 : _GEN_10109; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10111 = 10'h160 == _T_174[9:0] ? 4'h4 : _GEN_10110; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10112 = 10'h161 == _T_174[9:0] ? 4'h4 : _GEN_10111; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10113 = 10'h162 == _T_174[9:0] ? 4'h4 : _GEN_10112; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10114 = 10'h163 == _T_174[9:0] ? 4'h4 : _GEN_10113; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10115 = 10'h164 == _T_174[9:0] ? 4'h5 : _GEN_10114; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10116 = 10'h165 == _T_174[9:0] ? 4'ha : _GEN_10115; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10117 = 10'h166 == _T_174[9:0] ? 4'h9 : _GEN_10116; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10118 = 10'h167 == _T_174[9:0] ? 4'ha : _GEN_10117; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10119 = 10'h168 == _T_174[9:0] ? 4'ha : _GEN_10118; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10120 = 10'h169 == _T_174[9:0] ? 4'h6 : _GEN_10119; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10121 = 10'h16a == _T_174[9:0] ? 4'h3 : _GEN_10120; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10122 = 10'h16b == _T_174[9:0] ? 4'h3 : _GEN_10121; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10123 = 10'h16c == _T_174[9:0] ? 4'h3 : _GEN_10122; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10124 = 10'h16d == _T_174[9:0] ? 4'h4 : _GEN_10123; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10125 = 10'h16e == _T_174[9:0] ? 4'h3 : _GEN_10124; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10126 = 10'h16f == _T_174[9:0] ? 4'h3 : _GEN_10125; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10127 = 10'h170 == _T_174[9:0] ? 4'h3 : _GEN_10126; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10128 = 10'h171 == _T_174[9:0] ? 4'h7 : _GEN_10127; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10129 = 10'h172 == _T_174[9:0] ? 4'ha : _GEN_10128; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10130 = 10'h173 == _T_174[9:0] ? 4'h5 : _GEN_10129; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10131 = 10'h174 == _T_174[9:0] ? 4'h3 : _GEN_10130; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10132 = 10'h175 == _T_174[9:0] ? 4'h4 : _GEN_10131; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10133 = 10'h176 == _T_174[9:0] ? 4'h4 : _GEN_10132; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10134 = 10'h177 == _T_174[9:0] ? 4'h4 : _GEN_10133; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10135 = 10'h178 == _T_174[9:0] ? 4'h4 : _GEN_10134; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10136 = 10'h179 == _T_174[9:0] ? 4'h3 : _GEN_10135; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10137 = 10'h17a == _T_174[9:0] ? 4'h3 : _GEN_10136; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10138 = 10'h17b == _T_174[9:0] ? 4'h3 : _GEN_10137; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10139 = 10'h17c == _T_174[9:0] ? 4'h8 : _GEN_10138; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10140 = 10'h17d == _T_174[9:0] ? 4'h8 : _GEN_10139; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10141 = 10'h17e == _T_174[9:0] ? 4'h8 : _GEN_10140; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10142 = 10'h17f == _T_174[9:0] ? 4'h8 : _GEN_10141; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10143 = 10'h180 == _T_174[9:0] ? 4'h8 : _GEN_10142; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10144 = 10'h181 == _T_174[9:0] ? 4'h8 : _GEN_10143; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10145 = 10'h182 == _T_174[9:0] ? 4'h8 : _GEN_10144; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10146 = 10'h183 == _T_174[9:0] ? 4'h8 : _GEN_10145; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10147 = 10'h184 == _T_174[9:0] ? 4'h8 : _GEN_10146; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10148 = 10'h185 == _T_174[9:0] ? 4'h5 : _GEN_10147; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10149 = 10'h186 == _T_174[9:0] ? 4'h3 : _GEN_10148; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10150 = 10'h187 == _T_174[9:0] ? 4'h4 : _GEN_10149; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10151 = 10'h188 == _T_174[9:0] ? 4'h4 : _GEN_10150; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10152 = 10'h189 == _T_174[9:0] ? 4'h4 : _GEN_10151; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10153 = 10'h18a == _T_174[9:0] ? 4'h5 : _GEN_10152; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10154 = 10'h18b == _T_174[9:0] ? 4'ha : _GEN_10153; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10155 = 10'h18c == _T_174[9:0] ? 4'ha : _GEN_10154; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10156 = 10'h18d == _T_174[9:0] ? 4'h9 : _GEN_10155; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10157 = 10'h18e == _T_174[9:0] ? 4'ha : _GEN_10156; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10158 = 10'h18f == _T_174[9:0] ? 4'h4 : _GEN_10157; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10159 = 10'h190 == _T_174[9:0] ? 4'h3 : _GEN_10158; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10160 = 10'h191 == _T_174[9:0] ? 4'h3 : _GEN_10159; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10161 = 10'h192 == _T_174[9:0] ? 4'h5 : _GEN_10160; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10162 = 10'h193 == _T_174[9:0] ? 4'h6 : _GEN_10161; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10163 = 10'h194 == _T_174[9:0] ? 4'h5 : _GEN_10162; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10164 = 10'h195 == _T_174[9:0] ? 4'h3 : _GEN_10163; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10165 = 10'h196 == _T_174[9:0] ? 4'h3 : _GEN_10164; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10166 = 10'h197 == _T_174[9:0] ? 4'h5 : _GEN_10165; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10167 = 10'h198 == _T_174[9:0] ? 4'ha : _GEN_10166; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10168 = 10'h199 == _T_174[9:0] ? 4'h3 : _GEN_10167; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10169 = 10'h19a == _T_174[9:0] ? 4'h1 : _GEN_10168; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10170 = 10'h19b == _T_174[9:0] ? 4'h2 : _GEN_10169; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10171 = 10'h19c == _T_174[9:0] ? 4'h4 : _GEN_10170; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10172 = 10'h19d == _T_174[9:0] ? 4'h3 : _GEN_10171; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10173 = 10'h19e == _T_174[9:0] ? 4'h1 : _GEN_10172; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10174 = 10'h19f == _T_174[9:0] ? 4'h2 : _GEN_10173; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10175 = 10'h1a0 == _T_174[9:0] ? 4'h3 : _GEN_10174; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10176 = 10'h1a1 == _T_174[9:0] ? 4'h4 : _GEN_10175; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10177 = 10'h1a2 == _T_174[9:0] ? 4'h8 : _GEN_10176; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10178 = 10'h1a3 == _T_174[9:0] ? 4'h8 : _GEN_10177; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10179 = 10'h1a4 == _T_174[9:0] ? 4'h8 : _GEN_10178; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10180 = 10'h1a5 == _T_174[9:0] ? 4'h8 : _GEN_10179; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10181 = 10'h1a6 == _T_174[9:0] ? 4'h7 : _GEN_10180; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10182 = 10'h1a7 == _T_174[9:0] ? 4'h8 : _GEN_10181; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10183 = 10'h1a8 == _T_174[9:0] ? 4'h8 : _GEN_10182; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10184 = 10'h1a9 == _T_174[9:0] ? 4'h8 : _GEN_10183; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10185 = 10'h1aa == _T_174[9:0] ? 4'h7 : _GEN_10184; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10186 = 10'h1ab == _T_174[9:0] ? 4'h4 : _GEN_10185; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10187 = 10'h1ac == _T_174[9:0] ? 4'h4 : _GEN_10186; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10188 = 10'h1ad == _T_174[9:0] ? 4'h3 : _GEN_10187; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10189 = 10'h1ae == _T_174[9:0] ? 4'h3 : _GEN_10188; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10190 = 10'h1af == _T_174[9:0] ? 4'h4 : _GEN_10189; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10191 = 10'h1b0 == _T_174[9:0] ? 4'h6 : _GEN_10190; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10192 = 10'h1b1 == _T_174[9:0] ? 4'ha : _GEN_10191; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10193 = 10'h1b2 == _T_174[9:0] ? 4'ha : _GEN_10192; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10194 = 10'h1b3 == _T_174[9:0] ? 4'h9 : _GEN_10193; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10195 = 10'h1b4 == _T_174[9:0] ? 4'h9 : _GEN_10194; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10196 = 10'h1b5 == _T_174[9:0] ? 4'h3 : _GEN_10195; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10197 = 10'h1b6 == _T_174[9:0] ? 4'h3 : _GEN_10196; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10198 = 10'h1b7 == _T_174[9:0] ? 4'h4 : _GEN_10197; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10199 = 10'h1b8 == _T_174[9:0] ? 4'h5 : _GEN_10198; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10200 = 10'h1b9 == _T_174[9:0] ? 4'h6 : _GEN_10199; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10201 = 10'h1ba == _T_174[9:0] ? 4'h4 : _GEN_10200; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10202 = 10'h1bb == _T_174[9:0] ? 4'h3 : _GEN_10201; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10203 = 10'h1bc == _T_174[9:0] ? 4'h3 : _GEN_10202; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10204 = 10'h1bd == _T_174[9:0] ? 4'h4 : _GEN_10203; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10205 = 10'h1be == _T_174[9:0] ? 4'ha : _GEN_10204; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10206 = 10'h1bf == _T_174[9:0] ? 4'h4 : _GEN_10205; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10207 = 10'h1c0 == _T_174[9:0] ? 4'h5 : _GEN_10206; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10208 = 10'h1c1 == _T_174[9:0] ? 4'h5 : _GEN_10207; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10209 = 10'h1c2 == _T_174[9:0] ? 4'h4 : _GEN_10208; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10210 = 10'h1c3 == _T_174[9:0] ? 4'h5 : _GEN_10209; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10211 = 10'h1c4 == _T_174[9:0] ? 4'h4 : _GEN_10210; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10212 = 10'h1c5 == _T_174[9:0] ? 4'h3 : _GEN_10211; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10213 = 10'h1c6 == _T_174[9:0] ? 4'h4 : _GEN_10212; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10214 = 10'h1c7 == _T_174[9:0] ? 4'h3 : _GEN_10213; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10215 = 10'h1c8 == _T_174[9:0] ? 4'h8 : _GEN_10214; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10216 = 10'h1c9 == _T_174[9:0] ? 4'h8 : _GEN_10215; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10217 = 10'h1ca == _T_174[9:0] ? 4'h8 : _GEN_10216; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10218 = 10'h1cb == _T_174[9:0] ? 4'h8 : _GEN_10217; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10219 = 10'h1cc == _T_174[9:0] ? 4'h8 : _GEN_10218; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10220 = 10'h1cd == _T_174[9:0] ? 4'h8 : _GEN_10219; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10221 = 10'h1ce == _T_174[9:0] ? 4'h8 : _GEN_10220; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10222 = 10'h1cf == _T_174[9:0] ? 4'h8 : _GEN_10221; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10223 = 10'h1d0 == _T_174[9:0] ? 4'h5 : _GEN_10222; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10224 = 10'h1d1 == _T_174[9:0] ? 4'h4 : _GEN_10223; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10225 = 10'h1d2 == _T_174[9:0] ? 4'h6 : _GEN_10224; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10226 = 10'h1d3 == _T_174[9:0] ? 4'h6 : _GEN_10225; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10227 = 10'h1d4 == _T_174[9:0] ? 4'h6 : _GEN_10226; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10228 = 10'h1d5 == _T_174[9:0] ? 4'h5 : _GEN_10227; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10229 = 10'h1d6 == _T_174[9:0] ? 4'h8 : _GEN_10228; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10230 = 10'h1d7 == _T_174[9:0] ? 4'ha : _GEN_10229; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10231 = 10'h1d8 == _T_174[9:0] ? 4'ha : _GEN_10230; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10232 = 10'h1d9 == _T_174[9:0] ? 4'ha : _GEN_10231; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10233 = 10'h1da == _T_174[9:0] ? 4'h6 : _GEN_10232; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10234 = 10'h1db == _T_174[9:0] ? 4'h3 : _GEN_10233; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10235 = 10'h1dc == _T_174[9:0] ? 4'h5 : _GEN_10234; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10236 = 10'h1dd == _T_174[9:0] ? 4'h2 : _GEN_10235; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10237 = 10'h1de == _T_174[9:0] ? 4'h5 : _GEN_10236; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10238 = 10'h1df == _T_174[9:0] ? 4'h5 : _GEN_10237; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10239 = 10'h1e0 == _T_174[9:0] ? 4'h5 : _GEN_10238; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10240 = 10'h1e1 == _T_174[9:0] ? 4'h3 : _GEN_10239; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10241 = 10'h1e2 == _T_174[9:0] ? 4'h3 : _GEN_10240; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10242 = 10'h1e3 == _T_174[9:0] ? 4'h3 : _GEN_10241; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10243 = 10'h1e4 == _T_174[9:0] ? 4'h9 : _GEN_10242; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10244 = 10'h1e5 == _T_174[9:0] ? 4'h4 : _GEN_10243; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10245 = 10'h1e6 == _T_174[9:0] ? 4'h4 : _GEN_10244; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10246 = 10'h1e7 == _T_174[9:0] ? 4'h4 : _GEN_10245; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10247 = 10'h1e8 == _T_174[9:0] ? 4'h4 : _GEN_10246; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10248 = 10'h1e9 == _T_174[9:0] ? 4'h4 : _GEN_10247; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10249 = 10'h1ea == _T_174[9:0] ? 4'h4 : _GEN_10248; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10250 = 10'h1eb == _T_174[9:0] ? 4'h4 : _GEN_10249; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10251 = 10'h1ec == _T_174[9:0] ? 4'h4 : _GEN_10250; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10252 = 10'h1ed == _T_174[9:0] ? 4'h4 : _GEN_10251; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10253 = 10'h1ee == _T_174[9:0] ? 4'h8 : _GEN_10252; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10254 = 10'h1ef == _T_174[9:0] ? 4'h8 : _GEN_10253; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10255 = 10'h1f0 == _T_174[9:0] ? 4'h8 : _GEN_10254; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10256 = 10'h1f1 == _T_174[9:0] ? 4'h8 : _GEN_10255; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10257 = 10'h1f2 == _T_174[9:0] ? 4'h8 : _GEN_10256; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10258 = 10'h1f3 == _T_174[9:0] ? 4'h8 : _GEN_10257; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10259 = 10'h1f4 == _T_174[9:0] ? 4'h9 : _GEN_10258; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10260 = 10'h1f5 == _T_174[9:0] ? 4'h9 : _GEN_10259; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10261 = 10'h1f6 == _T_174[9:0] ? 4'ha : _GEN_10260; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10262 = 10'h1f7 == _T_174[9:0] ? 4'h5 : _GEN_10261; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10263 = 10'h1f8 == _T_174[9:0] ? 4'h5 : _GEN_10262; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10264 = 10'h1f9 == _T_174[9:0] ? 4'h7 : _GEN_10263; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10265 = 10'h1fa == _T_174[9:0] ? 4'h7 : _GEN_10264; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10266 = 10'h1fb == _T_174[9:0] ? 4'h5 : _GEN_10265; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10267 = 10'h1fc == _T_174[9:0] ? 4'ha : _GEN_10266; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10268 = 10'h1fd == _T_174[9:0] ? 4'hb : _GEN_10267; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10269 = 10'h1fe == _T_174[9:0] ? 4'hb : _GEN_10268; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10270 = 10'h1ff == _T_174[9:0] ? 4'ha : _GEN_10269; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10271 = 10'h200 == _T_174[9:0] ? 4'h4 : _GEN_10270; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10272 = 10'h201 == _T_174[9:0] ? 4'h3 : _GEN_10271; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10273 = 10'h202 == _T_174[9:0] ? 4'h2 : _GEN_10272; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10274 = 10'h203 == _T_174[9:0] ? 4'h2 : _GEN_10273; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10275 = 10'h204 == _T_174[9:0] ? 4'h2 : _GEN_10274; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10276 = 10'h205 == _T_174[9:0] ? 4'h2 : _GEN_10275; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10277 = 10'h206 == _T_174[9:0] ? 4'h2 : _GEN_10276; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10278 = 10'h207 == _T_174[9:0] ? 4'h2 : _GEN_10277; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10279 = 10'h208 == _T_174[9:0] ? 4'h3 : _GEN_10278; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10280 = 10'h209 == _T_174[9:0] ? 4'h3 : _GEN_10279; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10281 = 10'h20a == _T_174[9:0] ? 4'h8 : _GEN_10280; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10282 = 10'h20b == _T_174[9:0] ? 4'h4 : _GEN_10281; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10283 = 10'h20c == _T_174[9:0] ? 4'h4 : _GEN_10282; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10284 = 10'h20d == _T_174[9:0] ? 4'h4 : _GEN_10283; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10285 = 10'h20e == _T_174[9:0] ? 4'h4 : _GEN_10284; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10286 = 10'h20f == _T_174[9:0] ? 4'h4 : _GEN_10285; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10287 = 10'h210 == _T_174[9:0] ? 4'h4 : _GEN_10286; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10288 = 10'h211 == _T_174[9:0] ? 4'h4 : _GEN_10287; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10289 = 10'h212 == _T_174[9:0] ? 4'h4 : _GEN_10288; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10290 = 10'h213 == _T_174[9:0] ? 4'h6 : _GEN_10289; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10291 = 10'h214 == _T_174[9:0] ? 4'h7 : _GEN_10290; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10292 = 10'h215 == _T_174[9:0] ? 4'h8 : _GEN_10291; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10293 = 10'h216 == _T_174[9:0] ? 4'h8 : _GEN_10292; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10294 = 10'h217 == _T_174[9:0] ? 4'h8 : _GEN_10293; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10295 = 10'h218 == _T_174[9:0] ? 4'h8 : _GEN_10294; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10296 = 10'h219 == _T_174[9:0] ? 4'h8 : _GEN_10295; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10297 = 10'h21a == _T_174[9:0] ? 4'h8 : _GEN_10296; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10298 = 10'h21b == _T_174[9:0] ? 4'h8 : _GEN_10297; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10299 = 10'h21c == _T_174[9:0] ? 4'ha : _GEN_10298; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10300 = 10'h21d == _T_174[9:0] ? 4'h9 : _GEN_10299; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10301 = 10'h21e == _T_174[9:0] ? 4'h6 : _GEN_10300; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10302 = 10'h21f == _T_174[9:0] ? 4'h4 : _GEN_10301; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10303 = 10'h220 == _T_174[9:0] ? 4'h4 : _GEN_10302; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10304 = 10'h221 == _T_174[9:0] ? 4'h5 : _GEN_10303; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10305 = 10'h222 == _T_174[9:0] ? 4'ha : _GEN_10304; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10306 = 10'h223 == _T_174[9:0] ? 4'ha : _GEN_10305; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10307 = 10'h224 == _T_174[9:0] ? 4'ha : _GEN_10306; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10308 = 10'h225 == _T_174[9:0] ? 4'h8 : _GEN_10307; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10309 = 10'h226 == _T_174[9:0] ? 4'h4 : _GEN_10308; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10310 = 10'h227 == _T_174[9:0] ? 4'h2 : _GEN_10309; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10311 = 10'h228 == _T_174[9:0] ? 4'h2 : _GEN_10310; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10312 = 10'h229 == _T_174[9:0] ? 4'h2 : _GEN_10311; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10313 = 10'h22a == _T_174[9:0] ? 4'h2 : _GEN_10312; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10314 = 10'h22b == _T_174[9:0] ? 4'h2 : _GEN_10313; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10315 = 10'h22c == _T_174[9:0] ? 4'h2 : _GEN_10314; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10316 = 10'h22d == _T_174[9:0] ? 4'h2 : _GEN_10315; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10317 = 10'h22e == _T_174[9:0] ? 4'h2 : _GEN_10316; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10318 = 10'h22f == _T_174[9:0] ? 4'h3 : _GEN_10317; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10319 = 10'h230 == _T_174[9:0] ? 4'h3 : _GEN_10318; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10320 = 10'h231 == _T_174[9:0] ? 4'h3 : _GEN_10319; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10321 = 10'h232 == _T_174[9:0] ? 4'h4 : _GEN_10320; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10322 = 10'h233 == _T_174[9:0] ? 4'h6 : _GEN_10321; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10323 = 10'h234 == _T_174[9:0] ? 4'h6 : _GEN_10322; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10324 = 10'h235 == _T_174[9:0] ? 4'h4 : _GEN_10323; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10325 = 10'h236 == _T_174[9:0] ? 4'h4 : _GEN_10324; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10326 = 10'h237 == _T_174[9:0] ? 4'h4 : _GEN_10325; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10327 = 10'h238 == _T_174[9:0] ? 4'h4 : _GEN_10326; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10328 = 10'h239 == _T_174[9:0] ? 4'h3 : _GEN_10327; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10329 = 10'h23a == _T_174[9:0] ? 4'h7 : _GEN_10328; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10330 = 10'h23b == _T_174[9:0] ? 4'h7 : _GEN_10329; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10331 = 10'h23c == _T_174[9:0] ? 4'h7 : _GEN_10330; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10332 = 10'h23d == _T_174[9:0] ? 4'h7 : _GEN_10331; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10333 = 10'h23e == _T_174[9:0] ? 4'h7 : _GEN_10332; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10334 = 10'h23f == _T_174[9:0] ? 4'h7 : _GEN_10333; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10335 = 10'h240 == _T_174[9:0] ? 4'h7 : _GEN_10334; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10336 = 10'h241 == _T_174[9:0] ? 4'h8 : _GEN_10335; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10337 = 10'h242 == _T_174[9:0] ? 4'ha : _GEN_10336; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10338 = 10'h243 == _T_174[9:0] ? 4'ha : _GEN_10337; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10339 = 10'h244 == _T_174[9:0] ? 4'ha : _GEN_10338; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10340 = 10'h245 == _T_174[9:0] ? 4'h8 : _GEN_10339; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10341 = 10'h246 == _T_174[9:0] ? 4'h7 : _GEN_10340; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10342 = 10'h247 == _T_174[9:0] ? 4'h8 : _GEN_10341; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10343 = 10'h248 == _T_174[9:0] ? 4'ha : _GEN_10342; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10344 = 10'h249 == _T_174[9:0] ? 4'ha : _GEN_10343; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10345 = 10'h24a == _T_174[9:0] ? 4'ha : _GEN_10344; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10346 = 10'h24b == _T_174[9:0] ? 4'h4 : _GEN_10345; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10347 = 10'h24c == _T_174[9:0] ? 4'h4 : _GEN_10346; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10348 = 10'h24d == _T_174[9:0] ? 4'h2 : _GEN_10347; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10349 = 10'h24e == _T_174[9:0] ? 4'h2 : _GEN_10348; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10350 = 10'h24f == _T_174[9:0] ? 4'h2 : _GEN_10349; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10351 = 10'h250 == _T_174[9:0] ? 4'h2 : _GEN_10350; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10352 = 10'h251 == _T_174[9:0] ? 4'h2 : _GEN_10351; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10353 = 10'h252 == _T_174[9:0] ? 4'h2 : _GEN_10352; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10354 = 10'h253 == _T_174[9:0] ? 4'h2 : _GEN_10353; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10355 = 10'h254 == _T_174[9:0] ? 4'h2 : _GEN_10354; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10356 = 10'h255 == _T_174[9:0] ? 4'h3 : _GEN_10355; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10357 = 10'h256 == _T_174[9:0] ? 4'h4 : _GEN_10356; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10358 = 10'h257 == _T_174[9:0] ? 4'h3 : _GEN_10357; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10359 = 10'h258 == _T_174[9:0] ? 4'h4 : _GEN_10358; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10360 = 10'h259 == _T_174[9:0] ? 4'h4 : _GEN_10359; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10361 = 10'h25a == _T_174[9:0] ? 4'h4 : _GEN_10360; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10362 = 10'h25b == _T_174[9:0] ? 4'h3 : _GEN_10361; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10363 = 10'h25c == _T_174[9:0] ? 4'h4 : _GEN_10362; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10364 = 10'h25d == _T_174[9:0] ? 4'h4 : _GEN_10363; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10365 = 10'h25e == _T_174[9:0] ? 4'h3 : _GEN_10364; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10366 = 10'h25f == _T_174[9:0] ? 4'h3 : _GEN_10365; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10367 = 10'h260 == _T_174[9:0] ? 4'h8 : _GEN_10366; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10368 = 10'h261 == _T_174[9:0] ? 4'h7 : _GEN_10367; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10369 = 10'h262 == _T_174[9:0] ? 4'h6 : _GEN_10368; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10370 = 10'h263 == _T_174[9:0] ? 4'h5 : _GEN_10369; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10371 = 10'h264 == _T_174[9:0] ? 4'h6 : _GEN_10370; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10372 = 10'h265 == _T_174[9:0] ? 4'h5 : _GEN_10371; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10373 = 10'h266 == _T_174[9:0] ? 4'h5 : _GEN_10372; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10374 = 10'h267 == _T_174[9:0] ? 4'h7 : _GEN_10373; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10375 = 10'h268 == _T_174[9:0] ? 4'ha : _GEN_10374; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10376 = 10'h269 == _T_174[9:0] ? 4'ha : _GEN_10375; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10377 = 10'h26a == _T_174[9:0] ? 4'ha : _GEN_10376; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10378 = 10'h26b == _T_174[9:0] ? 4'ha : _GEN_10377; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10379 = 10'h26c == _T_174[9:0] ? 4'ha : _GEN_10378; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10380 = 10'h26d == _T_174[9:0] ? 4'ha : _GEN_10379; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10381 = 10'h26e == _T_174[9:0] ? 4'ha : _GEN_10380; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10382 = 10'h26f == _T_174[9:0] ? 4'ha : _GEN_10381; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10383 = 10'h270 == _T_174[9:0] ? 4'h5 : _GEN_10382; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10384 = 10'h271 == _T_174[9:0] ? 4'h4 : _GEN_10383; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10385 = 10'h272 == _T_174[9:0] ? 4'h3 : _GEN_10384; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10386 = 10'h273 == _T_174[9:0] ? 4'h2 : _GEN_10385; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10387 = 10'h274 == _T_174[9:0] ? 4'h2 : _GEN_10386; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10388 = 10'h275 == _T_174[9:0] ? 4'h2 : _GEN_10387; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10389 = 10'h276 == _T_174[9:0] ? 4'h2 : _GEN_10388; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10390 = 10'h277 == _T_174[9:0] ? 4'h2 : _GEN_10389; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10391 = 10'h278 == _T_174[9:0] ? 4'h2 : _GEN_10390; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10392 = 10'h279 == _T_174[9:0] ? 4'h2 : _GEN_10391; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10393 = 10'h27a == _T_174[9:0] ? 4'h2 : _GEN_10392; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10394 = 10'h27b == _T_174[9:0] ? 4'h4 : _GEN_10393; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10395 = 10'h27c == _T_174[9:0] ? 4'h3 : _GEN_10394; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10396 = 10'h27d == _T_174[9:0] ? 4'h4 : _GEN_10395; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10397 = 10'h27e == _T_174[9:0] ? 4'h5 : _GEN_10396; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10398 = 10'h27f == _T_174[9:0] ? 4'h4 : _GEN_10397; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10399 = 10'h280 == _T_174[9:0] ? 4'h4 : _GEN_10398; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10400 = 10'h281 == _T_174[9:0] ? 4'h4 : _GEN_10399; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10401 = 10'h282 == _T_174[9:0] ? 4'h4 : _GEN_10400; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10402 = 10'h283 == _T_174[9:0] ? 4'h3 : _GEN_10401; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10403 = 10'h284 == _T_174[9:0] ? 4'h3 : _GEN_10402; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10404 = 10'h285 == _T_174[9:0] ? 4'h3 : _GEN_10403; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10405 = 10'h286 == _T_174[9:0] ? 4'h8 : _GEN_10404; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10406 = 10'h287 == _T_174[9:0] ? 4'h6 : _GEN_10405; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10407 = 10'h288 == _T_174[9:0] ? 4'h6 : _GEN_10406; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10408 = 10'h289 == _T_174[9:0] ? 4'h6 : _GEN_10407; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10409 = 10'h28a == _T_174[9:0] ? 4'h7 : _GEN_10408; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10410 = 10'h28b == _T_174[9:0] ? 4'h7 : _GEN_10409; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10411 = 10'h28c == _T_174[9:0] ? 4'h6 : _GEN_10410; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10412 = 10'h28d == _T_174[9:0] ? 4'h6 : _GEN_10411; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10413 = 10'h28e == _T_174[9:0] ? 4'h4 : _GEN_10412; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10414 = 10'h28f == _T_174[9:0] ? 4'h7 : _GEN_10413; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10415 = 10'h290 == _T_174[9:0] ? 4'h9 : _GEN_10414; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10416 = 10'h291 == _T_174[9:0] ? 4'ha : _GEN_10415; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10417 = 10'h292 == _T_174[9:0] ? 4'ha : _GEN_10416; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10418 = 10'h293 == _T_174[9:0] ? 4'ha : _GEN_10417; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10419 = 10'h294 == _T_174[9:0] ? 4'h9 : _GEN_10418; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10420 = 10'h295 == _T_174[9:0] ? 4'h5 : _GEN_10419; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10421 = 10'h296 == _T_174[9:0] ? 4'h4 : _GEN_10420; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10422 = 10'h297 == _T_174[9:0] ? 4'h4 : _GEN_10421; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10423 = 10'h298 == _T_174[9:0] ? 4'h3 : _GEN_10422; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10424 = 10'h299 == _T_174[9:0] ? 4'h3 : _GEN_10423; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10425 = 10'h29a == _T_174[9:0] ? 4'h2 : _GEN_10424; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10426 = 10'h29b == _T_174[9:0] ? 4'h2 : _GEN_10425; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10427 = 10'h29c == _T_174[9:0] ? 4'h2 : _GEN_10426; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10428 = 10'h29d == _T_174[9:0] ? 4'h2 : _GEN_10427; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10429 = 10'h29e == _T_174[9:0] ? 4'h2 : _GEN_10428; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10430 = 10'h29f == _T_174[9:0] ? 4'h2 : _GEN_10429; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10431 = 10'h2a0 == _T_174[9:0] ? 4'h2 : _GEN_10430; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10432 = 10'h2a1 == _T_174[9:0] ? 4'h4 : _GEN_10431; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10433 = 10'h2a2 == _T_174[9:0] ? 4'h3 : _GEN_10432; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10434 = 10'h2a3 == _T_174[9:0] ? 4'h4 : _GEN_10433; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10435 = 10'h2a4 == _T_174[9:0] ? 4'h5 : _GEN_10434; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10436 = 10'h2a5 == _T_174[9:0] ? 4'h4 : _GEN_10435; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10437 = 10'h2a6 == _T_174[9:0] ? 4'h4 : _GEN_10436; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10438 = 10'h2a7 == _T_174[9:0] ? 4'h4 : _GEN_10437; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10439 = 10'h2a8 == _T_174[9:0] ? 4'h3 : _GEN_10438; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10440 = 10'h2a9 == _T_174[9:0] ? 4'h3 : _GEN_10439; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10441 = 10'h2aa == _T_174[9:0] ? 4'h3 : _GEN_10440; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10442 = 10'h2ab == _T_174[9:0] ? 4'h3 : _GEN_10441; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10443 = 10'h2ac == _T_174[9:0] ? 4'h8 : _GEN_10442; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10444 = 10'h2ad == _T_174[9:0] ? 4'h7 : _GEN_10443; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10445 = 10'h2ae == _T_174[9:0] ? 4'h5 : _GEN_10444; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10446 = 10'h2af == _T_174[9:0] ? 4'h6 : _GEN_10445; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10447 = 10'h2b0 == _T_174[9:0] ? 4'h7 : _GEN_10446; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10448 = 10'h2b1 == _T_174[9:0] ? 4'h6 : _GEN_10447; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10449 = 10'h2b2 == _T_174[9:0] ? 4'h6 : _GEN_10448; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10450 = 10'h2b3 == _T_174[9:0] ? 4'h6 : _GEN_10449; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10451 = 10'h2b4 == _T_174[9:0] ? 4'h3 : _GEN_10450; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10452 = 10'h2b5 == _T_174[9:0] ? 4'h3 : _GEN_10451; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10453 = 10'h2b6 == _T_174[9:0] ? 4'h3 : _GEN_10452; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10454 = 10'h2b7 == _T_174[9:0] ? 4'h4 : _GEN_10453; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10455 = 10'h2b8 == _T_174[9:0] ? 4'h6 : _GEN_10454; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10456 = 10'h2b9 == _T_174[9:0] ? 4'h9 : _GEN_10455; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10457 = 10'h2ba == _T_174[9:0] ? 4'h4 : _GEN_10456; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10458 = 10'h2bb == _T_174[9:0] ? 4'h3 : _GEN_10457; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10459 = 10'h2bc == _T_174[9:0] ? 4'h4 : _GEN_10458; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10460 = 10'h2bd == _T_174[9:0] ? 4'h3 : _GEN_10459; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10461 = 10'h2be == _T_174[9:0] ? 4'h3 : _GEN_10460; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10462 = 10'h2bf == _T_174[9:0] ? 4'h3 : _GEN_10461; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10463 = 10'h2c0 == _T_174[9:0] ? 4'h2 : _GEN_10462; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10464 = 10'h2c1 == _T_174[9:0] ? 4'h2 : _GEN_10463; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10465 = 10'h2c2 == _T_174[9:0] ? 4'h2 : _GEN_10464; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10466 = 10'h2c3 == _T_174[9:0] ? 4'h2 : _GEN_10465; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10467 = 10'h2c4 == _T_174[9:0] ? 4'h2 : _GEN_10466; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10468 = 10'h2c5 == _T_174[9:0] ? 4'h2 : _GEN_10467; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10469 = 10'h2c6 == _T_174[9:0] ? 4'h2 : _GEN_10468; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10470 = 10'h2c7 == _T_174[9:0] ? 4'h4 : _GEN_10469; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10471 = 10'h2c8 == _T_174[9:0] ? 4'h3 : _GEN_10470; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10472 = 10'h2c9 == _T_174[9:0] ? 4'h4 : _GEN_10471; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10473 = 10'h2ca == _T_174[9:0] ? 4'h5 : _GEN_10472; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10474 = 10'h2cb == _T_174[9:0] ? 4'h3 : _GEN_10473; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10475 = 10'h2cc == _T_174[9:0] ? 4'h3 : _GEN_10474; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10476 = 10'h2cd == _T_174[9:0] ? 4'h3 : _GEN_10475; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10477 = 10'h2ce == _T_174[9:0] ? 4'h3 : _GEN_10476; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10478 = 10'h2cf == _T_174[9:0] ? 4'h3 : _GEN_10477; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10479 = 10'h2d0 == _T_174[9:0] ? 4'h3 : _GEN_10478; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10480 = 10'h2d1 == _T_174[9:0] ? 4'h3 : _GEN_10479; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10481 = 10'h2d2 == _T_174[9:0] ? 4'h8 : _GEN_10480; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10482 = 10'h2d3 == _T_174[9:0] ? 4'h6 : _GEN_10481; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10483 = 10'h2d4 == _T_174[9:0] ? 4'h6 : _GEN_10482; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10484 = 10'h2d5 == _T_174[9:0] ? 4'h7 : _GEN_10483; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10485 = 10'h2d6 == _T_174[9:0] ? 4'h7 : _GEN_10484; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10486 = 10'h2d7 == _T_174[9:0] ? 4'h7 : _GEN_10485; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10487 = 10'h2d8 == _T_174[9:0] ? 4'h6 : _GEN_10486; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10488 = 10'h2d9 == _T_174[9:0] ? 4'h7 : _GEN_10487; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10489 = 10'h2da == _T_174[9:0] ? 4'h5 : _GEN_10488; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10490 = 10'h2db == _T_174[9:0] ? 4'h3 : _GEN_10489; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10491 = 10'h2dc == _T_174[9:0] ? 4'h3 : _GEN_10490; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10492 = 10'h2dd == _T_174[9:0] ? 4'h3 : _GEN_10491; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10493 = 10'h2de == _T_174[9:0] ? 4'h3 : _GEN_10492; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10494 = 10'h2df == _T_174[9:0] ? 4'h4 : _GEN_10493; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10495 = 10'h2e0 == _T_174[9:0] ? 4'h3 : _GEN_10494; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10496 = 10'h2e1 == _T_174[9:0] ? 4'h3 : _GEN_10495; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10497 = 10'h2e2 == _T_174[9:0] ? 4'h3 : _GEN_10496; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10498 = 10'h2e3 == _T_174[9:0] ? 4'h3 : _GEN_10497; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10499 = 10'h2e4 == _T_174[9:0] ? 4'h3 : _GEN_10498; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10500 = 10'h2e5 == _T_174[9:0] ? 4'h3 : _GEN_10499; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10501 = 10'h2e6 == _T_174[9:0] ? 4'h2 : _GEN_10500; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10502 = 10'h2e7 == _T_174[9:0] ? 4'h2 : _GEN_10501; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10503 = 10'h2e8 == _T_174[9:0] ? 4'h2 : _GEN_10502; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10504 = 10'h2e9 == _T_174[9:0] ? 4'h2 : _GEN_10503; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10505 = 10'h2ea == _T_174[9:0] ? 4'h2 : _GEN_10504; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10506 = 10'h2eb == _T_174[9:0] ? 4'h2 : _GEN_10505; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10507 = 10'h2ec == _T_174[9:0] ? 4'h3 : _GEN_10506; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10508 = 10'h2ed == _T_174[9:0] ? 4'h4 : _GEN_10507; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10509 = 10'h2ee == _T_174[9:0] ? 4'h3 : _GEN_10508; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10510 = 10'h2ef == _T_174[9:0] ? 4'h3 : _GEN_10509; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10511 = 10'h2f0 == _T_174[9:0] ? 4'h6 : _GEN_10510; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10512 = 10'h2f1 == _T_174[9:0] ? 4'h3 : _GEN_10511; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10513 = 10'h2f2 == _T_174[9:0] ? 4'h3 : _GEN_10512; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10514 = 10'h2f3 == _T_174[9:0] ? 4'h3 : _GEN_10513; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10515 = 10'h2f4 == _T_174[9:0] ? 4'h3 : _GEN_10514; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10516 = 10'h2f5 == _T_174[9:0] ? 4'h3 : _GEN_10515; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10517 = 10'h2f6 == _T_174[9:0] ? 4'h3 : _GEN_10516; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10518 = 10'h2f7 == _T_174[9:0] ? 4'h3 : _GEN_10517; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10519 = 10'h2f8 == _T_174[9:0] ? 4'h8 : _GEN_10518; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10520 = 10'h2f9 == _T_174[9:0] ? 4'h6 : _GEN_10519; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10521 = 10'h2fa == _T_174[9:0] ? 4'h7 : _GEN_10520; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10522 = 10'h2fb == _T_174[9:0] ? 4'h7 : _GEN_10521; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10523 = 10'h2fc == _T_174[9:0] ? 4'h6 : _GEN_10522; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10524 = 10'h2fd == _T_174[9:0] ? 4'h6 : _GEN_10523; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10525 = 10'h2fe == _T_174[9:0] ? 4'h6 : _GEN_10524; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10526 = 10'h2ff == _T_174[9:0] ? 4'h8 : _GEN_10525; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10527 = 10'h300 == _T_174[9:0] ? 4'h9 : _GEN_10526; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10528 = 10'h301 == _T_174[9:0] ? 4'h7 : _GEN_10527; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10529 = 10'h302 == _T_174[9:0] ? 4'h4 : _GEN_10528; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10530 = 10'h303 == _T_174[9:0] ? 4'h4 : _GEN_10529; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10531 = 10'h304 == _T_174[9:0] ? 4'h3 : _GEN_10530; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10532 = 10'h305 == _T_174[9:0] ? 4'h3 : _GEN_10531; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10533 = 10'h306 == _T_174[9:0] ? 4'h3 : _GEN_10532; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10534 = 10'h307 == _T_174[9:0] ? 4'h3 : _GEN_10533; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10535 = 10'h308 == _T_174[9:0] ? 4'h3 : _GEN_10534; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10536 = 10'h309 == _T_174[9:0] ? 4'h3 : _GEN_10535; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10537 = 10'h30a == _T_174[9:0] ? 4'h3 : _GEN_10536; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10538 = 10'h30b == _T_174[9:0] ? 4'h3 : _GEN_10537; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10539 = 10'h30c == _T_174[9:0] ? 4'h2 : _GEN_10538; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10540 = 10'h30d == _T_174[9:0] ? 4'h2 : _GEN_10539; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10541 = 10'h30e == _T_174[9:0] ? 4'h2 : _GEN_10540; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10542 = 10'h30f == _T_174[9:0] ? 4'h2 : _GEN_10541; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10543 = 10'h310 == _T_174[9:0] ? 4'h2 : _GEN_10542; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10544 = 10'h311 == _T_174[9:0] ? 4'h2 : _GEN_10543; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10545 = 10'h312 == _T_174[9:0] ? 4'h3 : _GEN_10544; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10546 = 10'h313 == _T_174[9:0] ? 4'h4 : _GEN_10545; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10547 = 10'h314 == _T_174[9:0] ? 4'h3 : _GEN_10546; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10548 = 10'h315 == _T_174[9:0] ? 4'h3 : _GEN_10547; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10549 = 10'h316 == _T_174[9:0] ? 4'h5 : _GEN_10548; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10550 = 10'h317 == _T_174[9:0] ? 4'h5 : _GEN_10549; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10551 = 10'h318 == _T_174[9:0] ? 4'h3 : _GEN_10550; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10552 = 10'h319 == _T_174[9:0] ? 4'h3 : _GEN_10551; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10553 = 10'h31a == _T_174[9:0] ? 4'h3 : _GEN_10552; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10554 = 10'h31b == _T_174[9:0] ? 4'h3 : _GEN_10553; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10555 = 10'h31c == _T_174[9:0] ? 4'h3 : _GEN_10554; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10556 = 10'h31d == _T_174[9:0] ? 4'h3 : _GEN_10555; // @[Filter.scala 230:62]
  wire [4:0] _GEN_38978 = {{1'd0}, _GEN_10556}; // @[Filter.scala 230:62]
  wire [8:0] _T_176 = _GEN_38978 * 5'h14; // @[Filter.scala 230:62]
  wire [3:0] _GEN_10580 = 10'h17 == _T_174[9:0] ? 4'hb : 4'he; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10581 = 10'h18 == _T_174[9:0] ? 4'hc : _GEN_10580; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10582 = 10'h19 == _T_174[9:0] ? 4'he : _GEN_10581; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10583 = 10'h1a == _T_174[9:0] ? 4'he : _GEN_10582; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10584 = 10'h1b == _T_174[9:0] ? 4'he : _GEN_10583; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10585 = 10'h1c == _T_174[9:0] ? 4'he : _GEN_10584; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10586 = 10'h1d == _T_174[9:0] ? 4'he : _GEN_10585; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10587 = 10'h1e == _T_174[9:0] ? 4'he : _GEN_10586; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10588 = 10'h1f == _T_174[9:0] ? 4'he : _GEN_10587; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10589 = 10'h20 == _T_174[9:0] ? 4'he : _GEN_10588; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10590 = 10'h21 == _T_174[9:0] ? 4'he : _GEN_10589; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10591 = 10'h22 == _T_174[9:0] ? 4'he : _GEN_10590; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10592 = 10'h23 == _T_174[9:0] ? 4'he : _GEN_10591; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10593 = 10'h24 == _T_174[9:0] ? 4'he : _GEN_10592; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10594 = 10'h25 == _T_174[9:0] ? 4'he : _GEN_10593; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10595 = 10'h26 == _T_174[9:0] ? 4'he : _GEN_10594; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10596 = 10'h27 == _T_174[9:0] ? 4'he : _GEN_10595; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10597 = 10'h28 == _T_174[9:0] ? 4'he : _GEN_10596; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10598 = 10'h29 == _T_174[9:0] ? 4'he : _GEN_10597; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10599 = 10'h2a == _T_174[9:0] ? 4'he : _GEN_10598; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10600 = 10'h2b == _T_174[9:0] ? 4'he : _GEN_10599; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10601 = 10'h2c == _T_174[9:0] ? 4'he : _GEN_10600; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10602 = 10'h2d == _T_174[9:0] ? 4'he : _GEN_10601; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10603 = 10'h2e == _T_174[9:0] ? 4'he : _GEN_10602; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10604 = 10'h2f == _T_174[9:0] ? 4'he : _GEN_10603; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10605 = 10'h30 == _T_174[9:0] ? 4'he : _GEN_10604; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10606 = 10'h31 == _T_174[9:0] ? 4'he : _GEN_10605; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10607 = 10'h32 == _T_174[9:0] ? 4'he : _GEN_10606; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10608 = 10'h33 == _T_174[9:0] ? 4'he : _GEN_10607; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10609 = 10'h34 == _T_174[9:0] ? 4'he : _GEN_10608; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10610 = 10'h35 == _T_174[9:0] ? 4'he : _GEN_10609; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10611 = 10'h36 == _T_174[9:0] ? 4'he : _GEN_10610; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10612 = 10'h37 == _T_174[9:0] ? 4'he : _GEN_10611; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10613 = 10'h38 == _T_174[9:0] ? 4'he : _GEN_10612; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10614 = 10'h39 == _T_174[9:0] ? 4'he : _GEN_10613; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10615 = 10'h3a == _T_174[9:0] ? 4'he : _GEN_10614; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10616 = 10'h3b == _T_174[9:0] ? 4'he : _GEN_10615; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10617 = 10'h3c == _T_174[9:0] ? 4'ha : _GEN_10616; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10618 = 10'h3d == _T_174[9:0] ? 4'hc : _GEN_10617; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10619 = 10'h3e == _T_174[9:0] ? 4'hb : _GEN_10618; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10620 = 10'h3f == _T_174[9:0] ? 4'he : _GEN_10619; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10621 = 10'h40 == _T_174[9:0] ? 4'he : _GEN_10620; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10622 = 10'h41 == _T_174[9:0] ? 4'he : _GEN_10621; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10623 = 10'h42 == _T_174[9:0] ? 4'he : _GEN_10622; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10624 = 10'h43 == _T_174[9:0] ? 4'he : _GEN_10623; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10625 = 10'h44 == _T_174[9:0] ? 4'he : _GEN_10624; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10626 = 10'h45 == _T_174[9:0] ? 4'he : _GEN_10625; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10627 = 10'h46 == _T_174[9:0] ? 4'he : _GEN_10626; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10628 = 10'h47 == _T_174[9:0] ? 4'he : _GEN_10627; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10629 = 10'h48 == _T_174[9:0] ? 4'he : _GEN_10628; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10630 = 10'h49 == _T_174[9:0] ? 4'he : _GEN_10629; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10631 = 10'h4a == _T_174[9:0] ? 4'he : _GEN_10630; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10632 = 10'h4b == _T_174[9:0] ? 4'he : _GEN_10631; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10633 = 10'h4c == _T_174[9:0] ? 4'he : _GEN_10632; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10634 = 10'h4d == _T_174[9:0] ? 4'he : _GEN_10633; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10635 = 10'h4e == _T_174[9:0] ? 4'he : _GEN_10634; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10636 = 10'h4f == _T_174[9:0] ? 4'he : _GEN_10635; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10637 = 10'h50 == _T_174[9:0] ? 4'he : _GEN_10636; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10638 = 10'h51 == _T_174[9:0] ? 4'he : _GEN_10637; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10639 = 10'h52 == _T_174[9:0] ? 4'he : _GEN_10638; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10640 = 10'h53 == _T_174[9:0] ? 4'he : _GEN_10639; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10641 = 10'h54 == _T_174[9:0] ? 4'he : _GEN_10640; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10642 = 10'h55 == _T_174[9:0] ? 4'he : _GEN_10641; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10643 = 10'h56 == _T_174[9:0] ? 4'he : _GEN_10642; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10644 = 10'h57 == _T_174[9:0] ? 4'he : _GEN_10643; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10645 = 10'h58 == _T_174[9:0] ? 4'he : _GEN_10644; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10646 = 10'h59 == _T_174[9:0] ? 4'he : _GEN_10645; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10647 = 10'h5a == _T_174[9:0] ? 4'hc : _GEN_10646; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10648 = 10'h5b == _T_174[9:0] ? 4'hd : _GEN_10647; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10649 = 10'h5c == _T_174[9:0] ? 4'he : _GEN_10648; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10650 = 10'h5d == _T_174[9:0] ? 4'he : _GEN_10649; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10651 = 10'h5e == _T_174[9:0] ? 4'he : _GEN_10650; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10652 = 10'h5f == _T_174[9:0] ? 4'he : _GEN_10651; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10653 = 10'h60 == _T_174[9:0] ? 4'he : _GEN_10652; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10654 = 10'h61 == _T_174[9:0] ? 4'hd : _GEN_10653; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10655 = 10'h62 == _T_174[9:0] ? 4'hb : _GEN_10654; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10656 = 10'h63 == _T_174[9:0] ? 4'hc : _GEN_10655; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10657 = 10'h64 == _T_174[9:0] ? 4'ha : _GEN_10656; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10658 = 10'h65 == _T_174[9:0] ? 4'hd : _GEN_10657; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10659 = 10'h66 == _T_174[9:0] ? 4'he : _GEN_10658; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10660 = 10'h67 == _T_174[9:0] ? 4'he : _GEN_10659; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10661 = 10'h68 == _T_174[9:0] ? 4'he : _GEN_10660; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10662 = 10'h69 == _T_174[9:0] ? 4'he : _GEN_10661; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10663 = 10'h6a == _T_174[9:0] ? 4'he : _GEN_10662; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10664 = 10'h6b == _T_174[9:0] ? 4'hd : _GEN_10663; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10665 = 10'h6c == _T_174[9:0] ? 4'hc : _GEN_10664; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10666 = 10'h6d == _T_174[9:0] ? 4'hc : _GEN_10665; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10667 = 10'h6e == _T_174[9:0] ? 4'he : _GEN_10666; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10668 = 10'h6f == _T_174[9:0] ? 4'he : _GEN_10667; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10669 = 10'h70 == _T_174[9:0] ? 4'he : _GEN_10668; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10670 = 10'h71 == _T_174[9:0] ? 4'he : _GEN_10669; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10671 = 10'h72 == _T_174[9:0] ? 4'he : _GEN_10670; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10672 = 10'h73 == _T_174[9:0] ? 4'he : _GEN_10671; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10673 = 10'h74 == _T_174[9:0] ? 4'he : _GEN_10672; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10674 = 10'h75 == _T_174[9:0] ? 4'he : _GEN_10673; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10675 = 10'h76 == _T_174[9:0] ? 4'he : _GEN_10674; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10676 = 10'h77 == _T_174[9:0] ? 4'he : _GEN_10675; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10677 = 10'h78 == _T_174[9:0] ? 4'he : _GEN_10676; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10678 = 10'h79 == _T_174[9:0] ? 4'he : _GEN_10677; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10679 = 10'h7a == _T_174[9:0] ? 4'he : _GEN_10678; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10680 = 10'h7b == _T_174[9:0] ? 4'he : _GEN_10679; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10681 = 10'h7c == _T_174[9:0] ? 4'he : _GEN_10680; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10682 = 10'h7d == _T_174[9:0] ? 4'he : _GEN_10681; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10683 = 10'h7e == _T_174[9:0] ? 4'he : _GEN_10682; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10684 = 10'h7f == _T_174[9:0] ? 4'he : _GEN_10683; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10685 = 10'h80 == _T_174[9:0] ? 4'he : _GEN_10684; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10686 = 10'h81 == _T_174[9:0] ? 4'hb : _GEN_10685; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10687 = 10'h82 == _T_174[9:0] ? 4'hc : _GEN_10686; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10688 = 10'h83 == _T_174[9:0] ? 4'hc : _GEN_10687; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10689 = 10'h84 == _T_174[9:0] ? 4'he : _GEN_10688; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10690 = 10'h85 == _T_174[9:0] ? 4'he : _GEN_10689; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10691 = 10'h86 == _T_174[9:0] ? 4'he : _GEN_10690; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10692 = 10'h87 == _T_174[9:0] ? 4'ha : _GEN_10691; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10693 = 10'h88 == _T_174[9:0] ? 4'hd : _GEN_10692; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10694 = 10'h89 == _T_174[9:0] ? 4'hd : _GEN_10693; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10695 = 10'h8a == _T_174[9:0] ? 4'hc : _GEN_10694; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10696 = 10'h8b == _T_174[9:0] ? 4'he : _GEN_10695; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10697 = 10'h8c == _T_174[9:0] ? 4'he : _GEN_10696; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10698 = 10'h8d == _T_174[9:0] ? 4'he : _GEN_10697; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10699 = 10'h8e == _T_174[9:0] ? 4'he : _GEN_10698; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10700 = 10'h8f == _T_174[9:0] ? 4'hb : _GEN_10699; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10701 = 10'h90 == _T_174[9:0] ? 4'hc : _GEN_10700; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10702 = 10'h91 == _T_174[9:0] ? 4'hc : _GEN_10701; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10703 = 10'h92 == _T_174[9:0] ? 4'hd : _GEN_10702; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10704 = 10'h93 == _T_174[9:0] ? 4'he : _GEN_10703; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10705 = 10'h94 == _T_174[9:0] ? 4'he : _GEN_10704; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10706 = 10'h95 == _T_174[9:0] ? 4'he : _GEN_10705; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10707 = 10'h96 == _T_174[9:0] ? 4'he : _GEN_10706; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10708 = 10'h97 == _T_174[9:0] ? 4'he : _GEN_10707; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10709 = 10'h98 == _T_174[9:0] ? 4'he : _GEN_10708; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10710 = 10'h99 == _T_174[9:0] ? 4'he : _GEN_10709; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10711 = 10'h9a == _T_174[9:0] ? 4'he : _GEN_10710; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10712 = 10'h9b == _T_174[9:0] ? 4'he : _GEN_10711; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10713 = 10'h9c == _T_174[9:0] ? 4'he : _GEN_10712; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10714 = 10'h9d == _T_174[9:0] ? 4'he : _GEN_10713; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10715 = 10'h9e == _T_174[9:0] ? 4'he : _GEN_10714; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10716 = 10'h9f == _T_174[9:0] ? 4'he : _GEN_10715; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10717 = 10'ha0 == _T_174[9:0] ? 4'he : _GEN_10716; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10718 = 10'ha1 == _T_174[9:0] ? 4'he : _GEN_10717; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10719 = 10'ha2 == _T_174[9:0] ? 4'he : _GEN_10718; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10720 = 10'ha3 == _T_174[9:0] ? 4'he : _GEN_10719; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10721 = 10'ha4 == _T_174[9:0] ? 4'he : _GEN_10720; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10722 = 10'ha5 == _T_174[9:0] ? 4'he : _GEN_10721; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10723 = 10'ha6 == _T_174[9:0] ? 4'he : _GEN_10722; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10724 = 10'ha7 == _T_174[9:0] ? 4'he : _GEN_10723; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10725 = 10'ha8 == _T_174[9:0] ? 4'hb : _GEN_10724; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10726 = 10'ha9 == _T_174[9:0] ? 4'hc : _GEN_10725; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10727 = 10'haa == _T_174[9:0] ? 4'hb : _GEN_10726; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10728 = 10'hab == _T_174[9:0] ? 4'hc : _GEN_10727; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10729 = 10'hac == _T_174[9:0] ? 4'hd : _GEN_10728; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10730 = 10'had == _T_174[9:0] ? 4'ha : _GEN_10729; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10731 = 10'hae == _T_174[9:0] ? 4'hd : _GEN_10730; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10732 = 10'haf == _T_174[9:0] ? 4'hd : _GEN_10731; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10733 = 10'hb0 == _T_174[9:0] ? 4'hb : _GEN_10732; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10734 = 10'hb1 == _T_174[9:0] ? 4'hc : _GEN_10733; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10735 = 10'hb2 == _T_174[9:0] ? 4'he : _GEN_10734; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10736 = 10'hb3 == _T_174[9:0] ? 4'hb : _GEN_10735; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10737 = 10'hb4 == _T_174[9:0] ? 4'hc : _GEN_10736; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10738 = 10'hb5 == _T_174[9:0] ? 4'hd : _GEN_10737; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10739 = 10'hb6 == _T_174[9:0] ? 4'hd : _GEN_10738; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10740 = 10'hb7 == _T_174[9:0] ? 4'hc : _GEN_10739; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10741 = 10'hb8 == _T_174[9:0] ? 4'he : _GEN_10740; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10742 = 10'hb9 == _T_174[9:0] ? 4'he : _GEN_10741; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10743 = 10'hba == _T_174[9:0] ? 4'he : _GEN_10742; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10744 = 10'hbb == _T_174[9:0] ? 4'he : _GEN_10743; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10745 = 10'hbc == _T_174[9:0] ? 4'he : _GEN_10744; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10746 = 10'hbd == _T_174[9:0] ? 4'he : _GEN_10745; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10747 = 10'hbe == _T_174[9:0] ? 4'he : _GEN_10746; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10748 = 10'hbf == _T_174[9:0] ? 4'he : _GEN_10747; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10749 = 10'hc0 == _T_174[9:0] ? 4'he : _GEN_10748; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10750 = 10'hc1 == _T_174[9:0] ? 4'he : _GEN_10749; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10751 = 10'hc2 == _T_174[9:0] ? 4'he : _GEN_10750; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10752 = 10'hc3 == _T_174[9:0] ? 4'he : _GEN_10751; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10753 = 10'hc4 == _T_174[9:0] ? 4'he : _GEN_10752; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10754 = 10'hc5 == _T_174[9:0] ? 4'he : _GEN_10753; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10755 = 10'hc6 == _T_174[9:0] ? 4'he : _GEN_10754; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10756 = 10'hc7 == _T_174[9:0] ? 4'hd : _GEN_10755; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10757 = 10'hc8 == _T_174[9:0] ? 4'hb : _GEN_10756; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10758 = 10'hc9 == _T_174[9:0] ? 4'hc : _GEN_10757; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10759 = 10'hca == _T_174[9:0] ? 4'he : _GEN_10758; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10760 = 10'hcb == _T_174[9:0] ? 4'he : _GEN_10759; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10761 = 10'hcc == _T_174[9:0] ? 4'he : _GEN_10760; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10762 = 10'hcd == _T_174[9:0] ? 4'he : _GEN_10761; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10763 = 10'hce == _T_174[9:0] ? 4'hd : _GEN_10762; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10764 = 10'hcf == _T_174[9:0] ? 4'hb : _GEN_10763; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10765 = 10'hd0 == _T_174[9:0] ? 4'hc : _GEN_10764; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10766 = 10'hd1 == _T_174[9:0] ? 4'hc : _GEN_10765; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10767 = 10'hd2 == _T_174[9:0] ? 4'hb : _GEN_10766; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10768 = 10'hd3 == _T_174[9:0] ? 4'hd : _GEN_10767; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10769 = 10'hd4 == _T_174[9:0] ? 4'hd : _GEN_10768; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10770 = 10'hd5 == _T_174[9:0] ? 4'hd : _GEN_10769; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10771 = 10'hd6 == _T_174[9:0] ? 4'hd : _GEN_10770; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10772 = 10'hd7 == _T_174[9:0] ? 4'hc : _GEN_10771; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10773 = 10'hd8 == _T_174[9:0] ? 4'hc : _GEN_10772; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10774 = 10'hd9 == _T_174[9:0] ? 4'hc : _GEN_10773; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10775 = 10'hda == _T_174[9:0] ? 4'hd : _GEN_10774; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10776 = 10'hdb == _T_174[9:0] ? 4'hc : _GEN_10775; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10777 = 10'hdc == _T_174[9:0] ? 4'h9 : _GEN_10776; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10778 = 10'hdd == _T_174[9:0] ? 4'he : _GEN_10777; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10779 = 10'hde == _T_174[9:0] ? 4'he : _GEN_10778; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10780 = 10'hdf == _T_174[9:0] ? 4'he : _GEN_10779; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10781 = 10'he0 == _T_174[9:0] ? 4'he : _GEN_10780; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10782 = 10'he1 == _T_174[9:0] ? 4'he : _GEN_10781; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10783 = 10'he2 == _T_174[9:0] ? 4'he : _GEN_10782; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10784 = 10'he3 == _T_174[9:0] ? 4'h9 : _GEN_10783; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10785 = 10'he4 == _T_174[9:0] ? 4'he : _GEN_10784; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10786 = 10'he5 == _T_174[9:0] ? 4'he : _GEN_10785; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10787 = 10'he6 == _T_174[9:0] ? 4'he : _GEN_10786; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10788 = 10'he7 == _T_174[9:0] ? 4'he : _GEN_10787; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10789 = 10'he8 == _T_174[9:0] ? 4'he : _GEN_10788; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10790 = 10'he9 == _T_174[9:0] ? 4'he : _GEN_10789; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10791 = 10'hea == _T_174[9:0] ? 4'he : _GEN_10790; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10792 = 10'heb == _T_174[9:0] ? 4'hc : _GEN_10791; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10793 = 10'hec == _T_174[9:0] ? 4'h7 : _GEN_10792; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10794 = 10'hed == _T_174[9:0] ? 4'h1 : _GEN_10793; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10795 = 10'hee == _T_174[9:0] ? 4'h0 : _GEN_10794; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10796 = 10'hef == _T_174[9:0] ? 4'h0 : _GEN_10795; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10797 = 10'hf0 == _T_174[9:0] ? 4'h2 : _GEN_10796; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10798 = 10'hf1 == _T_174[9:0] ? 4'h9 : _GEN_10797; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10799 = 10'hf2 == _T_174[9:0] ? 4'he : _GEN_10798; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10800 = 10'hf3 == _T_174[9:0] ? 4'he : _GEN_10799; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10801 = 10'hf4 == _T_174[9:0] ? 4'he : _GEN_10800; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10802 = 10'hf5 == _T_174[9:0] ? 4'hc : _GEN_10801; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10803 = 10'hf6 == _T_174[9:0] ? 4'hc : _GEN_10802; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10804 = 10'hf7 == _T_174[9:0] ? 4'hd : _GEN_10803; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10805 = 10'hf8 == _T_174[9:0] ? 4'hd : _GEN_10804; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10806 = 10'hf9 == _T_174[9:0] ? 4'hd : _GEN_10805; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10807 = 10'hfa == _T_174[9:0] ? 4'hd : _GEN_10806; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10808 = 10'hfb == _T_174[9:0] ? 4'hd : _GEN_10807; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10809 = 10'hfc == _T_174[9:0] ? 4'hd : _GEN_10808; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10810 = 10'hfd == _T_174[9:0] ? 4'hd : _GEN_10809; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10811 = 10'hfe == _T_174[9:0] ? 4'hd : _GEN_10810; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10812 = 10'hff == _T_174[9:0] ? 4'hd : _GEN_10811; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10813 = 10'h100 == _T_174[9:0] ? 4'hd : _GEN_10812; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10814 = 10'h101 == _T_174[9:0] ? 4'h9 : _GEN_10813; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10815 = 10'h102 == _T_174[9:0] ? 4'h9 : _GEN_10814; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10816 = 10'h103 == _T_174[9:0] ? 4'he : _GEN_10815; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10817 = 10'h104 == _T_174[9:0] ? 4'he : _GEN_10816; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10818 = 10'h105 == _T_174[9:0] ? 4'he : _GEN_10817; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10819 = 10'h106 == _T_174[9:0] ? 4'he : _GEN_10818; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10820 = 10'h107 == _T_174[9:0] ? 4'he : _GEN_10819; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10821 = 10'h108 == _T_174[9:0] ? 4'he : _GEN_10820; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10822 = 10'h109 == _T_174[9:0] ? 4'h6 : _GEN_10821; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10823 = 10'h10a == _T_174[9:0] ? 4'he : _GEN_10822; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10824 = 10'h10b == _T_174[9:0] ? 4'he : _GEN_10823; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10825 = 10'h10c == _T_174[9:0] ? 4'he : _GEN_10824; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10826 = 10'h10d == _T_174[9:0] ? 4'he : _GEN_10825; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10827 = 10'h10e == _T_174[9:0] ? 4'he : _GEN_10826; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10828 = 10'h10f == _T_174[9:0] ? 4'ha : _GEN_10827; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10829 = 10'h110 == _T_174[9:0] ? 4'hd : _GEN_10828; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10830 = 10'h111 == _T_174[9:0] ? 4'h4 : _GEN_10829; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10831 = 10'h112 == _T_174[9:0] ? 4'h7 : _GEN_10830; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10832 = 10'h113 == _T_174[9:0] ? 4'h0 : _GEN_10831; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10833 = 10'h114 == _T_174[9:0] ? 4'h0 : _GEN_10832; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10834 = 10'h115 == _T_174[9:0] ? 4'h0 : _GEN_10833; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10835 = 10'h116 == _T_174[9:0] ? 4'h0 : _GEN_10834; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10836 = 10'h117 == _T_174[9:0] ? 4'h0 : _GEN_10835; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10837 = 10'h118 == _T_174[9:0] ? 4'ha : _GEN_10836; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10838 = 10'h119 == _T_174[9:0] ? 4'he : _GEN_10837; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10839 = 10'h11a == _T_174[9:0] ? 4'he : _GEN_10838; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10840 = 10'h11b == _T_174[9:0] ? 4'he : _GEN_10839; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10841 = 10'h11c == _T_174[9:0] ? 4'hb : _GEN_10840; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10842 = 10'h11d == _T_174[9:0] ? 4'hc : _GEN_10841; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10843 = 10'h11e == _T_174[9:0] ? 4'hd : _GEN_10842; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10844 = 10'h11f == _T_174[9:0] ? 4'hb : _GEN_10843; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10845 = 10'h120 == _T_174[9:0] ? 4'ha : _GEN_10844; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10846 = 10'h121 == _T_174[9:0] ? 4'hc : _GEN_10845; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10847 = 10'h122 == _T_174[9:0] ? 4'ha : _GEN_10846; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10848 = 10'h123 == _T_174[9:0] ? 4'ha : _GEN_10847; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10849 = 10'h124 == _T_174[9:0] ? 4'hd : _GEN_10848; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10850 = 10'h125 == _T_174[9:0] ? 4'hd : _GEN_10849; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10851 = 10'h126 == _T_174[9:0] ? 4'hb : _GEN_10850; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10852 = 10'h127 == _T_174[9:0] ? 4'h9 : _GEN_10851; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10853 = 10'h128 == _T_174[9:0] ? 4'h7 : _GEN_10852; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10854 = 10'h129 == _T_174[9:0] ? 4'hd : _GEN_10853; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10855 = 10'h12a == _T_174[9:0] ? 4'hc : _GEN_10854; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10856 = 10'h12b == _T_174[9:0] ? 4'hb : _GEN_10855; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10857 = 10'h12c == _T_174[9:0] ? 4'hc : _GEN_10856; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10858 = 10'h12d == _T_174[9:0] ? 4'hb : _GEN_10857; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10859 = 10'h12e == _T_174[9:0] ? 4'ha : _GEN_10858; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10860 = 10'h12f == _T_174[9:0] ? 4'h6 : _GEN_10859; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10861 = 10'h130 == _T_174[9:0] ? 4'he : _GEN_10860; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10862 = 10'h131 == _T_174[9:0] ? 4'hc : _GEN_10861; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10863 = 10'h132 == _T_174[9:0] ? 4'ha : _GEN_10862; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10864 = 10'h133 == _T_174[9:0] ? 4'h9 : _GEN_10863; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10865 = 10'h134 == _T_174[9:0] ? 4'hb : _GEN_10864; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10866 = 10'h135 == _T_174[9:0] ? 4'h8 : _GEN_10865; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10867 = 10'h136 == _T_174[9:0] ? 4'h8 : _GEN_10866; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10868 = 10'h137 == _T_174[9:0] ? 4'h4 : _GEN_10867; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10869 = 10'h138 == _T_174[9:0] ? 4'h7 : _GEN_10868; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10870 = 10'h139 == _T_174[9:0] ? 4'h0 : _GEN_10869; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10871 = 10'h13a == _T_174[9:0] ? 4'h0 : _GEN_10870; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10872 = 10'h13b == _T_174[9:0] ? 4'h0 : _GEN_10871; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10873 = 10'h13c == _T_174[9:0] ? 4'h0 : _GEN_10872; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10874 = 10'h13d == _T_174[9:0] ? 4'h0 : _GEN_10873; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10875 = 10'h13e == _T_174[9:0] ? 4'h4 : _GEN_10874; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10876 = 10'h13f == _T_174[9:0] ? 4'hc : _GEN_10875; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10877 = 10'h140 == _T_174[9:0] ? 4'he : _GEN_10876; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10878 = 10'h141 == _T_174[9:0] ? 4'he : _GEN_10877; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10879 = 10'h142 == _T_174[9:0] ? 4'he : _GEN_10878; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10880 = 10'h143 == _T_174[9:0] ? 4'hc : _GEN_10879; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10881 = 10'h144 == _T_174[9:0] ? 4'hd : _GEN_10880; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10882 = 10'h145 == _T_174[9:0] ? 4'hb : _GEN_10881; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10883 = 10'h146 == _T_174[9:0] ? 4'hb : _GEN_10882; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10884 = 10'h147 == _T_174[9:0] ? 4'ha : _GEN_10883; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10885 = 10'h148 == _T_174[9:0] ? 4'ha : _GEN_10884; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10886 = 10'h149 == _T_174[9:0] ? 4'hc : _GEN_10885; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10887 = 10'h14a == _T_174[9:0] ? 4'hd : _GEN_10886; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10888 = 10'h14b == _T_174[9:0] ? 4'hc : _GEN_10887; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10889 = 10'h14c == _T_174[9:0] ? 4'hd : _GEN_10888; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10890 = 10'h14d == _T_174[9:0] ? 4'h9 : _GEN_10889; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10891 = 10'h14e == _T_174[9:0] ? 4'h7 : _GEN_10890; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10892 = 10'h14f == _T_174[9:0] ? 4'ha : _GEN_10891; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10893 = 10'h150 == _T_174[9:0] ? 4'ha : _GEN_10892; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10894 = 10'h151 == _T_174[9:0] ? 4'hb : _GEN_10893; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10895 = 10'h152 == _T_174[9:0] ? 4'hb : _GEN_10894; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10896 = 10'h153 == _T_174[9:0] ? 4'hc : _GEN_10895; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10897 = 10'h154 == _T_174[9:0] ? 4'hb : _GEN_10896; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10898 = 10'h155 == _T_174[9:0] ? 4'h6 : _GEN_10897; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10899 = 10'h156 == _T_174[9:0] ? 4'hb : _GEN_10898; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10900 = 10'h157 == _T_174[9:0] ? 4'h7 : _GEN_10899; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10901 = 10'h158 == _T_174[9:0] ? 4'h7 : _GEN_10900; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10902 = 10'h159 == _T_174[9:0] ? 4'h7 : _GEN_10901; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10903 = 10'h15a == _T_174[9:0] ? 4'h7 : _GEN_10902; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10904 = 10'h15b == _T_174[9:0] ? 4'h7 : _GEN_10903; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10905 = 10'h15c == _T_174[9:0] ? 4'h7 : _GEN_10904; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10906 = 10'h15d == _T_174[9:0] ? 4'h6 : _GEN_10905; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10907 = 10'h15e == _T_174[9:0] ? 4'h7 : _GEN_10906; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10908 = 10'h15f == _T_174[9:0] ? 4'h0 : _GEN_10907; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10909 = 10'h160 == _T_174[9:0] ? 4'h0 : _GEN_10908; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10910 = 10'h161 == _T_174[9:0] ? 4'h0 : _GEN_10909; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10911 = 10'h162 == _T_174[9:0] ? 4'h0 : _GEN_10910; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10912 = 10'h163 == _T_174[9:0] ? 4'h2 : _GEN_10911; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10913 = 10'h164 == _T_174[9:0] ? 4'h4 : _GEN_10912; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10914 = 10'h165 == _T_174[9:0] ? 4'hb : _GEN_10913; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10915 = 10'h166 == _T_174[9:0] ? 4'hb : _GEN_10914; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10916 = 10'h167 == _T_174[9:0] ? 4'he : _GEN_10915; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10917 = 10'h168 == _T_174[9:0] ? 4'he : _GEN_10916; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10918 = 10'h169 == _T_174[9:0] ? 4'hc : _GEN_10917; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10919 = 10'h16a == _T_174[9:0] ? 4'hd : _GEN_10918; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10920 = 10'h16b == _T_174[9:0] ? 4'hd : _GEN_10919; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10921 = 10'h16c == _T_174[9:0] ? 4'ha : _GEN_10920; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10922 = 10'h16d == _T_174[9:0] ? 4'ha : _GEN_10921; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10923 = 10'h16e == _T_174[9:0] ? 4'ha : _GEN_10922; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10924 = 10'h16f == _T_174[9:0] ? 4'hd : _GEN_10923; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10925 = 10'h170 == _T_174[9:0] ? 4'hd : _GEN_10924; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10926 = 10'h171 == _T_174[9:0] ? 4'hd : _GEN_10925; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10927 = 10'h172 == _T_174[9:0] ? 4'he : _GEN_10926; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10928 = 10'h173 == _T_174[9:0] ? 4'h8 : _GEN_10927; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10929 = 10'h174 == _T_174[9:0] ? 4'h5 : _GEN_10928; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10930 = 10'h175 == _T_174[9:0] ? 4'h6 : _GEN_10929; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10931 = 10'h176 == _T_174[9:0] ? 4'h6 : _GEN_10930; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10932 = 10'h177 == _T_174[9:0] ? 4'h6 : _GEN_10931; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10933 = 10'h178 == _T_174[9:0] ? 4'h7 : _GEN_10932; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10934 = 10'h179 == _T_174[9:0] ? 4'h9 : _GEN_10933; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10935 = 10'h17a == _T_174[9:0] ? 4'h9 : _GEN_10934; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10936 = 10'h17b == _T_174[9:0] ? 4'h6 : _GEN_10935; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10937 = 10'h17c == _T_174[9:0] ? 4'h7 : _GEN_10936; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10938 = 10'h17d == _T_174[9:0] ? 4'h7 : _GEN_10937; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10939 = 10'h17e == _T_174[9:0] ? 4'h7 : _GEN_10938; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10940 = 10'h17f == _T_174[9:0] ? 4'h7 : _GEN_10939; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10941 = 10'h180 == _T_174[9:0] ? 4'h7 : _GEN_10940; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10942 = 10'h181 == _T_174[9:0] ? 4'h7 : _GEN_10941; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10943 = 10'h182 == _T_174[9:0] ? 4'h8 : _GEN_10942; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10944 = 10'h183 == _T_174[9:0] ? 4'h8 : _GEN_10943; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10945 = 10'h184 == _T_174[9:0] ? 4'h8 : _GEN_10944; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10946 = 10'h185 == _T_174[9:0] ? 4'h7 : _GEN_10945; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10947 = 10'h186 == _T_174[9:0] ? 4'h1 : _GEN_10946; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10948 = 10'h187 == _T_174[9:0] ? 4'h0 : _GEN_10947; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10949 = 10'h188 == _T_174[9:0] ? 4'h0 : _GEN_10948; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10950 = 10'h189 == _T_174[9:0] ? 4'h4 : _GEN_10949; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10951 = 10'h18a == _T_174[9:0] ? 4'h4 : _GEN_10950; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10952 = 10'h18b == _T_174[9:0] ? 4'hb : _GEN_10951; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10953 = 10'h18c == _T_174[9:0] ? 4'hb : _GEN_10952; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10954 = 10'h18d == _T_174[9:0] ? 4'hc : _GEN_10953; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10955 = 10'h18e == _T_174[9:0] ? 4'he : _GEN_10954; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10956 = 10'h18f == _T_174[9:0] ? 4'hb : _GEN_10955; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10957 = 10'h190 == _T_174[9:0] ? 4'hd : _GEN_10956; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10958 = 10'h191 == _T_174[9:0] ? 4'hc : _GEN_10957; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10959 = 10'h192 == _T_174[9:0] ? 4'h9 : _GEN_10958; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10960 = 10'h193 == _T_174[9:0] ? 4'ha : _GEN_10959; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10961 = 10'h194 == _T_174[9:0] ? 4'h9 : _GEN_10960; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10962 = 10'h195 == _T_174[9:0] ? 4'hd : _GEN_10961; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10963 = 10'h196 == _T_174[9:0] ? 4'hd : _GEN_10962; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10964 = 10'h197 == _T_174[9:0] ? 4'hb : _GEN_10963; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10965 = 10'h198 == _T_174[9:0] ? 4'he : _GEN_10964; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10966 = 10'h199 == _T_174[9:0] ? 4'h5 : _GEN_10965; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10967 = 10'h19a == _T_174[9:0] ? 4'h1 : _GEN_10966; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10968 = 10'h19b == _T_174[9:0] ? 4'h3 : _GEN_10967; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10969 = 10'h19c == _T_174[9:0] ? 4'h6 : _GEN_10968; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10970 = 10'h19d == _T_174[9:0] ? 4'h4 : _GEN_10969; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10971 = 10'h19e == _T_174[9:0] ? 4'h1 : _GEN_10970; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10972 = 10'h19f == _T_174[9:0] ? 4'h3 : _GEN_10971; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10973 = 10'h1a0 == _T_174[9:0] ? 4'h6 : _GEN_10972; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10974 = 10'h1a1 == _T_174[9:0] ? 4'h6 : _GEN_10973; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10975 = 10'h1a2 == _T_174[9:0] ? 4'h7 : _GEN_10974; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10976 = 10'h1a3 == _T_174[9:0] ? 4'h7 : _GEN_10975; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10977 = 10'h1a4 == _T_174[9:0] ? 4'h7 : _GEN_10976; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10978 = 10'h1a5 == _T_174[9:0] ? 4'h7 : _GEN_10977; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10979 = 10'h1a6 == _T_174[9:0] ? 4'h7 : _GEN_10978; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10980 = 10'h1a7 == _T_174[9:0] ? 4'h7 : _GEN_10979; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10981 = 10'h1a8 == _T_174[9:0] ? 4'h8 : _GEN_10980; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10982 = 10'h1a9 == _T_174[9:0] ? 4'h8 : _GEN_10981; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10983 = 10'h1aa == _T_174[9:0] ? 4'h7 : _GEN_10982; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10984 = 10'h1ab == _T_174[9:0] ? 4'h8 : _GEN_10983; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10985 = 10'h1ac == _T_174[9:0] ? 4'h8 : _GEN_10984; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10986 = 10'h1ad == _T_174[9:0] ? 4'h3 : _GEN_10985; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10987 = 10'h1ae == _T_174[9:0] ? 4'h2 : _GEN_10986; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10988 = 10'h1af == _T_174[9:0] ? 4'h8 : _GEN_10987; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10989 = 10'h1b0 == _T_174[9:0] ? 4'h6 : _GEN_10988; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10990 = 10'h1b1 == _T_174[9:0] ? 4'hb : _GEN_10989; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10991 = 10'h1b2 == _T_174[9:0] ? 4'hb : _GEN_10990; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10992 = 10'h1b3 == _T_174[9:0] ? 4'ha : _GEN_10991; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10993 = 10'h1b4 == _T_174[9:0] ? 4'he : _GEN_10992; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10994 = 10'h1b5 == _T_174[9:0] ? 4'hb : _GEN_10993; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10995 = 10'h1b6 == _T_174[9:0] ? 4'hc : _GEN_10994; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10996 = 10'h1b7 == _T_174[9:0] ? 4'ha : _GEN_10995; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10997 = 10'h1b8 == _T_174[9:0] ? 4'h9 : _GEN_10996; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10998 = 10'h1b9 == _T_174[9:0] ? 4'h9 : _GEN_10997; // @[Filter.scala 230:102]
  wire [3:0] _GEN_10999 = 10'h1ba == _T_174[9:0] ? 4'h9 : _GEN_10998; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11000 = 10'h1bb == _T_174[9:0] ? 4'hb : _GEN_10999; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11001 = 10'h1bc == _T_174[9:0] ? 4'hd : _GEN_11000; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11002 = 10'h1bd == _T_174[9:0] ? 4'hd : _GEN_11001; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11003 = 10'h1be == _T_174[9:0] ? 4'he : _GEN_11002; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11004 = 10'h1bf == _T_174[9:0] ? 4'h7 : _GEN_11003; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11005 = 10'h1c0 == _T_174[9:0] ? 4'h6 : _GEN_11004; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11006 = 10'h1c1 == _T_174[9:0] ? 4'h6 : _GEN_11005; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11007 = 10'h1c2 == _T_174[9:0] ? 4'h5 : _GEN_11006; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11008 = 10'h1c3 == _T_174[9:0] ? 4'h5 : _GEN_11007; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11009 = 10'h1c4 == _T_174[9:0] ? 4'h4 : _GEN_11008; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11010 = 10'h1c5 == _T_174[9:0] ? 4'h5 : _GEN_11009; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11011 = 10'h1c6 == _T_174[9:0] ? 4'h6 : _GEN_11010; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11012 = 10'h1c7 == _T_174[9:0] ? 4'h6 : _GEN_11011; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11013 = 10'h1c8 == _T_174[9:0] ? 4'h7 : _GEN_11012; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11014 = 10'h1c9 == _T_174[9:0] ? 4'h7 : _GEN_11013; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11015 = 10'h1ca == _T_174[9:0] ? 4'h7 : _GEN_11014; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11016 = 10'h1cb == _T_174[9:0] ? 4'h7 : _GEN_11015; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11017 = 10'h1cc == _T_174[9:0] ? 4'h7 : _GEN_11016; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11018 = 10'h1cd == _T_174[9:0] ? 4'h8 : _GEN_11017; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11019 = 10'h1ce == _T_174[9:0] ? 4'h8 : _GEN_11018; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11020 = 10'h1cf == _T_174[9:0] ? 4'h8 : _GEN_11019; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11021 = 10'h1d0 == _T_174[9:0] ? 4'h5 : _GEN_11020; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11022 = 10'h1d1 == _T_174[9:0] ? 4'h8 : _GEN_11021; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11023 = 10'h1d2 == _T_174[9:0] ? 4'h8 : _GEN_11022; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11024 = 10'h1d3 == _T_174[9:0] ? 4'h8 : _GEN_11023; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11025 = 10'h1d4 == _T_174[9:0] ? 4'h8 : _GEN_11024; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11026 = 10'h1d5 == _T_174[9:0] ? 4'h7 : _GEN_11025; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11027 = 10'h1d6 == _T_174[9:0] ? 4'h9 : _GEN_11026; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11028 = 10'h1d7 == _T_174[9:0] ? 4'hb : _GEN_11027; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11029 = 10'h1d8 == _T_174[9:0] ? 4'hb : _GEN_11028; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11030 = 10'h1d9 == _T_174[9:0] ? 4'hb : _GEN_11029; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11031 = 10'h1da == _T_174[9:0] ? 4'ha : _GEN_11030; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11032 = 10'h1db == _T_174[9:0] ? 4'hc : _GEN_11031; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11033 = 10'h1dc == _T_174[9:0] ? 4'hb : _GEN_11032; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11034 = 10'h1dd == _T_174[9:0] ? 4'h5 : _GEN_11033; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11035 = 10'h1de == _T_174[9:0] ? 4'h9 : _GEN_11034; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11036 = 10'h1df == _T_174[9:0] ? 4'h9 : _GEN_11035; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11037 = 10'h1e0 == _T_174[9:0] ? 4'h9 : _GEN_11036; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11038 = 10'h1e1 == _T_174[9:0] ? 4'h7 : _GEN_11037; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11039 = 10'h1e2 == _T_174[9:0] ? 4'hc : _GEN_11038; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11040 = 10'h1e3 == _T_174[9:0] ? 4'hc : _GEN_11039; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11041 = 10'h1e4 == _T_174[9:0] ? 4'hd : _GEN_11040; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11042 = 10'h1e5 == _T_174[9:0] ? 4'h7 : _GEN_11041; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11043 = 10'h1e6 == _T_174[9:0] ? 4'h6 : _GEN_11042; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11044 = 10'h1e7 == _T_174[9:0] ? 4'h6 : _GEN_11043; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11045 = 10'h1e8 == _T_174[9:0] ? 4'h6 : _GEN_11044; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11046 = 10'h1e9 == _T_174[9:0] ? 4'h6 : _GEN_11045; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11047 = 10'h1ea == _T_174[9:0] ? 4'h6 : _GEN_11046; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11048 = 10'h1eb == _T_174[9:0] ? 4'h6 : _GEN_11047; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11049 = 10'h1ec == _T_174[9:0] ? 4'h6 : _GEN_11048; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11050 = 10'h1ed == _T_174[9:0] ? 4'h8 : _GEN_11049; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11051 = 10'h1ee == _T_174[9:0] ? 4'h7 : _GEN_11050; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11052 = 10'h1ef == _T_174[9:0] ? 4'h7 : _GEN_11051; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11053 = 10'h1f0 == _T_174[9:0] ? 4'h7 : _GEN_11052; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11054 = 10'h1f1 == _T_174[9:0] ? 4'h7 : _GEN_11053; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11055 = 10'h1f2 == _T_174[9:0] ? 4'h7 : _GEN_11054; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11056 = 10'h1f3 == _T_174[9:0] ? 4'h8 : _GEN_11055; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11057 = 10'h1f4 == _T_174[9:0] ? 4'h8 : _GEN_11056; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11058 = 10'h1f5 == _T_174[9:0] ? 4'h8 : _GEN_11057; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11059 = 10'h1f6 == _T_174[9:0] ? 4'ha : _GEN_11058; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11060 = 10'h1f7 == _T_174[9:0] ? 4'h8 : _GEN_11059; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11061 = 10'h1f8 == _T_174[9:0] ? 4'h8 : _GEN_11060; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11062 = 10'h1f9 == _T_174[9:0] ? 4'h9 : _GEN_11061; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11063 = 10'h1fa == _T_174[9:0] ? 4'h9 : _GEN_11062; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11064 = 10'h1fb == _T_174[9:0] ? 4'h8 : _GEN_11063; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11065 = 10'h1fc == _T_174[9:0] ? 4'hb : _GEN_11064; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11066 = 10'h1fd == _T_174[9:0] ? 4'hb : _GEN_11065; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11067 = 10'h1fe == _T_174[9:0] ? 4'hb : _GEN_11066; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11068 = 10'h1ff == _T_174[9:0] ? 4'ha : _GEN_11067; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11069 = 10'h200 == _T_174[9:0] ? 4'h3 : _GEN_11068; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11070 = 10'h201 == _T_174[9:0] ? 4'h9 : _GEN_11069; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11071 = 10'h202 == _T_174[9:0] ? 4'h5 : _GEN_11070; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11072 = 10'h203 == _T_174[9:0] ? 4'h3 : _GEN_11071; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11073 = 10'h204 == _T_174[9:0] ? 4'h4 : _GEN_11072; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11074 = 10'h205 == _T_174[9:0] ? 4'h4 : _GEN_11073; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11075 = 10'h206 == _T_174[9:0] ? 4'h4 : _GEN_11074; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11076 = 10'h207 == _T_174[9:0] ? 4'h4 : _GEN_11075; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11077 = 10'h208 == _T_174[9:0] ? 4'h8 : _GEN_11076; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11078 = 10'h209 == _T_174[9:0] ? 4'hc : _GEN_11077; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11079 = 10'h20a == _T_174[9:0] ? 4'hd : _GEN_11078; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11080 = 10'h20b == _T_174[9:0] ? 4'h7 : _GEN_11079; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11081 = 10'h20c == _T_174[9:0] ? 4'h6 : _GEN_11080; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11082 = 10'h20d == _T_174[9:0] ? 4'h6 : _GEN_11081; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11083 = 10'h20e == _T_174[9:0] ? 4'h6 : _GEN_11082; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11084 = 10'h20f == _T_174[9:0] ? 4'h5 : _GEN_11083; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11085 = 10'h210 == _T_174[9:0] ? 4'h6 : _GEN_11084; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11086 = 10'h211 == _T_174[9:0] ? 4'h6 : _GEN_11085; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11087 = 10'h212 == _T_174[9:0] ? 4'h7 : _GEN_11086; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11088 = 10'h213 == _T_174[9:0] ? 4'ha : _GEN_11087; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11089 = 10'h214 == _T_174[9:0] ? 4'h6 : _GEN_11088; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11090 = 10'h215 == _T_174[9:0] ? 4'h7 : _GEN_11089; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11091 = 10'h216 == _T_174[9:0] ? 4'h7 : _GEN_11090; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11092 = 10'h217 == _T_174[9:0] ? 4'h7 : _GEN_11091; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11093 = 10'h218 == _T_174[9:0] ? 4'h7 : _GEN_11092; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11094 = 10'h219 == _T_174[9:0] ? 4'h8 : _GEN_11093; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11095 = 10'h21a == _T_174[9:0] ? 4'h7 : _GEN_11094; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11096 = 10'h21b == _T_174[9:0] ? 4'h8 : _GEN_11095; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11097 = 10'h21c == _T_174[9:0] ? 4'hb : _GEN_11096; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11098 = 10'h21d == _T_174[9:0] ? 4'ha : _GEN_11097; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11099 = 10'h21e == _T_174[9:0] ? 4'h9 : _GEN_11098; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11100 = 10'h21f == _T_174[9:0] ? 4'h9 : _GEN_11099; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11101 = 10'h220 == _T_174[9:0] ? 4'h8 : _GEN_11100; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11102 = 10'h221 == _T_174[9:0] ? 4'h9 : _GEN_11101; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11103 = 10'h222 == _T_174[9:0] ? 4'hb : _GEN_11102; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11104 = 10'h223 == _T_174[9:0] ? 4'hb : _GEN_11103; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11105 = 10'h224 == _T_174[9:0] ? 4'hb : _GEN_11104; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11106 = 10'h225 == _T_174[9:0] ? 4'h8 : _GEN_11105; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11107 = 10'h226 == _T_174[9:0] ? 4'h1 : _GEN_11106; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11108 = 10'h227 == _T_174[9:0] ? 4'h3 : _GEN_11107; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11109 = 10'h228 == _T_174[9:0] ? 4'h3 : _GEN_11108; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11110 = 10'h229 == _T_174[9:0] ? 4'h3 : _GEN_11109; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11111 = 10'h22a == _T_174[9:0] ? 4'h3 : _GEN_11110; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11112 = 10'h22b == _T_174[9:0] ? 4'h3 : _GEN_11111; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11113 = 10'h22c == _T_174[9:0] ? 4'h3 : _GEN_11112; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11114 = 10'h22d == _T_174[9:0] ? 4'h3 : _GEN_11113; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11115 = 10'h22e == _T_174[9:0] ? 4'h3 : _GEN_11114; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11116 = 10'h22f == _T_174[9:0] ? 4'h9 : _GEN_11115; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11117 = 10'h230 == _T_174[9:0] ? 4'h6 : _GEN_11116; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11118 = 10'h231 == _T_174[9:0] ? 4'h7 : _GEN_11117; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11119 = 10'h232 == _T_174[9:0] ? 4'h6 : _GEN_11118; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11120 = 10'h233 == _T_174[9:0] ? 4'h7 : _GEN_11119; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11121 = 10'h234 == _T_174[9:0] ? 4'h7 : _GEN_11120; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11122 = 10'h235 == _T_174[9:0] ? 4'h6 : _GEN_11121; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11123 = 10'h236 == _T_174[9:0] ? 4'h6 : _GEN_11122; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11124 = 10'h237 == _T_174[9:0] ? 4'h6 : _GEN_11123; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11125 = 10'h238 == _T_174[9:0] ? 4'h6 : _GEN_11124; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11126 = 10'h239 == _T_174[9:0] ? 4'h8 : _GEN_11125; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11127 = 10'h23a == _T_174[9:0] ? 4'h6 : _GEN_11126; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11128 = 10'h23b == _T_174[9:0] ? 4'h7 : _GEN_11127; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11129 = 10'h23c == _T_174[9:0] ? 4'h7 : _GEN_11128; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11130 = 10'h23d == _T_174[9:0] ? 4'h7 : _GEN_11129; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11131 = 10'h23e == _T_174[9:0] ? 4'h7 : _GEN_11130; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11132 = 10'h23f == _T_174[9:0] ? 4'h7 : _GEN_11131; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11133 = 10'h240 == _T_174[9:0] ? 4'h7 : _GEN_11132; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11134 = 10'h241 == _T_174[9:0] ? 4'h8 : _GEN_11133; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11135 = 10'h242 == _T_174[9:0] ? 4'hb : _GEN_11134; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11136 = 10'h243 == _T_174[9:0] ? 4'hb : _GEN_11135; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11137 = 10'h244 == _T_174[9:0] ? 4'hb : _GEN_11136; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11138 = 10'h245 == _T_174[9:0] ? 4'ha : _GEN_11137; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11139 = 10'h246 == _T_174[9:0] ? 4'h9 : _GEN_11138; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11140 = 10'h247 == _T_174[9:0] ? 4'ha : _GEN_11139; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11141 = 10'h248 == _T_174[9:0] ? 4'hb : _GEN_11140; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11142 = 10'h249 == _T_174[9:0] ? 4'hb : _GEN_11141; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11143 = 10'h24a == _T_174[9:0] ? 4'ha : _GEN_11142; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11144 = 10'h24b == _T_174[9:0] ? 4'h2 : _GEN_11143; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11145 = 10'h24c == _T_174[9:0] ? 4'h0 : _GEN_11144; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11146 = 10'h24d == _T_174[9:0] ? 4'h2 : _GEN_11145; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11147 = 10'h24e == _T_174[9:0] ? 4'h3 : _GEN_11146; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11148 = 10'h24f == _T_174[9:0] ? 4'h3 : _GEN_11147; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11149 = 10'h250 == _T_174[9:0] ? 4'h3 : _GEN_11148; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11150 = 10'h251 == _T_174[9:0] ? 4'h3 : _GEN_11149; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11151 = 10'h252 == _T_174[9:0] ? 4'h3 : _GEN_11150; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11152 = 10'h253 == _T_174[9:0] ? 4'h3 : _GEN_11151; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11153 = 10'h254 == _T_174[9:0] ? 4'h3 : _GEN_11152; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11154 = 10'h255 == _T_174[9:0] ? 4'h5 : _GEN_11153; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11155 = 10'h256 == _T_174[9:0] ? 4'h6 : _GEN_11154; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11156 = 10'h257 == _T_174[9:0] ? 4'h8 : _GEN_11155; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11157 = 10'h258 == _T_174[9:0] ? 4'h5 : _GEN_11156; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11158 = 10'h259 == _T_174[9:0] ? 4'h6 : _GEN_11157; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11159 = 10'h25a == _T_174[9:0] ? 4'h6 : _GEN_11158; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11160 = 10'h25b == _T_174[9:0] ? 4'h5 : _GEN_11159; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11161 = 10'h25c == _T_174[9:0] ? 4'h6 : _GEN_11160; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11162 = 10'h25d == _T_174[9:0] ? 4'h6 : _GEN_11161; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11163 = 10'h25e == _T_174[9:0] ? 4'h9 : _GEN_11162; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11164 = 10'h25f == _T_174[9:0] ? 4'hc : _GEN_11163; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11165 = 10'h260 == _T_174[9:0] ? 4'h7 : _GEN_11164; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11166 = 10'h261 == _T_174[9:0] ? 4'h9 : _GEN_11165; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11167 = 10'h262 == _T_174[9:0] ? 4'ha : _GEN_11166; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11168 = 10'h263 == _T_174[9:0] ? 4'h8 : _GEN_11167; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11169 = 10'h264 == _T_174[9:0] ? 4'ha : _GEN_11168; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11170 = 10'h265 == _T_174[9:0] ? 4'h9 : _GEN_11169; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11171 = 10'h266 == _T_174[9:0] ? 4'h8 : _GEN_11170; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11172 = 10'h267 == _T_174[9:0] ? 4'h8 : _GEN_11171; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11173 = 10'h268 == _T_174[9:0] ? 4'ha : _GEN_11172; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11174 = 10'h269 == _T_174[9:0] ? 4'ha : _GEN_11173; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11175 = 10'h26a == _T_174[9:0] ? 4'hb : _GEN_11174; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11176 = 10'h26b == _T_174[9:0] ? 4'hb : _GEN_11175; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11177 = 10'h26c == _T_174[9:0] ? 4'hb : _GEN_11176; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11178 = 10'h26d == _T_174[9:0] ? 4'hb : _GEN_11177; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11179 = 10'h26e == _T_174[9:0] ? 4'hb : _GEN_11178; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11180 = 10'h26f == _T_174[9:0] ? 4'ha : _GEN_11179; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11181 = 10'h270 == _T_174[9:0] ? 4'h3 : _GEN_11180; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11182 = 10'h271 == _T_174[9:0] ? 4'h0 : _GEN_11181; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11183 = 10'h272 == _T_174[9:0] ? 4'h0 : _GEN_11182; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11184 = 10'h273 == _T_174[9:0] ? 4'h2 : _GEN_11183; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11185 = 10'h274 == _T_174[9:0] ? 4'h3 : _GEN_11184; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11186 = 10'h275 == _T_174[9:0] ? 4'h3 : _GEN_11185; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11187 = 10'h276 == _T_174[9:0] ? 4'h3 : _GEN_11186; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11188 = 10'h277 == _T_174[9:0] ? 4'h3 : _GEN_11187; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11189 = 10'h278 == _T_174[9:0] ? 4'h3 : _GEN_11188; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11190 = 10'h279 == _T_174[9:0] ? 4'h3 : _GEN_11189; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11191 = 10'h27a == _T_174[9:0] ? 4'h3 : _GEN_11190; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11192 = 10'h27b == _T_174[9:0] ? 4'h6 : _GEN_11191; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11193 = 10'h27c == _T_174[9:0] ? 4'h7 : _GEN_11192; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11194 = 10'h27d == _T_174[9:0] ? 4'h7 : _GEN_11193; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11195 = 10'h27e == _T_174[9:0] ? 4'h4 : _GEN_11194; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11196 = 10'h27f == _T_174[9:0] ? 4'h6 : _GEN_11195; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11197 = 10'h280 == _T_174[9:0] ? 4'h6 : _GEN_11196; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11198 = 10'h281 == _T_174[9:0] ? 4'h6 : _GEN_11197; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11199 = 10'h282 == _T_174[9:0] ? 4'h6 : _GEN_11198; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11200 = 10'h283 == _T_174[9:0] ? 4'ha : _GEN_11199; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11201 = 10'h284 == _T_174[9:0] ? 4'hc : _GEN_11200; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11202 = 10'h285 == _T_174[9:0] ? 4'hc : _GEN_11201; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11203 = 10'h286 == _T_174[9:0] ? 4'h8 : _GEN_11202; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11204 = 10'h287 == _T_174[9:0] ? 4'ha : _GEN_11203; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11205 = 10'h288 == _T_174[9:0] ? 4'ha : _GEN_11204; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11206 = 10'h289 == _T_174[9:0] ? 4'ha : _GEN_11205; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11207 = 10'h28a == _T_174[9:0] ? 4'hc : _GEN_11206; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11208 = 10'h28b == _T_174[9:0] ? 4'hb : _GEN_11207; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11209 = 10'h28c == _T_174[9:0] ? 4'ha : _GEN_11208; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11210 = 10'h28d == _T_174[9:0] ? 4'h7 : _GEN_11209; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11211 = 10'h28e == _T_174[9:0] ? 4'h2 : _GEN_11210; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11212 = 10'h28f == _T_174[9:0] ? 4'h5 : _GEN_11211; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11213 = 10'h290 == _T_174[9:0] ? 4'h8 : _GEN_11212; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11214 = 10'h291 == _T_174[9:0] ? 4'ha : _GEN_11213; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11215 = 10'h292 == _T_174[9:0] ? 4'ha : _GEN_11214; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11216 = 10'h293 == _T_174[9:0] ? 4'ha : _GEN_11215; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11217 = 10'h294 == _T_174[9:0] ? 4'h9 : _GEN_11216; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11218 = 10'h295 == _T_174[9:0] ? 4'h3 : _GEN_11217; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11219 = 10'h296 == _T_174[9:0] ? 4'h0 : _GEN_11218; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11220 = 10'h297 == _T_174[9:0] ? 4'h0 : _GEN_11219; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11221 = 10'h298 == _T_174[9:0] ? 4'h0 : _GEN_11220; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11222 = 10'h299 == _T_174[9:0] ? 4'h1 : _GEN_11221; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11223 = 10'h29a == _T_174[9:0] ? 4'h3 : _GEN_11222; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11224 = 10'h29b == _T_174[9:0] ? 4'h3 : _GEN_11223; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11225 = 10'h29c == _T_174[9:0] ? 4'h3 : _GEN_11224; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11226 = 10'h29d == _T_174[9:0] ? 4'h3 : _GEN_11225; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11227 = 10'h29e == _T_174[9:0] ? 4'h3 : _GEN_11226; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11228 = 10'h29f == _T_174[9:0] ? 4'h3 : _GEN_11227; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11229 = 10'h2a0 == _T_174[9:0] ? 4'h4 : _GEN_11228; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11230 = 10'h2a1 == _T_174[9:0] ? 4'h6 : _GEN_11229; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11231 = 10'h2a2 == _T_174[9:0] ? 4'h7 : _GEN_11230; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11232 = 10'h2a3 == _T_174[9:0] ? 4'h6 : _GEN_11231; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11233 = 10'h2a4 == _T_174[9:0] ? 4'h4 : _GEN_11232; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11234 = 10'h2a5 == _T_174[9:0] ? 4'h6 : _GEN_11233; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11235 = 10'h2a6 == _T_174[9:0] ? 4'h6 : _GEN_11234; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11236 = 10'h2a7 == _T_174[9:0] ? 4'h7 : _GEN_11235; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11237 = 10'h2a8 == _T_174[9:0] ? 4'ha : _GEN_11236; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11238 = 10'h2a9 == _T_174[9:0] ? 4'hb : _GEN_11237; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11239 = 10'h2aa == _T_174[9:0] ? 4'hb : _GEN_11238; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11240 = 10'h2ab == _T_174[9:0] ? 4'hb : _GEN_11239; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11241 = 10'h2ac == _T_174[9:0] ? 4'h8 : _GEN_11240; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11242 = 10'h2ad == _T_174[9:0] ? 4'hb : _GEN_11241; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11243 = 10'h2ae == _T_174[9:0] ? 4'ha : _GEN_11242; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11244 = 10'h2af == _T_174[9:0] ? 4'hb : _GEN_11243; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11245 = 10'h2b0 == _T_174[9:0] ? 4'hc : _GEN_11244; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11246 = 10'h2b1 == _T_174[9:0] ? 4'hb : _GEN_11245; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11247 = 10'h2b2 == _T_174[9:0] ? 4'ha : _GEN_11246; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11248 = 10'h2b3 == _T_174[9:0] ? 4'h6 : _GEN_11247; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11249 = 10'h2b4 == _T_174[9:0] ? 4'h0 : _GEN_11248; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11250 = 10'h2b5 == _T_174[9:0] ? 4'h0 : _GEN_11249; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11251 = 10'h2b6 == _T_174[9:0] ? 4'h0 : _GEN_11250; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11252 = 10'h2b7 == _T_174[9:0] ? 4'h1 : _GEN_11251; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11253 = 10'h2b8 == _T_174[9:0] ? 4'h5 : _GEN_11252; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11254 = 10'h2b9 == _T_174[9:0] ? 4'h9 : _GEN_11253; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11255 = 10'h2ba == _T_174[9:0] ? 4'h1 : _GEN_11254; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11256 = 10'h2bb == _T_174[9:0] ? 4'h0 : _GEN_11255; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11257 = 10'h2bc == _T_174[9:0] ? 4'h0 : _GEN_11256; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11258 = 10'h2bd == _T_174[9:0] ? 4'h0 : _GEN_11257; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11259 = 10'h2be == _T_174[9:0] ? 4'h0 : _GEN_11258; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11260 = 10'h2bf == _T_174[9:0] ? 4'h0 : _GEN_11259; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11261 = 10'h2c0 == _T_174[9:0] ? 4'h3 : _GEN_11260; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11262 = 10'h2c1 == _T_174[9:0] ? 4'h3 : _GEN_11261; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11263 = 10'h2c2 == _T_174[9:0] ? 4'h3 : _GEN_11262; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11264 = 10'h2c3 == _T_174[9:0] ? 4'h3 : _GEN_11263; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11265 = 10'h2c4 == _T_174[9:0] ? 4'h3 : _GEN_11264; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11266 = 10'h2c5 == _T_174[9:0] ? 4'h3 : _GEN_11265; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11267 = 10'h2c6 == _T_174[9:0] ? 4'h4 : _GEN_11266; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11268 = 10'h2c7 == _T_174[9:0] ? 4'h5 : _GEN_11267; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11269 = 10'h2c8 == _T_174[9:0] ? 4'h7 : _GEN_11268; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11270 = 10'h2c9 == _T_174[9:0] ? 4'h7 : _GEN_11269; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11271 = 10'h2ca == _T_174[9:0] ? 4'h4 : _GEN_11270; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11272 = 10'h2cb == _T_174[9:0] ? 4'h9 : _GEN_11271; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11273 = 10'h2cc == _T_174[9:0] ? 4'h9 : _GEN_11272; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11274 = 10'h2cd == _T_174[9:0] ? 4'hb : _GEN_11273; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11275 = 10'h2ce == _T_174[9:0] ? 4'hb : _GEN_11274; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11276 = 10'h2cf == _T_174[9:0] ? 4'hb : _GEN_11275; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11277 = 10'h2d0 == _T_174[9:0] ? 4'hb : _GEN_11276; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11278 = 10'h2d1 == _T_174[9:0] ? 4'hb : _GEN_11277; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11279 = 10'h2d2 == _T_174[9:0] ? 4'h8 : _GEN_11278; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11280 = 10'h2d3 == _T_174[9:0] ? 4'ha : _GEN_11279; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11281 = 10'h2d4 == _T_174[9:0] ? 4'hb : _GEN_11280; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11282 = 10'h2d5 == _T_174[9:0] ? 4'ha : _GEN_11281; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11283 = 10'h2d6 == _T_174[9:0] ? 4'ha : _GEN_11282; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11284 = 10'h2d7 == _T_174[9:0] ? 4'ha : _GEN_11283; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11285 = 10'h2d8 == _T_174[9:0] ? 4'ha : _GEN_11284; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11286 = 10'h2d9 == _T_174[9:0] ? 4'h7 : _GEN_11285; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11287 = 10'h2da == _T_174[9:0] ? 4'h2 : _GEN_11286; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11288 = 10'h2db == _T_174[9:0] ? 4'h0 : _GEN_11287; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11289 = 10'h2dc == _T_174[9:0] ? 4'h0 : _GEN_11288; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11290 = 10'h2dd == _T_174[9:0] ? 4'h0 : _GEN_11289; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11291 = 10'h2de == _T_174[9:0] ? 4'h0 : _GEN_11290; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11292 = 10'h2df == _T_174[9:0] ? 4'h2 : _GEN_11291; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11293 = 10'h2e0 == _T_174[9:0] ? 4'h0 : _GEN_11292; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11294 = 10'h2e1 == _T_174[9:0] ? 4'h0 : _GEN_11293; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11295 = 10'h2e2 == _T_174[9:0] ? 4'h0 : _GEN_11294; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11296 = 10'h2e3 == _T_174[9:0] ? 4'h0 : _GEN_11295; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11297 = 10'h2e4 == _T_174[9:0] ? 4'h0 : _GEN_11296; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11298 = 10'h2e5 == _T_174[9:0] ? 4'h0 : _GEN_11297; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11299 = 10'h2e6 == _T_174[9:0] ? 4'h2 : _GEN_11298; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11300 = 10'h2e7 == _T_174[9:0] ? 4'h3 : _GEN_11299; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11301 = 10'h2e8 == _T_174[9:0] ? 4'h3 : _GEN_11300; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11302 = 10'h2e9 == _T_174[9:0] ? 4'h3 : _GEN_11301; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11303 = 10'h2ea == _T_174[9:0] ? 4'h3 : _GEN_11302; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11304 = 10'h2eb == _T_174[9:0] ? 4'h3 : _GEN_11303; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11305 = 10'h2ec == _T_174[9:0] ? 4'h4 : _GEN_11304; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11306 = 10'h2ed == _T_174[9:0] ? 4'h5 : _GEN_11305; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11307 = 10'h2ee == _T_174[9:0] ? 4'h6 : _GEN_11306; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11308 = 10'h2ef == _T_174[9:0] ? 4'h8 : _GEN_11307; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11309 = 10'h2f0 == _T_174[9:0] ? 4'h4 : _GEN_11308; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11310 = 10'h2f1 == _T_174[9:0] ? 4'h9 : _GEN_11309; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11311 = 10'h2f2 == _T_174[9:0] ? 4'hb : _GEN_11310; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11312 = 10'h2f3 == _T_174[9:0] ? 4'hb : _GEN_11311; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11313 = 10'h2f4 == _T_174[9:0] ? 4'hb : _GEN_11312; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11314 = 10'h2f5 == _T_174[9:0] ? 4'hb : _GEN_11313; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11315 = 10'h2f6 == _T_174[9:0] ? 4'hb : _GEN_11314; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11316 = 10'h2f7 == _T_174[9:0] ? 4'hb : _GEN_11315; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11317 = 10'h2f8 == _T_174[9:0] ? 4'h8 : _GEN_11316; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11318 = 10'h2f9 == _T_174[9:0] ? 4'h9 : _GEN_11317; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11319 = 10'h2fa == _T_174[9:0] ? 4'hb : _GEN_11318; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11320 = 10'h2fb == _T_174[9:0] ? 4'hb : _GEN_11319; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11321 = 10'h2fc == _T_174[9:0] ? 4'ha : _GEN_11320; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11322 = 10'h2fd == _T_174[9:0] ? 4'ha : _GEN_11321; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11323 = 10'h2fe == _T_174[9:0] ? 4'h9 : _GEN_11322; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11324 = 10'h2ff == _T_174[9:0] ? 4'h8 : _GEN_11323; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11325 = 10'h300 == _T_174[9:0] ? 4'h8 : _GEN_11324; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11326 = 10'h301 == _T_174[9:0] ? 4'h6 : _GEN_11325; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11327 = 10'h302 == _T_174[9:0] ? 4'h1 : _GEN_11326; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11328 = 10'h303 == _T_174[9:0] ? 4'h0 : _GEN_11327; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11329 = 10'h304 == _T_174[9:0] ? 4'h0 : _GEN_11328; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11330 = 10'h305 == _T_174[9:0] ? 4'h0 : _GEN_11329; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11331 = 10'h306 == _T_174[9:0] ? 4'h0 : _GEN_11330; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11332 = 10'h307 == _T_174[9:0] ? 4'h0 : _GEN_11331; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11333 = 10'h308 == _T_174[9:0] ? 4'h0 : _GEN_11332; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11334 = 10'h309 == _T_174[9:0] ? 4'h0 : _GEN_11333; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11335 = 10'h30a == _T_174[9:0] ? 4'h0 : _GEN_11334; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11336 = 10'h30b == _T_174[9:0] ? 4'h0 : _GEN_11335; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11337 = 10'h30c == _T_174[9:0] ? 4'h2 : _GEN_11336; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11338 = 10'h30d == _T_174[9:0] ? 4'h3 : _GEN_11337; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11339 = 10'h30e == _T_174[9:0] ? 4'h3 : _GEN_11338; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11340 = 10'h30f == _T_174[9:0] ? 4'h3 : _GEN_11339; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11341 = 10'h310 == _T_174[9:0] ? 4'h3 : _GEN_11340; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11342 = 10'h311 == _T_174[9:0] ? 4'h3 : _GEN_11341; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11343 = 10'h312 == _T_174[9:0] ? 4'h4 : _GEN_11342; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11344 = 10'h313 == _T_174[9:0] ? 4'h5 : _GEN_11343; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11345 = 10'h314 == _T_174[9:0] ? 4'h5 : _GEN_11344; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11346 = 10'h315 == _T_174[9:0] ? 4'h8 : _GEN_11345; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11347 = 10'h316 == _T_174[9:0] ? 4'h4 : _GEN_11346; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11348 = 10'h317 == _T_174[9:0] ? 4'h6 : _GEN_11347; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11349 = 10'h318 == _T_174[9:0] ? 4'hb : _GEN_11348; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11350 = 10'h319 == _T_174[9:0] ? 4'hb : _GEN_11349; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11351 = 10'h31a == _T_174[9:0] ? 4'hb : _GEN_11350; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11352 = 10'h31b == _T_174[9:0] ? 4'hb : _GEN_11351; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11353 = 10'h31c == _T_174[9:0] ? 4'hb : _GEN_11352; // @[Filter.scala 230:102]
  wire [3:0] _GEN_11354 = 10'h31d == _T_174[9:0] ? 4'hb : _GEN_11353; // @[Filter.scala 230:102]
  wire [6:0] _GEN_38980 = {{3'd0}, _GEN_11354}; // @[Filter.scala 230:102]
  wire [10:0] _T_181 = _GEN_38980 * 7'h46; // @[Filter.scala 230:102]
  wire [10:0] _GEN_38981 = {{2'd0}, _T_176}; // @[Filter.scala 230:69]
  wire [10:0] _T_183 = _GEN_38981 + _T_181; // @[Filter.scala 230:69]
  wire [3:0] _GEN_11377 = 10'h16 == _T_174[9:0] ? 4'hb : 4'hc; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11378 = 10'h17 == _T_174[9:0] ? 4'h8 : _GEN_11377; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11379 = 10'h18 == _T_174[9:0] ? 4'ha : _GEN_11378; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11380 = 10'h19 == _T_174[9:0] ? 4'hc : _GEN_11379; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11381 = 10'h1a == _T_174[9:0] ? 4'hc : _GEN_11380; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11382 = 10'h1b == _T_174[9:0] ? 4'hc : _GEN_11381; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11383 = 10'h1c == _T_174[9:0] ? 4'hc : _GEN_11382; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11384 = 10'h1d == _T_174[9:0] ? 4'hc : _GEN_11383; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11385 = 10'h1e == _T_174[9:0] ? 4'hc : _GEN_11384; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11386 = 10'h1f == _T_174[9:0] ? 4'hc : _GEN_11385; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11387 = 10'h20 == _T_174[9:0] ? 4'hc : _GEN_11386; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11388 = 10'h21 == _T_174[9:0] ? 4'hc : _GEN_11387; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11389 = 10'h22 == _T_174[9:0] ? 4'hc : _GEN_11388; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11390 = 10'h23 == _T_174[9:0] ? 4'hc : _GEN_11389; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11391 = 10'h24 == _T_174[9:0] ? 4'hc : _GEN_11390; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11392 = 10'h25 == _T_174[9:0] ? 4'hc : _GEN_11391; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11393 = 10'h26 == _T_174[9:0] ? 4'hc : _GEN_11392; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11394 = 10'h27 == _T_174[9:0] ? 4'hc : _GEN_11393; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11395 = 10'h28 == _T_174[9:0] ? 4'hc : _GEN_11394; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11396 = 10'h29 == _T_174[9:0] ? 4'hc : _GEN_11395; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11397 = 10'h2a == _T_174[9:0] ? 4'hc : _GEN_11396; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11398 = 10'h2b == _T_174[9:0] ? 4'hc : _GEN_11397; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11399 = 10'h2c == _T_174[9:0] ? 4'hc : _GEN_11398; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11400 = 10'h2d == _T_174[9:0] ? 4'hc : _GEN_11399; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11401 = 10'h2e == _T_174[9:0] ? 4'hc : _GEN_11400; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11402 = 10'h2f == _T_174[9:0] ? 4'hc : _GEN_11401; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11403 = 10'h30 == _T_174[9:0] ? 4'hc : _GEN_11402; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11404 = 10'h31 == _T_174[9:0] ? 4'hc : _GEN_11403; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11405 = 10'h32 == _T_174[9:0] ? 4'hc : _GEN_11404; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11406 = 10'h33 == _T_174[9:0] ? 4'hc : _GEN_11405; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11407 = 10'h34 == _T_174[9:0] ? 4'hc : _GEN_11406; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11408 = 10'h35 == _T_174[9:0] ? 4'hc : _GEN_11407; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11409 = 10'h36 == _T_174[9:0] ? 4'hc : _GEN_11408; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11410 = 10'h37 == _T_174[9:0] ? 4'hc : _GEN_11409; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11411 = 10'h38 == _T_174[9:0] ? 4'hc : _GEN_11410; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11412 = 10'h39 == _T_174[9:0] ? 4'hc : _GEN_11411; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11413 = 10'h3a == _T_174[9:0] ? 4'hc : _GEN_11412; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11414 = 10'h3b == _T_174[9:0] ? 4'hc : _GEN_11413; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11415 = 10'h3c == _T_174[9:0] ? 4'h7 : _GEN_11414; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11416 = 10'h3d == _T_174[9:0] ? 4'h9 : _GEN_11415; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11417 = 10'h3e == _T_174[9:0] ? 4'h8 : _GEN_11416; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11418 = 10'h3f == _T_174[9:0] ? 4'hc : _GEN_11417; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11419 = 10'h40 == _T_174[9:0] ? 4'hc : _GEN_11418; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11420 = 10'h41 == _T_174[9:0] ? 4'hc : _GEN_11419; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11421 = 10'h42 == _T_174[9:0] ? 4'hc : _GEN_11420; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11422 = 10'h43 == _T_174[9:0] ? 4'hc : _GEN_11421; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11423 = 10'h44 == _T_174[9:0] ? 4'hc : _GEN_11422; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11424 = 10'h45 == _T_174[9:0] ? 4'hc : _GEN_11423; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11425 = 10'h46 == _T_174[9:0] ? 4'hc : _GEN_11424; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11426 = 10'h47 == _T_174[9:0] ? 4'hc : _GEN_11425; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11427 = 10'h48 == _T_174[9:0] ? 4'hc : _GEN_11426; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11428 = 10'h49 == _T_174[9:0] ? 4'hc : _GEN_11427; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11429 = 10'h4a == _T_174[9:0] ? 4'hc : _GEN_11428; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11430 = 10'h4b == _T_174[9:0] ? 4'hc : _GEN_11429; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11431 = 10'h4c == _T_174[9:0] ? 4'hc : _GEN_11430; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11432 = 10'h4d == _T_174[9:0] ? 4'hc : _GEN_11431; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11433 = 10'h4e == _T_174[9:0] ? 4'hc : _GEN_11432; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11434 = 10'h4f == _T_174[9:0] ? 4'hc : _GEN_11433; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11435 = 10'h50 == _T_174[9:0] ? 4'hc : _GEN_11434; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11436 = 10'h51 == _T_174[9:0] ? 4'hc : _GEN_11435; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11437 = 10'h52 == _T_174[9:0] ? 4'hc : _GEN_11436; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11438 = 10'h53 == _T_174[9:0] ? 4'hc : _GEN_11437; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11439 = 10'h54 == _T_174[9:0] ? 4'hc : _GEN_11438; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11440 = 10'h55 == _T_174[9:0] ? 4'hc : _GEN_11439; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11441 = 10'h56 == _T_174[9:0] ? 4'hc : _GEN_11440; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11442 = 10'h57 == _T_174[9:0] ? 4'hc : _GEN_11441; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11443 = 10'h58 == _T_174[9:0] ? 4'hc : _GEN_11442; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11444 = 10'h59 == _T_174[9:0] ? 4'hc : _GEN_11443; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11445 = 10'h5a == _T_174[9:0] ? 4'h9 : _GEN_11444; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11446 = 10'h5b == _T_174[9:0] ? 4'ha : _GEN_11445; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11447 = 10'h5c == _T_174[9:0] ? 4'hc : _GEN_11446; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11448 = 10'h5d == _T_174[9:0] ? 4'hc : _GEN_11447; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11449 = 10'h5e == _T_174[9:0] ? 4'hc : _GEN_11448; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11450 = 10'h5f == _T_174[9:0] ? 4'hc : _GEN_11449; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11451 = 10'h60 == _T_174[9:0] ? 4'hc : _GEN_11450; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11452 = 10'h61 == _T_174[9:0] ? 4'hb : _GEN_11451; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11453 = 10'h62 == _T_174[9:0] ? 4'h8 : _GEN_11452; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11454 = 10'h63 == _T_174[9:0] ? 4'h9 : _GEN_11453; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11455 = 10'h64 == _T_174[9:0] ? 4'h7 : _GEN_11454; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11456 = 10'h65 == _T_174[9:0] ? 4'hb : _GEN_11455; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11457 = 10'h66 == _T_174[9:0] ? 4'hc : _GEN_11456; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11458 = 10'h67 == _T_174[9:0] ? 4'hc : _GEN_11457; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11459 = 10'h68 == _T_174[9:0] ? 4'hc : _GEN_11458; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11460 = 10'h69 == _T_174[9:0] ? 4'hc : _GEN_11459; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11461 = 10'h6a == _T_174[9:0] ? 4'hc : _GEN_11460; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11462 = 10'h6b == _T_174[9:0] ? 4'hb : _GEN_11461; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11463 = 10'h6c == _T_174[9:0] ? 4'h9 : _GEN_11462; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11464 = 10'h6d == _T_174[9:0] ? 4'ha : _GEN_11463; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11465 = 10'h6e == _T_174[9:0] ? 4'hc : _GEN_11464; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11466 = 10'h6f == _T_174[9:0] ? 4'hc : _GEN_11465; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11467 = 10'h70 == _T_174[9:0] ? 4'hc : _GEN_11466; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11468 = 10'h71 == _T_174[9:0] ? 4'hc : _GEN_11467; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11469 = 10'h72 == _T_174[9:0] ? 4'hc : _GEN_11468; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11470 = 10'h73 == _T_174[9:0] ? 4'hc : _GEN_11469; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11471 = 10'h74 == _T_174[9:0] ? 4'hc : _GEN_11470; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11472 = 10'h75 == _T_174[9:0] ? 4'hc : _GEN_11471; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11473 = 10'h76 == _T_174[9:0] ? 4'hc : _GEN_11472; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11474 = 10'h77 == _T_174[9:0] ? 4'hc : _GEN_11473; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11475 = 10'h78 == _T_174[9:0] ? 4'hc : _GEN_11474; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11476 = 10'h79 == _T_174[9:0] ? 4'hc : _GEN_11475; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11477 = 10'h7a == _T_174[9:0] ? 4'hc : _GEN_11476; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11478 = 10'h7b == _T_174[9:0] ? 4'hc : _GEN_11477; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11479 = 10'h7c == _T_174[9:0] ? 4'hc : _GEN_11478; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11480 = 10'h7d == _T_174[9:0] ? 4'hc : _GEN_11479; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11481 = 10'h7e == _T_174[9:0] ? 4'hc : _GEN_11480; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11482 = 10'h7f == _T_174[9:0] ? 4'hc : _GEN_11481; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11483 = 10'h80 == _T_174[9:0] ? 4'hc : _GEN_11482; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11484 = 10'h81 == _T_174[9:0] ? 4'h9 : _GEN_11483; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11485 = 10'h82 == _T_174[9:0] ? 4'h9 : _GEN_11484; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11486 = 10'h83 == _T_174[9:0] ? 4'h9 : _GEN_11485; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11487 = 10'h84 == _T_174[9:0] ? 4'hc : _GEN_11486; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11488 = 10'h85 == _T_174[9:0] ? 4'hc : _GEN_11487; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11489 = 10'h86 == _T_174[9:0] ? 4'hc : _GEN_11488; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11490 = 10'h87 == _T_174[9:0] ? 4'h8 : _GEN_11489; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11491 = 10'h88 == _T_174[9:0] ? 4'h9 : _GEN_11490; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11492 = 10'h89 == _T_174[9:0] ? 4'h9 : _GEN_11491; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11493 = 10'h8a == _T_174[9:0] ? 4'h9 : _GEN_11492; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11494 = 10'h8b == _T_174[9:0] ? 4'hc : _GEN_11493; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11495 = 10'h8c == _T_174[9:0] ? 4'hc : _GEN_11494; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11496 = 10'h8d == _T_174[9:0] ? 4'hc : _GEN_11495; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11497 = 10'h8e == _T_174[9:0] ? 4'hc : _GEN_11496; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11498 = 10'h8f == _T_174[9:0] ? 4'h9 : _GEN_11497; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11499 = 10'h90 == _T_174[9:0] ? 4'h9 : _GEN_11498; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11500 = 10'h91 == _T_174[9:0] ? 4'h9 : _GEN_11499; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11501 = 10'h92 == _T_174[9:0] ? 4'ha : _GEN_11500; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11502 = 10'h93 == _T_174[9:0] ? 4'hc : _GEN_11501; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11503 = 10'h94 == _T_174[9:0] ? 4'hc : _GEN_11502; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11504 = 10'h95 == _T_174[9:0] ? 4'hc : _GEN_11503; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11505 = 10'h96 == _T_174[9:0] ? 4'hc : _GEN_11504; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11506 = 10'h97 == _T_174[9:0] ? 4'hc : _GEN_11505; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11507 = 10'h98 == _T_174[9:0] ? 4'hc : _GEN_11506; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11508 = 10'h99 == _T_174[9:0] ? 4'hc : _GEN_11507; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11509 = 10'h9a == _T_174[9:0] ? 4'hc : _GEN_11508; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11510 = 10'h9b == _T_174[9:0] ? 4'hc : _GEN_11509; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11511 = 10'h9c == _T_174[9:0] ? 4'hc : _GEN_11510; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11512 = 10'h9d == _T_174[9:0] ? 4'hc : _GEN_11511; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11513 = 10'h9e == _T_174[9:0] ? 4'hc : _GEN_11512; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11514 = 10'h9f == _T_174[9:0] ? 4'hc : _GEN_11513; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11515 = 10'ha0 == _T_174[9:0] ? 4'hc : _GEN_11514; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11516 = 10'ha1 == _T_174[9:0] ? 4'hc : _GEN_11515; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11517 = 10'ha2 == _T_174[9:0] ? 4'hc : _GEN_11516; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11518 = 10'ha3 == _T_174[9:0] ? 4'hc : _GEN_11517; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11519 = 10'ha4 == _T_174[9:0] ? 4'hc : _GEN_11518; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11520 = 10'ha5 == _T_174[9:0] ? 4'hc : _GEN_11519; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11521 = 10'ha6 == _T_174[9:0] ? 4'hc : _GEN_11520; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11522 = 10'ha7 == _T_174[9:0] ? 4'hc : _GEN_11521; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11523 = 10'ha8 == _T_174[9:0] ? 4'h9 : _GEN_11522; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11524 = 10'ha9 == _T_174[9:0] ? 4'h8 : _GEN_11523; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11525 = 10'haa == _T_174[9:0] ? 4'h8 : _GEN_11524; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11526 = 10'hab == _T_174[9:0] ? 4'ha : _GEN_11525; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11527 = 10'hac == _T_174[9:0] ? 4'hb : _GEN_11526; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11528 = 10'had == _T_174[9:0] ? 4'h7 : _GEN_11527; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11529 = 10'hae == _T_174[9:0] ? 4'h9 : _GEN_11528; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11530 = 10'haf == _T_174[9:0] ? 4'h9 : _GEN_11529; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11531 = 10'hb0 == _T_174[9:0] ? 4'h8 : _GEN_11530; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11532 = 10'hb1 == _T_174[9:0] ? 4'h9 : _GEN_11531; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11533 = 10'hb2 == _T_174[9:0] ? 4'hc : _GEN_11532; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11534 = 10'hb3 == _T_174[9:0] ? 4'h9 : _GEN_11533; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11535 = 10'hb4 == _T_174[9:0] ? 4'h9 : _GEN_11534; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11536 = 10'hb5 == _T_174[9:0] ? 4'h9 : _GEN_11535; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11537 = 10'hb6 == _T_174[9:0] ? 4'h9 : _GEN_11536; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11538 = 10'hb7 == _T_174[9:0] ? 4'ha : _GEN_11537; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11539 = 10'hb8 == _T_174[9:0] ? 4'hc : _GEN_11538; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11540 = 10'hb9 == _T_174[9:0] ? 4'hc : _GEN_11539; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11541 = 10'hba == _T_174[9:0] ? 4'hc : _GEN_11540; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11542 = 10'hbb == _T_174[9:0] ? 4'hc : _GEN_11541; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11543 = 10'hbc == _T_174[9:0] ? 4'hc : _GEN_11542; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11544 = 10'hbd == _T_174[9:0] ? 4'hb : _GEN_11543; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11545 = 10'hbe == _T_174[9:0] ? 4'hc : _GEN_11544; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11546 = 10'hbf == _T_174[9:0] ? 4'hc : _GEN_11545; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11547 = 10'hc0 == _T_174[9:0] ? 4'hc : _GEN_11546; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11548 = 10'hc1 == _T_174[9:0] ? 4'hc : _GEN_11547; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11549 = 10'hc2 == _T_174[9:0] ? 4'hc : _GEN_11548; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11550 = 10'hc3 == _T_174[9:0] ? 4'hc : _GEN_11549; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11551 = 10'hc4 == _T_174[9:0] ? 4'hc : _GEN_11550; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11552 = 10'hc5 == _T_174[9:0] ? 4'hc : _GEN_11551; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11553 = 10'hc6 == _T_174[9:0] ? 4'hb : _GEN_11552; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11554 = 10'hc7 == _T_174[9:0] ? 4'hb : _GEN_11553; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11555 = 10'hc8 == _T_174[9:0] ? 4'ha : _GEN_11554; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11556 = 10'hc9 == _T_174[9:0] ? 4'ha : _GEN_11555; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11557 = 10'hca == _T_174[9:0] ? 4'hb : _GEN_11556; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11558 = 10'hcb == _T_174[9:0] ? 4'hc : _GEN_11557; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11559 = 10'hcc == _T_174[9:0] ? 4'hc : _GEN_11558; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11560 = 10'hcd == _T_174[9:0] ? 4'hc : _GEN_11559; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11561 = 10'hce == _T_174[9:0] ? 4'ha : _GEN_11560; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11562 = 10'hcf == _T_174[9:0] ? 4'h8 : _GEN_11561; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11563 = 10'hd0 == _T_174[9:0] ? 4'h9 : _GEN_11562; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11564 = 10'hd1 == _T_174[9:0] ? 4'h8 : _GEN_11563; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11565 = 10'hd2 == _T_174[9:0] ? 4'h9 : _GEN_11564; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11566 = 10'hd3 == _T_174[9:0] ? 4'h9 : _GEN_11565; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11567 = 10'hd4 == _T_174[9:0] ? 4'h9 : _GEN_11566; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11568 = 10'hd5 == _T_174[9:0] ? 4'h9 : _GEN_11567; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11569 = 10'hd6 == _T_174[9:0] ? 4'ha : _GEN_11568; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11570 = 10'hd7 == _T_174[9:0] ? 4'h9 : _GEN_11569; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11571 = 10'hd8 == _T_174[9:0] ? 4'h9 : _GEN_11570; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11572 = 10'hd9 == _T_174[9:0] ? 4'h9 : _GEN_11571; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11573 = 10'hda == _T_174[9:0] ? 4'ha : _GEN_11572; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11574 = 10'hdb == _T_174[9:0] ? 4'h9 : _GEN_11573; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11575 = 10'hdc == _T_174[9:0] ? 4'h7 : _GEN_11574; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11576 = 10'hdd == _T_174[9:0] ? 4'hc : _GEN_11575; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11577 = 10'hde == _T_174[9:0] ? 4'hc : _GEN_11576; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11578 = 10'hdf == _T_174[9:0] ? 4'hc : _GEN_11577; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11579 = 10'he0 == _T_174[9:0] ? 4'hc : _GEN_11578; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11580 = 10'he1 == _T_174[9:0] ? 4'hc : _GEN_11579; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11581 = 10'he2 == _T_174[9:0] ? 4'hc : _GEN_11580; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11582 = 10'he3 == _T_174[9:0] ? 4'h8 : _GEN_11581; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11583 = 10'he4 == _T_174[9:0] ? 4'hc : _GEN_11582; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11584 = 10'he5 == _T_174[9:0] ? 4'hc : _GEN_11583; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11585 = 10'he6 == _T_174[9:0] ? 4'hc : _GEN_11584; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11586 = 10'he7 == _T_174[9:0] ? 4'hc : _GEN_11585; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11587 = 10'he8 == _T_174[9:0] ? 4'hc : _GEN_11586; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11588 = 10'he9 == _T_174[9:0] ? 4'hc : _GEN_11587; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11589 = 10'hea == _T_174[9:0] ? 4'hc : _GEN_11588; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11590 = 10'heb == _T_174[9:0] ? 4'ha : _GEN_11589; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11591 = 10'hec == _T_174[9:0] ? 4'h7 : _GEN_11590; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11592 = 10'hed == _T_174[9:0] ? 4'h3 : _GEN_11591; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11593 = 10'hee == _T_174[9:0] ? 4'h3 : _GEN_11592; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11594 = 10'hef == _T_174[9:0] ? 4'h3 : _GEN_11593; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11595 = 10'hf0 == _T_174[9:0] ? 4'h3 : _GEN_11594; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11596 = 10'hf1 == _T_174[9:0] ? 4'h8 : _GEN_11595; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11597 = 10'hf2 == _T_174[9:0] ? 4'hc : _GEN_11596; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11598 = 10'hf3 == _T_174[9:0] ? 4'hc : _GEN_11597; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11599 = 10'hf4 == _T_174[9:0] ? 4'hc : _GEN_11598; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11600 = 10'hf5 == _T_174[9:0] ? 4'h9 : _GEN_11599; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11601 = 10'hf6 == _T_174[9:0] ? 4'h9 : _GEN_11600; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11602 = 10'hf7 == _T_174[9:0] ? 4'h9 : _GEN_11601; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11603 = 10'hf8 == _T_174[9:0] ? 4'h9 : _GEN_11602; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11604 = 10'hf9 == _T_174[9:0] ? 4'ha : _GEN_11603; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11605 = 10'hfa == _T_174[9:0] ? 4'h9 : _GEN_11604; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11606 = 10'hfb == _T_174[9:0] ? 4'h9 : _GEN_11605; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11607 = 10'hfc == _T_174[9:0] ? 4'h9 : _GEN_11606; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11608 = 10'hfd == _T_174[9:0] ? 4'h9 : _GEN_11607; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11609 = 10'hfe == _T_174[9:0] ? 4'h9 : _GEN_11608; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11610 = 10'hff == _T_174[9:0] ? 4'ha : _GEN_11609; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11611 = 10'h100 == _T_174[9:0] ? 4'ha : _GEN_11610; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11612 = 10'h101 == _T_174[9:0] ? 4'h7 : _GEN_11611; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11613 = 10'h102 == _T_174[9:0] ? 4'h9 : _GEN_11612; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11614 = 10'h103 == _T_174[9:0] ? 4'hc : _GEN_11613; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11615 = 10'h104 == _T_174[9:0] ? 4'hc : _GEN_11614; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11616 = 10'h105 == _T_174[9:0] ? 4'hb : _GEN_11615; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11617 = 10'h106 == _T_174[9:0] ? 4'hb : _GEN_11616; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11618 = 10'h107 == _T_174[9:0] ? 4'hb : _GEN_11617; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11619 = 10'h108 == _T_174[9:0] ? 4'hb : _GEN_11618; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11620 = 10'h109 == _T_174[9:0] ? 4'h7 : _GEN_11619; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11621 = 10'h10a == _T_174[9:0] ? 4'hc : _GEN_11620; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11622 = 10'h10b == _T_174[9:0] ? 4'hc : _GEN_11621; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11623 = 10'h10c == _T_174[9:0] ? 4'hc : _GEN_11622; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11624 = 10'h10d == _T_174[9:0] ? 4'hc : _GEN_11623; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11625 = 10'h10e == _T_174[9:0] ? 4'hc : _GEN_11624; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11626 = 10'h10f == _T_174[9:0] ? 4'h9 : _GEN_11625; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11627 = 10'h110 == _T_174[9:0] ? 4'hb : _GEN_11626; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11628 = 10'h111 == _T_174[9:0] ? 4'h4 : _GEN_11627; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11629 = 10'h112 == _T_174[9:0] ? 4'h7 : _GEN_11628; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11630 = 10'h113 == _T_174[9:0] ? 4'h3 : _GEN_11629; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11631 = 10'h114 == _T_174[9:0] ? 4'h3 : _GEN_11630; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11632 = 10'h115 == _T_174[9:0] ? 4'h3 : _GEN_11631; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11633 = 10'h116 == _T_174[9:0] ? 4'h3 : _GEN_11632; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11634 = 10'h117 == _T_174[9:0] ? 4'h2 : _GEN_11633; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11635 = 10'h118 == _T_174[9:0] ? 4'h9 : _GEN_11634; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11636 = 10'h119 == _T_174[9:0] ? 4'hc : _GEN_11635; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11637 = 10'h11a == _T_174[9:0] ? 4'hc : _GEN_11636; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11638 = 10'h11b == _T_174[9:0] ? 4'hc : _GEN_11637; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11639 = 10'h11c == _T_174[9:0] ? 4'h9 : _GEN_11638; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11640 = 10'h11d == _T_174[9:0] ? 4'h9 : _GEN_11639; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11641 = 10'h11e == _T_174[9:0] ? 4'h9 : _GEN_11640; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11642 = 10'h11f == _T_174[9:0] ? 4'h8 : _GEN_11641; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11643 = 10'h120 == _T_174[9:0] ? 4'h7 : _GEN_11642; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11644 = 10'h121 == _T_174[9:0] ? 4'h9 : _GEN_11643; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11645 = 10'h122 == _T_174[9:0] ? 4'h7 : _GEN_11644; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11646 = 10'h123 == _T_174[9:0] ? 4'h7 : _GEN_11645; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11647 = 10'h124 == _T_174[9:0] ? 4'h9 : _GEN_11646; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11648 = 10'h125 == _T_174[9:0] ? 4'h9 : _GEN_11647; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11649 = 10'h126 == _T_174[9:0] ? 4'h8 : _GEN_11648; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11650 = 10'h127 == _T_174[9:0] ? 4'h9 : _GEN_11649; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11651 = 10'h128 == _T_174[9:0] ? 4'h8 : _GEN_11650; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11652 = 10'h129 == _T_174[9:0] ? 4'ha : _GEN_11651; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11653 = 10'h12a == _T_174[9:0] ? 4'h5 : _GEN_11652; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11654 = 10'h12b == _T_174[9:0] ? 4'h3 : _GEN_11653; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11655 = 10'h12c == _T_174[9:0] ? 4'h3 : _GEN_11654; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11656 = 10'h12d == _T_174[9:0] ? 4'h3 : _GEN_11655; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11657 = 10'h12e == _T_174[9:0] ? 4'h5 : _GEN_11656; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11658 = 10'h12f == _T_174[9:0] ? 4'h8 : _GEN_11657; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11659 = 10'h130 == _T_174[9:0] ? 4'hc : _GEN_11658; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11660 = 10'h131 == _T_174[9:0] ? 4'hb : _GEN_11659; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11661 = 10'h132 == _T_174[9:0] ? 4'h9 : _GEN_11660; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11662 = 10'h133 == _T_174[9:0] ? 4'h8 : _GEN_11661; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11663 = 10'h134 == _T_174[9:0] ? 4'h9 : _GEN_11662; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11664 = 10'h135 == _T_174[9:0] ? 4'h7 : _GEN_11663; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11665 = 10'h136 == _T_174[9:0] ? 4'h7 : _GEN_11664; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11666 = 10'h137 == _T_174[9:0] ? 4'h5 : _GEN_11665; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11667 = 10'h138 == _T_174[9:0] ? 4'h7 : _GEN_11666; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11668 = 10'h139 == _T_174[9:0] ? 4'h3 : _GEN_11667; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11669 = 10'h13a == _T_174[9:0] ? 4'h3 : _GEN_11668; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11670 = 10'h13b == _T_174[9:0] ? 4'h3 : _GEN_11669; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11671 = 10'h13c == _T_174[9:0] ? 4'h3 : _GEN_11670; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11672 = 10'h13d == _T_174[9:0] ? 4'h3 : _GEN_11671; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11673 = 10'h13e == _T_174[9:0] ? 4'h5 : _GEN_11672; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11674 = 10'h13f == _T_174[9:0] ? 4'ha : _GEN_11673; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11675 = 10'h140 == _T_174[9:0] ? 4'hc : _GEN_11674; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11676 = 10'h141 == _T_174[9:0] ? 4'hc : _GEN_11675; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11677 = 10'h142 == _T_174[9:0] ? 4'hc : _GEN_11676; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11678 = 10'h143 == _T_174[9:0] ? 4'h9 : _GEN_11677; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11679 = 10'h144 == _T_174[9:0] ? 4'h9 : _GEN_11678; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11680 = 10'h145 == _T_174[9:0] ? 4'h8 : _GEN_11679; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11681 = 10'h146 == _T_174[9:0] ? 4'h8 : _GEN_11680; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11682 = 10'h147 == _T_174[9:0] ? 4'h7 : _GEN_11681; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11683 = 10'h148 == _T_174[9:0] ? 4'h8 : _GEN_11682; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11684 = 10'h149 == _T_174[9:0] ? 4'h9 : _GEN_11683; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11685 = 10'h14a == _T_174[9:0] ? 4'ha : _GEN_11684; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11686 = 10'h14b == _T_174[9:0] ? 4'h9 : _GEN_11685; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11687 = 10'h14c == _T_174[9:0] ? 4'ha : _GEN_11686; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11688 = 10'h14d == _T_174[9:0] ? 4'h9 : _GEN_11687; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11689 = 10'h14e == _T_174[9:0] ? 4'h7 : _GEN_11688; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11690 = 10'h14f == _T_174[9:0] ? 4'h3 : _GEN_11689; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11691 = 10'h150 == _T_174[9:0] ? 4'h3 : _GEN_11690; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11692 = 10'h151 == _T_174[9:0] ? 4'h3 : _GEN_11691; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11693 = 10'h152 == _T_174[9:0] ? 4'h3 : _GEN_11692; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11694 = 10'h153 == _T_174[9:0] ? 4'h3 : _GEN_11693; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11695 = 10'h154 == _T_174[9:0] ? 4'h3 : _GEN_11694; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11696 = 10'h155 == _T_174[9:0] ? 4'h8 : _GEN_11695; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11697 = 10'h156 == _T_174[9:0] ? 4'ha : _GEN_11696; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11698 = 10'h157 == _T_174[9:0] ? 4'h7 : _GEN_11697; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11699 = 10'h158 == _T_174[9:0] ? 4'h7 : _GEN_11698; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11700 = 10'h159 == _T_174[9:0] ? 4'h7 : _GEN_11699; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11701 = 10'h15a == _T_174[9:0] ? 4'h7 : _GEN_11700; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11702 = 10'h15b == _T_174[9:0] ? 4'h7 : _GEN_11701; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11703 = 10'h15c == _T_174[9:0] ? 4'h7 : _GEN_11702; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11704 = 10'h15d == _T_174[9:0] ? 4'h7 : _GEN_11703; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11705 = 10'h15e == _T_174[9:0] ? 4'h7 : _GEN_11704; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11706 = 10'h15f == _T_174[9:0] ? 4'h3 : _GEN_11705; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11707 = 10'h160 == _T_174[9:0] ? 4'h3 : _GEN_11706; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11708 = 10'h161 == _T_174[9:0] ? 4'h3 : _GEN_11707; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11709 = 10'h162 == _T_174[9:0] ? 4'h3 : _GEN_11708; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11710 = 10'h163 == _T_174[9:0] ? 4'h3 : _GEN_11709; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11711 = 10'h164 == _T_174[9:0] ? 4'h4 : _GEN_11710; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11712 = 10'h165 == _T_174[9:0] ? 4'ha : _GEN_11711; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11713 = 10'h166 == _T_174[9:0] ? 4'ha : _GEN_11712; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11714 = 10'h167 == _T_174[9:0] ? 4'hc : _GEN_11713; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11715 = 10'h168 == _T_174[9:0] ? 4'hc : _GEN_11714; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11716 = 10'h169 == _T_174[9:0] ? 4'h9 : _GEN_11715; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11717 = 10'h16a == _T_174[9:0] ? 4'h9 : _GEN_11716; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11718 = 10'h16b == _T_174[9:0] ? 4'ha : _GEN_11717; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11719 = 10'h16c == _T_174[9:0] ? 4'h7 : _GEN_11718; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11720 = 10'h16d == _T_174[9:0] ? 4'h7 : _GEN_11719; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11721 = 10'h16e == _T_174[9:0] ? 4'h7 : _GEN_11720; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11722 = 10'h16f == _T_174[9:0] ? 4'ha : _GEN_11721; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11723 = 10'h170 == _T_174[9:0] ? 4'ha : _GEN_11722; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11724 = 10'h171 == _T_174[9:0] ? 4'ha : _GEN_11723; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11725 = 10'h172 == _T_174[9:0] ? 4'hc : _GEN_11724; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11726 = 10'h173 == _T_174[9:0] ? 4'h8 : _GEN_11725; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11727 = 10'h174 == _T_174[9:0] ? 4'h5 : _GEN_11726; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11728 = 10'h175 == _T_174[9:0] ? 4'h8 : _GEN_11727; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11729 = 10'h176 == _T_174[9:0] ? 4'h7 : _GEN_11728; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11730 = 10'h177 == _T_174[9:0] ? 4'h8 : _GEN_11729; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11731 = 10'h178 == _T_174[9:0] ? 4'h7 : _GEN_11730; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11732 = 10'h179 == _T_174[9:0] ? 4'h5 : _GEN_11731; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11733 = 10'h17a == _T_174[9:0] ? 4'h5 : _GEN_11732; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11734 = 10'h17b == _T_174[9:0] ? 4'h7 : _GEN_11733; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11735 = 10'h17c == _T_174[9:0] ? 4'h7 : _GEN_11734; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11736 = 10'h17d == _T_174[9:0] ? 4'h7 : _GEN_11735; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11737 = 10'h17e == _T_174[9:0] ? 4'h7 : _GEN_11736; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11738 = 10'h17f == _T_174[9:0] ? 4'h7 : _GEN_11737; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11739 = 10'h180 == _T_174[9:0] ? 4'h7 : _GEN_11738; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11740 = 10'h181 == _T_174[9:0] ? 4'h7 : _GEN_11739; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11741 = 10'h182 == _T_174[9:0] ? 4'h7 : _GEN_11740; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11742 = 10'h183 == _T_174[9:0] ? 4'h7 : _GEN_11741; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11743 = 10'h184 == _T_174[9:0] ? 4'h7 : _GEN_11742; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11744 = 10'h185 == _T_174[9:0] ? 4'h5 : _GEN_11743; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11745 = 10'h186 == _T_174[9:0] ? 4'h3 : _GEN_11744; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11746 = 10'h187 == _T_174[9:0] ? 4'h3 : _GEN_11745; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11747 = 10'h188 == _T_174[9:0] ? 4'h3 : _GEN_11746; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11748 = 10'h189 == _T_174[9:0] ? 4'h4 : _GEN_11747; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11749 = 10'h18a == _T_174[9:0] ? 4'h5 : _GEN_11748; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11750 = 10'h18b == _T_174[9:0] ? 4'ha : _GEN_11749; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11751 = 10'h18c == _T_174[9:0] ? 4'ha : _GEN_11750; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11752 = 10'h18d == _T_174[9:0] ? 4'ha : _GEN_11751; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11753 = 10'h18e == _T_174[9:0] ? 4'hc : _GEN_11752; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11754 = 10'h18f == _T_174[9:0] ? 4'h8 : _GEN_11753; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11755 = 10'h190 == _T_174[9:0] ? 4'h9 : _GEN_11754; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11756 = 10'h191 == _T_174[9:0] ? 4'h8 : _GEN_11755; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11757 = 10'h192 == _T_174[9:0] ? 4'h7 : _GEN_11756; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11758 = 10'h193 == _T_174[9:0] ? 4'h7 : _GEN_11757; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11759 = 10'h194 == _T_174[9:0] ? 4'h7 : _GEN_11758; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11760 = 10'h195 == _T_174[9:0] ? 4'h9 : _GEN_11759; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11761 = 10'h196 == _T_174[9:0] ? 4'ha : _GEN_11760; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11762 = 10'h197 == _T_174[9:0] ? 4'h8 : _GEN_11761; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11763 = 10'h198 == _T_174[9:0] ? 4'hc : _GEN_11762; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11764 = 10'h199 == _T_174[9:0] ? 4'h5 : _GEN_11763; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11765 = 10'h19a == _T_174[9:0] ? 4'h1 : _GEN_11764; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11766 = 10'h19b == _T_174[9:0] ? 4'h4 : _GEN_11765; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11767 = 10'h19c == _T_174[9:0] ? 4'h7 : _GEN_11766; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11768 = 10'h19d == _T_174[9:0] ? 4'h5 : _GEN_11767; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11769 = 10'h19e == _T_174[9:0] ? 4'h2 : _GEN_11768; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11770 = 10'h19f == _T_174[9:0] ? 4'h3 : _GEN_11769; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11771 = 10'h1a0 == _T_174[9:0] ? 4'h7 : _GEN_11770; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11772 = 10'h1a1 == _T_174[9:0] ? 4'h7 : _GEN_11771; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11773 = 10'h1a2 == _T_174[9:0] ? 4'h7 : _GEN_11772; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11774 = 10'h1a3 == _T_174[9:0] ? 4'h7 : _GEN_11773; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11775 = 10'h1a4 == _T_174[9:0] ? 4'h7 : _GEN_11774; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11776 = 10'h1a5 == _T_174[9:0] ? 4'h7 : _GEN_11775; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11777 = 10'h1a6 == _T_174[9:0] ? 4'h7 : _GEN_11776; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11778 = 10'h1a7 == _T_174[9:0] ? 4'h7 : _GEN_11777; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11779 = 10'h1a8 == _T_174[9:0] ? 4'h8 : _GEN_11778; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11780 = 10'h1a9 == _T_174[9:0] ? 4'h8 : _GEN_11779; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11781 = 10'h1aa == _T_174[9:0] ? 4'h6 : _GEN_11780; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11782 = 10'h1ab == _T_174[9:0] ? 4'h6 : _GEN_11781; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11783 = 10'h1ac == _T_174[9:0] ? 4'h5 : _GEN_11782; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11784 = 10'h1ad == _T_174[9:0] ? 4'h4 : _GEN_11783; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11785 = 10'h1ae == _T_174[9:0] ? 4'h3 : _GEN_11784; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11786 = 10'h1af == _T_174[9:0] ? 4'h6 : _GEN_11785; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11787 = 10'h1b0 == _T_174[9:0] ? 4'h6 : _GEN_11786; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11788 = 10'h1b1 == _T_174[9:0] ? 4'ha : _GEN_11787; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11789 = 10'h1b2 == _T_174[9:0] ? 4'ha : _GEN_11788; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11790 = 10'h1b3 == _T_174[9:0] ? 4'h9 : _GEN_11789; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11791 = 10'h1b4 == _T_174[9:0] ? 4'hb : _GEN_11790; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11792 = 10'h1b5 == _T_174[9:0] ? 4'h8 : _GEN_11791; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11793 = 10'h1b6 == _T_174[9:0] ? 4'h8 : _GEN_11792; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11794 = 10'h1b7 == _T_174[9:0] ? 4'h7 : _GEN_11793; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11795 = 10'h1b8 == _T_174[9:0] ? 4'h6 : _GEN_11794; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11796 = 10'h1b9 == _T_174[9:0] ? 4'h7 : _GEN_11795; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11797 = 10'h1ba == _T_174[9:0] ? 4'h6 : _GEN_11796; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11798 = 10'h1bb == _T_174[9:0] ? 4'h8 : _GEN_11797; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11799 = 10'h1bc == _T_174[9:0] ? 4'ha : _GEN_11798; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11800 = 10'h1bd == _T_174[9:0] ? 4'h9 : _GEN_11799; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11801 = 10'h1be == _T_174[9:0] ? 4'hc : _GEN_11800; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11802 = 10'h1bf == _T_174[9:0] ? 4'h7 : _GEN_11801; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11803 = 10'h1c0 == _T_174[9:0] ? 4'h6 : _GEN_11802; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11804 = 10'h1c1 == _T_174[9:0] ? 4'h7 : _GEN_11803; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11805 = 10'h1c2 == _T_174[9:0] ? 4'h7 : _GEN_11804; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11806 = 10'h1c3 == _T_174[9:0] ? 4'h6 : _GEN_11805; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11807 = 10'h1c4 == _T_174[9:0] ? 4'h5 : _GEN_11806; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11808 = 10'h1c5 == _T_174[9:0] ? 4'h6 : _GEN_11807; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11809 = 10'h1c6 == _T_174[9:0] ? 4'h8 : _GEN_11808; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11810 = 10'h1c7 == _T_174[9:0] ? 4'h7 : _GEN_11809; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11811 = 10'h1c8 == _T_174[9:0] ? 4'h7 : _GEN_11810; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11812 = 10'h1c9 == _T_174[9:0] ? 4'h7 : _GEN_11811; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11813 = 10'h1ca == _T_174[9:0] ? 4'h7 : _GEN_11812; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11814 = 10'h1cb == _T_174[9:0] ? 4'h7 : _GEN_11813; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11815 = 10'h1cc == _T_174[9:0] ? 4'h7 : _GEN_11814; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11816 = 10'h1cd == _T_174[9:0] ? 4'h8 : _GEN_11815; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11817 = 10'h1ce == _T_174[9:0] ? 4'h8 : _GEN_11816; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11818 = 10'h1cf == _T_174[9:0] ? 4'h8 : _GEN_11817; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11819 = 10'h1d0 == _T_174[9:0] ? 4'h5 : _GEN_11818; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11820 = 10'h1d1 == _T_174[9:0] ? 4'h6 : _GEN_11819; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11821 = 10'h1d2 == _T_174[9:0] ? 4'h7 : _GEN_11820; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11822 = 10'h1d3 == _T_174[9:0] ? 4'h7 : _GEN_11821; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11823 = 10'h1d4 == _T_174[9:0] ? 4'h7 : _GEN_11822; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11824 = 10'h1d5 == _T_174[9:0] ? 4'h6 : _GEN_11823; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11825 = 10'h1d6 == _T_174[9:0] ? 4'h8 : _GEN_11824; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11826 = 10'h1d7 == _T_174[9:0] ? 4'ha : _GEN_11825; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11827 = 10'h1d8 == _T_174[9:0] ? 4'ha : _GEN_11826; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11828 = 10'h1d9 == _T_174[9:0] ? 4'ha : _GEN_11827; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11829 = 10'h1da == _T_174[9:0] ? 4'h8 : _GEN_11828; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11830 = 10'h1db == _T_174[9:0] ? 4'h9 : _GEN_11829; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11831 = 10'h1dc == _T_174[9:0] ? 4'h9 : _GEN_11830; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11832 = 10'h1dd == _T_174[9:0] ? 4'h5 : _GEN_11831; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11833 = 10'h1de == _T_174[9:0] ? 4'h7 : _GEN_11832; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11834 = 10'h1df == _T_174[9:0] ? 4'h7 : _GEN_11833; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11835 = 10'h1e0 == _T_174[9:0] ? 4'h7 : _GEN_11834; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11836 = 10'h1e1 == _T_174[9:0] ? 4'h6 : _GEN_11835; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11837 = 10'h1e2 == _T_174[9:0] ? 4'h9 : _GEN_11836; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11838 = 10'h1e3 == _T_174[9:0] ? 4'h9 : _GEN_11837; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11839 = 10'h1e4 == _T_174[9:0] ? 4'hb : _GEN_11838; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11840 = 10'h1e5 == _T_174[9:0] ? 4'h8 : _GEN_11839; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11841 = 10'h1e6 == _T_174[9:0] ? 4'h7 : _GEN_11840; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11842 = 10'h1e7 == _T_174[9:0] ? 4'h8 : _GEN_11841; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11843 = 10'h1e8 == _T_174[9:0] ? 4'h8 : _GEN_11842; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11844 = 10'h1e9 == _T_174[9:0] ? 4'h8 : _GEN_11843; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11845 = 10'h1ea == _T_174[9:0] ? 4'h8 : _GEN_11844; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11846 = 10'h1eb == _T_174[9:0] ? 4'h8 : _GEN_11845; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11847 = 10'h1ec == _T_174[9:0] ? 4'h8 : _GEN_11846; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11848 = 10'h1ed == _T_174[9:0] ? 4'h6 : _GEN_11847; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11849 = 10'h1ee == _T_174[9:0] ? 4'h7 : _GEN_11848; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11850 = 10'h1ef == _T_174[9:0] ? 4'h7 : _GEN_11849; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11851 = 10'h1f0 == _T_174[9:0] ? 4'h7 : _GEN_11850; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11852 = 10'h1f1 == _T_174[9:0] ? 4'h7 : _GEN_11851; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11853 = 10'h1f2 == _T_174[9:0] ? 4'h7 : _GEN_11852; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11854 = 10'h1f3 == _T_174[9:0] ? 4'h8 : _GEN_11853; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11855 = 10'h1f4 == _T_174[9:0] ? 4'h8 : _GEN_11854; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11856 = 10'h1f5 == _T_174[9:0] ? 4'h8 : _GEN_11855; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11857 = 10'h1f6 == _T_174[9:0] ? 4'ha : _GEN_11856; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11858 = 10'h1f7 == _T_174[9:0] ? 4'h6 : _GEN_11857; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11859 = 10'h1f8 == _T_174[9:0] ? 4'h6 : _GEN_11858; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11860 = 10'h1f9 == _T_174[9:0] ? 4'h8 : _GEN_11859; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11861 = 10'h1fa == _T_174[9:0] ? 4'h8 : _GEN_11860; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11862 = 10'h1fb == _T_174[9:0] ? 4'h6 : _GEN_11861; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11863 = 10'h1fc == _T_174[9:0] ? 4'ha : _GEN_11862; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11864 = 10'h1fd == _T_174[9:0] ? 4'hb : _GEN_11863; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11865 = 10'h1fe == _T_174[9:0] ? 4'ha : _GEN_11864; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11866 = 10'h1ff == _T_174[9:0] ? 4'ha : _GEN_11865; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11867 = 10'h200 == _T_174[9:0] ? 4'h4 : _GEN_11866; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11868 = 10'h201 == _T_174[9:0] ? 4'h7 : _GEN_11867; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11869 = 10'h202 == _T_174[9:0] ? 4'h6 : _GEN_11868; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11870 = 10'h203 == _T_174[9:0] ? 4'h6 : _GEN_11869; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11871 = 10'h204 == _T_174[9:0] ? 4'h5 : _GEN_11870; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11872 = 10'h205 == _T_174[9:0] ? 4'h6 : _GEN_11871; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11873 = 10'h206 == _T_174[9:0] ? 4'h6 : _GEN_11872; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11874 = 10'h207 == _T_174[9:0] ? 4'h5 : _GEN_11873; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11875 = 10'h208 == _T_174[9:0] ? 4'h7 : _GEN_11874; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11876 = 10'h209 == _T_174[9:0] ? 4'h9 : _GEN_11875; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11877 = 10'h20a == _T_174[9:0] ? 4'hb : _GEN_11876; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11878 = 10'h20b == _T_174[9:0] ? 4'h7 : _GEN_11877; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11879 = 10'h20c == _T_174[9:0] ? 4'h7 : _GEN_11878; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11880 = 10'h20d == _T_174[9:0] ? 4'h7 : _GEN_11879; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11881 = 10'h20e == _T_174[9:0] ? 4'h7 : _GEN_11880; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11882 = 10'h20f == _T_174[9:0] ? 4'h7 : _GEN_11881; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11883 = 10'h210 == _T_174[9:0] ? 4'h7 : _GEN_11882; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11884 = 10'h211 == _T_174[9:0] ? 4'h8 : _GEN_11883; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11885 = 10'h212 == _T_174[9:0] ? 4'h8 : _GEN_11884; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11886 = 10'h213 == _T_174[9:0] ? 4'h9 : _GEN_11885; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11887 = 10'h214 == _T_174[9:0] ? 4'h6 : _GEN_11886; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11888 = 10'h215 == _T_174[9:0] ? 4'h7 : _GEN_11887; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11889 = 10'h216 == _T_174[9:0] ? 4'h7 : _GEN_11888; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11890 = 10'h217 == _T_174[9:0] ? 4'h7 : _GEN_11889; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11891 = 10'h218 == _T_174[9:0] ? 4'h7 : _GEN_11890; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11892 = 10'h219 == _T_174[9:0] ? 4'h8 : _GEN_11891; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11893 = 10'h21a == _T_174[9:0] ? 4'h7 : _GEN_11892; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11894 = 10'h21b == _T_174[9:0] ? 4'h8 : _GEN_11893; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11895 = 10'h21c == _T_174[9:0] ? 4'ha : _GEN_11894; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11896 = 10'h21d == _T_174[9:0] ? 4'ha : _GEN_11895; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11897 = 10'h21e == _T_174[9:0] ? 4'h7 : _GEN_11896; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11898 = 10'h21f == _T_174[9:0] ? 4'h6 : _GEN_11897; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11899 = 10'h220 == _T_174[9:0] ? 4'h6 : _GEN_11898; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11900 = 10'h221 == _T_174[9:0] ? 4'h7 : _GEN_11899; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11901 = 10'h222 == _T_174[9:0] ? 4'ha : _GEN_11900; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11902 = 10'h223 == _T_174[9:0] ? 4'ha : _GEN_11901; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11903 = 10'h224 == _T_174[9:0] ? 4'ha : _GEN_11902; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11904 = 10'h225 == _T_174[9:0] ? 4'h8 : _GEN_11903; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11905 = 10'h226 == _T_174[9:0] ? 4'h3 : _GEN_11904; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11906 = 10'h227 == _T_174[9:0] ? 4'h4 : _GEN_11905; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11907 = 10'h228 == _T_174[9:0] ? 4'h6 : _GEN_11906; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11908 = 10'h229 == _T_174[9:0] ? 4'h6 : _GEN_11907; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11909 = 10'h22a == _T_174[9:0] ? 4'h6 : _GEN_11908; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11910 = 10'h22b == _T_174[9:0] ? 4'h6 : _GEN_11909; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11911 = 10'h22c == _T_174[9:0] ? 4'h5 : _GEN_11910; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11912 = 10'h22d == _T_174[9:0] ? 4'h6 : _GEN_11911; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11913 = 10'h22e == _T_174[9:0] ? 4'h6 : _GEN_11912; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11914 = 10'h22f == _T_174[9:0] ? 4'h8 : _GEN_11913; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11915 = 10'h230 == _T_174[9:0] ? 4'h7 : _GEN_11914; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11916 = 10'h231 == _T_174[9:0] ? 4'h5 : _GEN_11915; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11917 = 10'h232 == _T_174[9:0] ? 4'h6 : _GEN_11916; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11918 = 10'h233 == _T_174[9:0] ? 4'h8 : _GEN_11917; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11919 = 10'h234 == _T_174[9:0] ? 4'h8 : _GEN_11918; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11920 = 10'h235 == _T_174[9:0] ? 4'h8 : _GEN_11919; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11921 = 10'h236 == _T_174[9:0] ? 4'h8 : _GEN_11920; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11922 = 10'h237 == _T_174[9:0] ? 4'h8 : _GEN_11921; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11923 = 10'h238 == _T_174[9:0] ? 4'h8 : _GEN_11922; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11924 = 10'h239 == _T_174[9:0] ? 4'h6 : _GEN_11923; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11925 = 10'h23a == _T_174[9:0] ? 4'h6 : _GEN_11924; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11926 = 10'h23b == _T_174[9:0] ? 4'h7 : _GEN_11925; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11927 = 10'h23c == _T_174[9:0] ? 4'h6 : _GEN_11926; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11928 = 10'h23d == _T_174[9:0] ? 4'h7 : _GEN_11927; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11929 = 10'h23e == _T_174[9:0] ? 4'h7 : _GEN_11928; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11930 = 10'h23f == _T_174[9:0] ? 4'h6 : _GEN_11929; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11931 = 10'h240 == _T_174[9:0] ? 4'h6 : _GEN_11930; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11932 = 10'h241 == _T_174[9:0] ? 4'h8 : _GEN_11931; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11933 = 10'h242 == _T_174[9:0] ? 4'ha : _GEN_11932; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11934 = 10'h243 == _T_174[9:0] ? 4'ha : _GEN_11933; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11935 = 10'h244 == _T_174[9:0] ? 4'ha : _GEN_11934; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11936 = 10'h245 == _T_174[9:0] ? 4'h8 : _GEN_11935; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11937 = 10'h246 == _T_174[9:0] ? 4'h8 : _GEN_11936; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11938 = 10'h247 == _T_174[9:0] ? 4'h9 : _GEN_11937; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11939 = 10'h248 == _T_174[9:0] ? 4'ha : _GEN_11938; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11940 = 10'h249 == _T_174[9:0] ? 4'ha : _GEN_11939; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11941 = 10'h24a == _T_174[9:0] ? 4'ha : _GEN_11940; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11942 = 10'h24b == _T_174[9:0] ? 4'h4 : _GEN_11941; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11943 = 10'h24c == _T_174[9:0] ? 4'h3 : _GEN_11942; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11944 = 10'h24d == _T_174[9:0] ? 4'h4 : _GEN_11943; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11945 = 10'h24e == _T_174[9:0] ? 4'h5 : _GEN_11944; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11946 = 10'h24f == _T_174[9:0] ? 4'h5 : _GEN_11945; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11947 = 10'h250 == _T_174[9:0] ? 4'h5 : _GEN_11946; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11948 = 10'h251 == _T_174[9:0] ? 4'h5 : _GEN_11947; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11949 = 10'h252 == _T_174[9:0] ? 4'h5 : _GEN_11948; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11950 = 10'h253 == _T_174[9:0] ? 4'h5 : _GEN_11949; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11951 = 10'h254 == _T_174[9:0] ? 4'h5 : _GEN_11950; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11952 = 10'h255 == _T_174[9:0] ? 4'h6 : _GEN_11951; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11953 = 10'h256 == _T_174[9:0] ? 4'h7 : _GEN_11952; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11954 = 10'h257 == _T_174[9:0] ? 4'h3 : _GEN_11953; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11955 = 10'h258 == _T_174[9:0] ? 4'h6 : _GEN_11954; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11956 = 10'h259 == _T_174[9:0] ? 4'h7 : _GEN_11955; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11957 = 10'h25a == _T_174[9:0] ? 4'h7 : _GEN_11956; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11958 = 10'h25b == _T_174[9:0] ? 4'h7 : _GEN_11957; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11959 = 10'h25c == _T_174[9:0] ? 4'h8 : _GEN_11958; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11960 = 10'h25d == _T_174[9:0] ? 4'h8 : _GEN_11959; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11961 = 10'h25e == _T_174[9:0] ? 4'h4 : _GEN_11960; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11962 = 10'h25f == _T_174[9:0] ? 4'h3 : _GEN_11961; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11963 = 10'h260 == _T_174[9:0] ? 4'h7 : _GEN_11962; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11964 = 10'h261 == _T_174[9:0] ? 4'h7 : _GEN_11963; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11965 = 10'h262 == _T_174[9:0] ? 4'h7 : _GEN_11964; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11966 = 10'h263 == _T_174[9:0] ? 4'h6 : _GEN_11965; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11967 = 10'h264 == _T_174[9:0] ? 4'h7 : _GEN_11966; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11968 = 10'h265 == _T_174[9:0] ? 4'h6 : _GEN_11967; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11969 = 10'h266 == _T_174[9:0] ? 4'h5 : _GEN_11968; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11970 = 10'h267 == _T_174[9:0] ? 4'h7 : _GEN_11969; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11971 = 10'h268 == _T_174[9:0] ? 4'ha : _GEN_11970; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11972 = 10'h269 == _T_174[9:0] ? 4'ha : _GEN_11971; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11973 = 10'h26a == _T_174[9:0] ? 4'ha : _GEN_11972; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11974 = 10'h26b == _T_174[9:0] ? 4'ha : _GEN_11973; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11975 = 10'h26c == _T_174[9:0] ? 4'ha : _GEN_11974; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11976 = 10'h26d == _T_174[9:0] ? 4'ha : _GEN_11975; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11977 = 10'h26e == _T_174[9:0] ? 4'ha : _GEN_11976; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11978 = 10'h26f == _T_174[9:0] ? 4'ha : _GEN_11977; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11979 = 10'h270 == _T_174[9:0] ? 4'h5 : _GEN_11978; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11980 = 10'h271 == _T_174[9:0] ? 4'h3 : _GEN_11979; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11981 = 10'h272 == _T_174[9:0] ? 4'h3 : _GEN_11980; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11982 = 10'h273 == _T_174[9:0] ? 4'h4 : _GEN_11981; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11983 = 10'h274 == _T_174[9:0] ? 4'h6 : _GEN_11982; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11984 = 10'h275 == _T_174[9:0] ? 4'h5 : _GEN_11983; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11985 = 10'h276 == _T_174[9:0] ? 4'h6 : _GEN_11984; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11986 = 10'h277 == _T_174[9:0] ? 4'h5 : _GEN_11985; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11987 = 10'h278 == _T_174[9:0] ? 4'h6 : _GEN_11986; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11988 = 10'h279 == _T_174[9:0] ? 4'h6 : _GEN_11987; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11989 = 10'h27a == _T_174[9:0] ? 4'h6 : _GEN_11988; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11990 = 10'h27b == _T_174[9:0] ? 4'h8 : _GEN_11989; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11991 = 10'h27c == _T_174[9:0] ? 4'h6 : _GEN_11990; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11992 = 10'h27d == _T_174[9:0] ? 4'h2 : _GEN_11991; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11993 = 10'h27e == _T_174[9:0] ? 4'h5 : _GEN_11992; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11994 = 10'h27f == _T_174[9:0] ? 4'h7 : _GEN_11993; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11995 = 10'h280 == _T_174[9:0] ? 4'h7 : _GEN_11994; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11996 = 10'h281 == _T_174[9:0] ? 4'h8 : _GEN_11995; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11997 = 10'h282 == _T_174[9:0] ? 4'h7 : _GEN_11996; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11998 = 10'h283 == _T_174[9:0] ? 4'h3 : _GEN_11997; // @[Filter.scala 230:142]
  wire [3:0] _GEN_11999 = 10'h284 == _T_174[9:0] ? 4'h3 : _GEN_11998; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12000 = 10'h285 == _T_174[9:0] ? 4'h3 : _GEN_11999; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12001 = 10'h286 == _T_174[9:0] ? 4'h7 : _GEN_12000; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12002 = 10'h287 == _T_174[9:0] ? 4'h7 : _GEN_12001; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12003 = 10'h288 == _T_174[9:0] ? 4'h7 : _GEN_12002; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12004 = 10'h289 == _T_174[9:0] ? 4'h7 : _GEN_12003; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12005 = 10'h28a == _T_174[9:0] ? 4'h8 : _GEN_12004; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12006 = 10'h28b == _T_174[9:0] ? 4'h8 : _GEN_12005; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12007 = 10'h28c == _T_174[9:0] ? 4'h7 : _GEN_12006; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12008 = 10'h28d == _T_174[9:0] ? 4'h6 : _GEN_12007; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12009 = 10'h28e == _T_174[9:0] ? 4'h3 : _GEN_12008; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12010 = 10'h28f == _T_174[9:0] ? 4'h6 : _GEN_12009; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12011 = 10'h290 == _T_174[9:0] ? 4'h8 : _GEN_12010; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12012 = 10'h291 == _T_174[9:0] ? 4'ha : _GEN_12011; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12013 = 10'h292 == _T_174[9:0] ? 4'ha : _GEN_12012; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12014 = 10'h293 == _T_174[9:0] ? 4'ha : _GEN_12013; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12015 = 10'h294 == _T_174[9:0] ? 4'h9 : _GEN_12014; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12016 = 10'h295 == _T_174[9:0] ? 4'h4 : _GEN_12015; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12017 = 10'h296 == _T_174[9:0] ? 4'h3 : _GEN_12016; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12018 = 10'h297 == _T_174[9:0] ? 4'h3 : _GEN_12017; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12019 = 10'h298 == _T_174[9:0] ? 4'h3 : _GEN_12018; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12020 = 10'h299 == _T_174[9:0] ? 4'h4 : _GEN_12019; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12021 = 10'h29a == _T_174[9:0] ? 4'h5 : _GEN_12020; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12022 = 10'h29b == _T_174[9:0] ? 4'h5 : _GEN_12021; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12023 = 10'h29c == _T_174[9:0] ? 4'h5 : _GEN_12022; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12024 = 10'h29d == _T_174[9:0] ? 4'h5 : _GEN_12023; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12025 = 10'h29e == _T_174[9:0] ? 4'h5 : _GEN_12024; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12026 = 10'h29f == _T_174[9:0] ? 4'h5 : _GEN_12025; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12027 = 10'h2a0 == _T_174[9:0] ? 4'h6 : _GEN_12026; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12028 = 10'h2a1 == _T_174[9:0] ? 4'h7 : _GEN_12027; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12029 = 10'h2a2 == _T_174[9:0] ? 4'h5 : _GEN_12028; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12030 = 10'h2a3 == _T_174[9:0] ? 4'h2 : _GEN_12029; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12031 = 10'h2a4 == _T_174[9:0] ? 4'h3 : _GEN_12030; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12032 = 10'h2a5 == _T_174[9:0] ? 4'h7 : _GEN_12031; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12033 = 10'h2a6 == _T_174[9:0] ? 4'h8 : _GEN_12032; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12034 = 10'h2a7 == _T_174[9:0] ? 4'h7 : _GEN_12033; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12035 = 10'h2a8 == _T_174[9:0] ? 4'h3 : _GEN_12034; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12036 = 10'h2a9 == _T_174[9:0] ? 4'h2 : _GEN_12035; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12037 = 10'h2aa == _T_174[9:0] ? 4'h3 : _GEN_12036; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12038 = 10'h2ab == _T_174[9:0] ? 4'h3 : _GEN_12037; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12039 = 10'h2ac == _T_174[9:0] ? 4'h7 : _GEN_12038; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12040 = 10'h2ad == _T_174[9:0] ? 4'h8 : _GEN_12039; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12041 = 10'h2ae == _T_174[9:0] ? 4'h7 : _GEN_12040; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12042 = 10'h2af == _T_174[9:0] ? 4'h8 : _GEN_12041; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12043 = 10'h2b0 == _T_174[9:0] ? 4'h8 : _GEN_12042; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12044 = 10'h2b1 == _T_174[9:0] ? 4'h8 : _GEN_12043; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12045 = 10'h2b2 == _T_174[9:0] ? 4'h7 : _GEN_12044; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12046 = 10'h2b3 == _T_174[9:0] ? 4'h6 : _GEN_12045; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12047 = 10'h2b4 == _T_174[9:0] ? 4'h2 : _GEN_12046; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12048 = 10'h2b5 == _T_174[9:0] ? 4'h2 : _GEN_12047; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12049 = 10'h2b6 == _T_174[9:0] ? 4'h3 : _GEN_12048; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12050 = 10'h2b7 == _T_174[9:0] ? 4'h3 : _GEN_12049; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12051 = 10'h2b8 == _T_174[9:0] ? 4'h6 : _GEN_12050; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12052 = 10'h2b9 == _T_174[9:0] ? 4'h9 : _GEN_12051; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12053 = 10'h2ba == _T_174[9:0] ? 4'h3 : _GEN_12052; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12054 = 10'h2bb == _T_174[9:0] ? 4'h3 : _GEN_12053; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12055 = 10'h2bc == _T_174[9:0] ? 4'h3 : _GEN_12054; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12056 = 10'h2bd == _T_174[9:0] ? 4'h2 : _GEN_12055; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12057 = 10'h2be == _T_174[9:0] ? 4'h3 : _GEN_12056; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12058 = 10'h2bf == _T_174[9:0] ? 4'h3 : _GEN_12057; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12059 = 10'h2c0 == _T_174[9:0] ? 4'h5 : _GEN_12058; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12060 = 10'h2c1 == _T_174[9:0] ? 4'h5 : _GEN_12059; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12061 = 10'h2c2 == _T_174[9:0] ? 4'h5 : _GEN_12060; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12062 = 10'h2c3 == _T_174[9:0] ? 4'h5 : _GEN_12061; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12063 = 10'h2c4 == _T_174[9:0] ? 4'h5 : _GEN_12062; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12064 = 10'h2c5 == _T_174[9:0] ? 4'h5 : _GEN_12063; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12065 = 10'h2c6 == _T_174[9:0] ? 4'h6 : _GEN_12064; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12066 = 10'h2c7 == _T_174[9:0] ? 4'h7 : _GEN_12065; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12067 = 10'h2c8 == _T_174[9:0] ? 4'h5 : _GEN_12066; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12068 = 10'h2c9 == _T_174[9:0] ? 4'h2 : _GEN_12067; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12069 = 10'h2ca == _T_174[9:0] ? 4'h2 : _GEN_12068; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12070 = 10'h2cb == _T_174[9:0] ? 4'h3 : _GEN_12069; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12071 = 10'h2cc == _T_174[9:0] ? 4'h3 : _GEN_12070; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12072 = 10'h2cd == _T_174[9:0] ? 4'h2 : _GEN_12071; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12073 = 10'h2ce == _T_174[9:0] ? 4'h2 : _GEN_12072; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12074 = 10'h2cf == _T_174[9:0] ? 4'h2 : _GEN_12073; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12075 = 10'h2d0 == _T_174[9:0] ? 4'h2 : _GEN_12074; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12076 = 10'h2d1 == _T_174[9:0] ? 4'h2 : _GEN_12075; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12077 = 10'h2d2 == _T_174[9:0] ? 4'h7 : _GEN_12076; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12078 = 10'h2d3 == _T_174[9:0] ? 4'h7 : _GEN_12077; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12079 = 10'h2d4 == _T_174[9:0] ? 4'h8 : _GEN_12078; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12080 = 10'h2d5 == _T_174[9:0] ? 4'h8 : _GEN_12079; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12081 = 10'h2d6 == _T_174[9:0] ? 4'h8 : _GEN_12080; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12082 = 10'h2d7 == _T_174[9:0] ? 4'h8 : _GEN_12081; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12083 = 10'h2d8 == _T_174[9:0] ? 4'h7 : _GEN_12082; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12084 = 10'h2d9 == _T_174[9:0] ? 4'h6 : _GEN_12083; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12085 = 10'h2da == _T_174[9:0] ? 4'h4 : _GEN_12084; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12086 = 10'h2db == _T_174[9:0] ? 4'h2 : _GEN_12085; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12087 = 10'h2dc == _T_174[9:0] ? 4'h2 : _GEN_12086; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12088 = 10'h2dd == _T_174[9:0] ? 4'h3 : _GEN_12087; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12089 = 10'h2de == _T_174[9:0] ? 4'h3 : _GEN_12088; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12090 = 10'h2df == _T_174[9:0] ? 4'h3 : _GEN_12089; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12091 = 10'h2e0 == _T_174[9:0] ? 4'h3 : _GEN_12090; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12092 = 10'h2e1 == _T_174[9:0] ? 4'h3 : _GEN_12091; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12093 = 10'h2e2 == _T_174[9:0] ? 4'h3 : _GEN_12092; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12094 = 10'h2e3 == _T_174[9:0] ? 4'h2 : _GEN_12093; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12095 = 10'h2e4 == _T_174[9:0] ? 4'h3 : _GEN_12094; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12096 = 10'h2e5 == _T_174[9:0] ? 4'h2 : _GEN_12095; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12097 = 10'h2e6 == _T_174[9:0] ? 4'h5 : _GEN_12096; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12098 = 10'h2e7 == _T_174[9:0] ? 4'h5 : _GEN_12097; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12099 = 10'h2e8 == _T_174[9:0] ? 4'h5 : _GEN_12098; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12100 = 10'h2e9 == _T_174[9:0] ? 4'h5 : _GEN_12099; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12101 = 10'h2ea == _T_174[9:0] ? 4'h5 : _GEN_12100; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12102 = 10'h2eb == _T_174[9:0] ? 4'h5 : _GEN_12101; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12103 = 10'h2ec == _T_174[9:0] ? 4'h6 : _GEN_12102; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12104 = 10'h2ed == _T_174[9:0] ? 4'h7 : _GEN_12103; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12105 = 10'h2ee == _T_174[9:0] ? 4'h6 : _GEN_12104; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12106 = 10'h2ef == _T_174[9:0] ? 4'h2 : _GEN_12105; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12107 = 10'h2f0 == _T_174[9:0] ? 4'h2 : _GEN_12106; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12108 = 10'h2f1 == _T_174[9:0] ? 4'h2 : _GEN_12107; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12109 = 10'h2f2 == _T_174[9:0] ? 4'h2 : _GEN_12108; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12110 = 10'h2f3 == _T_174[9:0] ? 4'h2 : _GEN_12109; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12111 = 10'h2f4 == _T_174[9:0] ? 4'h2 : _GEN_12110; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12112 = 10'h2f5 == _T_174[9:0] ? 4'h2 : _GEN_12111; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12113 = 10'h2f6 == _T_174[9:0] ? 4'h2 : _GEN_12112; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12114 = 10'h2f7 == _T_174[9:0] ? 4'h2 : _GEN_12113; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12115 = 10'h2f8 == _T_174[9:0] ? 4'h7 : _GEN_12114; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12116 = 10'h2f9 == _T_174[9:0] ? 4'h7 : _GEN_12115; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12117 = 10'h2fa == _T_174[9:0] ? 4'h8 : _GEN_12116; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12118 = 10'h2fb == _T_174[9:0] ? 4'h8 : _GEN_12117; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12119 = 10'h2fc == _T_174[9:0] ? 4'h7 : _GEN_12118; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12120 = 10'h2fd == _T_174[9:0] ? 4'h7 : _GEN_12119; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12121 = 10'h2fe == _T_174[9:0] ? 4'h7 : _GEN_12120; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12122 = 10'h2ff == _T_174[9:0] ? 4'h7 : _GEN_12121; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12123 = 10'h300 == _T_174[9:0] ? 4'h8 : _GEN_12122; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12124 = 10'h301 == _T_174[9:0] ? 4'h7 : _GEN_12123; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12125 = 10'h302 == _T_174[9:0] ? 4'h3 : _GEN_12124; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12126 = 10'h303 == _T_174[9:0] ? 4'h3 : _GEN_12125; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12127 = 10'h304 == _T_174[9:0] ? 4'h2 : _GEN_12126; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12128 = 10'h305 == _T_174[9:0] ? 4'h2 : _GEN_12127; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12129 = 10'h306 == _T_174[9:0] ? 4'h2 : _GEN_12128; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12130 = 10'h307 == _T_174[9:0] ? 4'h2 : _GEN_12129; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12131 = 10'h308 == _T_174[9:0] ? 4'h2 : _GEN_12130; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12132 = 10'h309 == _T_174[9:0] ? 4'h2 : _GEN_12131; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12133 = 10'h30a == _T_174[9:0] ? 4'h2 : _GEN_12132; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12134 = 10'h30b == _T_174[9:0] ? 4'h3 : _GEN_12133; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12135 = 10'h30c == _T_174[9:0] ? 4'h4 : _GEN_12134; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12136 = 10'h30d == _T_174[9:0] ? 4'h5 : _GEN_12135; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12137 = 10'h30e == _T_174[9:0] ? 4'h5 : _GEN_12136; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12138 = 10'h30f == _T_174[9:0] ? 4'h5 : _GEN_12137; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12139 = 10'h310 == _T_174[9:0] ? 4'h5 : _GEN_12138; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12140 = 10'h311 == _T_174[9:0] ? 4'h5 : _GEN_12139; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12141 = 10'h312 == _T_174[9:0] ? 4'h6 : _GEN_12140; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12142 = 10'h313 == _T_174[9:0] ? 4'h7 : _GEN_12141; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12143 = 10'h314 == _T_174[9:0] ? 4'h7 : _GEN_12142; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12144 = 10'h315 == _T_174[9:0] ? 4'h3 : _GEN_12143; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12145 = 10'h316 == _T_174[9:0] ? 4'h2 : _GEN_12144; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12146 = 10'h317 == _T_174[9:0] ? 4'h2 : _GEN_12145; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12147 = 10'h318 == _T_174[9:0] ? 4'h2 : _GEN_12146; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12148 = 10'h319 == _T_174[9:0] ? 4'h2 : _GEN_12147; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12149 = 10'h31a == _T_174[9:0] ? 4'h2 : _GEN_12148; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12150 = 10'h31b == _T_174[9:0] ? 4'h2 : _GEN_12149; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12151 = 10'h31c == _T_174[9:0] ? 4'h2 : _GEN_12150; // @[Filter.scala 230:142]
  wire [3:0] _GEN_12152 = 10'h31d == _T_174[9:0] ? 4'h2 : _GEN_12151; // @[Filter.scala 230:142]
  wire [7:0] _T_188 = _GEN_12152 * 4'ha; // @[Filter.scala 230:142]
  wire [10:0] _GEN_38983 = {{3'd0}, _T_188}; // @[Filter.scala 230:109]
  wire [10:0] _T_190 = _T_183 + _GEN_38983; // @[Filter.scala 230:109]
  wire [10:0] _T_191 = _T_190 / 11'h64; // @[Filter.scala 230:150]
  wire  _T_193 = _T_164 >= 6'h20; // @[Filter.scala 233:31]
  wire  _T_197 = _T_171 >= 32'h12; // @[Filter.scala 233:63]
  wire  _T_198 = _T_193 | _T_197; // @[Filter.scala 233:58]
  wire [10:0] _GEN_12951 = io_SPI_distort ? _T_191 : {{7'd0}, _GEN_10556}; // @[Filter.scala 235:35]
  wire [10:0] _GEN_12952 = _T_198 ? 11'h0 : _GEN_12951; // @[Filter.scala 233:80]
  wire [10:0] _GEN_13751 = io_SPI_distort ? _T_191 : {{7'd0}, _GEN_11354}; // @[Filter.scala 235:35]
  wire [10:0] _GEN_13752 = _T_198 ? 11'h0 : _GEN_13751; // @[Filter.scala 233:80]
  wire [10:0] _GEN_14551 = io_SPI_distort ? _T_191 : {{7'd0}, _GEN_12152}; // @[Filter.scala 235:35]
  wire [10:0] _GEN_14552 = _T_198 ? 11'h0 : _GEN_14551; // @[Filter.scala 233:80]
  wire [31:0] _T_226 = pixelIndex + 32'h3; // @[Filter.scala 228:31]
  wire [31:0] _GEN_3 = _T_226 % 32'h20; // @[Filter.scala 228:38]
  wire [5:0] _T_227 = _GEN_3[5:0]; // @[Filter.scala 228:38]
  wire [5:0] _T_229 = _T_227 + _GEN_38951; // @[Filter.scala 228:53]
  wire [5:0] _T_231 = _T_229 - 6'h1; // @[Filter.scala 228:69]
  wire [31:0] _T_234 = _T_226 / 32'h20; // @[Filter.scala 229:38]
  wire [31:0] _T_236 = _T_234 + _GEN_38952; // @[Filter.scala 229:53]
  wire [31:0] _T_238 = _T_236 - 32'h1; // @[Filter.scala 229:69]
  wire [37:0] _T_239 = _T_238 * 32'h20; // @[Filter.scala 230:42]
  wire [37:0] _GEN_38989 = {{32'd0}, _T_231}; // @[Filter.scala 230:57]
  wire [37:0] _T_241 = _T_239 + _GEN_38989; // @[Filter.scala 230:57]
  wire [3:0] _GEN_14575 = 10'h16 == _T_241[9:0] ? 4'h9 : 4'ha; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14576 = 10'h17 == _T_241[9:0] ? 4'h3 : _GEN_14575; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14577 = 10'h18 == _T_241[9:0] ? 4'h6 : _GEN_14576; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14578 = 10'h19 == _T_241[9:0] ? 4'ha : _GEN_14577; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14579 = 10'h1a == _T_241[9:0] ? 4'ha : _GEN_14578; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14580 = 10'h1b == _T_241[9:0] ? 4'ha : _GEN_14579; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14581 = 10'h1c == _T_241[9:0] ? 4'ha : _GEN_14580; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14582 = 10'h1d == _T_241[9:0] ? 4'ha : _GEN_14581; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14583 = 10'h1e == _T_241[9:0] ? 4'ha : _GEN_14582; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14584 = 10'h1f == _T_241[9:0] ? 4'ha : _GEN_14583; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14585 = 10'h20 == _T_241[9:0] ? 4'ha : _GEN_14584; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14586 = 10'h21 == _T_241[9:0] ? 4'ha : _GEN_14585; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14587 = 10'h22 == _T_241[9:0] ? 4'ha : _GEN_14586; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14588 = 10'h23 == _T_241[9:0] ? 4'ha : _GEN_14587; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14589 = 10'h24 == _T_241[9:0] ? 4'ha : _GEN_14588; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14590 = 10'h25 == _T_241[9:0] ? 4'ha : _GEN_14589; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14591 = 10'h26 == _T_241[9:0] ? 4'ha : _GEN_14590; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14592 = 10'h27 == _T_241[9:0] ? 4'ha : _GEN_14591; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14593 = 10'h28 == _T_241[9:0] ? 4'ha : _GEN_14592; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14594 = 10'h29 == _T_241[9:0] ? 4'ha : _GEN_14593; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14595 = 10'h2a == _T_241[9:0] ? 4'ha : _GEN_14594; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14596 = 10'h2b == _T_241[9:0] ? 4'ha : _GEN_14595; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14597 = 10'h2c == _T_241[9:0] ? 4'ha : _GEN_14596; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14598 = 10'h2d == _T_241[9:0] ? 4'ha : _GEN_14597; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14599 = 10'h2e == _T_241[9:0] ? 4'ha : _GEN_14598; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14600 = 10'h2f == _T_241[9:0] ? 4'ha : _GEN_14599; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14601 = 10'h30 == _T_241[9:0] ? 4'ha : _GEN_14600; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14602 = 10'h31 == _T_241[9:0] ? 4'ha : _GEN_14601; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14603 = 10'h32 == _T_241[9:0] ? 4'ha : _GEN_14602; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14604 = 10'h33 == _T_241[9:0] ? 4'ha : _GEN_14603; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14605 = 10'h34 == _T_241[9:0] ? 4'ha : _GEN_14604; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14606 = 10'h35 == _T_241[9:0] ? 4'ha : _GEN_14605; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14607 = 10'h36 == _T_241[9:0] ? 4'ha : _GEN_14606; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14608 = 10'h37 == _T_241[9:0] ? 4'ha : _GEN_14607; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14609 = 10'h38 == _T_241[9:0] ? 4'ha : _GEN_14608; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14610 = 10'h39 == _T_241[9:0] ? 4'ha : _GEN_14609; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14611 = 10'h3a == _T_241[9:0] ? 4'ha : _GEN_14610; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14612 = 10'h3b == _T_241[9:0] ? 4'h9 : _GEN_14611; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14613 = 10'h3c == _T_241[9:0] ? 4'h4 : _GEN_14612; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14614 = 10'h3d == _T_241[9:0] ? 4'h3 : _GEN_14613; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14615 = 10'h3e == _T_241[9:0] ? 4'h4 : _GEN_14614; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14616 = 10'h3f == _T_241[9:0] ? 4'ha : _GEN_14615; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14617 = 10'h40 == _T_241[9:0] ? 4'ha : _GEN_14616; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14618 = 10'h41 == _T_241[9:0] ? 4'ha : _GEN_14617; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14619 = 10'h42 == _T_241[9:0] ? 4'ha : _GEN_14618; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14620 = 10'h43 == _T_241[9:0] ? 4'ha : _GEN_14619; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14621 = 10'h44 == _T_241[9:0] ? 4'ha : _GEN_14620; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14622 = 10'h45 == _T_241[9:0] ? 4'ha : _GEN_14621; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14623 = 10'h46 == _T_241[9:0] ? 4'ha : _GEN_14622; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14624 = 10'h47 == _T_241[9:0] ? 4'ha : _GEN_14623; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14625 = 10'h48 == _T_241[9:0] ? 4'ha : _GEN_14624; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14626 = 10'h49 == _T_241[9:0] ? 4'ha : _GEN_14625; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14627 = 10'h4a == _T_241[9:0] ? 4'ha : _GEN_14626; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14628 = 10'h4b == _T_241[9:0] ? 4'ha : _GEN_14627; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14629 = 10'h4c == _T_241[9:0] ? 4'ha : _GEN_14628; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14630 = 10'h4d == _T_241[9:0] ? 4'ha : _GEN_14629; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14631 = 10'h4e == _T_241[9:0] ? 4'ha : _GEN_14630; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14632 = 10'h4f == _T_241[9:0] ? 4'ha : _GEN_14631; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14633 = 10'h50 == _T_241[9:0] ? 4'ha : _GEN_14632; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14634 = 10'h51 == _T_241[9:0] ? 4'ha : _GEN_14633; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14635 = 10'h52 == _T_241[9:0] ? 4'ha : _GEN_14634; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14636 = 10'h53 == _T_241[9:0] ? 4'ha : _GEN_14635; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14637 = 10'h54 == _T_241[9:0] ? 4'ha : _GEN_14636; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14638 = 10'h55 == _T_241[9:0] ? 4'ha : _GEN_14637; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14639 = 10'h56 == _T_241[9:0] ? 4'ha : _GEN_14638; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14640 = 10'h57 == _T_241[9:0] ? 4'ha : _GEN_14639; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14641 = 10'h58 == _T_241[9:0] ? 4'ha : _GEN_14640; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14642 = 10'h59 == _T_241[9:0] ? 4'ha : _GEN_14641; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14643 = 10'h5a == _T_241[9:0] ? 4'h7 : _GEN_14642; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14644 = 10'h5b == _T_241[9:0] ? 4'h7 : _GEN_14643; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14645 = 10'h5c == _T_241[9:0] ? 4'ha : _GEN_14644; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14646 = 10'h5d == _T_241[9:0] ? 4'ha : _GEN_14645; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14647 = 10'h5e == _T_241[9:0] ? 4'ha : _GEN_14646; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14648 = 10'h5f == _T_241[9:0] ? 4'ha : _GEN_14647; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14649 = 10'h60 == _T_241[9:0] ? 4'ha : _GEN_14648; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14650 = 10'h61 == _T_241[9:0] ? 4'h8 : _GEN_14649; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14651 = 10'h62 == _T_241[9:0] ? 4'h3 : _GEN_14650; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14652 = 10'h63 == _T_241[9:0] ? 4'h3 : _GEN_14651; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14653 = 10'h64 == _T_241[9:0] ? 4'h3 : _GEN_14652; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14654 = 10'h65 == _T_241[9:0] ? 4'h9 : _GEN_14653; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14655 = 10'h66 == _T_241[9:0] ? 4'ha : _GEN_14654; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14656 = 10'h67 == _T_241[9:0] ? 4'ha : _GEN_14655; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14657 = 10'h68 == _T_241[9:0] ? 4'ha : _GEN_14656; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14658 = 10'h69 == _T_241[9:0] ? 4'ha : _GEN_14657; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14659 = 10'h6a == _T_241[9:0] ? 4'ha : _GEN_14658; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14660 = 10'h6b == _T_241[9:0] ? 4'h8 : _GEN_14659; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14661 = 10'h6c == _T_241[9:0] ? 4'h5 : _GEN_14660; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14662 = 10'h6d == _T_241[9:0] ? 4'h8 : _GEN_14661; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14663 = 10'h6e == _T_241[9:0] ? 4'ha : _GEN_14662; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14664 = 10'h6f == _T_241[9:0] ? 4'ha : _GEN_14663; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14665 = 10'h70 == _T_241[9:0] ? 4'ha : _GEN_14664; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14666 = 10'h71 == _T_241[9:0] ? 4'ha : _GEN_14665; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14667 = 10'h72 == _T_241[9:0] ? 4'ha : _GEN_14666; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14668 = 10'h73 == _T_241[9:0] ? 4'ha : _GEN_14667; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14669 = 10'h74 == _T_241[9:0] ? 4'ha : _GEN_14668; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14670 = 10'h75 == _T_241[9:0] ? 4'ha : _GEN_14669; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14671 = 10'h76 == _T_241[9:0] ? 4'ha : _GEN_14670; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14672 = 10'h77 == _T_241[9:0] ? 4'ha : _GEN_14671; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14673 = 10'h78 == _T_241[9:0] ? 4'ha : _GEN_14672; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14674 = 10'h79 == _T_241[9:0] ? 4'ha : _GEN_14673; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14675 = 10'h7a == _T_241[9:0] ? 4'ha : _GEN_14674; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14676 = 10'h7b == _T_241[9:0] ? 4'ha : _GEN_14675; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14677 = 10'h7c == _T_241[9:0] ? 4'ha : _GEN_14676; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14678 = 10'h7d == _T_241[9:0] ? 4'ha : _GEN_14677; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14679 = 10'h7e == _T_241[9:0] ? 4'ha : _GEN_14678; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14680 = 10'h7f == _T_241[9:0] ? 4'ha : _GEN_14679; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14681 = 10'h80 == _T_241[9:0] ? 4'ha : _GEN_14680; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14682 = 10'h81 == _T_241[9:0] ? 4'h5 : _GEN_14681; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14683 = 10'h82 == _T_241[9:0] ? 4'h5 : _GEN_14682; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14684 = 10'h83 == _T_241[9:0] ? 4'h7 : _GEN_14683; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14685 = 10'h84 == _T_241[9:0] ? 4'ha : _GEN_14684; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14686 = 10'h85 == _T_241[9:0] ? 4'ha : _GEN_14685; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14687 = 10'h86 == _T_241[9:0] ? 4'ha : _GEN_14686; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14688 = 10'h87 == _T_241[9:0] ? 4'h5 : _GEN_14687; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14689 = 10'h88 == _T_241[9:0] ? 4'h3 : _GEN_14688; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14690 = 10'h89 == _T_241[9:0] ? 4'h3 : _GEN_14689; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14691 = 10'h8a == _T_241[9:0] ? 4'h4 : _GEN_14690; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14692 = 10'h8b == _T_241[9:0] ? 4'h9 : _GEN_14691; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14693 = 10'h8c == _T_241[9:0] ? 4'ha : _GEN_14692; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14694 = 10'h8d == _T_241[9:0] ? 4'ha : _GEN_14693; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14695 = 10'h8e == _T_241[9:0] ? 4'ha : _GEN_14694; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14696 = 10'h8f == _T_241[9:0] ? 4'h6 : _GEN_14695; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14697 = 10'h90 == _T_241[9:0] ? 4'h4 : _GEN_14696; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14698 = 10'h91 == _T_241[9:0] ? 4'h3 : _GEN_14697; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14699 = 10'h92 == _T_241[9:0] ? 4'h7 : _GEN_14698; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14700 = 10'h93 == _T_241[9:0] ? 4'ha : _GEN_14699; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14701 = 10'h94 == _T_241[9:0] ? 4'ha : _GEN_14700; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14702 = 10'h95 == _T_241[9:0] ? 4'ha : _GEN_14701; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14703 = 10'h96 == _T_241[9:0] ? 4'ha : _GEN_14702; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14704 = 10'h97 == _T_241[9:0] ? 4'ha : _GEN_14703; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14705 = 10'h98 == _T_241[9:0] ? 4'ha : _GEN_14704; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14706 = 10'h99 == _T_241[9:0] ? 4'ha : _GEN_14705; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14707 = 10'h9a == _T_241[9:0] ? 4'ha : _GEN_14706; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14708 = 10'h9b == _T_241[9:0] ? 4'ha : _GEN_14707; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14709 = 10'h9c == _T_241[9:0] ? 4'ha : _GEN_14708; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14710 = 10'h9d == _T_241[9:0] ? 4'ha : _GEN_14709; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14711 = 10'h9e == _T_241[9:0] ? 4'ha : _GEN_14710; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14712 = 10'h9f == _T_241[9:0] ? 4'ha : _GEN_14711; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14713 = 10'ha0 == _T_241[9:0] ? 4'ha : _GEN_14712; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14714 = 10'ha1 == _T_241[9:0] ? 4'ha : _GEN_14713; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14715 = 10'ha2 == _T_241[9:0] ? 4'ha : _GEN_14714; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14716 = 10'ha3 == _T_241[9:0] ? 4'ha : _GEN_14715; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14717 = 10'ha4 == _T_241[9:0] ? 4'ha : _GEN_14716; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14718 = 10'ha5 == _T_241[9:0] ? 4'ha : _GEN_14717; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14719 = 10'ha6 == _T_241[9:0] ? 4'ha : _GEN_14718; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14720 = 10'ha7 == _T_241[9:0] ? 4'h9 : _GEN_14719; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14721 = 10'ha8 == _T_241[9:0] ? 4'h4 : _GEN_14720; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14722 = 10'ha9 == _T_241[9:0] ? 4'h3 : _GEN_14721; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14723 = 10'haa == _T_241[9:0] ? 4'h4 : _GEN_14722; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14724 = 10'hab == _T_241[9:0] ? 4'h7 : _GEN_14723; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14725 = 10'hac == _T_241[9:0] ? 4'h8 : _GEN_14724; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14726 = 10'had == _T_241[9:0] ? 4'h3 : _GEN_14725; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14727 = 10'hae == _T_241[9:0] ? 4'h3 : _GEN_14726; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14728 = 10'haf == _T_241[9:0] ? 4'h3 : _GEN_14727; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14729 = 10'hb0 == _T_241[9:0] ? 4'h3 : _GEN_14728; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14730 = 10'hb1 == _T_241[9:0] ? 4'h7 : _GEN_14729; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14731 = 10'hb2 == _T_241[9:0] ? 4'h9 : _GEN_14730; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14732 = 10'hb3 == _T_241[9:0] ? 4'h6 : _GEN_14731; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14733 = 10'hb4 == _T_241[9:0] ? 4'h4 : _GEN_14732; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14734 = 10'hb5 == _T_241[9:0] ? 4'h3 : _GEN_14733; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14735 = 10'hb6 == _T_241[9:0] ? 4'h3 : _GEN_14734; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14736 = 10'hb7 == _T_241[9:0] ? 4'h6 : _GEN_14735; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14737 = 10'hb8 == _T_241[9:0] ? 4'ha : _GEN_14736; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14738 = 10'hb9 == _T_241[9:0] ? 4'ha : _GEN_14737; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14739 = 10'hba == _T_241[9:0] ? 4'ha : _GEN_14738; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14740 = 10'hbb == _T_241[9:0] ? 4'ha : _GEN_14739; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14741 = 10'hbc == _T_241[9:0] ? 4'ha : _GEN_14740; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14742 = 10'hbd == _T_241[9:0] ? 4'h9 : _GEN_14741; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14743 = 10'hbe == _T_241[9:0] ? 4'ha : _GEN_14742; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14744 = 10'hbf == _T_241[9:0] ? 4'ha : _GEN_14743; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14745 = 10'hc0 == _T_241[9:0] ? 4'ha : _GEN_14744; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14746 = 10'hc1 == _T_241[9:0] ? 4'ha : _GEN_14745; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14747 = 10'hc2 == _T_241[9:0] ? 4'ha : _GEN_14746; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14748 = 10'hc3 == _T_241[9:0] ? 4'ha : _GEN_14747; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14749 = 10'hc4 == _T_241[9:0] ? 4'ha : _GEN_14748; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14750 = 10'hc5 == _T_241[9:0] ? 4'ha : _GEN_14749; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14751 = 10'hc6 == _T_241[9:0] ? 4'ha : _GEN_14750; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14752 = 10'hc7 == _T_241[9:0] ? 4'h9 : _GEN_14751; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14753 = 10'hc8 == _T_241[9:0] ? 4'h8 : _GEN_14752; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14754 = 10'hc9 == _T_241[9:0] ? 4'h8 : _GEN_14753; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14755 = 10'hca == _T_241[9:0] ? 4'h9 : _GEN_14754; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14756 = 10'hcb == _T_241[9:0] ? 4'ha : _GEN_14755; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14757 = 10'hcc == _T_241[9:0] ? 4'ha : _GEN_14756; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14758 = 10'hcd == _T_241[9:0] ? 4'ha : _GEN_14757; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14759 = 10'hce == _T_241[9:0] ? 4'h8 : _GEN_14758; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14760 = 10'hcf == _T_241[9:0] ? 4'h3 : _GEN_14759; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14761 = 10'hd0 == _T_241[9:0] ? 4'h3 : _GEN_14760; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14762 = 10'hd1 == _T_241[9:0] ? 4'h3 : _GEN_14761; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14763 = 10'hd2 == _T_241[9:0] ? 4'h4 : _GEN_14762; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14764 = 10'hd3 == _T_241[9:0] ? 4'h3 : _GEN_14763; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14765 = 10'hd4 == _T_241[9:0] ? 4'h3 : _GEN_14764; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14766 = 10'hd5 == _T_241[9:0] ? 4'h3 : _GEN_14765; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14767 = 10'hd6 == _T_241[9:0] ? 4'h3 : _GEN_14766; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14768 = 10'hd7 == _T_241[9:0] ? 4'h5 : _GEN_14767; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14769 = 10'hd8 == _T_241[9:0] ? 4'h4 : _GEN_14768; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14770 = 10'hd9 == _T_241[9:0] ? 4'h3 : _GEN_14769; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14771 = 10'hda == _T_241[9:0] ? 4'h3 : _GEN_14770; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14772 = 10'hdb == _T_241[9:0] ? 4'h3 : _GEN_14771; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14773 = 10'hdc == _T_241[9:0] ? 4'h4 : _GEN_14772; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14774 = 10'hdd == _T_241[9:0] ? 4'ha : _GEN_14773; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14775 = 10'hde == _T_241[9:0] ? 4'ha : _GEN_14774; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14776 = 10'hdf == _T_241[9:0] ? 4'ha : _GEN_14775; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14777 = 10'he0 == _T_241[9:0] ? 4'ha : _GEN_14776; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14778 = 10'he1 == _T_241[9:0] ? 4'ha : _GEN_14777; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14779 = 10'he2 == _T_241[9:0] ? 4'ha : _GEN_14778; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14780 = 10'he3 == _T_241[9:0] ? 4'h5 : _GEN_14779; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14781 = 10'he4 == _T_241[9:0] ? 4'ha : _GEN_14780; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14782 = 10'he5 == _T_241[9:0] ? 4'ha : _GEN_14781; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14783 = 10'he6 == _T_241[9:0] ? 4'ha : _GEN_14782; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14784 = 10'he7 == _T_241[9:0] ? 4'ha : _GEN_14783; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14785 = 10'he8 == _T_241[9:0] ? 4'ha : _GEN_14784; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14786 = 10'he9 == _T_241[9:0] ? 4'ha : _GEN_14785; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14787 = 10'hea == _T_241[9:0] ? 4'ha : _GEN_14786; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14788 = 10'heb == _T_241[9:0] ? 4'h9 : _GEN_14787; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14789 = 10'hec == _T_241[9:0] ? 4'h7 : _GEN_14788; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14790 = 10'hed == _T_241[9:0] ? 4'h3 : _GEN_14789; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14791 = 10'hee == _T_241[9:0] ? 4'h3 : _GEN_14790; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14792 = 10'hef == _T_241[9:0] ? 4'h3 : _GEN_14791; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14793 = 10'hf0 == _T_241[9:0] ? 4'h4 : _GEN_14792; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14794 = 10'hf1 == _T_241[9:0] ? 4'h7 : _GEN_14793; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14795 = 10'hf2 == _T_241[9:0] ? 4'ha : _GEN_14794; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14796 = 10'hf3 == _T_241[9:0] ? 4'ha : _GEN_14795; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14797 = 10'hf4 == _T_241[9:0] ? 4'ha : _GEN_14796; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14798 = 10'hf5 == _T_241[9:0] ? 4'h7 : _GEN_14797; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14799 = 10'hf6 == _T_241[9:0] ? 4'h3 : _GEN_14798; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14800 = 10'hf7 == _T_241[9:0] ? 4'h3 : _GEN_14799; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14801 = 10'hf8 == _T_241[9:0] ? 4'h3 : _GEN_14800; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14802 = 10'hf9 == _T_241[9:0] ? 4'h3 : _GEN_14801; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14803 = 10'hfa == _T_241[9:0] ? 4'h3 : _GEN_14802; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14804 = 10'hfb == _T_241[9:0] ? 4'h3 : _GEN_14803; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14805 = 10'hfc == _T_241[9:0] ? 4'h3 : _GEN_14804; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14806 = 10'hfd == _T_241[9:0] ? 4'h3 : _GEN_14805; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14807 = 10'hfe == _T_241[9:0] ? 4'h3 : _GEN_14806; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14808 = 10'hff == _T_241[9:0] ? 4'h3 : _GEN_14807; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14809 = 10'h100 == _T_241[9:0] ? 4'h3 : _GEN_14808; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14810 = 10'h101 == _T_241[9:0] ? 4'h4 : _GEN_14809; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14811 = 10'h102 == _T_241[9:0] ? 4'h6 : _GEN_14810; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14812 = 10'h103 == _T_241[9:0] ? 4'ha : _GEN_14811; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14813 = 10'h104 == _T_241[9:0] ? 4'ha : _GEN_14812; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14814 = 10'h105 == _T_241[9:0] ? 4'h9 : _GEN_14813; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14815 = 10'h106 == _T_241[9:0] ? 4'h9 : _GEN_14814; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14816 = 10'h107 == _T_241[9:0] ? 4'h9 : _GEN_14815; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14817 = 10'h108 == _T_241[9:0] ? 4'h9 : _GEN_14816; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14818 = 10'h109 == _T_241[9:0] ? 4'h3 : _GEN_14817; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14819 = 10'h10a == _T_241[9:0] ? 4'ha : _GEN_14818; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14820 = 10'h10b == _T_241[9:0] ? 4'ha : _GEN_14819; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14821 = 10'h10c == _T_241[9:0] ? 4'ha : _GEN_14820; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14822 = 10'h10d == _T_241[9:0] ? 4'ha : _GEN_14821; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14823 = 10'h10e == _T_241[9:0] ? 4'ha : _GEN_14822; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14824 = 10'h10f == _T_241[9:0] ? 4'h9 : _GEN_14823; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14825 = 10'h110 == _T_241[9:0] ? 4'h9 : _GEN_14824; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14826 = 10'h111 == _T_241[9:0] ? 4'h4 : _GEN_14825; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14827 = 10'h112 == _T_241[9:0] ? 4'h8 : _GEN_14826; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14828 = 10'h113 == _T_241[9:0] ? 4'h3 : _GEN_14827; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14829 = 10'h114 == _T_241[9:0] ? 4'h3 : _GEN_14828; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14830 = 10'h115 == _T_241[9:0] ? 4'h4 : _GEN_14829; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14831 = 10'h116 == _T_241[9:0] ? 4'h4 : _GEN_14830; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14832 = 10'h117 == _T_241[9:0] ? 4'h3 : _GEN_14831; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14833 = 10'h118 == _T_241[9:0] ? 4'h8 : _GEN_14832; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14834 = 10'h119 == _T_241[9:0] ? 4'ha : _GEN_14833; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14835 = 10'h11a == _T_241[9:0] ? 4'ha : _GEN_14834; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14836 = 10'h11b == _T_241[9:0] ? 4'ha : _GEN_14835; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14837 = 10'h11c == _T_241[9:0] ? 4'h6 : _GEN_14836; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14838 = 10'h11d == _T_241[9:0] ? 4'h3 : _GEN_14837; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14839 = 10'h11e == _T_241[9:0] ? 4'h3 : _GEN_14838; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14840 = 10'h11f == _T_241[9:0] ? 4'h3 : _GEN_14839; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14841 = 10'h120 == _T_241[9:0] ? 4'h3 : _GEN_14840; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14842 = 10'h121 == _T_241[9:0] ? 4'h3 : _GEN_14841; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14843 = 10'h122 == _T_241[9:0] ? 4'h3 : _GEN_14842; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14844 = 10'h123 == _T_241[9:0] ? 4'h3 : _GEN_14843; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14845 = 10'h124 == _T_241[9:0] ? 4'h3 : _GEN_14844; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14846 = 10'h125 == _T_241[9:0] ? 4'h3 : _GEN_14845; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14847 = 10'h126 == _T_241[9:0] ? 4'h4 : _GEN_14846; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14848 = 10'h127 == _T_241[9:0] ? 4'h6 : _GEN_14847; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14849 = 10'h128 == _T_241[9:0] ? 4'h5 : _GEN_14848; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14850 = 10'h129 == _T_241[9:0] ? 4'h8 : _GEN_14849; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14851 = 10'h12a == _T_241[9:0] ? 4'h5 : _GEN_14850; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14852 = 10'h12b == _T_241[9:0] ? 4'h3 : _GEN_14851; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14853 = 10'h12c == _T_241[9:0] ? 4'h3 : _GEN_14852; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14854 = 10'h12d == _T_241[9:0] ? 4'h3 : _GEN_14853; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14855 = 10'h12e == _T_241[9:0] ? 4'h4 : _GEN_14854; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14856 = 10'h12f == _T_241[9:0] ? 4'h4 : _GEN_14855; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14857 = 10'h130 == _T_241[9:0] ? 4'ha : _GEN_14856; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14858 = 10'h131 == _T_241[9:0] ? 4'h9 : _GEN_14857; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14859 = 10'h132 == _T_241[9:0] ? 4'h9 : _GEN_14858; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14860 = 10'h133 == _T_241[9:0] ? 4'h8 : _GEN_14859; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14861 = 10'h134 == _T_241[9:0] ? 4'h9 : _GEN_14860; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14862 = 10'h135 == _T_241[9:0] ? 4'h8 : _GEN_14861; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14863 = 10'h136 == _T_241[9:0] ? 4'h7 : _GEN_14862; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14864 = 10'h137 == _T_241[9:0] ? 4'h6 : _GEN_14863; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14865 = 10'h138 == _T_241[9:0] ? 4'h8 : _GEN_14864; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14866 = 10'h139 == _T_241[9:0] ? 4'h3 : _GEN_14865; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14867 = 10'h13a == _T_241[9:0] ? 4'h3 : _GEN_14866; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14868 = 10'h13b == _T_241[9:0] ? 4'h4 : _GEN_14867; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14869 = 10'h13c == _T_241[9:0] ? 4'h4 : _GEN_14868; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14870 = 10'h13d == _T_241[9:0] ? 4'h3 : _GEN_14869; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14871 = 10'h13e == _T_241[9:0] ? 4'h5 : _GEN_14870; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14872 = 10'h13f == _T_241[9:0] ? 4'h9 : _GEN_14871; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14873 = 10'h140 == _T_241[9:0] ? 4'ha : _GEN_14872; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14874 = 10'h141 == _T_241[9:0] ? 4'ha : _GEN_14873; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14875 = 10'h142 == _T_241[9:0] ? 4'ha : _GEN_14874; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14876 = 10'h143 == _T_241[9:0] ? 4'h5 : _GEN_14875; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14877 = 10'h144 == _T_241[9:0] ? 4'h3 : _GEN_14876; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14878 = 10'h145 == _T_241[9:0] ? 4'h3 : _GEN_14877; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14879 = 10'h146 == _T_241[9:0] ? 4'h3 : _GEN_14878; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14880 = 10'h147 == _T_241[9:0] ? 4'h4 : _GEN_14879; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14881 = 10'h148 == _T_241[9:0] ? 4'h3 : _GEN_14880; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14882 = 10'h149 == _T_241[9:0] ? 4'h3 : _GEN_14881; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14883 = 10'h14a == _T_241[9:0] ? 4'h3 : _GEN_14882; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14884 = 10'h14b == _T_241[9:0] ? 4'h6 : _GEN_14883; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14885 = 10'h14c == _T_241[9:0] ? 4'h8 : _GEN_14884; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14886 = 10'h14d == _T_241[9:0] ? 4'h5 : _GEN_14885; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14887 = 10'h14e == _T_241[9:0] ? 4'h4 : _GEN_14886; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14888 = 10'h14f == _T_241[9:0] ? 4'h3 : _GEN_14887; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14889 = 10'h150 == _T_241[9:0] ? 4'h3 : _GEN_14888; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14890 = 10'h151 == _T_241[9:0] ? 4'h3 : _GEN_14889; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14891 = 10'h152 == _T_241[9:0] ? 4'h3 : _GEN_14890; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14892 = 10'h153 == _T_241[9:0] ? 4'h3 : _GEN_14891; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14893 = 10'h154 == _T_241[9:0] ? 4'h3 : _GEN_14892; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14894 = 10'h155 == _T_241[9:0] ? 4'h4 : _GEN_14893; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14895 = 10'h156 == _T_241[9:0] ? 4'h9 : _GEN_14894; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14896 = 10'h157 == _T_241[9:0] ? 4'h8 : _GEN_14895; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14897 = 10'h158 == _T_241[9:0] ? 4'h8 : _GEN_14896; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14898 = 10'h159 == _T_241[9:0] ? 4'h8 : _GEN_14897; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14899 = 10'h15a == _T_241[9:0] ? 4'h8 : _GEN_14898; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14900 = 10'h15b == _T_241[9:0] ? 4'h8 : _GEN_14899; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14901 = 10'h15c == _T_241[9:0] ? 4'h7 : _GEN_14900; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14902 = 10'h15d == _T_241[9:0] ? 4'h7 : _GEN_14901; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14903 = 10'h15e == _T_241[9:0] ? 4'h8 : _GEN_14902; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14904 = 10'h15f == _T_241[9:0] ? 4'h3 : _GEN_14903; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14905 = 10'h160 == _T_241[9:0] ? 4'h4 : _GEN_14904; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14906 = 10'h161 == _T_241[9:0] ? 4'h4 : _GEN_14905; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14907 = 10'h162 == _T_241[9:0] ? 4'h4 : _GEN_14906; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14908 = 10'h163 == _T_241[9:0] ? 4'h4 : _GEN_14907; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14909 = 10'h164 == _T_241[9:0] ? 4'h5 : _GEN_14908; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14910 = 10'h165 == _T_241[9:0] ? 4'ha : _GEN_14909; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14911 = 10'h166 == _T_241[9:0] ? 4'h9 : _GEN_14910; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14912 = 10'h167 == _T_241[9:0] ? 4'ha : _GEN_14911; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14913 = 10'h168 == _T_241[9:0] ? 4'ha : _GEN_14912; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14914 = 10'h169 == _T_241[9:0] ? 4'h6 : _GEN_14913; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14915 = 10'h16a == _T_241[9:0] ? 4'h3 : _GEN_14914; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14916 = 10'h16b == _T_241[9:0] ? 4'h3 : _GEN_14915; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14917 = 10'h16c == _T_241[9:0] ? 4'h3 : _GEN_14916; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14918 = 10'h16d == _T_241[9:0] ? 4'h4 : _GEN_14917; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14919 = 10'h16e == _T_241[9:0] ? 4'h3 : _GEN_14918; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14920 = 10'h16f == _T_241[9:0] ? 4'h3 : _GEN_14919; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14921 = 10'h170 == _T_241[9:0] ? 4'h3 : _GEN_14920; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14922 = 10'h171 == _T_241[9:0] ? 4'h7 : _GEN_14921; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14923 = 10'h172 == _T_241[9:0] ? 4'ha : _GEN_14922; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14924 = 10'h173 == _T_241[9:0] ? 4'h5 : _GEN_14923; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14925 = 10'h174 == _T_241[9:0] ? 4'h3 : _GEN_14924; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14926 = 10'h175 == _T_241[9:0] ? 4'h4 : _GEN_14925; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14927 = 10'h176 == _T_241[9:0] ? 4'h4 : _GEN_14926; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14928 = 10'h177 == _T_241[9:0] ? 4'h4 : _GEN_14927; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14929 = 10'h178 == _T_241[9:0] ? 4'h4 : _GEN_14928; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14930 = 10'h179 == _T_241[9:0] ? 4'h3 : _GEN_14929; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14931 = 10'h17a == _T_241[9:0] ? 4'h3 : _GEN_14930; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14932 = 10'h17b == _T_241[9:0] ? 4'h3 : _GEN_14931; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14933 = 10'h17c == _T_241[9:0] ? 4'h8 : _GEN_14932; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14934 = 10'h17d == _T_241[9:0] ? 4'h8 : _GEN_14933; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14935 = 10'h17e == _T_241[9:0] ? 4'h8 : _GEN_14934; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14936 = 10'h17f == _T_241[9:0] ? 4'h8 : _GEN_14935; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14937 = 10'h180 == _T_241[9:0] ? 4'h8 : _GEN_14936; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14938 = 10'h181 == _T_241[9:0] ? 4'h8 : _GEN_14937; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14939 = 10'h182 == _T_241[9:0] ? 4'h8 : _GEN_14938; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14940 = 10'h183 == _T_241[9:0] ? 4'h8 : _GEN_14939; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14941 = 10'h184 == _T_241[9:0] ? 4'h8 : _GEN_14940; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14942 = 10'h185 == _T_241[9:0] ? 4'h5 : _GEN_14941; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14943 = 10'h186 == _T_241[9:0] ? 4'h3 : _GEN_14942; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14944 = 10'h187 == _T_241[9:0] ? 4'h4 : _GEN_14943; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14945 = 10'h188 == _T_241[9:0] ? 4'h4 : _GEN_14944; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14946 = 10'h189 == _T_241[9:0] ? 4'h4 : _GEN_14945; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14947 = 10'h18a == _T_241[9:0] ? 4'h5 : _GEN_14946; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14948 = 10'h18b == _T_241[9:0] ? 4'ha : _GEN_14947; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14949 = 10'h18c == _T_241[9:0] ? 4'ha : _GEN_14948; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14950 = 10'h18d == _T_241[9:0] ? 4'h9 : _GEN_14949; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14951 = 10'h18e == _T_241[9:0] ? 4'ha : _GEN_14950; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14952 = 10'h18f == _T_241[9:0] ? 4'h4 : _GEN_14951; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14953 = 10'h190 == _T_241[9:0] ? 4'h3 : _GEN_14952; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14954 = 10'h191 == _T_241[9:0] ? 4'h3 : _GEN_14953; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14955 = 10'h192 == _T_241[9:0] ? 4'h5 : _GEN_14954; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14956 = 10'h193 == _T_241[9:0] ? 4'h6 : _GEN_14955; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14957 = 10'h194 == _T_241[9:0] ? 4'h5 : _GEN_14956; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14958 = 10'h195 == _T_241[9:0] ? 4'h3 : _GEN_14957; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14959 = 10'h196 == _T_241[9:0] ? 4'h3 : _GEN_14958; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14960 = 10'h197 == _T_241[9:0] ? 4'h5 : _GEN_14959; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14961 = 10'h198 == _T_241[9:0] ? 4'ha : _GEN_14960; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14962 = 10'h199 == _T_241[9:0] ? 4'h3 : _GEN_14961; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14963 = 10'h19a == _T_241[9:0] ? 4'h1 : _GEN_14962; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14964 = 10'h19b == _T_241[9:0] ? 4'h2 : _GEN_14963; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14965 = 10'h19c == _T_241[9:0] ? 4'h4 : _GEN_14964; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14966 = 10'h19d == _T_241[9:0] ? 4'h3 : _GEN_14965; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14967 = 10'h19e == _T_241[9:0] ? 4'h1 : _GEN_14966; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14968 = 10'h19f == _T_241[9:0] ? 4'h2 : _GEN_14967; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14969 = 10'h1a0 == _T_241[9:0] ? 4'h3 : _GEN_14968; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14970 = 10'h1a1 == _T_241[9:0] ? 4'h4 : _GEN_14969; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14971 = 10'h1a2 == _T_241[9:0] ? 4'h8 : _GEN_14970; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14972 = 10'h1a3 == _T_241[9:0] ? 4'h8 : _GEN_14971; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14973 = 10'h1a4 == _T_241[9:0] ? 4'h8 : _GEN_14972; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14974 = 10'h1a5 == _T_241[9:0] ? 4'h8 : _GEN_14973; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14975 = 10'h1a6 == _T_241[9:0] ? 4'h7 : _GEN_14974; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14976 = 10'h1a7 == _T_241[9:0] ? 4'h8 : _GEN_14975; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14977 = 10'h1a8 == _T_241[9:0] ? 4'h8 : _GEN_14976; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14978 = 10'h1a9 == _T_241[9:0] ? 4'h8 : _GEN_14977; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14979 = 10'h1aa == _T_241[9:0] ? 4'h7 : _GEN_14978; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14980 = 10'h1ab == _T_241[9:0] ? 4'h4 : _GEN_14979; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14981 = 10'h1ac == _T_241[9:0] ? 4'h4 : _GEN_14980; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14982 = 10'h1ad == _T_241[9:0] ? 4'h3 : _GEN_14981; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14983 = 10'h1ae == _T_241[9:0] ? 4'h3 : _GEN_14982; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14984 = 10'h1af == _T_241[9:0] ? 4'h4 : _GEN_14983; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14985 = 10'h1b0 == _T_241[9:0] ? 4'h6 : _GEN_14984; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14986 = 10'h1b1 == _T_241[9:0] ? 4'ha : _GEN_14985; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14987 = 10'h1b2 == _T_241[9:0] ? 4'ha : _GEN_14986; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14988 = 10'h1b3 == _T_241[9:0] ? 4'h9 : _GEN_14987; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14989 = 10'h1b4 == _T_241[9:0] ? 4'h9 : _GEN_14988; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14990 = 10'h1b5 == _T_241[9:0] ? 4'h3 : _GEN_14989; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14991 = 10'h1b6 == _T_241[9:0] ? 4'h3 : _GEN_14990; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14992 = 10'h1b7 == _T_241[9:0] ? 4'h4 : _GEN_14991; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14993 = 10'h1b8 == _T_241[9:0] ? 4'h5 : _GEN_14992; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14994 = 10'h1b9 == _T_241[9:0] ? 4'h6 : _GEN_14993; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14995 = 10'h1ba == _T_241[9:0] ? 4'h4 : _GEN_14994; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14996 = 10'h1bb == _T_241[9:0] ? 4'h3 : _GEN_14995; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14997 = 10'h1bc == _T_241[9:0] ? 4'h3 : _GEN_14996; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14998 = 10'h1bd == _T_241[9:0] ? 4'h4 : _GEN_14997; // @[Filter.scala 230:62]
  wire [3:0] _GEN_14999 = 10'h1be == _T_241[9:0] ? 4'ha : _GEN_14998; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15000 = 10'h1bf == _T_241[9:0] ? 4'h4 : _GEN_14999; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15001 = 10'h1c0 == _T_241[9:0] ? 4'h5 : _GEN_15000; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15002 = 10'h1c1 == _T_241[9:0] ? 4'h5 : _GEN_15001; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15003 = 10'h1c2 == _T_241[9:0] ? 4'h4 : _GEN_15002; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15004 = 10'h1c3 == _T_241[9:0] ? 4'h5 : _GEN_15003; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15005 = 10'h1c4 == _T_241[9:0] ? 4'h4 : _GEN_15004; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15006 = 10'h1c5 == _T_241[9:0] ? 4'h3 : _GEN_15005; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15007 = 10'h1c6 == _T_241[9:0] ? 4'h4 : _GEN_15006; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15008 = 10'h1c7 == _T_241[9:0] ? 4'h3 : _GEN_15007; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15009 = 10'h1c8 == _T_241[9:0] ? 4'h8 : _GEN_15008; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15010 = 10'h1c9 == _T_241[9:0] ? 4'h8 : _GEN_15009; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15011 = 10'h1ca == _T_241[9:0] ? 4'h8 : _GEN_15010; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15012 = 10'h1cb == _T_241[9:0] ? 4'h8 : _GEN_15011; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15013 = 10'h1cc == _T_241[9:0] ? 4'h8 : _GEN_15012; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15014 = 10'h1cd == _T_241[9:0] ? 4'h8 : _GEN_15013; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15015 = 10'h1ce == _T_241[9:0] ? 4'h8 : _GEN_15014; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15016 = 10'h1cf == _T_241[9:0] ? 4'h8 : _GEN_15015; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15017 = 10'h1d0 == _T_241[9:0] ? 4'h5 : _GEN_15016; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15018 = 10'h1d1 == _T_241[9:0] ? 4'h4 : _GEN_15017; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15019 = 10'h1d2 == _T_241[9:0] ? 4'h6 : _GEN_15018; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15020 = 10'h1d3 == _T_241[9:0] ? 4'h6 : _GEN_15019; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15021 = 10'h1d4 == _T_241[9:0] ? 4'h6 : _GEN_15020; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15022 = 10'h1d5 == _T_241[9:0] ? 4'h5 : _GEN_15021; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15023 = 10'h1d6 == _T_241[9:0] ? 4'h8 : _GEN_15022; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15024 = 10'h1d7 == _T_241[9:0] ? 4'ha : _GEN_15023; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15025 = 10'h1d8 == _T_241[9:0] ? 4'ha : _GEN_15024; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15026 = 10'h1d9 == _T_241[9:0] ? 4'ha : _GEN_15025; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15027 = 10'h1da == _T_241[9:0] ? 4'h6 : _GEN_15026; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15028 = 10'h1db == _T_241[9:0] ? 4'h3 : _GEN_15027; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15029 = 10'h1dc == _T_241[9:0] ? 4'h5 : _GEN_15028; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15030 = 10'h1dd == _T_241[9:0] ? 4'h2 : _GEN_15029; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15031 = 10'h1de == _T_241[9:0] ? 4'h5 : _GEN_15030; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15032 = 10'h1df == _T_241[9:0] ? 4'h5 : _GEN_15031; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15033 = 10'h1e0 == _T_241[9:0] ? 4'h5 : _GEN_15032; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15034 = 10'h1e1 == _T_241[9:0] ? 4'h3 : _GEN_15033; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15035 = 10'h1e2 == _T_241[9:0] ? 4'h3 : _GEN_15034; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15036 = 10'h1e3 == _T_241[9:0] ? 4'h3 : _GEN_15035; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15037 = 10'h1e4 == _T_241[9:0] ? 4'h9 : _GEN_15036; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15038 = 10'h1e5 == _T_241[9:0] ? 4'h4 : _GEN_15037; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15039 = 10'h1e6 == _T_241[9:0] ? 4'h4 : _GEN_15038; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15040 = 10'h1e7 == _T_241[9:0] ? 4'h4 : _GEN_15039; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15041 = 10'h1e8 == _T_241[9:0] ? 4'h4 : _GEN_15040; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15042 = 10'h1e9 == _T_241[9:0] ? 4'h4 : _GEN_15041; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15043 = 10'h1ea == _T_241[9:0] ? 4'h4 : _GEN_15042; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15044 = 10'h1eb == _T_241[9:0] ? 4'h4 : _GEN_15043; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15045 = 10'h1ec == _T_241[9:0] ? 4'h4 : _GEN_15044; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15046 = 10'h1ed == _T_241[9:0] ? 4'h4 : _GEN_15045; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15047 = 10'h1ee == _T_241[9:0] ? 4'h8 : _GEN_15046; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15048 = 10'h1ef == _T_241[9:0] ? 4'h8 : _GEN_15047; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15049 = 10'h1f0 == _T_241[9:0] ? 4'h8 : _GEN_15048; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15050 = 10'h1f1 == _T_241[9:0] ? 4'h8 : _GEN_15049; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15051 = 10'h1f2 == _T_241[9:0] ? 4'h8 : _GEN_15050; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15052 = 10'h1f3 == _T_241[9:0] ? 4'h8 : _GEN_15051; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15053 = 10'h1f4 == _T_241[9:0] ? 4'h9 : _GEN_15052; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15054 = 10'h1f5 == _T_241[9:0] ? 4'h9 : _GEN_15053; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15055 = 10'h1f6 == _T_241[9:0] ? 4'ha : _GEN_15054; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15056 = 10'h1f7 == _T_241[9:0] ? 4'h5 : _GEN_15055; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15057 = 10'h1f8 == _T_241[9:0] ? 4'h5 : _GEN_15056; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15058 = 10'h1f9 == _T_241[9:0] ? 4'h7 : _GEN_15057; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15059 = 10'h1fa == _T_241[9:0] ? 4'h7 : _GEN_15058; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15060 = 10'h1fb == _T_241[9:0] ? 4'h5 : _GEN_15059; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15061 = 10'h1fc == _T_241[9:0] ? 4'ha : _GEN_15060; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15062 = 10'h1fd == _T_241[9:0] ? 4'hb : _GEN_15061; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15063 = 10'h1fe == _T_241[9:0] ? 4'hb : _GEN_15062; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15064 = 10'h1ff == _T_241[9:0] ? 4'ha : _GEN_15063; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15065 = 10'h200 == _T_241[9:0] ? 4'h4 : _GEN_15064; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15066 = 10'h201 == _T_241[9:0] ? 4'h3 : _GEN_15065; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15067 = 10'h202 == _T_241[9:0] ? 4'h2 : _GEN_15066; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15068 = 10'h203 == _T_241[9:0] ? 4'h2 : _GEN_15067; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15069 = 10'h204 == _T_241[9:0] ? 4'h2 : _GEN_15068; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15070 = 10'h205 == _T_241[9:0] ? 4'h2 : _GEN_15069; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15071 = 10'h206 == _T_241[9:0] ? 4'h2 : _GEN_15070; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15072 = 10'h207 == _T_241[9:0] ? 4'h2 : _GEN_15071; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15073 = 10'h208 == _T_241[9:0] ? 4'h3 : _GEN_15072; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15074 = 10'h209 == _T_241[9:0] ? 4'h3 : _GEN_15073; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15075 = 10'h20a == _T_241[9:0] ? 4'h8 : _GEN_15074; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15076 = 10'h20b == _T_241[9:0] ? 4'h4 : _GEN_15075; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15077 = 10'h20c == _T_241[9:0] ? 4'h4 : _GEN_15076; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15078 = 10'h20d == _T_241[9:0] ? 4'h4 : _GEN_15077; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15079 = 10'h20e == _T_241[9:0] ? 4'h4 : _GEN_15078; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15080 = 10'h20f == _T_241[9:0] ? 4'h4 : _GEN_15079; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15081 = 10'h210 == _T_241[9:0] ? 4'h4 : _GEN_15080; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15082 = 10'h211 == _T_241[9:0] ? 4'h4 : _GEN_15081; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15083 = 10'h212 == _T_241[9:0] ? 4'h4 : _GEN_15082; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15084 = 10'h213 == _T_241[9:0] ? 4'h6 : _GEN_15083; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15085 = 10'h214 == _T_241[9:0] ? 4'h7 : _GEN_15084; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15086 = 10'h215 == _T_241[9:0] ? 4'h8 : _GEN_15085; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15087 = 10'h216 == _T_241[9:0] ? 4'h8 : _GEN_15086; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15088 = 10'h217 == _T_241[9:0] ? 4'h8 : _GEN_15087; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15089 = 10'h218 == _T_241[9:0] ? 4'h8 : _GEN_15088; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15090 = 10'h219 == _T_241[9:0] ? 4'h8 : _GEN_15089; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15091 = 10'h21a == _T_241[9:0] ? 4'h8 : _GEN_15090; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15092 = 10'h21b == _T_241[9:0] ? 4'h8 : _GEN_15091; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15093 = 10'h21c == _T_241[9:0] ? 4'ha : _GEN_15092; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15094 = 10'h21d == _T_241[9:0] ? 4'h9 : _GEN_15093; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15095 = 10'h21e == _T_241[9:0] ? 4'h6 : _GEN_15094; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15096 = 10'h21f == _T_241[9:0] ? 4'h4 : _GEN_15095; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15097 = 10'h220 == _T_241[9:0] ? 4'h4 : _GEN_15096; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15098 = 10'h221 == _T_241[9:0] ? 4'h5 : _GEN_15097; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15099 = 10'h222 == _T_241[9:0] ? 4'ha : _GEN_15098; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15100 = 10'h223 == _T_241[9:0] ? 4'ha : _GEN_15099; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15101 = 10'h224 == _T_241[9:0] ? 4'ha : _GEN_15100; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15102 = 10'h225 == _T_241[9:0] ? 4'h8 : _GEN_15101; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15103 = 10'h226 == _T_241[9:0] ? 4'h4 : _GEN_15102; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15104 = 10'h227 == _T_241[9:0] ? 4'h2 : _GEN_15103; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15105 = 10'h228 == _T_241[9:0] ? 4'h2 : _GEN_15104; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15106 = 10'h229 == _T_241[9:0] ? 4'h2 : _GEN_15105; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15107 = 10'h22a == _T_241[9:0] ? 4'h2 : _GEN_15106; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15108 = 10'h22b == _T_241[9:0] ? 4'h2 : _GEN_15107; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15109 = 10'h22c == _T_241[9:0] ? 4'h2 : _GEN_15108; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15110 = 10'h22d == _T_241[9:0] ? 4'h2 : _GEN_15109; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15111 = 10'h22e == _T_241[9:0] ? 4'h2 : _GEN_15110; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15112 = 10'h22f == _T_241[9:0] ? 4'h3 : _GEN_15111; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15113 = 10'h230 == _T_241[9:0] ? 4'h3 : _GEN_15112; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15114 = 10'h231 == _T_241[9:0] ? 4'h3 : _GEN_15113; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15115 = 10'h232 == _T_241[9:0] ? 4'h4 : _GEN_15114; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15116 = 10'h233 == _T_241[9:0] ? 4'h6 : _GEN_15115; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15117 = 10'h234 == _T_241[9:0] ? 4'h6 : _GEN_15116; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15118 = 10'h235 == _T_241[9:0] ? 4'h4 : _GEN_15117; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15119 = 10'h236 == _T_241[9:0] ? 4'h4 : _GEN_15118; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15120 = 10'h237 == _T_241[9:0] ? 4'h4 : _GEN_15119; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15121 = 10'h238 == _T_241[9:0] ? 4'h4 : _GEN_15120; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15122 = 10'h239 == _T_241[9:0] ? 4'h3 : _GEN_15121; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15123 = 10'h23a == _T_241[9:0] ? 4'h7 : _GEN_15122; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15124 = 10'h23b == _T_241[9:0] ? 4'h7 : _GEN_15123; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15125 = 10'h23c == _T_241[9:0] ? 4'h7 : _GEN_15124; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15126 = 10'h23d == _T_241[9:0] ? 4'h7 : _GEN_15125; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15127 = 10'h23e == _T_241[9:0] ? 4'h7 : _GEN_15126; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15128 = 10'h23f == _T_241[9:0] ? 4'h7 : _GEN_15127; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15129 = 10'h240 == _T_241[9:0] ? 4'h7 : _GEN_15128; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15130 = 10'h241 == _T_241[9:0] ? 4'h8 : _GEN_15129; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15131 = 10'h242 == _T_241[9:0] ? 4'ha : _GEN_15130; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15132 = 10'h243 == _T_241[9:0] ? 4'ha : _GEN_15131; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15133 = 10'h244 == _T_241[9:0] ? 4'ha : _GEN_15132; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15134 = 10'h245 == _T_241[9:0] ? 4'h8 : _GEN_15133; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15135 = 10'h246 == _T_241[9:0] ? 4'h7 : _GEN_15134; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15136 = 10'h247 == _T_241[9:0] ? 4'h8 : _GEN_15135; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15137 = 10'h248 == _T_241[9:0] ? 4'ha : _GEN_15136; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15138 = 10'h249 == _T_241[9:0] ? 4'ha : _GEN_15137; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15139 = 10'h24a == _T_241[9:0] ? 4'ha : _GEN_15138; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15140 = 10'h24b == _T_241[9:0] ? 4'h4 : _GEN_15139; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15141 = 10'h24c == _T_241[9:0] ? 4'h4 : _GEN_15140; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15142 = 10'h24d == _T_241[9:0] ? 4'h2 : _GEN_15141; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15143 = 10'h24e == _T_241[9:0] ? 4'h2 : _GEN_15142; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15144 = 10'h24f == _T_241[9:0] ? 4'h2 : _GEN_15143; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15145 = 10'h250 == _T_241[9:0] ? 4'h2 : _GEN_15144; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15146 = 10'h251 == _T_241[9:0] ? 4'h2 : _GEN_15145; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15147 = 10'h252 == _T_241[9:0] ? 4'h2 : _GEN_15146; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15148 = 10'h253 == _T_241[9:0] ? 4'h2 : _GEN_15147; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15149 = 10'h254 == _T_241[9:0] ? 4'h2 : _GEN_15148; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15150 = 10'h255 == _T_241[9:0] ? 4'h3 : _GEN_15149; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15151 = 10'h256 == _T_241[9:0] ? 4'h4 : _GEN_15150; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15152 = 10'h257 == _T_241[9:0] ? 4'h3 : _GEN_15151; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15153 = 10'h258 == _T_241[9:0] ? 4'h4 : _GEN_15152; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15154 = 10'h259 == _T_241[9:0] ? 4'h4 : _GEN_15153; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15155 = 10'h25a == _T_241[9:0] ? 4'h4 : _GEN_15154; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15156 = 10'h25b == _T_241[9:0] ? 4'h3 : _GEN_15155; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15157 = 10'h25c == _T_241[9:0] ? 4'h4 : _GEN_15156; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15158 = 10'h25d == _T_241[9:0] ? 4'h4 : _GEN_15157; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15159 = 10'h25e == _T_241[9:0] ? 4'h3 : _GEN_15158; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15160 = 10'h25f == _T_241[9:0] ? 4'h3 : _GEN_15159; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15161 = 10'h260 == _T_241[9:0] ? 4'h8 : _GEN_15160; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15162 = 10'h261 == _T_241[9:0] ? 4'h7 : _GEN_15161; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15163 = 10'h262 == _T_241[9:0] ? 4'h6 : _GEN_15162; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15164 = 10'h263 == _T_241[9:0] ? 4'h5 : _GEN_15163; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15165 = 10'h264 == _T_241[9:0] ? 4'h6 : _GEN_15164; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15166 = 10'h265 == _T_241[9:0] ? 4'h5 : _GEN_15165; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15167 = 10'h266 == _T_241[9:0] ? 4'h5 : _GEN_15166; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15168 = 10'h267 == _T_241[9:0] ? 4'h7 : _GEN_15167; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15169 = 10'h268 == _T_241[9:0] ? 4'ha : _GEN_15168; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15170 = 10'h269 == _T_241[9:0] ? 4'ha : _GEN_15169; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15171 = 10'h26a == _T_241[9:0] ? 4'ha : _GEN_15170; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15172 = 10'h26b == _T_241[9:0] ? 4'ha : _GEN_15171; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15173 = 10'h26c == _T_241[9:0] ? 4'ha : _GEN_15172; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15174 = 10'h26d == _T_241[9:0] ? 4'ha : _GEN_15173; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15175 = 10'h26e == _T_241[9:0] ? 4'ha : _GEN_15174; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15176 = 10'h26f == _T_241[9:0] ? 4'ha : _GEN_15175; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15177 = 10'h270 == _T_241[9:0] ? 4'h5 : _GEN_15176; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15178 = 10'h271 == _T_241[9:0] ? 4'h4 : _GEN_15177; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15179 = 10'h272 == _T_241[9:0] ? 4'h3 : _GEN_15178; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15180 = 10'h273 == _T_241[9:0] ? 4'h2 : _GEN_15179; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15181 = 10'h274 == _T_241[9:0] ? 4'h2 : _GEN_15180; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15182 = 10'h275 == _T_241[9:0] ? 4'h2 : _GEN_15181; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15183 = 10'h276 == _T_241[9:0] ? 4'h2 : _GEN_15182; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15184 = 10'h277 == _T_241[9:0] ? 4'h2 : _GEN_15183; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15185 = 10'h278 == _T_241[9:0] ? 4'h2 : _GEN_15184; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15186 = 10'h279 == _T_241[9:0] ? 4'h2 : _GEN_15185; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15187 = 10'h27a == _T_241[9:0] ? 4'h2 : _GEN_15186; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15188 = 10'h27b == _T_241[9:0] ? 4'h4 : _GEN_15187; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15189 = 10'h27c == _T_241[9:0] ? 4'h3 : _GEN_15188; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15190 = 10'h27d == _T_241[9:0] ? 4'h4 : _GEN_15189; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15191 = 10'h27e == _T_241[9:0] ? 4'h5 : _GEN_15190; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15192 = 10'h27f == _T_241[9:0] ? 4'h4 : _GEN_15191; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15193 = 10'h280 == _T_241[9:0] ? 4'h4 : _GEN_15192; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15194 = 10'h281 == _T_241[9:0] ? 4'h4 : _GEN_15193; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15195 = 10'h282 == _T_241[9:0] ? 4'h4 : _GEN_15194; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15196 = 10'h283 == _T_241[9:0] ? 4'h3 : _GEN_15195; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15197 = 10'h284 == _T_241[9:0] ? 4'h3 : _GEN_15196; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15198 = 10'h285 == _T_241[9:0] ? 4'h3 : _GEN_15197; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15199 = 10'h286 == _T_241[9:0] ? 4'h8 : _GEN_15198; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15200 = 10'h287 == _T_241[9:0] ? 4'h6 : _GEN_15199; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15201 = 10'h288 == _T_241[9:0] ? 4'h6 : _GEN_15200; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15202 = 10'h289 == _T_241[9:0] ? 4'h6 : _GEN_15201; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15203 = 10'h28a == _T_241[9:0] ? 4'h7 : _GEN_15202; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15204 = 10'h28b == _T_241[9:0] ? 4'h7 : _GEN_15203; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15205 = 10'h28c == _T_241[9:0] ? 4'h6 : _GEN_15204; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15206 = 10'h28d == _T_241[9:0] ? 4'h6 : _GEN_15205; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15207 = 10'h28e == _T_241[9:0] ? 4'h4 : _GEN_15206; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15208 = 10'h28f == _T_241[9:0] ? 4'h7 : _GEN_15207; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15209 = 10'h290 == _T_241[9:0] ? 4'h9 : _GEN_15208; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15210 = 10'h291 == _T_241[9:0] ? 4'ha : _GEN_15209; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15211 = 10'h292 == _T_241[9:0] ? 4'ha : _GEN_15210; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15212 = 10'h293 == _T_241[9:0] ? 4'ha : _GEN_15211; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15213 = 10'h294 == _T_241[9:0] ? 4'h9 : _GEN_15212; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15214 = 10'h295 == _T_241[9:0] ? 4'h5 : _GEN_15213; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15215 = 10'h296 == _T_241[9:0] ? 4'h4 : _GEN_15214; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15216 = 10'h297 == _T_241[9:0] ? 4'h4 : _GEN_15215; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15217 = 10'h298 == _T_241[9:0] ? 4'h3 : _GEN_15216; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15218 = 10'h299 == _T_241[9:0] ? 4'h3 : _GEN_15217; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15219 = 10'h29a == _T_241[9:0] ? 4'h2 : _GEN_15218; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15220 = 10'h29b == _T_241[9:0] ? 4'h2 : _GEN_15219; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15221 = 10'h29c == _T_241[9:0] ? 4'h2 : _GEN_15220; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15222 = 10'h29d == _T_241[9:0] ? 4'h2 : _GEN_15221; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15223 = 10'h29e == _T_241[9:0] ? 4'h2 : _GEN_15222; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15224 = 10'h29f == _T_241[9:0] ? 4'h2 : _GEN_15223; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15225 = 10'h2a0 == _T_241[9:0] ? 4'h2 : _GEN_15224; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15226 = 10'h2a1 == _T_241[9:0] ? 4'h4 : _GEN_15225; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15227 = 10'h2a2 == _T_241[9:0] ? 4'h3 : _GEN_15226; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15228 = 10'h2a3 == _T_241[9:0] ? 4'h4 : _GEN_15227; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15229 = 10'h2a4 == _T_241[9:0] ? 4'h5 : _GEN_15228; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15230 = 10'h2a5 == _T_241[9:0] ? 4'h4 : _GEN_15229; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15231 = 10'h2a6 == _T_241[9:0] ? 4'h4 : _GEN_15230; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15232 = 10'h2a7 == _T_241[9:0] ? 4'h4 : _GEN_15231; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15233 = 10'h2a8 == _T_241[9:0] ? 4'h3 : _GEN_15232; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15234 = 10'h2a9 == _T_241[9:0] ? 4'h3 : _GEN_15233; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15235 = 10'h2aa == _T_241[9:0] ? 4'h3 : _GEN_15234; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15236 = 10'h2ab == _T_241[9:0] ? 4'h3 : _GEN_15235; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15237 = 10'h2ac == _T_241[9:0] ? 4'h8 : _GEN_15236; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15238 = 10'h2ad == _T_241[9:0] ? 4'h7 : _GEN_15237; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15239 = 10'h2ae == _T_241[9:0] ? 4'h5 : _GEN_15238; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15240 = 10'h2af == _T_241[9:0] ? 4'h6 : _GEN_15239; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15241 = 10'h2b0 == _T_241[9:0] ? 4'h7 : _GEN_15240; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15242 = 10'h2b1 == _T_241[9:0] ? 4'h6 : _GEN_15241; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15243 = 10'h2b2 == _T_241[9:0] ? 4'h6 : _GEN_15242; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15244 = 10'h2b3 == _T_241[9:0] ? 4'h6 : _GEN_15243; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15245 = 10'h2b4 == _T_241[9:0] ? 4'h3 : _GEN_15244; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15246 = 10'h2b5 == _T_241[9:0] ? 4'h3 : _GEN_15245; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15247 = 10'h2b6 == _T_241[9:0] ? 4'h3 : _GEN_15246; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15248 = 10'h2b7 == _T_241[9:0] ? 4'h4 : _GEN_15247; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15249 = 10'h2b8 == _T_241[9:0] ? 4'h6 : _GEN_15248; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15250 = 10'h2b9 == _T_241[9:0] ? 4'h9 : _GEN_15249; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15251 = 10'h2ba == _T_241[9:0] ? 4'h4 : _GEN_15250; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15252 = 10'h2bb == _T_241[9:0] ? 4'h3 : _GEN_15251; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15253 = 10'h2bc == _T_241[9:0] ? 4'h4 : _GEN_15252; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15254 = 10'h2bd == _T_241[9:0] ? 4'h3 : _GEN_15253; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15255 = 10'h2be == _T_241[9:0] ? 4'h3 : _GEN_15254; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15256 = 10'h2bf == _T_241[9:0] ? 4'h3 : _GEN_15255; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15257 = 10'h2c0 == _T_241[9:0] ? 4'h2 : _GEN_15256; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15258 = 10'h2c1 == _T_241[9:0] ? 4'h2 : _GEN_15257; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15259 = 10'h2c2 == _T_241[9:0] ? 4'h2 : _GEN_15258; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15260 = 10'h2c3 == _T_241[9:0] ? 4'h2 : _GEN_15259; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15261 = 10'h2c4 == _T_241[9:0] ? 4'h2 : _GEN_15260; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15262 = 10'h2c5 == _T_241[9:0] ? 4'h2 : _GEN_15261; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15263 = 10'h2c6 == _T_241[9:0] ? 4'h2 : _GEN_15262; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15264 = 10'h2c7 == _T_241[9:0] ? 4'h4 : _GEN_15263; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15265 = 10'h2c8 == _T_241[9:0] ? 4'h3 : _GEN_15264; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15266 = 10'h2c9 == _T_241[9:0] ? 4'h4 : _GEN_15265; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15267 = 10'h2ca == _T_241[9:0] ? 4'h5 : _GEN_15266; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15268 = 10'h2cb == _T_241[9:0] ? 4'h3 : _GEN_15267; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15269 = 10'h2cc == _T_241[9:0] ? 4'h3 : _GEN_15268; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15270 = 10'h2cd == _T_241[9:0] ? 4'h3 : _GEN_15269; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15271 = 10'h2ce == _T_241[9:0] ? 4'h3 : _GEN_15270; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15272 = 10'h2cf == _T_241[9:0] ? 4'h3 : _GEN_15271; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15273 = 10'h2d0 == _T_241[9:0] ? 4'h3 : _GEN_15272; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15274 = 10'h2d1 == _T_241[9:0] ? 4'h3 : _GEN_15273; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15275 = 10'h2d2 == _T_241[9:0] ? 4'h8 : _GEN_15274; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15276 = 10'h2d3 == _T_241[9:0] ? 4'h6 : _GEN_15275; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15277 = 10'h2d4 == _T_241[9:0] ? 4'h6 : _GEN_15276; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15278 = 10'h2d5 == _T_241[9:0] ? 4'h7 : _GEN_15277; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15279 = 10'h2d6 == _T_241[9:0] ? 4'h7 : _GEN_15278; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15280 = 10'h2d7 == _T_241[9:0] ? 4'h7 : _GEN_15279; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15281 = 10'h2d8 == _T_241[9:0] ? 4'h6 : _GEN_15280; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15282 = 10'h2d9 == _T_241[9:0] ? 4'h7 : _GEN_15281; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15283 = 10'h2da == _T_241[9:0] ? 4'h5 : _GEN_15282; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15284 = 10'h2db == _T_241[9:0] ? 4'h3 : _GEN_15283; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15285 = 10'h2dc == _T_241[9:0] ? 4'h3 : _GEN_15284; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15286 = 10'h2dd == _T_241[9:0] ? 4'h3 : _GEN_15285; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15287 = 10'h2de == _T_241[9:0] ? 4'h3 : _GEN_15286; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15288 = 10'h2df == _T_241[9:0] ? 4'h4 : _GEN_15287; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15289 = 10'h2e0 == _T_241[9:0] ? 4'h3 : _GEN_15288; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15290 = 10'h2e1 == _T_241[9:0] ? 4'h3 : _GEN_15289; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15291 = 10'h2e2 == _T_241[9:0] ? 4'h3 : _GEN_15290; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15292 = 10'h2e3 == _T_241[9:0] ? 4'h3 : _GEN_15291; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15293 = 10'h2e4 == _T_241[9:0] ? 4'h3 : _GEN_15292; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15294 = 10'h2e5 == _T_241[9:0] ? 4'h3 : _GEN_15293; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15295 = 10'h2e6 == _T_241[9:0] ? 4'h2 : _GEN_15294; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15296 = 10'h2e7 == _T_241[9:0] ? 4'h2 : _GEN_15295; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15297 = 10'h2e8 == _T_241[9:0] ? 4'h2 : _GEN_15296; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15298 = 10'h2e9 == _T_241[9:0] ? 4'h2 : _GEN_15297; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15299 = 10'h2ea == _T_241[9:0] ? 4'h2 : _GEN_15298; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15300 = 10'h2eb == _T_241[9:0] ? 4'h2 : _GEN_15299; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15301 = 10'h2ec == _T_241[9:0] ? 4'h3 : _GEN_15300; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15302 = 10'h2ed == _T_241[9:0] ? 4'h4 : _GEN_15301; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15303 = 10'h2ee == _T_241[9:0] ? 4'h3 : _GEN_15302; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15304 = 10'h2ef == _T_241[9:0] ? 4'h3 : _GEN_15303; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15305 = 10'h2f0 == _T_241[9:0] ? 4'h6 : _GEN_15304; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15306 = 10'h2f1 == _T_241[9:0] ? 4'h3 : _GEN_15305; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15307 = 10'h2f2 == _T_241[9:0] ? 4'h3 : _GEN_15306; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15308 = 10'h2f3 == _T_241[9:0] ? 4'h3 : _GEN_15307; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15309 = 10'h2f4 == _T_241[9:0] ? 4'h3 : _GEN_15308; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15310 = 10'h2f5 == _T_241[9:0] ? 4'h3 : _GEN_15309; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15311 = 10'h2f6 == _T_241[9:0] ? 4'h3 : _GEN_15310; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15312 = 10'h2f7 == _T_241[9:0] ? 4'h3 : _GEN_15311; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15313 = 10'h2f8 == _T_241[9:0] ? 4'h8 : _GEN_15312; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15314 = 10'h2f9 == _T_241[9:0] ? 4'h6 : _GEN_15313; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15315 = 10'h2fa == _T_241[9:0] ? 4'h7 : _GEN_15314; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15316 = 10'h2fb == _T_241[9:0] ? 4'h7 : _GEN_15315; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15317 = 10'h2fc == _T_241[9:0] ? 4'h6 : _GEN_15316; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15318 = 10'h2fd == _T_241[9:0] ? 4'h6 : _GEN_15317; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15319 = 10'h2fe == _T_241[9:0] ? 4'h6 : _GEN_15318; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15320 = 10'h2ff == _T_241[9:0] ? 4'h8 : _GEN_15319; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15321 = 10'h300 == _T_241[9:0] ? 4'h9 : _GEN_15320; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15322 = 10'h301 == _T_241[9:0] ? 4'h7 : _GEN_15321; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15323 = 10'h302 == _T_241[9:0] ? 4'h4 : _GEN_15322; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15324 = 10'h303 == _T_241[9:0] ? 4'h4 : _GEN_15323; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15325 = 10'h304 == _T_241[9:0] ? 4'h3 : _GEN_15324; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15326 = 10'h305 == _T_241[9:0] ? 4'h3 : _GEN_15325; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15327 = 10'h306 == _T_241[9:0] ? 4'h3 : _GEN_15326; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15328 = 10'h307 == _T_241[9:0] ? 4'h3 : _GEN_15327; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15329 = 10'h308 == _T_241[9:0] ? 4'h3 : _GEN_15328; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15330 = 10'h309 == _T_241[9:0] ? 4'h3 : _GEN_15329; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15331 = 10'h30a == _T_241[9:0] ? 4'h3 : _GEN_15330; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15332 = 10'h30b == _T_241[9:0] ? 4'h3 : _GEN_15331; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15333 = 10'h30c == _T_241[9:0] ? 4'h2 : _GEN_15332; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15334 = 10'h30d == _T_241[9:0] ? 4'h2 : _GEN_15333; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15335 = 10'h30e == _T_241[9:0] ? 4'h2 : _GEN_15334; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15336 = 10'h30f == _T_241[9:0] ? 4'h2 : _GEN_15335; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15337 = 10'h310 == _T_241[9:0] ? 4'h2 : _GEN_15336; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15338 = 10'h311 == _T_241[9:0] ? 4'h2 : _GEN_15337; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15339 = 10'h312 == _T_241[9:0] ? 4'h3 : _GEN_15338; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15340 = 10'h313 == _T_241[9:0] ? 4'h4 : _GEN_15339; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15341 = 10'h314 == _T_241[9:0] ? 4'h3 : _GEN_15340; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15342 = 10'h315 == _T_241[9:0] ? 4'h3 : _GEN_15341; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15343 = 10'h316 == _T_241[9:0] ? 4'h5 : _GEN_15342; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15344 = 10'h317 == _T_241[9:0] ? 4'h5 : _GEN_15343; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15345 = 10'h318 == _T_241[9:0] ? 4'h3 : _GEN_15344; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15346 = 10'h319 == _T_241[9:0] ? 4'h3 : _GEN_15345; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15347 = 10'h31a == _T_241[9:0] ? 4'h3 : _GEN_15346; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15348 = 10'h31b == _T_241[9:0] ? 4'h3 : _GEN_15347; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15349 = 10'h31c == _T_241[9:0] ? 4'h3 : _GEN_15348; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15350 = 10'h31d == _T_241[9:0] ? 4'h3 : _GEN_15349; // @[Filter.scala 230:62]
  wire [4:0] _GEN_38990 = {{1'd0}, _GEN_15350}; // @[Filter.scala 230:62]
  wire [8:0] _T_243 = _GEN_38990 * 5'h14; // @[Filter.scala 230:62]
  wire [3:0] _GEN_15374 = 10'h17 == _T_241[9:0] ? 4'hb : 4'he; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15375 = 10'h18 == _T_241[9:0] ? 4'hc : _GEN_15374; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15376 = 10'h19 == _T_241[9:0] ? 4'he : _GEN_15375; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15377 = 10'h1a == _T_241[9:0] ? 4'he : _GEN_15376; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15378 = 10'h1b == _T_241[9:0] ? 4'he : _GEN_15377; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15379 = 10'h1c == _T_241[9:0] ? 4'he : _GEN_15378; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15380 = 10'h1d == _T_241[9:0] ? 4'he : _GEN_15379; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15381 = 10'h1e == _T_241[9:0] ? 4'he : _GEN_15380; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15382 = 10'h1f == _T_241[9:0] ? 4'he : _GEN_15381; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15383 = 10'h20 == _T_241[9:0] ? 4'he : _GEN_15382; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15384 = 10'h21 == _T_241[9:0] ? 4'he : _GEN_15383; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15385 = 10'h22 == _T_241[9:0] ? 4'he : _GEN_15384; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15386 = 10'h23 == _T_241[9:0] ? 4'he : _GEN_15385; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15387 = 10'h24 == _T_241[9:0] ? 4'he : _GEN_15386; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15388 = 10'h25 == _T_241[9:0] ? 4'he : _GEN_15387; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15389 = 10'h26 == _T_241[9:0] ? 4'he : _GEN_15388; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15390 = 10'h27 == _T_241[9:0] ? 4'he : _GEN_15389; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15391 = 10'h28 == _T_241[9:0] ? 4'he : _GEN_15390; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15392 = 10'h29 == _T_241[9:0] ? 4'he : _GEN_15391; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15393 = 10'h2a == _T_241[9:0] ? 4'he : _GEN_15392; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15394 = 10'h2b == _T_241[9:0] ? 4'he : _GEN_15393; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15395 = 10'h2c == _T_241[9:0] ? 4'he : _GEN_15394; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15396 = 10'h2d == _T_241[9:0] ? 4'he : _GEN_15395; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15397 = 10'h2e == _T_241[9:0] ? 4'he : _GEN_15396; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15398 = 10'h2f == _T_241[9:0] ? 4'he : _GEN_15397; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15399 = 10'h30 == _T_241[9:0] ? 4'he : _GEN_15398; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15400 = 10'h31 == _T_241[9:0] ? 4'he : _GEN_15399; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15401 = 10'h32 == _T_241[9:0] ? 4'he : _GEN_15400; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15402 = 10'h33 == _T_241[9:0] ? 4'he : _GEN_15401; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15403 = 10'h34 == _T_241[9:0] ? 4'he : _GEN_15402; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15404 = 10'h35 == _T_241[9:0] ? 4'he : _GEN_15403; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15405 = 10'h36 == _T_241[9:0] ? 4'he : _GEN_15404; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15406 = 10'h37 == _T_241[9:0] ? 4'he : _GEN_15405; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15407 = 10'h38 == _T_241[9:0] ? 4'he : _GEN_15406; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15408 = 10'h39 == _T_241[9:0] ? 4'he : _GEN_15407; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15409 = 10'h3a == _T_241[9:0] ? 4'he : _GEN_15408; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15410 = 10'h3b == _T_241[9:0] ? 4'he : _GEN_15409; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15411 = 10'h3c == _T_241[9:0] ? 4'ha : _GEN_15410; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15412 = 10'h3d == _T_241[9:0] ? 4'hc : _GEN_15411; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15413 = 10'h3e == _T_241[9:0] ? 4'hb : _GEN_15412; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15414 = 10'h3f == _T_241[9:0] ? 4'he : _GEN_15413; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15415 = 10'h40 == _T_241[9:0] ? 4'he : _GEN_15414; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15416 = 10'h41 == _T_241[9:0] ? 4'he : _GEN_15415; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15417 = 10'h42 == _T_241[9:0] ? 4'he : _GEN_15416; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15418 = 10'h43 == _T_241[9:0] ? 4'he : _GEN_15417; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15419 = 10'h44 == _T_241[9:0] ? 4'he : _GEN_15418; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15420 = 10'h45 == _T_241[9:0] ? 4'he : _GEN_15419; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15421 = 10'h46 == _T_241[9:0] ? 4'he : _GEN_15420; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15422 = 10'h47 == _T_241[9:0] ? 4'he : _GEN_15421; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15423 = 10'h48 == _T_241[9:0] ? 4'he : _GEN_15422; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15424 = 10'h49 == _T_241[9:0] ? 4'he : _GEN_15423; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15425 = 10'h4a == _T_241[9:0] ? 4'he : _GEN_15424; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15426 = 10'h4b == _T_241[9:0] ? 4'he : _GEN_15425; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15427 = 10'h4c == _T_241[9:0] ? 4'he : _GEN_15426; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15428 = 10'h4d == _T_241[9:0] ? 4'he : _GEN_15427; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15429 = 10'h4e == _T_241[9:0] ? 4'he : _GEN_15428; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15430 = 10'h4f == _T_241[9:0] ? 4'he : _GEN_15429; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15431 = 10'h50 == _T_241[9:0] ? 4'he : _GEN_15430; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15432 = 10'h51 == _T_241[9:0] ? 4'he : _GEN_15431; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15433 = 10'h52 == _T_241[9:0] ? 4'he : _GEN_15432; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15434 = 10'h53 == _T_241[9:0] ? 4'he : _GEN_15433; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15435 = 10'h54 == _T_241[9:0] ? 4'he : _GEN_15434; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15436 = 10'h55 == _T_241[9:0] ? 4'he : _GEN_15435; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15437 = 10'h56 == _T_241[9:0] ? 4'he : _GEN_15436; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15438 = 10'h57 == _T_241[9:0] ? 4'he : _GEN_15437; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15439 = 10'h58 == _T_241[9:0] ? 4'he : _GEN_15438; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15440 = 10'h59 == _T_241[9:0] ? 4'he : _GEN_15439; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15441 = 10'h5a == _T_241[9:0] ? 4'hc : _GEN_15440; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15442 = 10'h5b == _T_241[9:0] ? 4'hd : _GEN_15441; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15443 = 10'h5c == _T_241[9:0] ? 4'he : _GEN_15442; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15444 = 10'h5d == _T_241[9:0] ? 4'he : _GEN_15443; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15445 = 10'h5e == _T_241[9:0] ? 4'he : _GEN_15444; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15446 = 10'h5f == _T_241[9:0] ? 4'he : _GEN_15445; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15447 = 10'h60 == _T_241[9:0] ? 4'he : _GEN_15446; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15448 = 10'h61 == _T_241[9:0] ? 4'hd : _GEN_15447; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15449 = 10'h62 == _T_241[9:0] ? 4'hb : _GEN_15448; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15450 = 10'h63 == _T_241[9:0] ? 4'hc : _GEN_15449; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15451 = 10'h64 == _T_241[9:0] ? 4'ha : _GEN_15450; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15452 = 10'h65 == _T_241[9:0] ? 4'hd : _GEN_15451; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15453 = 10'h66 == _T_241[9:0] ? 4'he : _GEN_15452; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15454 = 10'h67 == _T_241[9:0] ? 4'he : _GEN_15453; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15455 = 10'h68 == _T_241[9:0] ? 4'he : _GEN_15454; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15456 = 10'h69 == _T_241[9:0] ? 4'he : _GEN_15455; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15457 = 10'h6a == _T_241[9:0] ? 4'he : _GEN_15456; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15458 = 10'h6b == _T_241[9:0] ? 4'hd : _GEN_15457; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15459 = 10'h6c == _T_241[9:0] ? 4'hc : _GEN_15458; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15460 = 10'h6d == _T_241[9:0] ? 4'hc : _GEN_15459; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15461 = 10'h6e == _T_241[9:0] ? 4'he : _GEN_15460; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15462 = 10'h6f == _T_241[9:0] ? 4'he : _GEN_15461; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15463 = 10'h70 == _T_241[9:0] ? 4'he : _GEN_15462; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15464 = 10'h71 == _T_241[9:0] ? 4'he : _GEN_15463; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15465 = 10'h72 == _T_241[9:0] ? 4'he : _GEN_15464; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15466 = 10'h73 == _T_241[9:0] ? 4'he : _GEN_15465; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15467 = 10'h74 == _T_241[9:0] ? 4'he : _GEN_15466; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15468 = 10'h75 == _T_241[9:0] ? 4'he : _GEN_15467; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15469 = 10'h76 == _T_241[9:0] ? 4'he : _GEN_15468; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15470 = 10'h77 == _T_241[9:0] ? 4'he : _GEN_15469; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15471 = 10'h78 == _T_241[9:0] ? 4'he : _GEN_15470; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15472 = 10'h79 == _T_241[9:0] ? 4'he : _GEN_15471; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15473 = 10'h7a == _T_241[9:0] ? 4'he : _GEN_15472; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15474 = 10'h7b == _T_241[9:0] ? 4'he : _GEN_15473; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15475 = 10'h7c == _T_241[9:0] ? 4'he : _GEN_15474; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15476 = 10'h7d == _T_241[9:0] ? 4'he : _GEN_15475; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15477 = 10'h7e == _T_241[9:0] ? 4'he : _GEN_15476; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15478 = 10'h7f == _T_241[9:0] ? 4'he : _GEN_15477; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15479 = 10'h80 == _T_241[9:0] ? 4'he : _GEN_15478; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15480 = 10'h81 == _T_241[9:0] ? 4'hb : _GEN_15479; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15481 = 10'h82 == _T_241[9:0] ? 4'hc : _GEN_15480; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15482 = 10'h83 == _T_241[9:0] ? 4'hc : _GEN_15481; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15483 = 10'h84 == _T_241[9:0] ? 4'he : _GEN_15482; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15484 = 10'h85 == _T_241[9:0] ? 4'he : _GEN_15483; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15485 = 10'h86 == _T_241[9:0] ? 4'he : _GEN_15484; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15486 = 10'h87 == _T_241[9:0] ? 4'ha : _GEN_15485; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15487 = 10'h88 == _T_241[9:0] ? 4'hd : _GEN_15486; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15488 = 10'h89 == _T_241[9:0] ? 4'hd : _GEN_15487; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15489 = 10'h8a == _T_241[9:0] ? 4'hc : _GEN_15488; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15490 = 10'h8b == _T_241[9:0] ? 4'he : _GEN_15489; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15491 = 10'h8c == _T_241[9:0] ? 4'he : _GEN_15490; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15492 = 10'h8d == _T_241[9:0] ? 4'he : _GEN_15491; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15493 = 10'h8e == _T_241[9:0] ? 4'he : _GEN_15492; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15494 = 10'h8f == _T_241[9:0] ? 4'hb : _GEN_15493; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15495 = 10'h90 == _T_241[9:0] ? 4'hc : _GEN_15494; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15496 = 10'h91 == _T_241[9:0] ? 4'hc : _GEN_15495; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15497 = 10'h92 == _T_241[9:0] ? 4'hd : _GEN_15496; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15498 = 10'h93 == _T_241[9:0] ? 4'he : _GEN_15497; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15499 = 10'h94 == _T_241[9:0] ? 4'he : _GEN_15498; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15500 = 10'h95 == _T_241[9:0] ? 4'he : _GEN_15499; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15501 = 10'h96 == _T_241[9:0] ? 4'he : _GEN_15500; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15502 = 10'h97 == _T_241[9:0] ? 4'he : _GEN_15501; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15503 = 10'h98 == _T_241[9:0] ? 4'he : _GEN_15502; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15504 = 10'h99 == _T_241[9:0] ? 4'he : _GEN_15503; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15505 = 10'h9a == _T_241[9:0] ? 4'he : _GEN_15504; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15506 = 10'h9b == _T_241[9:0] ? 4'he : _GEN_15505; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15507 = 10'h9c == _T_241[9:0] ? 4'he : _GEN_15506; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15508 = 10'h9d == _T_241[9:0] ? 4'he : _GEN_15507; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15509 = 10'h9e == _T_241[9:0] ? 4'he : _GEN_15508; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15510 = 10'h9f == _T_241[9:0] ? 4'he : _GEN_15509; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15511 = 10'ha0 == _T_241[9:0] ? 4'he : _GEN_15510; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15512 = 10'ha1 == _T_241[9:0] ? 4'he : _GEN_15511; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15513 = 10'ha2 == _T_241[9:0] ? 4'he : _GEN_15512; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15514 = 10'ha3 == _T_241[9:0] ? 4'he : _GEN_15513; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15515 = 10'ha4 == _T_241[9:0] ? 4'he : _GEN_15514; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15516 = 10'ha5 == _T_241[9:0] ? 4'he : _GEN_15515; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15517 = 10'ha6 == _T_241[9:0] ? 4'he : _GEN_15516; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15518 = 10'ha7 == _T_241[9:0] ? 4'he : _GEN_15517; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15519 = 10'ha8 == _T_241[9:0] ? 4'hb : _GEN_15518; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15520 = 10'ha9 == _T_241[9:0] ? 4'hc : _GEN_15519; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15521 = 10'haa == _T_241[9:0] ? 4'hb : _GEN_15520; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15522 = 10'hab == _T_241[9:0] ? 4'hc : _GEN_15521; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15523 = 10'hac == _T_241[9:0] ? 4'hd : _GEN_15522; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15524 = 10'had == _T_241[9:0] ? 4'ha : _GEN_15523; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15525 = 10'hae == _T_241[9:0] ? 4'hd : _GEN_15524; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15526 = 10'haf == _T_241[9:0] ? 4'hd : _GEN_15525; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15527 = 10'hb0 == _T_241[9:0] ? 4'hb : _GEN_15526; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15528 = 10'hb1 == _T_241[9:0] ? 4'hc : _GEN_15527; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15529 = 10'hb2 == _T_241[9:0] ? 4'he : _GEN_15528; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15530 = 10'hb3 == _T_241[9:0] ? 4'hb : _GEN_15529; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15531 = 10'hb4 == _T_241[9:0] ? 4'hc : _GEN_15530; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15532 = 10'hb5 == _T_241[9:0] ? 4'hd : _GEN_15531; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15533 = 10'hb6 == _T_241[9:0] ? 4'hd : _GEN_15532; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15534 = 10'hb7 == _T_241[9:0] ? 4'hc : _GEN_15533; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15535 = 10'hb8 == _T_241[9:0] ? 4'he : _GEN_15534; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15536 = 10'hb9 == _T_241[9:0] ? 4'he : _GEN_15535; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15537 = 10'hba == _T_241[9:0] ? 4'he : _GEN_15536; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15538 = 10'hbb == _T_241[9:0] ? 4'he : _GEN_15537; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15539 = 10'hbc == _T_241[9:0] ? 4'he : _GEN_15538; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15540 = 10'hbd == _T_241[9:0] ? 4'he : _GEN_15539; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15541 = 10'hbe == _T_241[9:0] ? 4'he : _GEN_15540; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15542 = 10'hbf == _T_241[9:0] ? 4'he : _GEN_15541; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15543 = 10'hc0 == _T_241[9:0] ? 4'he : _GEN_15542; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15544 = 10'hc1 == _T_241[9:0] ? 4'he : _GEN_15543; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15545 = 10'hc2 == _T_241[9:0] ? 4'he : _GEN_15544; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15546 = 10'hc3 == _T_241[9:0] ? 4'he : _GEN_15545; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15547 = 10'hc4 == _T_241[9:0] ? 4'he : _GEN_15546; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15548 = 10'hc5 == _T_241[9:0] ? 4'he : _GEN_15547; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15549 = 10'hc6 == _T_241[9:0] ? 4'he : _GEN_15548; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15550 = 10'hc7 == _T_241[9:0] ? 4'hd : _GEN_15549; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15551 = 10'hc8 == _T_241[9:0] ? 4'hb : _GEN_15550; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15552 = 10'hc9 == _T_241[9:0] ? 4'hc : _GEN_15551; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15553 = 10'hca == _T_241[9:0] ? 4'he : _GEN_15552; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15554 = 10'hcb == _T_241[9:0] ? 4'he : _GEN_15553; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15555 = 10'hcc == _T_241[9:0] ? 4'he : _GEN_15554; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15556 = 10'hcd == _T_241[9:0] ? 4'he : _GEN_15555; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15557 = 10'hce == _T_241[9:0] ? 4'hd : _GEN_15556; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15558 = 10'hcf == _T_241[9:0] ? 4'hb : _GEN_15557; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15559 = 10'hd0 == _T_241[9:0] ? 4'hc : _GEN_15558; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15560 = 10'hd1 == _T_241[9:0] ? 4'hc : _GEN_15559; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15561 = 10'hd2 == _T_241[9:0] ? 4'hb : _GEN_15560; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15562 = 10'hd3 == _T_241[9:0] ? 4'hd : _GEN_15561; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15563 = 10'hd4 == _T_241[9:0] ? 4'hd : _GEN_15562; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15564 = 10'hd5 == _T_241[9:0] ? 4'hd : _GEN_15563; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15565 = 10'hd6 == _T_241[9:0] ? 4'hd : _GEN_15564; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15566 = 10'hd7 == _T_241[9:0] ? 4'hc : _GEN_15565; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15567 = 10'hd8 == _T_241[9:0] ? 4'hc : _GEN_15566; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15568 = 10'hd9 == _T_241[9:0] ? 4'hc : _GEN_15567; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15569 = 10'hda == _T_241[9:0] ? 4'hd : _GEN_15568; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15570 = 10'hdb == _T_241[9:0] ? 4'hc : _GEN_15569; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15571 = 10'hdc == _T_241[9:0] ? 4'h9 : _GEN_15570; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15572 = 10'hdd == _T_241[9:0] ? 4'he : _GEN_15571; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15573 = 10'hde == _T_241[9:0] ? 4'he : _GEN_15572; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15574 = 10'hdf == _T_241[9:0] ? 4'he : _GEN_15573; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15575 = 10'he0 == _T_241[9:0] ? 4'he : _GEN_15574; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15576 = 10'he1 == _T_241[9:0] ? 4'he : _GEN_15575; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15577 = 10'he2 == _T_241[9:0] ? 4'he : _GEN_15576; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15578 = 10'he3 == _T_241[9:0] ? 4'h9 : _GEN_15577; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15579 = 10'he4 == _T_241[9:0] ? 4'he : _GEN_15578; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15580 = 10'he5 == _T_241[9:0] ? 4'he : _GEN_15579; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15581 = 10'he6 == _T_241[9:0] ? 4'he : _GEN_15580; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15582 = 10'he7 == _T_241[9:0] ? 4'he : _GEN_15581; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15583 = 10'he8 == _T_241[9:0] ? 4'he : _GEN_15582; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15584 = 10'he9 == _T_241[9:0] ? 4'he : _GEN_15583; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15585 = 10'hea == _T_241[9:0] ? 4'he : _GEN_15584; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15586 = 10'heb == _T_241[9:0] ? 4'hc : _GEN_15585; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15587 = 10'hec == _T_241[9:0] ? 4'h7 : _GEN_15586; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15588 = 10'hed == _T_241[9:0] ? 4'h1 : _GEN_15587; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15589 = 10'hee == _T_241[9:0] ? 4'h0 : _GEN_15588; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15590 = 10'hef == _T_241[9:0] ? 4'h0 : _GEN_15589; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15591 = 10'hf0 == _T_241[9:0] ? 4'h2 : _GEN_15590; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15592 = 10'hf1 == _T_241[9:0] ? 4'h9 : _GEN_15591; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15593 = 10'hf2 == _T_241[9:0] ? 4'he : _GEN_15592; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15594 = 10'hf3 == _T_241[9:0] ? 4'he : _GEN_15593; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15595 = 10'hf4 == _T_241[9:0] ? 4'he : _GEN_15594; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15596 = 10'hf5 == _T_241[9:0] ? 4'hc : _GEN_15595; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15597 = 10'hf6 == _T_241[9:0] ? 4'hc : _GEN_15596; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15598 = 10'hf7 == _T_241[9:0] ? 4'hd : _GEN_15597; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15599 = 10'hf8 == _T_241[9:0] ? 4'hd : _GEN_15598; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15600 = 10'hf9 == _T_241[9:0] ? 4'hd : _GEN_15599; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15601 = 10'hfa == _T_241[9:0] ? 4'hd : _GEN_15600; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15602 = 10'hfb == _T_241[9:0] ? 4'hd : _GEN_15601; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15603 = 10'hfc == _T_241[9:0] ? 4'hd : _GEN_15602; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15604 = 10'hfd == _T_241[9:0] ? 4'hd : _GEN_15603; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15605 = 10'hfe == _T_241[9:0] ? 4'hd : _GEN_15604; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15606 = 10'hff == _T_241[9:0] ? 4'hd : _GEN_15605; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15607 = 10'h100 == _T_241[9:0] ? 4'hd : _GEN_15606; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15608 = 10'h101 == _T_241[9:0] ? 4'h9 : _GEN_15607; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15609 = 10'h102 == _T_241[9:0] ? 4'h9 : _GEN_15608; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15610 = 10'h103 == _T_241[9:0] ? 4'he : _GEN_15609; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15611 = 10'h104 == _T_241[9:0] ? 4'he : _GEN_15610; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15612 = 10'h105 == _T_241[9:0] ? 4'he : _GEN_15611; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15613 = 10'h106 == _T_241[9:0] ? 4'he : _GEN_15612; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15614 = 10'h107 == _T_241[9:0] ? 4'he : _GEN_15613; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15615 = 10'h108 == _T_241[9:0] ? 4'he : _GEN_15614; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15616 = 10'h109 == _T_241[9:0] ? 4'h6 : _GEN_15615; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15617 = 10'h10a == _T_241[9:0] ? 4'he : _GEN_15616; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15618 = 10'h10b == _T_241[9:0] ? 4'he : _GEN_15617; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15619 = 10'h10c == _T_241[9:0] ? 4'he : _GEN_15618; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15620 = 10'h10d == _T_241[9:0] ? 4'he : _GEN_15619; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15621 = 10'h10e == _T_241[9:0] ? 4'he : _GEN_15620; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15622 = 10'h10f == _T_241[9:0] ? 4'ha : _GEN_15621; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15623 = 10'h110 == _T_241[9:0] ? 4'hd : _GEN_15622; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15624 = 10'h111 == _T_241[9:0] ? 4'h4 : _GEN_15623; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15625 = 10'h112 == _T_241[9:0] ? 4'h7 : _GEN_15624; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15626 = 10'h113 == _T_241[9:0] ? 4'h0 : _GEN_15625; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15627 = 10'h114 == _T_241[9:0] ? 4'h0 : _GEN_15626; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15628 = 10'h115 == _T_241[9:0] ? 4'h0 : _GEN_15627; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15629 = 10'h116 == _T_241[9:0] ? 4'h0 : _GEN_15628; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15630 = 10'h117 == _T_241[9:0] ? 4'h0 : _GEN_15629; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15631 = 10'h118 == _T_241[9:0] ? 4'ha : _GEN_15630; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15632 = 10'h119 == _T_241[9:0] ? 4'he : _GEN_15631; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15633 = 10'h11a == _T_241[9:0] ? 4'he : _GEN_15632; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15634 = 10'h11b == _T_241[9:0] ? 4'he : _GEN_15633; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15635 = 10'h11c == _T_241[9:0] ? 4'hb : _GEN_15634; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15636 = 10'h11d == _T_241[9:0] ? 4'hc : _GEN_15635; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15637 = 10'h11e == _T_241[9:0] ? 4'hd : _GEN_15636; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15638 = 10'h11f == _T_241[9:0] ? 4'hb : _GEN_15637; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15639 = 10'h120 == _T_241[9:0] ? 4'ha : _GEN_15638; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15640 = 10'h121 == _T_241[9:0] ? 4'hc : _GEN_15639; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15641 = 10'h122 == _T_241[9:0] ? 4'ha : _GEN_15640; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15642 = 10'h123 == _T_241[9:0] ? 4'ha : _GEN_15641; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15643 = 10'h124 == _T_241[9:0] ? 4'hd : _GEN_15642; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15644 = 10'h125 == _T_241[9:0] ? 4'hd : _GEN_15643; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15645 = 10'h126 == _T_241[9:0] ? 4'hb : _GEN_15644; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15646 = 10'h127 == _T_241[9:0] ? 4'h9 : _GEN_15645; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15647 = 10'h128 == _T_241[9:0] ? 4'h7 : _GEN_15646; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15648 = 10'h129 == _T_241[9:0] ? 4'hd : _GEN_15647; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15649 = 10'h12a == _T_241[9:0] ? 4'hc : _GEN_15648; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15650 = 10'h12b == _T_241[9:0] ? 4'hb : _GEN_15649; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15651 = 10'h12c == _T_241[9:0] ? 4'hc : _GEN_15650; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15652 = 10'h12d == _T_241[9:0] ? 4'hb : _GEN_15651; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15653 = 10'h12e == _T_241[9:0] ? 4'ha : _GEN_15652; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15654 = 10'h12f == _T_241[9:0] ? 4'h6 : _GEN_15653; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15655 = 10'h130 == _T_241[9:0] ? 4'he : _GEN_15654; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15656 = 10'h131 == _T_241[9:0] ? 4'hc : _GEN_15655; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15657 = 10'h132 == _T_241[9:0] ? 4'ha : _GEN_15656; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15658 = 10'h133 == _T_241[9:0] ? 4'h9 : _GEN_15657; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15659 = 10'h134 == _T_241[9:0] ? 4'hb : _GEN_15658; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15660 = 10'h135 == _T_241[9:0] ? 4'h8 : _GEN_15659; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15661 = 10'h136 == _T_241[9:0] ? 4'h8 : _GEN_15660; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15662 = 10'h137 == _T_241[9:0] ? 4'h4 : _GEN_15661; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15663 = 10'h138 == _T_241[9:0] ? 4'h7 : _GEN_15662; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15664 = 10'h139 == _T_241[9:0] ? 4'h0 : _GEN_15663; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15665 = 10'h13a == _T_241[9:0] ? 4'h0 : _GEN_15664; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15666 = 10'h13b == _T_241[9:0] ? 4'h0 : _GEN_15665; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15667 = 10'h13c == _T_241[9:0] ? 4'h0 : _GEN_15666; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15668 = 10'h13d == _T_241[9:0] ? 4'h0 : _GEN_15667; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15669 = 10'h13e == _T_241[9:0] ? 4'h4 : _GEN_15668; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15670 = 10'h13f == _T_241[9:0] ? 4'hc : _GEN_15669; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15671 = 10'h140 == _T_241[9:0] ? 4'he : _GEN_15670; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15672 = 10'h141 == _T_241[9:0] ? 4'he : _GEN_15671; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15673 = 10'h142 == _T_241[9:0] ? 4'he : _GEN_15672; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15674 = 10'h143 == _T_241[9:0] ? 4'hc : _GEN_15673; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15675 = 10'h144 == _T_241[9:0] ? 4'hd : _GEN_15674; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15676 = 10'h145 == _T_241[9:0] ? 4'hb : _GEN_15675; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15677 = 10'h146 == _T_241[9:0] ? 4'hb : _GEN_15676; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15678 = 10'h147 == _T_241[9:0] ? 4'ha : _GEN_15677; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15679 = 10'h148 == _T_241[9:0] ? 4'ha : _GEN_15678; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15680 = 10'h149 == _T_241[9:0] ? 4'hc : _GEN_15679; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15681 = 10'h14a == _T_241[9:0] ? 4'hd : _GEN_15680; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15682 = 10'h14b == _T_241[9:0] ? 4'hc : _GEN_15681; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15683 = 10'h14c == _T_241[9:0] ? 4'hd : _GEN_15682; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15684 = 10'h14d == _T_241[9:0] ? 4'h9 : _GEN_15683; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15685 = 10'h14e == _T_241[9:0] ? 4'h7 : _GEN_15684; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15686 = 10'h14f == _T_241[9:0] ? 4'ha : _GEN_15685; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15687 = 10'h150 == _T_241[9:0] ? 4'ha : _GEN_15686; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15688 = 10'h151 == _T_241[9:0] ? 4'hb : _GEN_15687; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15689 = 10'h152 == _T_241[9:0] ? 4'hb : _GEN_15688; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15690 = 10'h153 == _T_241[9:0] ? 4'hc : _GEN_15689; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15691 = 10'h154 == _T_241[9:0] ? 4'hb : _GEN_15690; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15692 = 10'h155 == _T_241[9:0] ? 4'h6 : _GEN_15691; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15693 = 10'h156 == _T_241[9:0] ? 4'hb : _GEN_15692; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15694 = 10'h157 == _T_241[9:0] ? 4'h7 : _GEN_15693; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15695 = 10'h158 == _T_241[9:0] ? 4'h7 : _GEN_15694; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15696 = 10'h159 == _T_241[9:0] ? 4'h7 : _GEN_15695; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15697 = 10'h15a == _T_241[9:0] ? 4'h7 : _GEN_15696; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15698 = 10'h15b == _T_241[9:0] ? 4'h7 : _GEN_15697; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15699 = 10'h15c == _T_241[9:0] ? 4'h7 : _GEN_15698; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15700 = 10'h15d == _T_241[9:0] ? 4'h6 : _GEN_15699; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15701 = 10'h15e == _T_241[9:0] ? 4'h7 : _GEN_15700; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15702 = 10'h15f == _T_241[9:0] ? 4'h0 : _GEN_15701; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15703 = 10'h160 == _T_241[9:0] ? 4'h0 : _GEN_15702; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15704 = 10'h161 == _T_241[9:0] ? 4'h0 : _GEN_15703; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15705 = 10'h162 == _T_241[9:0] ? 4'h0 : _GEN_15704; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15706 = 10'h163 == _T_241[9:0] ? 4'h2 : _GEN_15705; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15707 = 10'h164 == _T_241[9:0] ? 4'h4 : _GEN_15706; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15708 = 10'h165 == _T_241[9:0] ? 4'hb : _GEN_15707; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15709 = 10'h166 == _T_241[9:0] ? 4'hb : _GEN_15708; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15710 = 10'h167 == _T_241[9:0] ? 4'he : _GEN_15709; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15711 = 10'h168 == _T_241[9:0] ? 4'he : _GEN_15710; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15712 = 10'h169 == _T_241[9:0] ? 4'hc : _GEN_15711; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15713 = 10'h16a == _T_241[9:0] ? 4'hd : _GEN_15712; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15714 = 10'h16b == _T_241[9:0] ? 4'hd : _GEN_15713; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15715 = 10'h16c == _T_241[9:0] ? 4'ha : _GEN_15714; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15716 = 10'h16d == _T_241[9:0] ? 4'ha : _GEN_15715; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15717 = 10'h16e == _T_241[9:0] ? 4'ha : _GEN_15716; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15718 = 10'h16f == _T_241[9:0] ? 4'hd : _GEN_15717; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15719 = 10'h170 == _T_241[9:0] ? 4'hd : _GEN_15718; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15720 = 10'h171 == _T_241[9:0] ? 4'hd : _GEN_15719; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15721 = 10'h172 == _T_241[9:0] ? 4'he : _GEN_15720; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15722 = 10'h173 == _T_241[9:0] ? 4'h8 : _GEN_15721; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15723 = 10'h174 == _T_241[9:0] ? 4'h5 : _GEN_15722; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15724 = 10'h175 == _T_241[9:0] ? 4'h6 : _GEN_15723; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15725 = 10'h176 == _T_241[9:0] ? 4'h6 : _GEN_15724; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15726 = 10'h177 == _T_241[9:0] ? 4'h6 : _GEN_15725; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15727 = 10'h178 == _T_241[9:0] ? 4'h7 : _GEN_15726; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15728 = 10'h179 == _T_241[9:0] ? 4'h9 : _GEN_15727; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15729 = 10'h17a == _T_241[9:0] ? 4'h9 : _GEN_15728; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15730 = 10'h17b == _T_241[9:0] ? 4'h6 : _GEN_15729; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15731 = 10'h17c == _T_241[9:0] ? 4'h7 : _GEN_15730; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15732 = 10'h17d == _T_241[9:0] ? 4'h7 : _GEN_15731; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15733 = 10'h17e == _T_241[9:0] ? 4'h7 : _GEN_15732; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15734 = 10'h17f == _T_241[9:0] ? 4'h7 : _GEN_15733; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15735 = 10'h180 == _T_241[9:0] ? 4'h7 : _GEN_15734; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15736 = 10'h181 == _T_241[9:0] ? 4'h7 : _GEN_15735; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15737 = 10'h182 == _T_241[9:0] ? 4'h8 : _GEN_15736; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15738 = 10'h183 == _T_241[9:0] ? 4'h8 : _GEN_15737; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15739 = 10'h184 == _T_241[9:0] ? 4'h8 : _GEN_15738; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15740 = 10'h185 == _T_241[9:0] ? 4'h7 : _GEN_15739; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15741 = 10'h186 == _T_241[9:0] ? 4'h1 : _GEN_15740; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15742 = 10'h187 == _T_241[9:0] ? 4'h0 : _GEN_15741; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15743 = 10'h188 == _T_241[9:0] ? 4'h0 : _GEN_15742; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15744 = 10'h189 == _T_241[9:0] ? 4'h4 : _GEN_15743; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15745 = 10'h18a == _T_241[9:0] ? 4'h4 : _GEN_15744; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15746 = 10'h18b == _T_241[9:0] ? 4'hb : _GEN_15745; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15747 = 10'h18c == _T_241[9:0] ? 4'hb : _GEN_15746; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15748 = 10'h18d == _T_241[9:0] ? 4'hc : _GEN_15747; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15749 = 10'h18e == _T_241[9:0] ? 4'he : _GEN_15748; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15750 = 10'h18f == _T_241[9:0] ? 4'hb : _GEN_15749; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15751 = 10'h190 == _T_241[9:0] ? 4'hd : _GEN_15750; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15752 = 10'h191 == _T_241[9:0] ? 4'hc : _GEN_15751; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15753 = 10'h192 == _T_241[9:0] ? 4'h9 : _GEN_15752; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15754 = 10'h193 == _T_241[9:0] ? 4'ha : _GEN_15753; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15755 = 10'h194 == _T_241[9:0] ? 4'h9 : _GEN_15754; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15756 = 10'h195 == _T_241[9:0] ? 4'hd : _GEN_15755; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15757 = 10'h196 == _T_241[9:0] ? 4'hd : _GEN_15756; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15758 = 10'h197 == _T_241[9:0] ? 4'hb : _GEN_15757; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15759 = 10'h198 == _T_241[9:0] ? 4'he : _GEN_15758; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15760 = 10'h199 == _T_241[9:0] ? 4'h5 : _GEN_15759; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15761 = 10'h19a == _T_241[9:0] ? 4'h1 : _GEN_15760; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15762 = 10'h19b == _T_241[9:0] ? 4'h3 : _GEN_15761; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15763 = 10'h19c == _T_241[9:0] ? 4'h6 : _GEN_15762; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15764 = 10'h19d == _T_241[9:0] ? 4'h4 : _GEN_15763; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15765 = 10'h19e == _T_241[9:0] ? 4'h1 : _GEN_15764; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15766 = 10'h19f == _T_241[9:0] ? 4'h3 : _GEN_15765; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15767 = 10'h1a0 == _T_241[9:0] ? 4'h6 : _GEN_15766; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15768 = 10'h1a1 == _T_241[9:0] ? 4'h6 : _GEN_15767; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15769 = 10'h1a2 == _T_241[9:0] ? 4'h7 : _GEN_15768; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15770 = 10'h1a3 == _T_241[9:0] ? 4'h7 : _GEN_15769; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15771 = 10'h1a4 == _T_241[9:0] ? 4'h7 : _GEN_15770; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15772 = 10'h1a5 == _T_241[9:0] ? 4'h7 : _GEN_15771; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15773 = 10'h1a6 == _T_241[9:0] ? 4'h7 : _GEN_15772; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15774 = 10'h1a7 == _T_241[9:0] ? 4'h7 : _GEN_15773; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15775 = 10'h1a8 == _T_241[9:0] ? 4'h8 : _GEN_15774; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15776 = 10'h1a9 == _T_241[9:0] ? 4'h8 : _GEN_15775; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15777 = 10'h1aa == _T_241[9:0] ? 4'h7 : _GEN_15776; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15778 = 10'h1ab == _T_241[9:0] ? 4'h8 : _GEN_15777; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15779 = 10'h1ac == _T_241[9:0] ? 4'h8 : _GEN_15778; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15780 = 10'h1ad == _T_241[9:0] ? 4'h3 : _GEN_15779; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15781 = 10'h1ae == _T_241[9:0] ? 4'h2 : _GEN_15780; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15782 = 10'h1af == _T_241[9:0] ? 4'h8 : _GEN_15781; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15783 = 10'h1b0 == _T_241[9:0] ? 4'h6 : _GEN_15782; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15784 = 10'h1b1 == _T_241[9:0] ? 4'hb : _GEN_15783; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15785 = 10'h1b2 == _T_241[9:0] ? 4'hb : _GEN_15784; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15786 = 10'h1b3 == _T_241[9:0] ? 4'ha : _GEN_15785; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15787 = 10'h1b4 == _T_241[9:0] ? 4'he : _GEN_15786; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15788 = 10'h1b5 == _T_241[9:0] ? 4'hb : _GEN_15787; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15789 = 10'h1b6 == _T_241[9:0] ? 4'hc : _GEN_15788; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15790 = 10'h1b7 == _T_241[9:0] ? 4'ha : _GEN_15789; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15791 = 10'h1b8 == _T_241[9:0] ? 4'h9 : _GEN_15790; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15792 = 10'h1b9 == _T_241[9:0] ? 4'h9 : _GEN_15791; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15793 = 10'h1ba == _T_241[9:0] ? 4'h9 : _GEN_15792; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15794 = 10'h1bb == _T_241[9:0] ? 4'hb : _GEN_15793; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15795 = 10'h1bc == _T_241[9:0] ? 4'hd : _GEN_15794; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15796 = 10'h1bd == _T_241[9:0] ? 4'hd : _GEN_15795; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15797 = 10'h1be == _T_241[9:0] ? 4'he : _GEN_15796; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15798 = 10'h1bf == _T_241[9:0] ? 4'h7 : _GEN_15797; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15799 = 10'h1c0 == _T_241[9:0] ? 4'h6 : _GEN_15798; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15800 = 10'h1c1 == _T_241[9:0] ? 4'h6 : _GEN_15799; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15801 = 10'h1c2 == _T_241[9:0] ? 4'h5 : _GEN_15800; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15802 = 10'h1c3 == _T_241[9:0] ? 4'h5 : _GEN_15801; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15803 = 10'h1c4 == _T_241[9:0] ? 4'h4 : _GEN_15802; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15804 = 10'h1c5 == _T_241[9:0] ? 4'h5 : _GEN_15803; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15805 = 10'h1c6 == _T_241[9:0] ? 4'h6 : _GEN_15804; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15806 = 10'h1c7 == _T_241[9:0] ? 4'h6 : _GEN_15805; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15807 = 10'h1c8 == _T_241[9:0] ? 4'h7 : _GEN_15806; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15808 = 10'h1c9 == _T_241[9:0] ? 4'h7 : _GEN_15807; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15809 = 10'h1ca == _T_241[9:0] ? 4'h7 : _GEN_15808; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15810 = 10'h1cb == _T_241[9:0] ? 4'h7 : _GEN_15809; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15811 = 10'h1cc == _T_241[9:0] ? 4'h7 : _GEN_15810; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15812 = 10'h1cd == _T_241[9:0] ? 4'h8 : _GEN_15811; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15813 = 10'h1ce == _T_241[9:0] ? 4'h8 : _GEN_15812; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15814 = 10'h1cf == _T_241[9:0] ? 4'h8 : _GEN_15813; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15815 = 10'h1d0 == _T_241[9:0] ? 4'h5 : _GEN_15814; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15816 = 10'h1d1 == _T_241[9:0] ? 4'h8 : _GEN_15815; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15817 = 10'h1d2 == _T_241[9:0] ? 4'h8 : _GEN_15816; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15818 = 10'h1d3 == _T_241[9:0] ? 4'h8 : _GEN_15817; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15819 = 10'h1d4 == _T_241[9:0] ? 4'h8 : _GEN_15818; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15820 = 10'h1d5 == _T_241[9:0] ? 4'h7 : _GEN_15819; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15821 = 10'h1d6 == _T_241[9:0] ? 4'h9 : _GEN_15820; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15822 = 10'h1d7 == _T_241[9:0] ? 4'hb : _GEN_15821; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15823 = 10'h1d8 == _T_241[9:0] ? 4'hb : _GEN_15822; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15824 = 10'h1d9 == _T_241[9:0] ? 4'hb : _GEN_15823; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15825 = 10'h1da == _T_241[9:0] ? 4'ha : _GEN_15824; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15826 = 10'h1db == _T_241[9:0] ? 4'hc : _GEN_15825; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15827 = 10'h1dc == _T_241[9:0] ? 4'hb : _GEN_15826; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15828 = 10'h1dd == _T_241[9:0] ? 4'h5 : _GEN_15827; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15829 = 10'h1de == _T_241[9:0] ? 4'h9 : _GEN_15828; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15830 = 10'h1df == _T_241[9:0] ? 4'h9 : _GEN_15829; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15831 = 10'h1e0 == _T_241[9:0] ? 4'h9 : _GEN_15830; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15832 = 10'h1e1 == _T_241[9:0] ? 4'h7 : _GEN_15831; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15833 = 10'h1e2 == _T_241[9:0] ? 4'hc : _GEN_15832; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15834 = 10'h1e3 == _T_241[9:0] ? 4'hc : _GEN_15833; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15835 = 10'h1e4 == _T_241[9:0] ? 4'hd : _GEN_15834; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15836 = 10'h1e5 == _T_241[9:0] ? 4'h7 : _GEN_15835; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15837 = 10'h1e6 == _T_241[9:0] ? 4'h6 : _GEN_15836; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15838 = 10'h1e7 == _T_241[9:0] ? 4'h6 : _GEN_15837; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15839 = 10'h1e8 == _T_241[9:0] ? 4'h6 : _GEN_15838; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15840 = 10'h1e9 == _T_241[9:0] ? 4'h6 : _GEN_15839; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15841 = 10'h1ea == _T_241[9:0] ? 4'h6 : _GEN_15840; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15842 = 10'h1eb == _T_241[9:0] ? 4'h6 : _GEN_15841; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15843 = 10'h1ec == _T_241[9:0] ? 4'h6 : _GEN_15842; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15844 = 10'h1ed == _T_241[9:0] ? 4'h8 : _GEN_15843; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15845 = 10'h1ee == _T_241[9:0] ? 4'h7 : _GEN_15844; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15846 = 10'h1ef == _T_241[9:0] ? 4'h7 : _GEN_15845; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15847 = 10'h1f0 == _T_241[9:0] ? 4'h7 : _GEN_15846; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15848 = 10'h1f1 == _T_241[9:0] ? 4'h7 : _GEN_15847; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15849 = 10'h1f2 == _T_241[9:0] ? 4'h7 : _GEN_15848; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15850 = 10'h1f3 == _T_241[9:0] ? 4'h8 : _GEN_15849; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15851 = 10'h1f4 == _T_241[9:0] ? 4'h8 : _GEN_15850; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15852 = 10'h1f5 == _T_241[9:0] ? 4'h8 : _GEN_15851; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15853 = 10'h1f6 == _T_241[9:0] ? 4'ha : _GEN_15852; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15854 = 10'h1f7 == _T_241[9:0] ? 4'h8 : _GEN_15853; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15855 = 10'h1f8 == _T_241[9:0] ? 4'h8 : _GEN_15854; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15856 = 10'h1f9 == _T_241[9:0] ? 4'h9 : _GEN_15855; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15857 = 10'h1fa == _T_241[9:0] ? 4'h9 : _GEN_15856; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15858 = 10'h1fb == _T_241[9:0] ? 4'h8 : _GEN_15857; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15859 = 10'h1fc == _T_241[9:0] ? 4'hb : _GEN_15858; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15860 = 10'h1fd == _T_241[9:0] ? 4'hb : _GEN_15859; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15861 = 10'h1fe == _T_241[9:0] ? 4'hb : _GEN_15860; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15862 = 10'h1ff == _T_241[9:0] ? 4'ha : _GEN_15861; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15863 = 10'h200 == _T_241[9:0] ? 4'h3 : _GEN_15862; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15864 = 10'h201 == _T_241[9:0] ? 4'h9 : _GEN_15863; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15865 = 10'h202 == _T_241[9:0] ? 4'h5 : _GEN_15864; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15866 = 10'h203 == _T_241[9:0] ? 4'h3 : _GEN_15865; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15867 = 10'h204 == _T_241[9:0] ? 4'h4 : _GEN_15866; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15868 = 10'h205 == _T_241[9:0] ? 4'h4 : _GEN_15867; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15869 = 10'h206 == _T_241[9:0] ? 4'h4 : _GEN_15868; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15870 = 10'h207 == _T_241[9:0] ? 4'h4 : _GEN_15869; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15871 = 10'h208 == _T_241[9:0] ? 4'h8 : _GEN_15870; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15872 = 10'h209 == _T_241[9:0] ? 4'hc : _GEN_15871; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15873 = 10'h20a == _T_241[9:0] ? 4'hd : _GEN_15872; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15874 = 10'h20b == _T_241[9:0] ? 4'h7 : _GEN_15873; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15875 = 10'h20c == _T_241[9:0] ? 4'h6 : _GEN_15874; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15876 = 10'h20d == _T_241[9:0] ? 4'h6 : _GEN_15875; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15877 = 10'h20e == _T_241[9:0] ? 4'h6 : _GEN_15876; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15878 = 10'h20f == _T_241[9:0] ? 4'h5 : _GEN_15877; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15879 = 10'h210 == _T_241[9:0] ? 4'h6 : _GEN_15878; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15880 = 10'h211 == _T_241[9:0] ? 4'h6 : _GEN_15879; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15881 = 10'h212 == _T_241[9:0] ? 4'h7 : _GEN_15880; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15882 = 10'h213 == _T_241[9:0] ? 4'ha : _GEN_15881; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15883 = 10'h214 == _T_241[9:0] ? 4'h6 : _GEN_15882; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15884 = 10'h215 == _T_241[9:0] ? 4'h7 : _GEN_15883; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15885 = 10'h216 == _T_241[9:0] ? 4'h7 : _GEN_15884; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15886 = 10'h217 == _T_241[9:0] ? 4'h7 : _GEN_15885; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15887 = 10'h218 == _T_241[9:0] ? 4'h7 : _GEN_15886; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15888 = 10'h219 == _T_241[9:0] ? 4'h8 : _GEN_15887; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15889 = 10'h21a == _T_241[9:0] ? 4'h7 : _GEN_15888; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15890 = 10'h21b == _T_241[9:0] ? 4'h8 : _GEN_15889; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15891 = 10'h21c == _T_241[9:0] ? 4'hb : _GEN_15890; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15892 = 10'h21d == _T_241[9:0] ? 4'ha : _GEN_15891; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15893 = 10'h21e == _T_241[9:0] ? 4'h9 : _GEN_15892; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15894 = 10'h21f == _T_241[9:0] ? 4'h9 : _GEN_15893; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15895 = 10'h220 == _T_241[9:0] ? 4'h8 : _GEN_15894; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15896 = 10'h221 == _T_241[9:0] ? 4'h9 : _GEN_15895; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15897 = 10'h222 == _T_241[9:0] ? 4'hb : _GEN_15896; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15898 = 10'h223 == _T_241[9:0] ? 4'hb : _GEN_15897; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15899 = 10'h224 == _T_241[9:0] ? 4'hb : _GEN_15898; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15900 = 10'h225 == _T_241[9:0] ? 4'h8 : _GEN_15899; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15901 = 10'h226 == _T_241[9:0] ? 4'h1 : _GEN_15900; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15902 = 10'h227 == _T_241[9:0] ? 4'h3 : _GEN_15901; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15903 = 10'h228 == _T_241[9:0] ? 4'h3 : _GEN_15902; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15904 = 10'h229 == _T_241[9:0] ? 4'h3 : _GEN_15903; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15905 = 10'h22a == _T_241[9:0] ? 4'h3 : _GEN_15904; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15906 = 10'h22b == _T_241[9:0] ? 4'h3 : _GEN_15905; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15907 = 10'h22c == _T_241[9:0] ? 4'h3 : _GEN_15906; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15908 = 10'h22d == _T_241[9:0] ? 4'h3 : _GEN_15907; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15909 = 10'h22e == _T_241[9:0] ? 4'h3 : _GEN_15908; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15910 = 10'h22f == _T_241[9:0] ? 4'h9 : _GEN_15909; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15911 = 10'h230 == _T_241[9:0] ? 4'h6 : _GEN_15910; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15912 = 10'h231 == _T_241[9:0] ? 4'h7 : _GEN_15911; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15913 = 10'h232 == _T_241[9:0] ? 4'h6 : _GEN_15912; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15914 = 10'h233 == _T_241[9:0] ? 4'h7 : _GEN_15913; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15915 = 10'h234 == _T_241[9:0] ? 4'h7 : _GEN_15914; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15916 = 10'h235 == _T_241[9:0] ? 4'h6 : _GEN_15915; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15917 = 10'h236 == _T_241[9:0] ? 4'h6 : _GEN_15916; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15918 = 10'h237 == _T_241[9:0] ? 4'h6 : _GEN_15917; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15919 = 10'h238 == _T_241[9:0] ? 4'h6 : _GEN_15918; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15920 = 10'h239 == _T_241[9:0] ? 4'h8 : _GEN_15919; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15921 = 10'h23a == _T_241[9:0] ? 4'h6 : _GEN_15920; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15922 = 10'h23b == _T_241[9:0] ? 4'h7 : _GEN_15921; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15923 = 10'h23c == _T_241[9:0] ? 4'h7 : _GEN_15922; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15924 = 10'h23d == _T_241[9:0] ? 4'h7 : _GEN_15923; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15925 = 10'h23e == _T_241[9:0] ? 4'h7 : _GEN_15924; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15926 = 10'h23f == _T_241[9:0] ? 4'h7 : _GEN_15925; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15927 = 10'h240 == _T_241[9:0] ? 4'h7 : _GEN_15926; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15928 = 10'h241 == _T_241[9:0] ? 4'h8 : _GEN_15927; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15929 = 10'h242 == _T_241[9:0] ? 4'hb : _GEN_15928; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15930 = 10'h243 == _T_241[9:0] ? 4'hb : _GEN_15929; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15931 = 10'h244 == _T_241[9:0] ? 4'hb : _GEN_15930; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15932 = 10'h245 == _T_241[9:0] ? 4'ha : _GEN_15931; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15933 = 10'h246 == _T_241[9:0] ? 4'h9 : _GEN_15932; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15934 = 10'h247 == _T_241[9:0] ? 4'ha : _GEN_15933; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15935 = 10'h248 == _T_241[9:0] ? 4'hb : _GEN_15934; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15936 = 10'h249 == _T_241[9:0] ? 4'hb : _GEN_15935; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15937 = 10'h24a == _T_241[9:0] ? 4'ha : _GEN_15936; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15938 = 10'h24b == _T_241[9:0] ? 4'h2 : _GEN_15937; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15939 = 10'h24c == _T_241[9:0] ? 4'h0 : _GEN_15938; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15940 = 10'h24d == _T_241[9:0] ? 4'h2 : _GEN_15939; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15941 = 10'h24e == _T_241[9:0] ? 4'h3 : _GEN_15940; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15942 = 10'h24f == _T_241[9:0] ? 4'h3 : _GEN_15941; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15943 = 10'h250 == _T_241[9:0] ? 4'h3 : _GEN_15942; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15944 = 10'h251 == _T_241[9:0] ? 4'h3 : _GEN_15943; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15945 = 10'h252 == _T_241[9:0] ? 4'h3 : _GEN_15944; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15946 = 10'h253 == _T_241[9:0] ? 4'h3 : _GEN_15945; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15947 = 10'h254 == _T_241[9:0] ? 4'h3 : _GEN_15946; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15948 = 10'h255 == _T_241[9:0] ? 4'h5 : _GEN_15947; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15949 = 10'h256 == _T_241[9:0] ? 4'h6 : _GEN_15948; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15950 = 10'h257 == _T_241[9:0] ? 4'h8 : _GEN_15949; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15951 = 10'h258 == _T_241[9:0] ? 4'h5 : _GEN_15950; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15952 = 10'h259 == _T_241[9:0] ? 4'h6 : _GEN_15951; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15953 = 10'h25a == _T_241[9:0] ? 4'h6 : _GEN_15952; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15954 = 10'h25b == _T_241[9:0] ? 4'h5 : _GEN_15953; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15955 = 10'h25c == _T_241[9:0] ? 4'h6 : _GEN_15954; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15956 = 10'h25d == _T_241[9:0] ? 4'h6 : _GEN_15955; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15957 = 10'h25e == _T_241[9:0] ? 4'h9 : _GEN_15956; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15958 = 10'h25f == _T_241[9:0] ? 4'hc : _GEN_15957; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15959 = 10'h260 == _T_241[9:0] ? 4'h7 : _GEN_15958; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15960 = 10'h261 == _T_241[9:0] ? 4'h9 : _GEN_15959; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15961 = 10'h262 == _T_241[9:0] ? 4'ha : _GEN_15960; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15962 = 10'h263 == _T_241[9:0] ? 4'h8 : _GEN_15961; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15963 = 10'h264 == _T_241[9:0] ? 4'ha : _GEN_15962; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15964 = 10'h265 == _T_241[9:0] ? 4'h9 : _GEN_15963; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15965 = 10'h266 == _T_241[9:0] ? 4'h8 : _GEN_15964; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15966 = 10'h267 == _T_241[9:0] ? 4'h8 : _GEN_15965; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15967 = 10'h268 == _T_241[9:0] ? 4'ha : _GEN_15966; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15968 = 10'h269 == _T_241[9:0] ? 4'ha : _GEN_15967; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15969 = 10'h26a == _T_241[9:0] ? 4'hb : _GEN_15968; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15970 = 10'h26b == _T_241[9:0] ? 4'hb : _GEN_15969; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15971 = 10'h26c == _T_241[9:0] ? 4'hb : _GEN_15970; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15972 = 10'h26d == _T_241[9:0] ? 4'hb : _GEN_15971; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15973 = 10'h26e == _T_241[9:0] ? 4'hb : _GEN_15972; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15974 = 10'h26f == _T_241[9:0] ? 4'ha : _GEN_15973; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15975 = 10'h270 == _T_241[9:0] ? 4'h3 : _GEN_15974; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15976 = 10'h271 == _T_241[9:0] ? 4'h0 : _GEN_15975; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15977 = 10'h272 == _T_241[9:0] ? 4'h0 : _GEN_15976; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15978 = 10'h273 == _T_241[9:0] ? 4'h2 : _GEN_15977; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15979 = 10'h274 == _T_241[9:0] ? 4'h3 : _GEN_15978; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15980 = 10'h275 == _T_241[9:0] ? 4'h3 : _GEN_15979; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15981 = 10'h276 == _T_241[9:0] ? 4'h3 : _GEN_15980; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15982 = 10'h277 == _T_241[9:0] ? 4'h3 : _GEN_15981; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15983 = 10'h278 == _T_241[9:0] ? 4'h3 : _GEN_15982; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15984 = 10'h279 == _T_241[9:0] ? 4'h3 : _GEN_15983; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15985 = 10'h27a == _T_241[9:0] ? 4'h3 : _GEN_15984; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15986 = 10'h27b == _T_241[9:0] ? 4'h6 : _GEN_15985; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15987 = 10'h27c == _T_241[9:0] ? 4'h7 : _GEN_15986; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15988 = 10'h27d == _T_241[9:0] ? 4'h7 : _GEN_15987; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15989 = 10'h27e == _T_241[9:0] ? 4'h4 : _GEN_15988; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15990 = 10'h27f == _T_241[9:0] ? 4'h6 : _GEN_15989; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15991 = 10'h280 == _T_241[9:0] ? 4'h6 : _GEN_15990; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15992 = 10'h281 == _T_241[9:0] ? 4'h6 : _GEN_15991; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15993 = 10'h282 == _T_241[9:0] ? 4'h6 : _GEN_15992; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15994 = 10'h283 == _T_241[9:0] ? 4'ha : _GEN_15993; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15995 = 10'h284 == _T_241[9:0] ? 4'hc : _GEN_15994; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15996 = 10'h285 == _T_241[9:0] ? 4'hc : _GEN_15995; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15997 = 10'h286 == _T_241[9:0] ? 4'h8 : _GEN_15996; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15998 = 10'h287 == _T_241[9:0] ? 4'ha : _GEN_15997; // @[Filter.scala 230:102]
  wire [3:0] _GEN_15999 = 10'h288 == _T_241[9:0] ? 4'ha : _GEN_15998; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16000 = 10'h289 == _T_241[9:0] ? 4'ha : _GEN_15999; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16001 = 10'h28a == _T_241[9:0] ? 4'hc : _GEN_16000; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16002 = 10'h28b == _T_241[9:0] ? 4'hb : _GEN_16001; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16003 = 10'h28c == _T_241[9:0] ? 4'ha : _GEN_16002; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16004 = 10'h28d == _T_241[9:0] ? 4'h7 : _GEN_16003; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16005 = 10'h28e == _T_241[9:0] ? 4'h2 : _GEN_16004; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16006 = 10'h28f == _T_241[9:0] ? 4'h5 : _GEN_16005; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16007 = 10'h290 == _T_241[9:0] ? 4'h8 : _GEN_16006; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16008 = 10'h291 == _T_241[9:0] ? 4'ha : _GEN_16007; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16009 = 10'h292 == _T_241[9:0] ? 4'ha : _GEN_16008; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16010 = 10'h293 == _T_241[9:0] ? 4'ha : _GEN_16009; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16011 = 10'h294 == _T_241[9:0] ? 4'h9 : _GEN_16010; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16012 = 10'h295 == _T_241[9:0] ? 4'h3 : _GEN_16011; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16013 = 10'h296 == _T_241[9:0] ? 4'h0 : _GEN_16012; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16014 = 10'h297 == _T_241[9:0] ? 4'h0 : _GEN_16013; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16015 = 10'h298 == _T_241[9:0] ? 4'h0 : _GEN_16014; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16016 = 10'h299 == _T_241[9:0] ? 4'h1 : _GEN_16015; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16017 = 10'h29a == _T_241[9:0] ? 4'h3 : _GEN_16016; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16018 = 10'h29b == _T_241[9:0] ? 4'h3 : _GEN_16017; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16019 = 10'h29c == _T_241[9:0] ? 4'h3 : _GEN_16018; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16020 = 10'h29d == _T_241[9:0] ? 4'h3 : _GEN_16019; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16021 = 10'h29e == _T_241[9:0] ? 4'h3 : _GEN_16020; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16022 = 10'h29f == _T_241[9:0] ? 4'h3 : _GEN_16021; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16023 = 10'h2a0 == _T_241[9:0] ? 4'h4 : _GEN_16022; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16024 = 10'h2a1 == _T_241[9:0] ? 4'h6 : _GEN_16023; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16025 = 10'h2a2 == _T_241[9:0] ? 4'h7 : _GEN_16024; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16026 = 10'h2a3 == _T_241[9:0] ? 4'h6 : _GEN_16025; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16027 = 10'h2a4 == _T_241[9:0] ? 4'h4 : _GEN_16026; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16028 = 10'h2a5 == _T_241[9:0] ? 4'h6 : _GEN_16027; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16029 = 10'h2a6 == _T_241[9:0] ? 4'h6 : _GEN_16028; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16030 = 10'h2a7 == _T_241[9:0] ? 4'h7 : _GEN_16029; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16031 = 10'h2a8 == _T_241[9:0] ? 4'ha : _GEN_16030; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16032 = 10'h2a9 == _T_241[9:0] ? 4'hb : _GEN_16031; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16033 = 10'h2aa == _T_241[9:0] ? 4'hb : _GEN_16032; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16034 = 10'h2ab == _T_241[9:0] ? 4'hb : _GEN_16033; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16035 = 10'h2ac == _T_241[9:0] ? 4'h8 : _GEN_16034; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16036 = 10'h2ad == _T_241[9:0] ? 4'hb : _GEN_16035; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16037 = 10'h2ae == _T_241[9:0] ? 4'ha : _GEN_16036; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16038 = 10'h2af == _T_241[9:0] ? 4'hb : _GEN_16037; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16039 = 10'h2b0 == _T_241[9:0] ? 4'hc : _GEN_16038; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16040 = 10'h2b1 == _T_241[9:0] ? 4'hb : _GEN_16039; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16041 = 10'h2b2 == _T_241[9:0] ? 4'ha : _GEN_16040; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16042 = 10'h2b3 == _T_241[9:0] ? 4'h6 : _GEN_16041; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16043 = 10'h2b4 == _T_241[9:0] ? 4'h0 : _GEN_16042; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16044 = 10'h2b5 == _T_241[9:0] ? 4'h0 : _GEN_16043; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16045 = 10'h2b6 == _T_241[9:0] ? 4'h0 : _GEN_16044; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16046 = 10'h2b7 == _T_241[9:0] ? 4'h1 : _GEN_16045; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16047 = 10'h2b8 == _T_241[9:0] ? 4'h5 : _GEN_16046; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16048 = 10'h2b9 == _T_241[9:0] ? 4'h9 : _GEN_16047; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16049 = 10'h2ba == _T_241[9:0] ? 4'h1 : _GEN_16048; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16050 = 10'h2bb == _T_241[9:0] ? 4'h0 : _GEN_16049; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16051 = 10'h2bc == _T_241[9:0] ? 4'h0 : _GEN_16050; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16052 = 10'h2bd == _T_241[9:0] ? 4'h0 : _GEN_16051; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16053 = 10'h2be == _T_241[9:0] ? 4'h0 : _GEN_16052; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16054 = 10'h2bf == _T_241[9:0] ? 4'h0 : _GEN_16053; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16055 = 10'h2c0 == _T_241[9:0] ? 4'h3 : _GEN_16054; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16056 = 10'h2c1 == _T_241[9:0] ? 4'h3 : _GEN_16055; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16057 = 10'h2c2 == _T_241[9:0] ? 4'h3 : _GEN_16056; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16058 = 10'h2c3 == _T_241[9:0] ? 4'h3 : _GEN_16057; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16059 = 10'h2c4 == _T_241[9:0] ? 4'h3 : _GEN_16058; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16060 = 10'h2c5 == _T_241[9:0] ? 4'h3 : _GEN_16059; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16061 = 10'h2c6 == _T_241[9:0] ? 4'h4 : _GEN_16060; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16062 = 10'h2c7 == _T_241[9:0] ? 4'h5 : _GEN_16061; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16063 = 10'h2c8 == _T_241[9:0] ? 4'h7 : _GEN_16062; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16064 = 10'h2c9 == _T_241[9:0] ? 4'h7 : _GEN_16063; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16065 = 10'h2ca == _T_241[9:0] ? 4'h4 : _GEN_16064; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16066 = 10'h2cb == _T_241[9:0] ? 4'h9 : _GEN_16065; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16067 = 10'h2cc == _T_241[9:0] ? 4'h9 : _GEN_16066; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16068 = 10'h2cd == _T_241[9:0] ? 4'hb : _GEN_16067; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16069 = 10'h2ce == _T_241[9:0] ? 4'hb : _GEN_16068; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16070 = 10'h2cf == _T_241[9:0] ? 4'hb : _GEN_16069; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16071 = 10'h2d0 == _T_241[9:0] ? 4'hb : _GEN_16070; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16072 = 10'h2d1 == _T_241[9:0] ? 4'hb : _GEN_16071; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16073 = 10'h2d2 == _T_241[9:0] ? 4'h8 : _GEN_16072; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16074 = 10'h2d3 == _T_241[9:0] ? 4'ha : _GEN_16073; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16075 = 10'h2d4 == _T_241[9:0] ? 4'hb : _GEN_16074; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16076 = 10'h2d5 == _T_241[9:0] ? 4'ha : _GEN_16075; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16077 = 10'h2d6 == _T_241[9:0] ? 4'ha : _GEN_16076; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16078 = 10'h2d7 == _T_241[9:0] ? 4'ha : _GEN_16077; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16079 = 10'h2d8 == _T_241[9:0] ? 4'ha : _GEN_16078; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16080 = 10'h2d9 == _T_241[9:0] ? 4'h7 : _GEN_16079; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16081 = 10'h2da == _T_241[9:0] ? 4'h2 : _GEN_16080; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16082 = 10'h2db == _T_241[9:0] ? 4'h0 : _GEN_16081; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16083 = 10'h2dc == _T_241[9:0] ? 4'h0 : _GEN_16082; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16084 = 10'h2dd == _T_241[9:0] ? 4'h0 : _GEN_16083; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16085 = 10'h2de == _T_241[9:0] ? 4'h0 : _GEN_16084; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16086 = 10'h2df == _T_241[9:0] ? 4'h2 : _GEN_16085; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16087 = 10'h2e0 == _T_241[9:0] ? 4'h0 : _GEN_16086; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16088 = 10'h2e1 == _T_241[9:0] ? 4'h0 : _GEN_16087; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16089 = 10'h2e2 == _T_241[9:0] ? 4'h0 : _GEN_16088; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16090 = 10'h2e3 == _T_241[9:0] ? 4'h0 : _GEN_16089; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16091 = 10'h2e4 == _T_241[9:0] ? 4'h0 : _GEN_16090; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16092 = 10'h2e5 == _T_241[9:0] ? 4'h0 : _GEN_16091; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16093 = 10'h2e6 == _T_241[9:0] ? 4'h2 : _GEN_16092; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16094 = 10'h2e7 == _T_241[9:0] ? 4'h3 : _GEN_16093; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16095 = 10'h2e8 == _T_241[9:0] ? 4'h3 : _GEN_16094; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16096 = 10'h2e9 == _T_241[9:0] ? 4'h3 : _GEN_16095; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16097 = 10'h2ea == _T_241[9:0] ? 4'h3 : _GEN_16096; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16098 = 10'h2eb == _T_241[9:0] ? 4'h3 : _GEN_16097; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16099 = 10'h2ec == _T_241[9:0] ? 4'h4 : _GEN_16098; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16100 = 10'h2ed == _T_241[9:0] ? 4'h5 : _GEN_16099; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16101 = 10'h2ee == _T_241[9:0] ? 4'h6 : _GEN_16100; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16102 = 10'h2ef == _T_241[9:0] ? 4'h8 : _GEN_16101; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16103 = 10'h2f0 == _T_241[9:0] ? 4'h4 : _GEN_16102; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16104 = 10'h2f1 == _T_241[9:0] ? 4'h9 : _GEN_16103; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16105 = 10'h2f2 == _T_241[9:0] ? 4'hb : _GEN_16104; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16106 = 10'h2f3 == _T_241[9:0] ? 4'hb : _GEN_16105; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16107 = 10'h2f4 == _T_241[9:0] ? 4'hb : _GEN_16106; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16108 = 10'h2f5 == _T_241[9:0] ? 4'hb : _GEN_16107; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16109 = 10'h2f6 == _T_241[9:0] ? 4'hb : _GEN_16108; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16110 = 10'h2f7 == _T_241[9:0] ? 4'hb : _GEN_16109; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16111 = 10'h2f8 == _T_241[9:0] ? 4'h8 : _GEN_16110; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16112 = 10'h2f9 == _T_241[9:0] ? 4'h9 : _GEN_16111; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16113 = 10'h2fa == _T_241[9:0] ? 4'hb : _GEN_16112; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16114 = 10'h2fb == _T_241[9:0] ? 4'hb : _GEN_16113; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16115 = 10'h2fc == _T_241[9:0] ? 4'ha : _GEN_16114; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16116 = 10'h2fd == _T_241[9:0] ? 4'ha : _GEN_16115; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16117 = 10'h2fe == _T_241[9:0] ? 4'h9 : _GEN_16116; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16118 = 10'h2ff == _T_241[9:0] ? 4'h8 : _GEN_16117; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16119 = 10'h300 == _T_241[9:0] ? 4'h8 : _GEN_16118; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16120 = 10'h301 == _T_241[9:0] ? 4'h6 : _GEN_16119; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16121 = 10'h302 == _T_241[9:0] ? 4'h1 : _GEN_16120; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16122 = 10'h303 == _T_241[9:0] ? 4'h0 : _GEN_16121; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16123 = 10'h304 == _T_241[9:0] ? 4'h0 : _GEN_16122; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16124 = 10'h305 == _T_241[9:0] ? 4'h0 : _GEN_16123; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16125 = 10'h306 == _T_241[9:0] ? 4'h0 : _GEN_16124; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16126 = 10'h307 == _T_241[9:0] ? 4'h0 : _GEN_16125; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16127 = 10'h308 == _T_241[9:0] ? 4'h0 : _GEN_16126; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16128 = 10'h309 == _T_241[9:0] ? 4'h0 : _GEN_16127; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16129 = 10'h30a == _T_241[9:0] ? 4'h0 : _GEN_16128; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16130 = 10'h30b == _T_241[9:0] ? 4'h0 : _GEN_16129; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16131 = 10'h30c == _T_241[9:0] ? 4'h2 : _GEN_16130; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16132 = 10'h30d == _T_241[9:0] ? 4'h3 : _GEN_16131; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16133 = 10'h30e == _T_241[9:0] ? 4'h3 : _GEN_16132; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16134 = 10'h30f == _T_241[9:0] ? 4'h3 : _GEN_16133; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16135 = 10'h310 == _T_241[9:0] ? 4'h3 : _GEN_16134; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16136 = 10'h311 == _T_241[9:0] ? 4'h3 : _GEN_16135; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16137 = 10'h312 == _T_241[9:0] ? 4'h4 : _GEN_16136; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16138 = 10'h313 == _T_241[9:0] ? 4'h5 : _GEN_16137; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16139 = 10'h314 == _T_241[9:0] ? 4'h5 : _GEN_16138; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16140 = 10'h315 == _T_241[9:0] ? 4'h8 : _GEN_16139; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16141 = 10'h316 == _T_241[9:0] ? 4'h4 : _GEN_16140; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16142 = 10'h317 == _T_241[9:0] ? 4'h6 : _GEN_16141; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16143 = 10'h318 == _T_241[9:0] ? 4'hb : _GEN_16142; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16144 = 10'h319 == _T_241[9:0] ? 4'hb : _GEN_16143; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16145 = 10'h31a == _T_241[9:0] ? 4'hb : _GEN_16144; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16146 = 10'h31b == _T_241[9:0] ? 4'hb : _GEN_16145; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16147 = 10'h31c == _T_241[9:0] ? 4'hb : _GEN_16146; // @[Filter.scala 230:102]
  wire [3:0] _GEN_16148 = 10'h31d == _T_241[9:0] ? 4'hb : _GEN_16147; // @[Filter.scala 230:102]
  wire [6:0] _GEN_38992 = {{3'd0}, _GEN_16148}; // @[Filter.scala 230:102]
  wire [10:0] _T_248 = _GEN_38992 * 7'h46; // @[Filter.scala 230:102]
  wire [10:0] _GEN_38993 = {{2'd0}, _T_243}; // @[Filter.scala 230:69]
  wire [10:0] _T_250 = _GEN_38993 + _T_248; // @[Filter.scala 230:69]
  wire [3:0] _GEN_16171 = 10'h16 == _T_241[9:0] ? 4'hb : 4'hc; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16172 = 10'h17 == _T_241[9:0] ? 4'h8 : _GEN_16171; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16173 = 10'h18 == _T_241[9:0] ? 4'ha : _GEN_16172; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16174 = 10'h19 == _T_241[9:0] ? 4'hc : _GEN_16173; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16175 = 10'h1a == _T_241[9:0] ? 4'hc : _GEN_16174; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16176 = 10'h1b == _T_241[9:0] ? 4'hc : _GEN_16175; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16177 = 10'h1c == _T_241[9:0] ? 4'hc : _GEN_16176; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16178 = 10'h1d == _T_241[9:0] ? 4'hc : _GEN_16177; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16179 = 10'h1e == _T_241[9:0] ? 4'hc : _GEN_16178; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16180 = 10'h1f == _T_241[9:0] ? 4'hc : _GEN_16179; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16181 = 10'h20 == _T_241[9:0] ? 4'hc : _GEN_16180; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16182 = 10'h21 == _T_241[9:0] ? 4'hc : _GEN_16181; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16183 = 10'h22 == _T_241[9:0] ? 4'hc : _GEN_16182; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16184 = 10'h23 == _T_241[9:0] ? 4'hc : _GEN_16183; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16185 = 10'h24 == _T_241[9:0] ? 4'hc : _GEN_16184; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16186 = 10'h25 == _T_241[9:0] ? 4'hc : _GEN_16185; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16187 = 10'h26 == _T_241[9:0] ? 4'hc : _GEN_16186; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16188 = 10'h27 == _T_241[9:0] ? 4'hc : _GEN_16187; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16189 = 10'h28 == _T_241[9:0] ? 4'hc : _GEN_16188; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16190 = 10'h29 == _T_241[9:0] ? 4'hc : _GEN_16189; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16191 = 10'h2a == _T_241[9:0] ? 4'hc : _GEN_16190; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16192 = 10'h2b == _T_241[9:0] ? 4'hc : _GEN_16191; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16193 = 10'h2c == _T_241[9:0] ? 4'hc : _GEN_16192; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16194 = 10'h2d == _T_241[9:0] ? 4'hc : _GEN_16193; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16195 = 10'h2e == _T_241[9:0] ? 4'hc : _GEN_16194; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16196 = 10'h2f == _T_241[9:0] ? 4'hc : _GEN_16195; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16197 = 10'h30 == _T_241[9:0] ? 4'hc : _GEN_16196; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16198 = 10'h31 == _T_241[9:0] ? 4'hc : _GEN_16197; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16199 = 10'h32 == _T_241[9:0] ? 4'hc : _GEN_16198; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16200 = 10'h33 == _T_241[9:0] ? 4'hc : _GEN_16199; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16201 = 10'h34 == _T_241[9:0] ? 4'hc : _GEN_16200; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16202 = 10'h35 == _T_241[9:0] ? 4'hc : _GEN_16201; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16203 = 10'h36 == _T_241[9:0] ? 4'hc : _GEN_16202; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16204 = 10'h37 == _T_241[9:0] ? 4'hc : _GEN_16203; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16205 = 10'h38 == _T_241[9:0] ? 4'hc : _GEN_16204; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16206 = 10'h39 == _T_241[9:0] ? 4'hc : _GEN_16205; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16207 = 10'h3a == _T_241[9:0] ? 4'hc : _GEN_16206; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16208 = 10'h3b == _T_241[9:0] ? 4'hc : _GEN_16207; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16209 = 10'h3c == _T_241[9:0] ? 4'h7 : _GEN_16208; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16210 = 10'h3d == _T_241[9:0] ? 4'h9 : _GEN_16209; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16211 = 10'h3e == _T_241[9:0] ? 4'h8 : _GEN_16210; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16212 = 10'h3f == _T_241[9:0] ? 4'hc : _GEN_16211; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16213 = 10'h40 == _T_241[9:0] ? 4'hc : _GEN_16212; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16214 = 10'h41 == _T_241[9:0] ? 4'hc : _GEN_16213; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16215 = 10'h42 == _T_241[9:0] ? 4'hc : _GEN_16214; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16216 = 10'h43 == _T_241[9:0] ? 4'hc : _GEN_16215; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16217 = 10'h44 == _T_241[9:0] ? 4'hc : _GEN_16216; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16218 = 10'h45 == _T_241[9:0] ? 4'hc : _GEN_16217; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16219 = 10'h46 == _T_241[9:0] ? 4'hc : _GEN_16218; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16220 = 10'h47 == _T_241[9:0] ? 4'hc : _GEN_16219; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16221 = 10'h48 == _T_241[9:0] ? 4'hc : _GEN_16220; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16222 = 10'h49 == _T_241[9:0] ? 4'hc : _GEN_16221; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16223 = 10'h4a == _T_241[9:0] ? 4'hc : _GEN_16222; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16224 = 10'h4b == _T_241[9:0] ? 4'hc : _GEN_16223; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16225 = 10'h4c == _T_241[9:0] ? 4'hc : _GEN_16224; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16226 = 10'h4d == _T_241[9:0] ? 4'hc : _GEN_16225; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16227 = 10'h4e == _T_241[9:0] ? 4'hc : _GEN_16226; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16228 = 10'h4f == _T_241[9:0] ? 4'hc : _GEN_16227; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16229 = 10'h50 == _T_241[9:0] ? 4'hc : _GEN_16228; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16230 = 10'h51 == _T_241[9:0] ? 4'hc : _GEN_16229; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16231 = 10'h52 == _T_241[9:0] ? 4'hc : _GEN_16230; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16232 = 10'h53 == _T_241[9:0] ? 4'hc : _GEN_16231; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16233 = 10'h54 == _T_241[9:0] ? 4'hc : _GEN_16232; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16234 = 10'h55 == _T_241[9:0] ? 4'hc : _GEN_16233; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16235 = 10'h56 == _T_241[9:0] ? 4'hc : _GEN_16234; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16236 = 10'h57 == _T_241[9:0] ? 4'hc : _GEN_16235; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16237 = 10'h58 == _T_241[9:0] ? 4'hc : _GEN_16236; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16238 = 10'h59 == _T_241[9:0] ? 4'hc : _GEN_16237; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16239 = 10'h5a == _T_241[9:0] ? 4'h9 : _GEN_16238; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16240 = 10'h5b == _T_241[9:0] ? 4'ha : _GEN_16239; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16241 = 10'h5c == _T_241[9:0] ? 4'hc : _GEN_16240; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16242 = 10'h5d == _T_241[9:0] ? 4'hc : _GEN_16241; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16243 = 10'h5e == _T_241[9:0] ? 4'hc : _GEN_16242; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16244 = 10'h5f == _T_241[9:0] ? 4'hc : _GEN_16243; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16245 = 10'h60 == _T_241[9:0] ? 4'hc : _GEN_16244; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16246 = 10'h61 == _T_241[9:0] ? 4'hb : _GEN_16245; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16247 = 10'h62 == _T_241[9:0] ? 4'h8 : _GEN_16246; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16248 = 10'h63 == _T_241[9:0] ? 4'h9 : _GEN_16247; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16249 = 10'h64 == _T_241[9:0] ? 4'h7 : _GEN_16248; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16250 = 10'h65 == _T_241[9:0] ? 4'hb : _GEN_16249; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16251 = 10'h66 == _T_241[9:0] ? 4'hc : _GEN_16250; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16252 = 10'h67 == _T_241[9:0] ? 4'hc : _GEN_16251; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16253 = 10'h68 == _T_241[9:0] ? 4'hc : _GEN_16252; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16254 = 10'h69 == _T_241[9:0] ? 4'hc : _GEN_16253; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16255 = 10'h6a == _T_241[9:0] ? 4'hc : _GEN_16254; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16256 = 10'h6b == _T_241[9:0] ? 4'hb : _GEN_16255; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16257 = 10'h6c == _T_241[9:0] ? 4'h9 : _GEN_16256; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16258 = 10'h6d == _T_241[9:0] ? 4'ha : _GEN_16257; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16259 = 10'h6e == _T_241[9:0] ? 4'hc : _GEN_16258; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16260 = 10'h6f == _T_241[9:0] ? 4'hc : _GEN_16259; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16261 = 10'h70 == _T_241[9:0] ? 4'hc : _GEN_16260; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16262 = 10'h71 == _T_241[9:0] ? 4'hc : _GEN_16261; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16263 = 10'h72 == _T_241[9:0] ? 4'hc : _GEN_16262; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16264 = 10'h73 == _T_241[9:0] ? 4'hc : _GEN_16263; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16265 = 10'h74 == _T_241[9:0] ? 4'hc : _GEN_16264; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16266 = 10'h75 == _T_241[9:0] ? 4'hc : _GEN_16265; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16267 = 10'h76 == _T_241[9:0] ? 4'hc : _GEN_16266; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16268 = 10'h77 == _T_241[9:0] ? 4'hc : _GEN_16267; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16269 = 10'h78 == _T_241[9:0] ? 4'hc : _GEN_16268; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16270 = 10'h79 == _T_241[9:0] ? 4'hc : _GEN_16269; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16271 = 10'h7a == _T_241[9:0] ? 4'hc : _GEN_16270; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16272 = 10'h7b == _T_241[9:0] ? 4'hc : _GEN_16271; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16273 = 10'h7c == _T_241[9:0] ? 4'hc : _GEN_16272; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16274 = 10'h7d == _T_241[9:0] ? 4'hc : _GEN_16273; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16275 = 10'h7e == _T_241[9:0] ? 4'hc : _GEN_16274; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16276 = 10'h7f == _T_241[9:0] ? 4'hc : _GEN_16275; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16277 = 10'h80 == _T_241[9:0] ? 4'hc : _GEN_16276; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16278 = 10'h81 == _T_241[9:0] ? 4'h9 : _GEN_16277; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16279 = 10'h82 == _T_241[9:0] ? 4'h9 : _GEN_16278; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16280 = 10'h83 == _T_241[9:0] ? 4'h9 : _GEN_16279; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16281 = 10'h84 == _T_241[9:0] ? 4'hc : _GEN_16280; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16282 = 10'h85 == _T_241[9:0] ? 4'hc : _GEN_16281; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16283 = 10'h86 == _T_241[9:0] ? 4'hc : _GEN_16282; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16284 = 10'h87 == _T_241[9:0] ? 4'h8 : _GEN_16283; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16285 = 10'h88 == _T_241[9:0] ? 4'h9 : _GEN_16284; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16286 = 10'h89 == _T_241[9:0] ? 4'h9 : _GEN_16285; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16287 = 10'h8a == _T_241[9:0] ? 4'h9 : _GEN_16286; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16288 = 10'h8b == _T_241[9:0] ? 4'hc : _GEN_16287; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16289 = 10'h8c == _T_241[9:0] ? 4'hc : _GEN_16288; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16290 = 10'h8d == _T_241[9:0] ? 4'hc : _GEN_16289; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16291 = 10'h8e == _T_241[9:0] ? 4'hc : _GEN_16290; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16292 = 10'h8f == _T_241[9:0] ? 4'h9 : _GEN_16291; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16293 = 10'h90 == _T_241[9:0] ? 4'h9 : _GEN_16292; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16294 = 10'h91 == _T_241[9:0] ? 4'h9 : _GEN_16293; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16295 = 10'h92 == _T_241[9:0] ? 4'ha : _GEN_16294; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16296 = 10'h93 == _T_241[9:0] ? 4'hc : _GEN_16295; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16297 = 10'h94 == _T_241[9:0] ? 4'hc : _GEN_16296; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16298 = 10'h95 == _T_241[9:0] ? 4'hc : _GEN_16297; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16299 = 10'h96 == _T_241[9:0] ? 4'hc : _GEN_16298; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16300 = 10'h97 == _T_241[9:0] ? 4'hc : _GEN_16299; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16301 = 10'h98 == _T_241[9:0] ? 4'hc : _GEN_16300; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16302 = 10'h99 == _T_241[9:0] ? 4'hc : _GEN_16301; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16303 = 10'h9a == _T_241[9:0] ? 4'hc : _GEN_16302; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16304 = 10'h9b == _T_241[9:0] ? 4'hc : _GEN_16303; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16305 = 10'h9c == _T_241[9:0] ? 4'hc : _GEN_16304; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16306 = 10'h9d == _T_241[9:0] ? 4'hc : _GEN_16305; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16307 = 10'h9e == _T_241[9:0] ? 4'hc : _GEN_16306; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16308 = 10'h9f == _T_241[9:0] ? 4'hc : _GEN_16307; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16309 = 10'ha0 == _T_241[9:0] ? 4'hc : _GEN_16308; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16310 = 10'ha1 == _T_241[9:0] ? 4'hc : _GEN_16309; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16311 = 10'ha2 == _T_241[9:0] ? 4'hc : _GEN_16310; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16312 = 10'ha3 == _T_241[9:0] ? 4'hc : _GEN_16311; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16313 = 10'ha4 == _T_241[9:0] ? 4'hc : _GEN_16312; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16314 = 10'ha5 == _T_241[9:0] ? 4'hc : _GEN_16313; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16315 = 10'ha6 == _T_241[9:0] ? 4'hc : _GEN_16314; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16316 = 10'ha7 == _T_241[9:0] ? 4'hc : _GEN_16315; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16317 = 10'ha8 == _T_241[9:0] ? 4'h9 : _GEN_16316; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16318 = 10'ha9 == _T_241[9:0] ? 4'h8 : _GEN_16317; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16319 = 10'haa == _T_241[9:0] ? 4'h8 : _GEN_16318; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16320 = 10'hab == _T_241[9:0] ? 4'ha : _GEN_16319; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16321 = 10'hac == _T_241[9:0] ? 4'hb : _GEN_16320; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16322 = 10'had == _T_241[9:0] ? 4'h7 : _GEN_16321; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16323 = 10'hae == _T_241[9:0] ? 4'h9 : _GEN_16322; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16324 = 10'haf == _T_241[9:0] ? 4'h9 : _GEN_16323; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16325 = 10'hb0 == _T_241[9:0] ? 4'h8 : _GEN_16324; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16326 = 10'hb1 == _T_241[9:0] ? 4'h9 : _GEN_16325; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16327 = 10'hb2 == _T_241[9:0] ? 4'hc : _GEN_16326; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16328 = 10'hb3 == _T_241[9:0] ? 4'h9 : _GEN_16327; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16329 = 10'hb4 == _T_241[9:0] ? 4'h9 : _GEN_16328; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16330 = 10'hb5 == _T_241[9:0] ? 4'h9 : _GEN_16329; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16331 = 10'hb6 == _T_241[9:0] ? 4'h9 : _GEN_16330; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16332 = 10'hb7 == _T_241[9:0] ? 4'ha : _GEN_16331; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16333 = 10'hb8 == _T_241[9:0] ? 4'hc : _GEN_16332; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16334 = 10'hb9 == _T_241[9:0] ? 4'hc : _GEN_16333; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16335 = 10'hba == _T_241[9:0] ? 4'hc : _GEN_16334; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16336 = 10'hbb == _T_241[9:0] ? 4'hc : _GEN_16335; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16337 = 10'hbc == _T_241[9:0] ? 4'hc : _GEN_16336; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16338 = 10'hbd == _T_241[9:0] ? 4'hb : _GEN_16337; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16339 = 10'hbe == _T_241[9:0] ? 4'hc : _GEN_16338; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16340 = 10'hbf == _T_241[9:0] ? 4'hc : _GEN_16339; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16341 = 10'hc0 == _T_241[9:0] ? 4'hc : _GEN_16340; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16342 = 10'hc1 == _T_241[9:0] ? 4'hc : _GEN_16341; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16343 = 10'hc2 == _T_241[9:0] ? 4'hc : _GEN_16342; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16344 = 10'hc3 == _T_241[9:0] ? 4'hc : _GEN_16343; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16345 = 10'hc4 == _T_241[9:0] ? 4'hc : _GEN_16344; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16346 = 10'hc5 == _T_241[9:0] ? 4'hc : _GEN_16345; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16347 = 10'hc6 == _T_241[9:0] ? 4'hb : _GEN_16346; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16348 = 10'hc7 == _T_241[9:0] ? 4'hb : _GEN_16347; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16349 = 10'hc8 == _T_241[9:0] ? 4'ha : _GEN_16348; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16350 = 10'hc9 == _T_241[9:0] ? 4'ha : _GEN_16349; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16351 = 10'hca == _T_241[9:0] ? 4'hb : _GEN_16350; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16352 = 10'hcb == _T_241[9:0] ? 4'hc : _GEN_16351; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16353 = 10'hcc == _T_241[9:0] ? 4'hc : _GEN_16352; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16354 = 10'hcd == _T_241[9:0] ? 4'hc : _GEN_16353; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16355 = 10'hce == _T_241[9:0] ? 4'ha : _GEN_16354; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16356 = 10'hcf == _T_241[9:0] ? 4'h8 : _GEN_16355; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16357 = 10'hd0 == _T_241[9:0] ? 4'h9 : _GEN_16356; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16358 = 10'hd1 == _T_241[9:0] ? 4'h8 : _GEN_16357; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16359 = 10'hd2 == _T_241[9:0] ? 4'h9 : _GEN_16358; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16360 = 10'hd3 == _T_241[9:0] ? 4'h9 : _GEN_16359; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16361 = 10'hd4 == _T_241[9:0] ? 4'h9 : _GEN_16360; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16362 = 10'hd5 == _T_241[9:0] ? 4'h9 : _GEN_16361; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16363 = 10'hd6 == _T_241[9:0] ? 4'ha : _GEN_16362; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16364 = 10'hd7 == _T_241[9:0] ? 4'h9 : _GEN_16363; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16365 = 10'hd8 == _T_241[9:0] ? 4'h9 : _GEN_16364; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16366 = 10'hd9 == _T_241[9:0] ? 4'h9 : _GEN_16365; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16367 = 10'hda == _T_241[9:0] ? 4'ha : _GEN_16366; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16368 = 10'hdb == _T_241[9:0] ? 4'h9 : _GEN_16367; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16369 = 10'hdc == _T_241[9:0] ? 4'h7 : _GEN_16368; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16370 = 10'hdd == _T_241[9:0] ? 4'hc : _GEN_16369; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16371 = 10'hde == _T_241[9:0] ? 4'hc : _GEN_16370; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16372 = 10'hdf == _T_241[9:0] ? 4'hc : _GEN_16371; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16373 = 10'he0 == _T_241[9:0] ? 4'hc : _GEN_16372; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16374 = 10'he1 == _T_241[9:0] ? 4'hc : _GEN_16373; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16375 = 10'he2 == _T_241[9:0] ? 4'hc : _GEN_16374; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16376 = 10'he3 == _T_241[9:0] ? 4'h8 : _GEN_16375; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16377 = 10'he4 == _T_241[9:0] ? 4'hc : _GEN_16376; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16378 = 10'he5 == _T_241[9:0] ? 4'hc : _GEN_16377; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16379 = 10'he6 == _T_241[9:0] ? 4'hc : _GEN_16378; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16380 = 10'he7 == _T_241[9:0] ? 4'hc : _GEN_16379; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16381 = 10'he8 == _T_241[9:0] ? 4'hc : _GEN_16380; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16382 = 10'he9 == _T_241[9:0] ? 4'hc : _GEN_16381; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16383 = 10'hea == _T_241[9:0] ? 4'hc : _GEN_16382; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16384 = 10'heb == _T_241[9:0] ? 4'ha : _GEN_16383; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16385 = 10'hec == _T_241[9:0] ? 4'h7 : _GEN_16384; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16386 = 10'hed == _T_241[9:0] ? 4'h3 : _GEN_16385; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16387 = 10'hee == _T_241[9:0] ? 4'h3 : _GEN_16386; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16388 = 10'hef == _T_241[9:0] ? 4'h3 : _GEN_16387; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16389 = 10'hf0 == _T_241[9:0] ? 4'h3 : _GEN_16388; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16390 = 10'hf1 == _T_241[9:0] ? 4'h8 : _GEN_16389; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16391 = 10'hf2 == _T_241[9:0] ? 4'hc : _GEN_16390; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16392 = 10'hf3 == _T_241[9:0] ? 4'hc : _GEN_16391; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16393 = 10'hf4 == _T_241[9:0] ? 4'hc : _GEN_16392; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16394 = 10'hf5 == _T_241[9:0] ? 4'h9 : _GEN_16393; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16395 = 10'hf6 == _T_241[9:0] ? 4'h9 : _GEN_16394; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16396 = 10'hf7 == _T_241[9:0] ? 4'h9 : _GEN_16395; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16397 = 10'hf8 == _T_241[9:0] ? 4'h9 : _GEN_16396; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16398 = 10'hf9 == _T_241[9:0] ? 4'ha : _GEN_16397; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16399 = 10'hfa == _T_241[9:0] ? 4'h9 : _GEN_16398; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16400 = 10'hfb == _T_241[9:0] ? 4'h9 : _GEN_16399; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16401 = 10'hfc == _T_241[9:0] ? 4'h9 : _GEN_16400; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16402 = 10'hfd == _T_241[9:0] ? 4'h9 : _GEN_16401; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16403 = 10'hfe == _T_241[9:0] ? 4'h9 : _GEN_16402; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16404 = 10'hff == _T_241[9:0] ? 4'ha : _GEN_16403; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16405 = 10'h100 == _T_241[9:0] ? 4'ha : _GEN_16404; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16406 = 10'h101 == _T_241[9:0] ? 4'h7 : _GEN_16405; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16407 = 10'h102 == _T_241[9:0] ? 4'h9 : _GEN_16406; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16408 = 10'h103 == _T_241[9:0] ? 4'hc : _GEN_16407; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16409 = 10'h104 == _T_241[9:0] ? 4'hc : _GEN_16408; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16410 = 10'h105 == _T_241[9:0] ? 4'hb : _GEN_16409; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16411 = 10'h106 == _T_241[9:0] ? 4'hb : _GEN_16410; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16412 = 10'h107 == _T_241[9:0] ? 4'hb : _GEN_16411; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16413 = 10'h108 == _T_241[9:0] ? 4'hb : _GEN_16412; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16414 = 10'h109 == _T_241[9:0] ? 4'h7 : _GEN_16413; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16415 = 10'h10a == _T_241[9:0] ? 4'hc : _GEN_16414; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16416 = 10'h10b == _T_241[9:0] ? 4'hc : _GEN_16415; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16417 = 10'h10c == _T_241[9:0] ? 4'hc : _GEN_16416; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16418 = 10'h10d == _T_241[9:0] ? 4'hc : _GEN_16417; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16419 = 10'h10e == _T_241[9:0] ? 4'hc : _GEN_16418; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16420 = 10'h10f == _T_241[9:0] ? 4'h9 : _GEN_16419; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16421 = 10'h110 == _T_241[9:0] ? 4'hb : _GEN_16420; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16422 = 10'h111 == _T_241[9:0] ? 4'h4 : _GEN_16421; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16423 = 10'h112 == _T_241[9:0] ? 4'h7 : _GEN_16422; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16424 = 10'h113 == _T_241[9:0] ? 4'h3 : _GEN_16423; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16425 = 10'h114 == _T_241[9:0] ? 4'h3 : _GEN_16424; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16426 = 10'h115 == _T_241[9:0] ? 4'h3 : _GEN_16425; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16427 = 10'h116 == _T_241[9:0] ? 4'h3 : _GEN_16426; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16428 = 10'h117 == _T_241[9:0] ? 4'h2 : _GEN_16427; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16429 = 10'h118 == _T_241[9:0] ? 4'h9 : _GEN_16428; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16430 = 10'h119 == _T_241[9:0] ? 4'hc : _GEN_16429; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16431 = 10'h11a == _T_241[9:0] ? 4'hc : _GEN_16430; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16432 = 10'h11b == _T_241[9:0] ? 4'hc : _GEN_16431; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16433 = 10'h11c == _T_241[9:0] ? 4'h9 : _GEN_16432; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16434 = 10'h11d == _T_241[9:0] ? 4'h9 : _GEN_16433; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16435 = 10'h11e == _T_241[9:0] ? 4'h9 : _GEN_16434; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16436 = 10'h11f == _T_241[9:0] ? 4'h8 : _GEN_16435; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16437 = 10'h120 == _T_241[9:0] ? 4'h7 : _GEN_16436; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16438 = 10'h121 == _T_241[9:0] ? 4'h9 : _GEN_16437; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16439 = 10'h122 == _T_241[9:0] ? 4'h7 : _GEN_16438; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16440 = 10'h123 == _T_241[9:0] ? 4'h7 : _GEN_16439; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16441 = 10'h124 == _T_241[9:0] ? 4'h9 : _GEN_16440; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16442 = 10'h125 == _T_241[9:0] ? 4'h9 : _GEN_16441; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16443 = 10'h126 == _T_241[9:0] ? 4'h8 : _GEN_16442; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16444 = 10'h127 == _T_241[9:0] ? 4'h9 : _GEN_16443; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16445 = 10'h128 == _T_241[9:0] ? 4'h8 : _GEN_16444; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16446 = 10'h129 == _T_241[9:0] ? 4'ha : _GEN_16445; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16447 = 10'h12a == _T_241[9:0] ? 4'h5 : _GEN_16446; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16448 = 10'h12b == _T_241[9:0] ? 4'h3 : _GEN_16447; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16449 = 10'h12c == _T_241[9:0] ? 4'h3 : _GEN_16448; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16450 = 10'h12d == _T_241[9:0] ? 4'h3 : _GEN_16449; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16451 = 10'h12e == _T_241[9:0] ? 4'h5 : _GEN_16450; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16452 = 10'h12f == _T_241[9:0] ? 4'h8 : _GEN_16451; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16453 = 10'h130 == _T_241[9:0] ? 4'hc : _GEN_16452; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16454 = 10'h131 == _T_241[9:0] ? 4'hb : _GEN_16453; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16455 = 10'h132 == _T_241[9:0] ? 4'h9 : _GEN_16454; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16456 = 10'h133 == _T_241[9:0] ? 4'h8 : _GEN_16455; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16457 = 10'h134 == _T_241[9:0] ? 4'h9 : _GEN_16456; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16458 = 10'h135 == _T_241[9:0] ? 4'h7 : _GEN_16457; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16459 = 10'h136 == _T_241[9:0] ? 4'h7 : _GEN_16458; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16460 = 10'h137 == _T_241[9:0] ? 4'h5 : _GEN_16459; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16461 = 10'h138 == _T_241[9:0] ? 4'h7 : _GEN_16460; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16462 = 10'h139 == _T_241[9:0] ? 4'h3 : _GEN_16461; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16463 = 10'h13a == _T_241[9:0] ? 4'h3 : _GEN_16462; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16464 = 10'h13b == _T_241[9:0] ? 4'h3 : _GEN_16463; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16465 = 10'h13c == _T_241[9:0] ? 4'h3 : _GEN_16464; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16466 = 10'h13d == _T_241[9:0] ? 4'h3 : _GEN_16465; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16467 = 10'h13e == _T_241[9:0] ? 4'h5 : _GEN_16466; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16468 = 10'h13f == _T_241[9:0] ? 4'ha : _GEN_16467; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16469 = 10'h140 == _T_241[9:0] ? 4'hc : _GEN_16468; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16470 = 10'h141 == _T_241[9:0] ? 4'hc : _GEN_16469; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16471 = 10'h142 == _T_241[9:0] ? 4'hc : _GEN_16470; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16472 = 10'h143 == _T_241[9:0] ? 4'h9 : _GEN_16471; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16473 = 10'h144 == _T_241[9:0] ? 4'h9 : _GEN_16472; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16474 = 10'h145 == _T_241[9:0] ? 4'h8 : _GEN_16473; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16475 = 10'h146 == _T_241[9:0] ? 4'h8 : _GEN_16474; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16476 = 10'h147 == _T_241[9:0] ? 4'h7 : _GEN_16475; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16477 = 10'h148 == _T_241[9:0] ? 4'h8 : _GEN_16476; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16478 = 10'h149 == _T_241[9:0] ? 4'h9 : _GEN_16477; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16479 = 10'h14a == _T_241[9:0] ? 4'ha : _GEN_16478; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16480 = 10'h14b == _T_241[9:0] ? 4'h9 : _GEN_16479; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16481 = 10'h14c == _T_241[9:0] ? 4'ha : _GEN_16480; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16482 = 10'h14d == _T_241[9:0] ? 4'h9 : _GEN_16481; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16483 = 10'h14e == _T_241[9:0] ? 4'h7 : _GEN_16482; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16484 = 10'h14f == _T_241[9:0] ? 4'h3 : _GEN_16483; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16485 = 10'h150 == _T_241[9:0] ? 4'h3 : _GEN_16484; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16486 = 10'h151 == _T_241[9:0] ? 4'h3 : _GEN_16485; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16487 = 10'h152 == _T_241[9:0] ? 4'h3 : _GEN_16486; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16488 = 10'h153 == _T_241[9:0] ? 4'h3 : _GEN_16487; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16489 = 10'h154 == _T_241[9:0] ? 4'h3 : _GEN_16488; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16490 = 10'h155 == _T_241[9:0] ? 4'h8 : _GEN_16489; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16491 = 10'h156 == _T_241[9:0] ? 4'ha : _GEN_16490; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16492 = 10'h157 == _T_241[9:0] ? 4'h7 : _GEN_16491; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16493 = 10'h158 == _T_241[9:0] ? 4'h7 : _GEN_16492; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16494 = 10'h159 == _T_241[9:0] ? 4'h7 : _GEN_16493; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16495 = 10'h15a == _T_241[9:0] ? 4'h7 : _GEN_16494; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16496 = 10'h15b == _T_241[9:0] ? 4'h7 : _GEN_16495; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16497 = 10'h15c == _T_241[9:0] ? 4'h7 : _GEN_16496; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16498 = 10'h15d == _T_241[9:0] ? 4'h7 : _GEN_16497; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16499 = 10'h15e == _T_241[9:0] ? 4'h7 : _GEN_16498; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16500 = 10'h15f == _T_241[9:0] ? 4'h3 : _GEN_16499; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16501 = 10'h160 == _T_241[9:0] ? 4'h3 : _GEN_16500; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16502 = 10'h161 == _T_241[9:0] ? 4'h3 : _GEN_16501; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16503 = 10'h162 == _T_241[9:0] ? 4'h3 : _GEN_16502; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16504 = 10'h163 == _T_241[9:0] ? 4'h3 : _GEN_16503; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16505 = 10'h164 == _T_241[9:0] ? 4'h4 : _GEN_16504; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16506 = 10'h165 == _T_241[9:0] ? 4'ha : _GEN_16505; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16507 = 10'h166 == _T_241[9:0] ? 4'ha : _GEN_16506; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16508 = 10'h167 == _T_241[9:0] ? 4'hc : _GEN_16507; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16509 = 10'h168 == _T_241[9:0] ? 4'hc : _GEN_16508; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16510 = 10'h169 == _T_241[9:0] ? 4'h9 : _GEN_16509; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16511 = 10'h16a == _T_241[9:0] ? 4'h9 : _GEN_16510; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16512 = 10'h16b == _T_241[9:0] ? 4'ha : _GEN_16511; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16513 = 10'h16c == _T_241[9:0] ? 4'h7 : _GEN_16512; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16514 = 10'h16d == _T_241[9:0] ? 4'h7 : _GEN_16513; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16515 = 10'h16e == _T_241[9:0] ? 4'h7 : _GEN_16514; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16516 = 10'h16f == _T_241[9:0] ? 4'ha : _GEN_16515; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16517 = 10'h170 == _T_241[9:0] ? 4'ha : _GEN_16516; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16518 = 10'h171 == _T_241[9:0] ? 4'ha : _GEN_16517; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16519 = 10'h172 == _T_241[9:0] ? 4'hc : _GEN_16518; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16520 = 10'h173 == _T_241[9:0] ? 4'h8 : _GEN_16519; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16521 = 10'h174 == _T_241[9:0] ? 4'h5 : _GEN_16520; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16522 = 10'h175 == _T_241[9:0] ? 4'h8 : _GEN_16521; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16523 = 10'h176 == _T_241[9:0] ? 4'h7 : _GEN_16522; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16524 = 10'h177 == _T_241[9:0] ? 4'h8 : _GEN_16523; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16525 = 10'h178 == _T_241[9:0] ? 4'h7 : _GEN_16524; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16526 = 10'h179 == _T_241[9:0] ? 4'h5 : _GEN_16525; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16527 = 10'h17a == _T_241[9:0] ? 4'h5 : _GEN_16526; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16528 = 10'h17b == _T_241[9:0] ? 4'h7 : _GEN_16527; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16529 = 10'h17c == _T_241[9:0] ? 4'h7 : _GEN_16528; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16530 = 10'h17d == _T_241[9:0] ? 4'h7 : _GEN_16529; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16531 = 10'h17e == _T_241[9:0] ? 4'h7 : _GEN_16530; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16532 = 10'h17f == _T_241[9:0] ? 4'h7 : _GEN_16531; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16533 = 10'h180 == _T_241[9:0] ? 4'h7 : _GEN_16532; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16534 = 10'h181 == _T_241[9:0] ? 4'h7 : _GEN_16533; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16535 = 10'h182 == _T_241[9:0] ? 4'h7 : _GEN_16534; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16536 = 10'h183 == _T_241[9:0] ? 4'h7 : _GEN_16535; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16537 = 10'h184 == _T_241[9:0] ? 4'h7 : _GEN_16536; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16538 = 10'h185 == _T_241[9:0] ? 4'h5 : _GEN_16537; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16539 = 10'h186 == _T_241[9:0] ? 4'h3 : _GEN_16538; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16540 = 10'h187 == _T_241[9:0] ? 4'h3 : _GEN_16539; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16541 = 10'h188 == _T_241[9:0] ? 4'h3 : _GEN_16540; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16542 = 10'h189 == _T_241[9:0] ? 4'h4 : _GEN_16541; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16543 = 10'h18a == _T_241[9:0] ? 4'h5 : _GEN_16542; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16544 = 10'h18b == _T_241[9:0] ? 4'ha : _GEN_16543; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16545 = 10'h18c == _T_241[9:0] ? 4'ha : _GEN_16544; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16546 = 10'h18d == _T_241[9:0] ? 4'ha : _GEN_16545; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16547 = 10'h18e == _T_241[9:0] ? 4'hc : _GEN_16546; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16548 = 10'h18f == _T_241[9:0] ? 4'h8 : _GEN_16547; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16549 = 10'h190 == _T_241[9:0] ? 4'h9 : _GEN_16548; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16550 = 10'h191 == _T_241[9:0] ? 4'h8 : _GEN_16549; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16551 = 10'h192 == _T_241[9:0] ? 4'h7 : _GEN_16550; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16552 = 10'h193 == _T_241[9:0] ? 4'h7 : _GEN_16551; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16553 = 10'h194 == _T_241[9:0] ? 4'h7 : _GEN_16552; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16554 = 10'h195 == _T_241[9:0] ? 4'h9 : _GEN_16553; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16555 = 10'h196 == _T_241[9:0] ? 4'ha : _GEN_16554; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16556 = 10'h197 == _T_241[9:0] ? 4'h8 : _GEN_16555; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16557 = 10'h198 == _T_241[9:0] ? 4'hc : _GEN_16556; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16558 = 10'h199 == _T_241[9:0] ? 4'h5 : _GEN_16557; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16559 = 10'h19a == _T_241[9:0] ? 4'h1 : _GEN_16558; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16560 = 10'h19b == _T_241[9:0] ? 4'h4 : _GEN_16559; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16561 = 10'h19c == _T_241[9:0] ? 4'h7 : _GEN_16560; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16562 = 10'h19d == _T_241[9:0] ? 4'h5 : _GEN_16561; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16563 = 10'h19e == _T_241[9:0] ? 4'h2 : _GEN_16562; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16564 = 10'h19f == _T_241[9:0] ? 4'h3 : _GEN_16563; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16565 = 10'h1a0 == _T_241[9:0] ? 4'h7 : _GEN_16564; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16566 = 10'h1a1 == _T_241[9:0] ? 4'h7 : _GEN_16565; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16567 = 10'h1a2 == _T_241[9:0] ? 4'h7 : _GEN_16566; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16568 = 10'h1a3 == _T_241[9:0] ? 4'h7 : _GEN_16567; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16569 = 10'h1a4 == _T_241[9:0] ? 4'h7 : _GEN_16568; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16570 = 10'h1a5 == _T_241[9:0] ? 4'h7 : _GEN_16569; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16571 = 10'h1a6 == _T_241[9:0] ? 4'h7 : _GEN_16570; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16572 = 10'h1a7 == _T_241[9:0] ? 4'h7 : _GEN_16571; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16573 = 10'h1a8 == _T_241[9:0] ? 4'h8 : _GEN_16572; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16574 = 10'h1a9 == _T_241[9:0] ? 4'h8 : _GEN_16573; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16575 = 10'h1aa == _T_241[9:0] ? 4'h6 : _GEN_16574; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16576 = 10'h1ab == _T_241[9:0] ? 4'h6 : _GEN_16575; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16577 = 10'h1ac == _T_241[9:0] ? 4'h5 : _GEN_16576; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16578 = 10'h1ad == _T_241[9:0] ? 4'h4 : _GEN_16577; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16579 = 10'h1ae == _T_241[9:0] ? 4'h3 : _GEN_16578; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16580 = 10'h1af == _T_241[9:0] ? 4'h6 : _GEN_16579; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16581 = 10'h1b0 == _T_241[9:0] ? 4'h6 : _GEN_16580; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16582 = 10'h1b1 == _T_241[9:0] ? 4'ha : _GEN_16581; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16583 = 10'h1b2 == _T_241[9:0] ? 4'ha : _GEN_16582; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16584 = 10'h1b3 == _T_241[9:0] ? 4'h9 : _GEN_16583; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16585 = 10'h1b4 == _T_241[9:0] ? 4'hb : _GEN_16584; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16586 = 10'h1b5 == _T_241[9:0] ? 4'h8 : _GEN_16585; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16587 = 10'h1b6 == _T_241[9:0] ? 4'h8 : _GEN_16586; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16588 = 10'h1b7 == _T_241[9:0] ? 4'h7 : _GEN_16587; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16589 = 10'h1b8 == _T_241[9:0] ? 4'h6 : _GEN_16588; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16590 = 10'h1b9 == _T_241[9:0] ? 4'h7 : _GEN_16589; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16591 = 10'h1ba == _T_241[9:0] ? 4'h6 : _GEN_16590; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16592 = 10'h1bb == _T_241[9:0] ? 4'h8 : _GEN_16591; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16593 = 10'h1bc == _T_241[9:0] ? 4'ha : _GEN_16592; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16594 = 10'h1bd == _T_241[9:0] ? 4'h9 : _GEN_16593; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16595 = 10'h1be == _T_241[9:0] ? 4'hc : _GEN_16594; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16596 = 10'h1bf == _T_241[9:0] ? 4'h7 : _GEN_16595; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16597 = 10'h1c0 == _T_241[9:0] ? 4'h6 : _GEN_16596; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16598 = 10'h1c1 == _T_241[9:0] ? 4'h7 : _GEN_16597; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16599 = 10'h1c2 == _T_241[9:0] ? 4'h7 : _GEN_16598; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16600 = 10'h1c3 == _T_241[9:0] ? 4'h6 : _GEN_16599; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16601 = 10'h1c4 == _T_241[9:0] ? 4'h5 : _GEN_16600; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16602 = 10'h1c5 == _T_241[9:0] ? 4'h6 : _GEN_16601; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16603 = 10'h1c6 == _T_241[9:0] ? 4'h8 : _GEN_16602; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16604 = 10'h1c7 == _T_241[9:0] ? 4'h7 : _GEN_16603; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16605 = 10'h1c8 == _T_241[9:0] ? 4'h7 : _GEN_16604; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16606 = 10'h1c9 == _T_241[9:0] ? 4'h7 : _GEN_16605; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16607 = 10'h1ca == _T_241[9:0] ? 4'h7 : _GEN_16606; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16608 = 10'h1cb == _T_241[9:0] ? 4'h7 : _GEN_16607; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16609 = 10'h1cc == _T_241[9:0] ? 4'h7 : _GEN_16608; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16610 = 10'h1cd == _T_241[9:0] ? 4'h8 : _GEN_16609; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16611 = 10'h1ce == _T_241[9:0] ? 4'h8 : _GEN_16610; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16612 = 10'h1cf == _T_241[9:0] ? 4'h8 : _GEN_16611; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16613 = 10'h1d0 == _T_241[9:0] ? 4'h5 : _GEN_16612; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16614 = 10'h1d1 == _T_241[9:0] ? 4'h6 : _GEN_16613; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16615 = 10'h1d2 == _T_241[9:0] ? 4'h7 : _GEN_16614; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16616 = 10'h1d3 == _T_241[9:0] ? 4'h7 : _GEN_16615; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16617 = 10'h1d4 == _T_241[9:0] ? 4'h7 : _GEN_16616; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16618 = 10'h1d5 == _T_241[9:0] ? 4'h6 : _GEN_16617; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16619 = 10'h1d6 == _T_241[9:0] ? 4'h8 : _GEN_16618; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16620 = 10'h1d7 == _T_241[9:0] ? 4'ha : _GEN_16619; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16621 = 10'h1d8 == _T_241[9:0] ? 4'ha : _GEN_16620; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16622 = 10'h1d9 == _T_241[9:0] ? 4'ha : _GEN_16621; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16623 = 10'h1da == _T_241[9:0] ? 4'h8 : _GEN_16622; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16624 = 10'h1db == _T_241[9:0] ? 4'h9 : _GEN_16623; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16625 = 10'h1dc == _T_241[9:0] ? 4'h9 : _GEN_16624; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16626 = 10'h1dd == _T_241[9:0] ? 4'h5 : _GEN_16625; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16627 = 10'h1de == _T_241[9:0] ? 4'h7 : _GEN_16626; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16628 = 10'h1df == _T_241[9:0] ? 4'h7 : _GEN_16627; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16629 = 10'h1e0 == _T_241[9:0] ? 4'h7 : _GEN_16628; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16630 = 10'h1e1 == _T_241[9:0] ? 4'h6 : _GEN_16629; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16631 = 10'h1e2 == _T_241[9:0] ? 4'h9 : _GEN_16630; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16632 = 10'h1e3 == _T_241[9:0] ? 4'h9 : _GEN_16631; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16633 = 10'h1e4 == _T_241[9:0] ? 4'hb : _GEN_16632; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16634 = 10'h1e5 == _T_241[9:0] ? 4'h8 : _GEN_16633; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16635 = 10'h1e6 == _T_241[9:0] ? 4'h7 : _GEN_16634; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16636 = 10'h1e7 == _T_241[9:0] ? 4'h8 : _GEN_16635; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16637 = 10'h1e8 == _T_241[9:0] ? 4'h8 : _GEN_16636; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16638 = 10'h1e9 == _T_241[9:0] ? 4'h8 : _GEN_16637; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16639 = 10'h1ea == _T_241[9:0] ? 4'h8 : _GEN_16638; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16640 = 10'h1eb == _T_241[9:0] ? 4'h8 : _GEN_16639; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16641 = 10'h1ec == _T_241[9:0] ? 4'h8 : _GEN_16640; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16642 = 10'h1ed == _T_241[9:0] ? 4'h6 : _GEN_16641; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16643 = 10'h1ee == _T_241[9:0] ? 4'h7 : _GEN_16642; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16644 = 10'h1ef == _T_241[9:0] ? 4'h7 : _GEN_16643; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16645 = 10'h1f0 == _T_241[9:0] ? 4'h7 : _GEN_16644; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16646 = 10'h1f1 == _T_241[9:0] ? 4'h7 : _GEN_16645; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16647 = 10'h1f2 == _T_241[9:0] ? 4'h7 : _GEN_16646; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16648 = 10'h1f3 == _T_241[9:0] ? 4'h8 : _GEN_16647; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16649 = 10'h1f4 == _T_241[9:0] ? 4'h8 : _GEN_16648; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16650 = 10'h1f5 == _T_241[9:0] ? 4'h8 : _GEN_16649; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16651 = 10'h1f6 == _T_241[9:0] ? 4'ha : _GEN_16650; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16652 = 10'h1f7 == _T_241[9:0] ? 4'h6 : _GEN_16651; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16653 = 10'h1f8 == _T_241[9:0] ? 4'h6 : _GEN_16652; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16654 = 10'h1f9 == _T_241[9:0] ? 4'h8 : _GEN_16653; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16655 = 10'h1fa == _T_241[9:0] ? 4'h8 : _GEN_16654; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16656 = 10'h1fb == _T_241[9:0] ? 4'h6 : _GEN_16655; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16657 = 10'h1fc == _T_241[9:0] ? 4'ha : _GEN_16656; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16658 = 10'h1fd == _T_241[9:0] ? 4'hb : _GEN_16657; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16659 = 10'h1fe == _T_241[9:0] ? 4'ha : _GEN_16658; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16660 = 10'h1ff == _T_241[9:0] ? 4'ha : _GEN_16659; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16661 = 10'h200 == _T_241[9:0] ? 4'h4 : _GEN_16660; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16662 = 10'h201 == _T_241[9:0] ? 4'h7 : _GEN_16661; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16663 = 10'h202 == _T_241[9:0] ? 4'h6 : _GEN_16662; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16664 = 10'h203 == _T_241[9:0] ? 4'h6 : _GEN_16663; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16665 = 10'h204 == _T_241[9:0] ? 4'h5 : _GEN_16664; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16666 = 10'h205 == _T_241[9:0] ? 4'h6 : _GEN_16665; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16667 = 10'h206 == _T_241[9:0] ? 4'h6 : _GEN_16666; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16668 = 10'h207 == _T_241[9:0] ? 4'h5 : _GEN_16667; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16669 = 10'h208 == _T_241[9:0] ? 4'h7 : _GEN_16668; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16670 = 10'h209 == _T_241[9:0] ? 4'h9 : _GEN_16669; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16671 = 10'h20a == _T_241[9:0] ? 4'hb : _GEN_16670; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16672 = 10'h20b == _T_241[9:0] ? 4'h7 : _GEN_16671; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16673 = 10'h20c == _T_241[9:0] ? 4'h7 : _GEN_16672; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16674 = 10'h20d == _T_241[9:0] ? 4'h7 : _GEN_16673; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16675 = 10'h20e == _T_241[9:0] ? 4'h7 : _GEN_16674; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16676 = 10'h20f == _T_241[9:0] ? 4'h7 : _GEN_16675; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16677 = 10'h210 == _T_241[9:0] ? 4'h7 : _GEN_16676; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16678 = 10'h211 == _T_241[9:0] ? 4'h8 : _GEN_16677; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16679 = 10'h212 == _T_241[9:0] ? 4'h8 : _GEN_16678; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16680 = 10'h213 == _T_241[9:0] ? 4'h9 : _GEN_16679; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16681 = 10'h214 == _T_241[9:0] ? 4'h6 : _GEN_16680; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16682 = 10'h215 == _T_241[9:0] ? 4'h7 : _GEN_16681; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16683 = 10'h216 == _T_241[9:0] ? 4'h7 : _GEN_16682; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16684 = 10'h217 == _T_241[9:0] ? 4'h7 : _GEN_16683; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16685 = 10'h218 == _T_241[9:0] ? 4'h7 : _GEN_16684; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16686 = 10'h219 == _T_241[9:0] ? 4'h8 : _GEN_16685; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16687 = 10'h21a == _T_241[9:0] ? 4'h7 : _GEN_16686; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16688 = 10'h21b == _T_241[9:0] ? 4'h8 : _GEN_16687; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16689 = 10'h21c == _T_241[9:0] ? 4'ha : _GEN_16688; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16690 = 10'h21d == _T_241[9:0] ? 4'ha : _GEN_16689; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16691 = 10'h21e == _T_241[9:0] ? 4'h7 : _GEN_16690; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16692 = 10'h21f == _T_241[9:0] ? 4'h6 : _GEN_16691; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16693 = 10'h220 == _T_241[9:0] ? 4'h6 : _GEN_16692; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16694 = 10'h221 == _T_241[9:0] ? 4'h7 : _GEN_16693; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16695 = 10'h222 == _T_241[9:0] ? 4'ha : _GEN_16694; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16696 = 10'h223 == _T_241[9:0] ? 4'ha : _GEN_16695; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16697 = 10'h224 == _T_241[9:0] ? 4'ha : _GEN_16696; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16698 = 10'h225 == _T_241[9:0] ? 4'h8 : _GEN_16697; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16699 = 10'h226 == _T_241[9:0] ? 4'h3 : _GEN_16698; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16700 = 10'h227 == _T_241[9:0] ? 4'h4 : _GEN_16699; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16701 = 10'h228 == _T_241[9:0] ? 4'h6 : _GEN_16700; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16702 = 10'h229 == _T_241[9:0] ? 4'h6 : _GEN_16701; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16703 = 10'h22a == _T_241[9:0] ? 4'h6 : _GEN_16702; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16704 = 10'h22b == _T_241[9:0] ? 4'h6 : _GEN_16703; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16705 = 10'h22c == _T_241[9:0] ? 4'h5 : _GEN_16704; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16706 = 10'h22d == _T_241[9:0] ? 4'h6 : _GEN_16705; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16707 = 10'h22e == _T_241[9:0] ? 4'h6 : _GEN_16706; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16708 = 10'h22f == _T_241[9:0] ? 4'h8 : _GEN_16707; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16709 = 10'h230 == _T_241[9:0] ? 4'h7 : _GEN_16708; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16710 = 10'h231 == _T_241[9:0] ? 4'h5 : _GEN_16709; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16711 = 10'h232 == _T_241[9:0] ? 4'h6 : _GEN_16710; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16712 = 10'h233 == _T_241[9:0] ? 4'h8 : _GEN_16711; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16713 = 10'h234 == _T_241[9:0] ? 4'h8 : _GEN_16712; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16714 = 10'h235 == _T_241[9:0] ? 4'h8 : _GEN_16713; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16715 = 10'h236 == _T_241[9:0] ? 4'h8 : _GEN_16714; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16716 = 10'h237 == _T_241[9:0] ? 4'h8 : _GEN_16715; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16717 = 10'h238 == _T_241[9:0] ? 4'h8 : _GEN_16716; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16718 = 10'h239 == _T_241[9:0] ? 4'h6 : _GEN_16717; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16719 = 10'h23a == _T_241[9:0] ? 4'h6 : _GEN_16718; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16720 = 10'h23b == _T_241[9:0] ? 4'h7 : _GEN_16719; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16721 = 10'h23c == _T_241[9:0] ? 4'h6 : _GEN_16720; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16722 = 10'h23d == _T_241[9:0] ? 4'h7 : _GEN_16721; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16723 = 10'h23e == _T_241[9:0] ? 4'h7 : _GEN_16722; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16724 = 10'h23f == _T_241[9:0] ? 4'h6 : _GEN_16723; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16725 = 10'h240 == _T_241[9:0] ? 4'h6 : _GEN_16724; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16726 = 10'h241 == _T_241[9:0] ? 4'h8 : _GEN_16725; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16727 = 10'h242 == _T_241[9:0] ? 4'ha : _GEN_16726; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16728 = 10'h243 == _T_241[9:0] ? 4'ha : _GEN_16727; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16729 = 10'h244 == _T_241[9:0] ? 4'ha : _GEN_16728; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16730 = 10'h245 == _T_241[9:0] ? 4'h8 : _GEN_16729; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16731 = 10'h246 == _T_241[9:0] ? 4'h8 : _GEN_16730; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16732 = 10'h247 == _T_241[9:0] ? 4'h9 : _GEN_16731; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16733 = 10'h248 == _T_241[9:0] ? 4'ha : _GEN_16732; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16734 = 10'h249 == _T_241[9:0] ? 4'ha : _GEN_16733; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16735 = 10'h24a == _T_241[9:0] ? 4'ha : _GEN_16734; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16736 = 10'h24b == _T_241[9:0] ? 4'h4 : _GEN_16735; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16737 = 10'h24c == _T_241[9:0] ? 4'h3 : _GEN_16736; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16738 = 10'h24d == _T_241[9:0] ? 4'h4 : _GEN_16737; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16739 = 10'h24e == _T_241[9:0] ? 4'h5 : _GEN_16738; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16740 = 10'h24f == _T_241[9:0] ? 4'h5 : _GEN_16739; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16741 = 10'h250 == _T_241[9:0] ? 4'h5 : _GEN_16740; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16742 = 10'h251 == _T_241[9:0] ? 4'h5 : _GEN_16741; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16743 = 10'h252 == _T_241[9:0] ? 4'h5 : _GEN_16742; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16744 = 10'h253 == _T_241[9:0] ? 4'h5 : _GEN_16743; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16745 = 10'h254 == _T_241[9:0] ? 4'h5 : _GEN_16744; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16746 = 10'h255 == _T_241[9:0] ? 4'h6 : _GEN_16745; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16747 = 10'h256 == _T_241[9:0] ? 4'h7 : _GEN_16746; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16748 = 10'h257 == _T_241[9:0] ? 4'h3 : _GEN_16747; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16749 = 10'h258 == _T_241[9:0] ? 4'h6 : _GEN_16748; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16750 = 10'h259 == _T_241[9:0] ? 4'h7 : _GEN_16749; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16751 = 10'h25a == _T_241[9:0] ? 4'h7 : _GEN_16750; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16752 = 10'h25b == _T_241[9:0] ? 4'h7 : _GEN_16751; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16753 = 10'h25c == _T_241[9:0] ? 4'h8 : _GEN_16752; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16754 = 10'h25d == _T_241[9:0] ? 4'h8 : _GEN_16753; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16755 = 10'h25e == _T_241[9:0] ? 4'h4 : _GEN_16754; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16756 = 10'h25f == _T_241[9:0] ? 4'h3 : _GEN_16755; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16757 = 10'h260 == _T_241[9:0] ? 4'h7 : _GEN_16756; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16758 = 10'h261 == _T_241[9:0] ? 4'h7 : _GEN_16757; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16759 = 10'h262 == _T_241[9:0] ? 4'h7 : _GEN_16758; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16760 = 10'h263 == _T_241[9:0] ? 4'h6 : _GEN_16759; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16761 = 10'h264 == _T_241[9:0] ? 4'h7 : _GEN_16760; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16762 = 10'h265 == _T_241[9:0] ? 4'h6 : _GEN_16761; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16763 = 10'h266 == _T_241[9:0] ? 4'h5 : _GEN_16762; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16764 = 10'h267 == _T_241[9:0] ? 4'h7 : _GEN_16763; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16765 = 10'h268 == _T_241[9:0] ? 4'ha : _GEN_16764; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16766 = 10'h269 == _T_241[9:0] ? 4'ha : _GEN_16765; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16767 = 10'h26a == _T_241[9:0] ? 4'ha : _GEN_16766; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16768 = 10'h26b == _T_241[9:0] ? 4'ha : _GEN_16767; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16769 = 10'h26c == _T_241[9:0] ? 4'ha : _GEN_16768; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16770 = 10'h26d == _T_241[9:0] ? 4'ha : _GEN_16769; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16771 = 10'h26e == _T_241[9:0] ? 4'ha : _GEN_16770; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16772 = 10'h26f == _T_241[9:0] ? 4'ha : _GEN_16771; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16773 = 10'h270 == _T_241[9:0] ? 4'h5 : _GEN_16772; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16774 = 10'h271 == _T_241[9:0] ? 4'h3 : _GEN_16773; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16775 = 10'h272 == _T_241[9:0] ? 4'h3 : _GEN_16774; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16776 = 10'h273 == _T_241[9:0] ? 4'h4 : _GEN_16775; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16777 = 10'h274 == _T_241[9:0] ? 4'h6 : _GEN_16776; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16778 = 10'h275 == _T_241[9:0] ? 4'h5 : _GEN_16777; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16779 = 10'h276 == _T_241[9:0] ? 4'h6 : _GEN_16778; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16780 = 10'h277 == _T_241[9:0] ? 4'h5 : _GEN_16779; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16781 = 10'h278 == _T_241[9:0] ? 4'h6 : _GEN_16780; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16782 = 10'h279 == _T_241[9:0] ? 4'h6 : _GEN_16781; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16783 = 10'h27a == _T_241[9:0] ? 4'h6 : _GEN_16782; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16784 = 10'h27b == _T_241[9:0] ? 4'h8 : _GEN_16783; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16785 = 10'h27c == _T_241[9:0] ? 4'h6 : _GEN_16784; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16786 = 10'h27d == _T_241[9:0] ? 4'h2 : _GEN_16785; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16787 = 10'h27e == _T_241[9:0] ? 4'h5 : _GEN_16786; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16788 = 10'h27f == _T_241[9:0] ? 4'h7 : _GEN_16787; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16789 = 10'h280 == _T_241[9:0] ? 4'h7 : _GEN_16788; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16790 = 10'h281 == _T_241[9:0] ? 4'h8 : _GEN_16789; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16791 = 10'h282 == _T_241[9:0] ? 4'h7 : _GEN_16790; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16792 = 10'h283 == _T_241[9:0] ? 4'h3 : _GEN_16791; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16793 = 10'h284 == _T_241[9:0] ? 4'h3 : _GEN_16792; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16794 = 10'h285 == _T_241[9:0] ? 4'h3 : _GEN_16793; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16795 = 10'h286 == _T_241[9:0] ? 4'h7 : _GEN_16794; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16796 = 10'h287 == _T_241[9:0] ? 4'h7 : _GEN_16795; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16797 = 10'h288 == _T_241[9:0] ? 4'h7 : _GEN_16796; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16798 = 10'h289 == _T_241[9:0] ? 4'h7 : _GEN_16797; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16799 = 10'h28a == _T_241[9:0] ? 4'h8 : _GEN_16798; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16800 = 10'h28b == _T_241[9:0] ? 4'h8 : _GEN_16799; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16801 = 10'h28c == _T_241[9:0] ? 4'h7 : _GEN_16800; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16802 = 10'h28d == _T_241[9:0] ? 4'h6 : _GEN_16801; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16803 = 10'h28e == _T_241[9:0] ? 4'h3 : _GEN_16802; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16804 = 10'h28f == _T_241[9:0] ? 4'h6 : _GEN_16803; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16805 = 10'h290 == _T_241[9:0] ? 4'h8 : _GEN_16804; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16806 = 10'h291 == _T_241[9:0] ? 4'ha : _GEN_16805; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16807 = 10'h292 == _T_241[9:0] ? 4'ha : _GEN_16806; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16808 = 10'h293 == _T_241[9:0] ? 4'ha : _GEN_16807; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16809 = 10'h294 == _T_241[9:0] ? 4'h9 : _GEN_16808; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16810 = 10'h295 == _T_241[9:0] ? 4'h4 : _GEN_16809; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16811 = 10'h296 == _T_241[9:0] ? 4'h3 : _GEN_16810; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16812 = 10'h297 == _T_241[9:0] ? 4'h3 : _GEN_16811; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16813 = 10'h298 == _T_241[9:0] ? 4'h3 : _GEN_16812; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16814 = 10'h299 == _T_241[9:0] ? 4'h4 : _GEN_16813; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16815 = 10'h29a == _T_241[9:0] ? 4'h5 : _GEN_16814; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16816 = 10'h29b == _T_241[9:0] ? 4'h5 : _GEN_16815; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16817 = 10'h29c == _T_241[9:0] ? 4'h5 : _GEN_16816; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16818 = 10'h29d == _T_241[9:0] ? 4'h5 : _GEN_16817; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16819 = 10'h29e == _T_241[9:0] ? 4'h5 : _GEN_16818; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16820 = 10'h29f == _T_241[9:0] ? 4'h5 : _GEN_16819; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16821 = 10'h2a0 == _T_241[9:0] ? 4'h6 : _GEN_16820; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16822 = 10'h2a1 == _T_241[9:0] ? 4'h7 : _GEN_16821; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16823 = 10'h2a2 == _T_241[9:0] ? 4'h5 : _GEN_16822; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16824 = 10'h2a3 == _T_241[9:0] ? 4'h2 : _GEN_16823; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16825 = 10'h2a4 == _T_241[9:0] ? 4'h3 : _GEN_16824; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16826 = 10'h2a5 == _T_241[9:0] ? 4'h7 : _GEN_16825; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16827 = 10'h2a6 == _T_241[9:0] ? 4'h8 : _GEN_16826; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16828 = 10'h2a7 == _T_241[9:0] ? 4'h7 : _GEN_16827; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16829 = 10'h2a8 == _T_241[9:0] ? 4'h3 : _GEN_16828; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16830 = 10'h2a9 == _T_241[9:0] ? 4'h2 : _GEN_16829; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16831 = 10'h2aa == _T_241[9:0] ? 4'h3 : _GEN_16830; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16832 = 10'h2ab == _T_241[9:0] ? 4'h3 : _GEN_16831; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16833 = 10'h2ac == _T_241[9:0] ? 4'h7 : _GEN_16832; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16834 = 10'h2ad == _T_241[9:0] ? 4'h8 : _GEN_16833; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16835 = 10'h2ae == _T_241[9:0] ? 4'h7 : _GEN_16834; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16836 = 10'h2af == _T_241[9:0] ? 4'h8 : _GEN_16835; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16837 = 10'h2b0 == _T_241[9:0] ? 4'h8 : _GEN_16836; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16838 = 10'h2b1 == _T_241[9:0] ? 4'h8 : _GEN_16837; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16839 = 10'h2b2 == _T_241[9:0] ? 4'h7 : _GEN_16838; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16840 = 10'h2b3 == _T_241[9:0] ? 4'h6 : _GEN_16839; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16841 = 10'h2b4 == _T_241[9:0] ? 4'h2 : _GEN_16840; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16842 = 10'h2b5 == _T_241[9:0] ? 4'h2 : _GEN_16841; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16843 = 10'h2b6 == _T_241[9:0] ? 4'h3 : _GEN_16842; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16844 = 10'h2b7 == _T_241[9:0] ? 4'h3 : _GEN_16843; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16845 = 10'h2b8 == _T_241[9:0] ? 4'h6 : _GEN_16844; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16846 = 10'h2b9 == _T_241[9:0] ? 4'h9 : _GEN_16845; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16847 = 10'h2ba == _T_241[9:0] ? 4'h3 : _GEN_16846; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16848 = 10'h2bb == _T_241[9:0] ? 4'h3 : _GEN_16847; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16849 = 10'h2bc == _T_241[9:0] ? 4'h3 : _GEN_16848; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16850 = 10'h2bd == _T_241[9:0] ? 4'h2 : _GEN_16849; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16851 = 10'h2be == _T_241[9:0] ? 4'h3 : _GEN_16850; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16852 = 10'h2bf == _T_241[9:0] ? 4'h3 : _GEN_16851; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16853 = 10'h2c0 == _T_241[9:0] ? 4'h5 : _GEN_16852; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16854 = 10'h2c1 == _T_241[9:0] ? 4'h5 : _GEN_16853; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16855 = 10'h2c2 == _T_241[9:0] ? 4'h5 : _GEN_16854; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16856 = 10'h2c3 == _T_241[9:0] ? 4'h5 : _GEN_16855; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16857 = 10'h2c4 == _T_241[9:0] ? 4'h5 : _GEN_16856; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16858 = 10'h2c5 == _T_241[9:0] ? 4'h5 : _GEN_16857; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16859 = 10'h2c6 == _T_241[9:0] ? 4'h6 : _GEN_16858; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16860 = 10'h2c7 == _T_241[9:0] ? 4'h7 : _GEN_16859; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16861 = 10'h2c8 == _T_241[9:0] ? 4'h5 : _GEN_16860; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16862 = 10'h2c9 == _T_241[9:0] ? 4'h2 : _GEN_16861; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16863 = 10'h2ca == _T_241[9:0] ? 4'h2 : _GEN_16862; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16864 = 10'h2cb == _T_241[9:0] ? 4'h3 : _GEN_16863; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16865 = 10'h2cc == _T_241[9:0] ? 4'h3 : _GEN_16864; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16866 = 10'h2cd == _T_241[9:0] ? 4'h2 : _GEN_16865; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16867 = 10'h2ce == _T_241[9:0] ? 4'h2 : _GEN_16866; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16868 = 10'h2cf == _T_241[9:0] ? 4'h2 : _GEN_16867; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16869 = 10'h2d0 == _T_241[9:0] ? 4'h2 : _GEN_16868; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16870 = 10'h2d1 == _T_241[9:0] ? 4'h2 : _GEN_16869; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16871 = 10'h2d2 == _T_241[9:0] ? 4'h7 : _GEN_16870; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16872 = 10'h2d3 == _T_241[9:0] ? 4'h7 : _GEN_16871; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16873 = 10'h2d4 == _T_241[9:0] ? 4'h8 : _GEN_16872; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16874 = 10'h2d5 == _T_241[9:0] ? 4'h8 : _GEN_16873; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16875 = 10'h2d6 == _T_241[9:0] ? 4'h8 : _GEN_16874; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16876 = 10'h2d7 == _T_241[9:0] ? 4'h8 : _GEN_16875; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16877 = 10'h2d8 == _T_241[9:0] ? 4'h7 : _GEN_16876; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16878 = 10'h2d9 == _T_241[9:0] ? 4'h6 : _GEN_16877; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16879 = 10'h2da == _T_241[9:0] ? 4'h4 : _GEN_16878; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16880 = 10'h2db == _T_241[9:0] ? 4'h2 : _GEN_16879; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16881 = 10'h2dc == _T_241[9:0] ? 4'h2 : _GEN_16880; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16882 = 10'h2dd == _T_241[9:0] ? 4'h3 : _GEN_16881; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16883 = 10'h2de == _T_241[9:0] ? 4'h3 : _GEN_16882; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16884 = 10'h2df == _T_241[9:0] ? 4'h3 : _GEN_16883; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16885 = 10'h2e0 == _T_241[9:0] ? 4'h3 : _GEN_16884; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16886 = 10'h2e1 == _T_241[9:0] ? 4'h3 : _GEN_16885; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16887 = 10'h2e2 == _T_241[9:0] ? 4'h3 : _GEN_16886; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16888 = 10'h2e3 == _T_241[9:0] ? 4'h2 : _GEN_16887; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16889 = 10'h2e4 == _T_241[9:0] ? 4'h3 : _GEN_16888; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16890 = 10'h2e5 == _T_241[9:0] ? 4'h2 : _GEN_16889; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16891 = 10'h2e6 == _T_241[9:0] ? 4'h5 : _GEN_16890; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16892 = 10'h2e7 == _T_241[9:0] ? 4'h5 : _GEN_16891; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16893 = 10'h2e8 == _T_241[9:0] ? 4'h5 : _GEN_16892; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16894 = 10'h2e9 == _T_241[9:0] ? 4'h5 : _GEN_16893; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16895 = 10'h2ea == _T_241[9:0] ? 4'h5 : _GEN_16894; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16896 = 10'h2eb == _T_241[9:0] ? 4'h5 : _GEN_16895; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16897 = 10'h2ec == _T_241[9:0] ? 4'h6 : _GEN_16896; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16898 = 10'h2ed == _T_241[9:0] ? 4'h7 : _GEN_16897; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16899 = 10'h2ee == _T_241[9:0] ? 4'h6 : _GEN_16898; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16900 = 10'h2ef == _T_241[9:0] ? 4'h2 : _GEN_16899; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16901 = 10'h2f0 == _T_241[9:0] ? 4'h2 : _GEN_16900; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16902 = 10'h2f1 == _T_241[9:0] ? 4'h2 : _GEN_16901; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16903 = 10'h2f2 == _T_241[9:0] ? 4'h2 : _GEN_16902; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16904 = 10'h2f3 == _T_241[9:0] ? 4'h2 : _GEN_16903; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16905 = 10'h2f4 == _T_241[9:0] ? 4'h2 : _GEN_16904; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16906 = 10'h2f5 == _T_241[9:0] ? 4'h2 : _GEN_16905; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16907 = 10'h2f6 == _T_241[9:0] ? 4'h2 : _GEN_16906; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16908 = 10'h2f7 == _T_241[9:0] ? 4'h2 : _GEN_16907; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16909 = 10'h2f8 == _T_241[9:0] ? 4'h7 : _GEN_16908; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16910 = 10'h2f9 == _T_241[9:0] ? 4'h7 : _GEN_16909; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16911 = 10'h2fa == _T_241[9:0] ? 4'h8 : _GEN_16910; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16912 = 10'h2fb == _T_241[9:0] ? 4'h8 : _GEN_16911; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16913 = 10'h2fc == _T_241[9:0] ? 4'h7 : _GEN_16912; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16914 = 10'h2fd == _T_241[9:0] ? 4'h7 : _GEN_16913; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16915 = 10'h2fe == _T_241[9:0] ? 4'h7 : _GEN_16914; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16916 = 10'h2ff == _T_241[9:0] ? 4'h7 : _GEN_16915; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16917 = 10'h300 == _T_241[9:0] ? 4'h8 : _GEN_16916; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16918 = 10'h301 == _T_241[9:0] ? 4'h7 : _GEN_16917; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16919 = 10'h302 == _T_241[9:0] ? 4'h3 : _GEN_16918; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16920 = 10'h303 == _T_241[9:0] ? 4'h3 : _GEN_16919; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16921 = 10'h304 == _T_241[9:0] ? 4'h2 : _GEN_16920; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16922 = 10'h305 == _T_241[9:0] ? 4'h2 : _GEN_16921; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16923 = 10'h306 == _T_241[9:0] ? 4'h2 : _GEN_16922; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16924 = 10'h307 == _T_241[9:0] ? 4'h2 : _GEN_16923; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16925 = 10'h308 == _T_241[9:0] ? 4'h2 : _GEN_16924; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16926 = 10'h309 == _T_241[9:0] ? 4'h2 : _GEN_16925; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16927 = 10'h30a == _T_241[9:0] ? 4'h2 : _GEN_16926; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16928 = 10'h30b == _T_241[9:0] ? 4'h3 : _GEN_16927; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16929 = 10'h30c == _T_241[9:0] ? 4'h4 : _GEN_16928; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16930 = 10'h30d == _T_241[9:0] ? 4'h5 : _GEN_16929; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16931 = 10'h30e == _T_241[9:0] ? 4'h5 : _GEN_16930; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16932 = 10'h30f == _T_241[9:0] ? 4'h5 : _GEN_16931; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16933 = 10'h310 == _T_241[9:0] ? 4'h5 : _GEN_16932; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16934 = 10'h311 == _T_241[9:0] ? 4'h5 : _GEN_16933; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16935 = 10'h312 == _T_241[9:0] ? 4'h6 : _GEN_16934; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16936 = 10'h313 == _T_241[9:0] ? 4'h7 : _GEN_16935; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16937 = 10'h314 == _T_241[9:0] ? 4'h7 : _GEN_16936; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16938 = 10'h315 == _T_241[9:0] ? 4'h3 : _GEN_16937; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16939 = 10'h316 == _T_241[9:0] ? 4'h2 : _GEN_16938; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16940 = 10'h317 == _T_241[9:0] ? 4'h2 : _GEN_16939; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16941 = 10'h318 == _T_241[9:0] ? 4'h2 : _GEN_16940; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16942 = 10'h319 == _T_241[9:0] ? 4'h2 : _GEN_16941; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16943 = 10'h31a == _T_241[9:0] ? 4'h2 : _GEN_16942; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16944 = 10'h31b == _T_241[9:0] ? 4'h2 : _GEN_16943; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16945 = 10'h31c == _T_241[9:0] ? 4'h2 : _GEN_16944; // @[Filter.scala 230:142]
  wire [3:0] _GEN_16946 = 10'h31d == _T_241[9:0] ? 4'h2 : _GEN_16945; // @[Filter.scala 230:142]
  wire [7:0] _T_255 = _GEN_16946 * 4'ha; // @[Filter.scala 230:142]
  wire [10:0] _GEN_38995 = {{3'd0}, _T_255}; // @[Filter.scala 230:109]
  wire [10:0] _T_257 = _T_250 + _GEN_38995; // @[Filter.scala 230:109]
  wire [10:0] _T_258 = _T_257 / 11'h64; // @[Filter.scala 230:150]
  wire  _T_260 = _T_231 >= 6'h20; // @[Filter.scala 233:31]
  wire  _T_264 = _T_238 >= 32'h12; // @[Filter.scala 233:63]
  wire  _T_265 = _T_260 | _T_264; // @[Filter.scala 233:58]
  wire [10:0] _GEN_17745 = io_SPI_distort ? _T_258 : {{7'd0}, _GEN_15350}; // @[Filter.scala 235:35]
  wire [10:0] _GEN_17746 = _T_265 ? 11'h0 : _GEN_17745; // @[Filter.scala 233:80]
  wire [10:0] _GEN_18545 = io_SPI_distort ? _T_258 : {{7'd0}, _GEN_16148}; // @[Filter.scala 235:35]
  wire [10:0] _GEN_18546 = _T_265 ? 11'h0 : _GEN_18545; // @[Filter.scala 233:80]
  wire [10:0] _GEN_19345 = io_SPI_distort ? _T_258 : {{7'd0}, _GEN_16946}; // @[Filter.scala 235:35]
  wire [10:0] _GEN_19346 = _T_265 ? 11'h0 : _GEN_19345; // @[Filter.scala 233:80]
  wire [31:0] _T_293 = pixelIndex + 32'h4; // @[Filter.scala 228:31]
  wire [31:0] _GEN_4 = _T_293 % 32'h20; // @[Filter.scala 228:38]
  wire [5:0] _T_294 = _GEN_4[5:0]; // @[Filter.scala 228:38]
  wire [5:0] _T_296 = _T_294 + _GEN_38951; // @[Filter.scala 228:53]
  wire [5:0] _T_298 = _T_296 - 6'h1; // @[Filter.scala 228:69]
  wire [31:0] _T_301 = _T_293 / 32'h20; // @[Filter.scala 229:38]
  wire [31:0] _T_303 = _T_301 + _GEN_38952; // @[Filter.scala 229:53]
  wire [31:0] _T_305 = _T_303 - 32'h1; // @[Filter.scala 229:69]
  wire [37:0] _T_306 = _T_305 * 32'h20; // @[Filter.scala 230:42]
  wire [37:0] _GEN_39001 = {{32'd0}, _T_298}; // @[Filter.scala 230:57]
  wire [37:0] _T_308 = _T_306 + _GEN_39001; // @[Filter.scala 230:57]
  wire [3:0] _GEN_19369 = 10'h16 == _T_308[9:0] ? 4'h9 : 4'ha; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19370 = 10'h17 == _T_308[9:0] ? 4'h3 : _GEN_19369; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19371 = 10'h18 == _T_308[9:0] ? 4'h6 : _GEN_19370; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19372 = 10'h19 == _T_308[9:0] ? 4'ha : _GEN_19371; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19373 = 10'h1a == _T_308[9:0] ? 4'ha : _GEN_19372; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19374 = 10'h1b == _T_308[9:0] ? 4'ha : _GEN_19373; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19375 = 10'h1c == _T_308[9:0] ? 4'ha : _GEN_19374; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19376 = 10'h1d == _T_308[9:0] ? 4'ha : _GEN_19375; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19377 = 10'h1e == _T_308[9:0] ? 4'ha : _GEN_19376; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19378 = 10'h1f == _T_308[9:0] ? 4'ha : _GEN_19377; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19379 = 10'h20 == _T_308[9:0] ? 4'ha : _GEN_19378; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19380 = 10'h21 == _T_308[9:0] ? 4'ha : _GEN_19379; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19381 = 10'h22 == _T_308[9:0] ? 4'ha : _GEN_19380; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19382 = 10'h23 == _T_308[9:0] ? 4'ha : _GEN_19381; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19383 = 10'h24 == _T_308[9:0] ? 4'ha : _GEN_19382; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19384 = 10'h25 == _T_308[9:0] ? 4'ha : _GEN_19383; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19385 = 10'h26 == _T_308[9:0] ? 4'ha : _GEN_19384; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19386 = 10'h27 == _T_308[9:0] ? 4'ha : _GEN_19385; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19387 = 10'h28 == _T_308[9:0] ? 4'ha : _GEN_19386; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19388 = 10'h29 == _T_308[9:0] ? 4'ha : _GEN_19387; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19389 = 10'h2a == _T_308[9:0] ? 4'ha : _GEN_19388; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19390 = 10'h2b == _T_308[9:0] ? 4'ha : _GEN_19389; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19391 = 10'h2c == _T_308[9:0] ? 4'ha : _GEN_19390; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19392 = 10'h2d == _T_308[9:0] ? 4'ha : _GEN_19391; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19393 = 10'h2e == _T_308[9:0] ? 4'ha : _GEN_19392; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19394 = 10'h2f == _T_308[9:0] ? 4'ha : _GEN_19393; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19395 = 10'h30 == _T_308[9:0] ? 4'ha : _GEN_19394; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19396 = 10'h31 == _T_308[9:0] ? 4'ha : _GEN_19395; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19397 = 10'h32 == _T_308[9:0] ? 4'ha : _GEN_19396; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19398 = 10'h33 == _T_308[9:0] ? 4'ha : _GEN_19397; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19399 = 10'h34 == _T_308[9:0] ? 4'ha : _GEN_19398; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19400 = 10'h35 == _T_308[9:0] ? 4'ha : _GEN_19399; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19401 = 10'h36 == _T_308[9:0] ? 4'ha : _GEN_19400; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19402 = 10'h37 == _T_308[9:0] ? 4'ha : _GEN_19401; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19403 = 10'h38 == _T_308[9:0] ? 4'ha : _GEN_19402; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19404 = 10'h39 == _T_308[9:0] ? 4'ha : _GEN_19403; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19405 = 10'h3a == _T_308[9:0] ? 4'ha : _GEN_19404; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19406 = 10'h3b == _T_308[9:0] ? 4'h9 : _GEN_19405; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19407 = 10'h3c == _T_308[9:0] ? 4'h4 : _GEN_19406; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19408 = 10'h3d == _T_308[9:0] ? 4'h3 : _GEN_19407; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19409 = 10'h3e == _T_308[9:0] ? 4'h4 : _GEN_19408; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19410 = 10'h3f == _T_308[9:0] ? 4'ha : _GEN_19409; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19411 = 10'h40 == _T_308[9:0] ? 4'ha : _GEN_19410; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19412 = 10'h41 == _T_308[9:0] ? 4'ha : _GEN_19411; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19413 = 10'h42 == _T_308[9:0] ? 4'ha : _GEN_19412; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19414 = 10'h43 == _T_308[9:0] ? 4'ha : _GEN_19413; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19415 = 10'h44 == _T_308[9:0] ? 4'ha : _GEN_19414; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19416 = 10'h45 == _T_308[9:0] ? 4'ha : _GEN_19415; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19417 = 10'h46 == _T_308[9:0] ? 4'ha : _GEN_19416; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19418 = 10'h47 == _T_308[9:0] ? 4'ha : _GEN_19417; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19419 = 10'h48 == _T_308[9:0] ? 4'ha : _GEN_19418; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19420 = 10'h49 == _T_308[9:0] ? 4'ha : _GEN_19419; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19421 = 10'h4a == _T_308[9:0] ? 4'ha : _GEN_19420; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19422 = 10'h4b == _T_308[9:0] ? 4'ha : _GEN_19421; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19423 = 10'h4c == _T_308[9:0] ? 4'ha : _GEN_19422; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19424 = 10'h4d == _T_308[9:0] ? 4'ha : _GEN_19423; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19425 = 10'h4e == _T_308[9:0] ? 4'ha : _GEN_19424; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19426 = 10'h4f == _T_308[9:0] ? 4'ha : _GEN_19425; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19427 = 10'h50 == _T_308[9:0] ? 4'ha : _GEN_19426; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19428 = 10'h51 == _T_308[9:0] ? 4'ha : _GEN_19427; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19429 = 10'h52 == _T_308[9:0] ? 4'ha : _GEN_19428; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19430 = 10'h53 == _T_308[9:0] ? 4'ha : _GEN_19429; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19431 = 10'h54 == _T_308[9:0] ? 4'ha : _GEN_19430; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19432 = 10'h55 == _T_308[9:0] ? 4'ha : _GEN_19431; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19433 = 10'h56 == _T_308[9:0] ? 4'ha : _GEN_19432; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19434 = 10'h57 == _T_308[9:0] ? 4'ha : _GEN_19433; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19435 = 10'h58 == _T_308[9:0] ? 4'ha : _GEN_19434; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19436 = 10'h59 == _T_308[9:0] ? 4'ha : _GEN_19435; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19437 = 10'h5a == _T_308[9:0] ? 4'h7 : _GEN_19436; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19438 = 10'h5b == _T_308[9:0] ? 4'h7 : _GEN_19437; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19439 = 10'h5c == _T_308[9:0] ? 4'ha : _GEN_19438; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19440 = 10'h5d == _T_308[9:0] ? 4'ha : _GEN_19439; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19441 = 10'h5e == _T_308[9:0] ? 4'ha : _GEN_19440; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19442 = 10'h5f == _T_308[9:0] ? 4'ha : _GEN_19441; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19443 = 10'h60 == _T_308[9:0] ? 4'ha : _GEN_19442; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19444 = 10'h61 == _T_308[9:0] ? 4'h8 : _GEN_19443; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19445 = 10'h62 == _T_308[9:0] ? 4'h3 : _GEN_19444; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19446 = 10'h63 == _T_308[9:0] ? 4'h3 : _GEN_19445; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19447 = 10'h64 == _T_308[9:0] ? 4'h3 : _GEN_19446; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19448 = 10'h65 == _T_308[9:0] ? 4'h9 : _GEN_19447; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19449 = 10'h66 == _T_308[9:0] ? 4'ha : _GEN_19448; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19450 = 10'h67 == _T_308[9:0] ? 4'ha : _GEN_19449; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19451 = 10'h68 == _T_308[9:0] ? 4'ha : _GEN_19450; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19452 = 10'h69 == _T_308[9:0] ? 4'ha : _GEN_19451; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19453 = 10'h6a == _T_308[9:0] ? 4'ha : _GEN_19452; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19454 = 10'h6b == _T_308[9:0] ? 4'h8 : _GEN_19453; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19455 = 10'h6c == _T_308[9:0] ? 4'h5 : _GEN_19454; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19456 = 10'h6d == _T_308[9:0] ? 4'h8 : _GEN_19455; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19457 = 10'h6e == _T_308[9:0] ? 4'ha : _GEN_19456; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19458 = 10'h6f == _T_308[9:0] ? 4'ha : _GEN_19457; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19459 = 10'h70 == _T_308[9:0] ? 4'ha : _GEN_19458; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19460 = 10'h71 == _T_308[9:0] ? 4'ha : _GEN_19459; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19461 = 10'h72 == _T_308[9:0] ? 4'ha : _GEN_19460; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19462 = 10'h73 == _T_308[9:0] ? 4'ha : _GEN_19461; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19463 = 10'h74 == _T_308[9:0] ? 4'ha : _GEN_19462; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19464 = 10'h75 == _T_308[9:0] ? 4'ha : _GEN_19463; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19465 = 10'h76 == _T_308[9:0] ? 4'ha : _GEN_19464; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19466 = 10'h77 == _T_308[9:0] ? 4'ha : _GEN_19465; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19467 = 10'h78 == _T_308[9:0] ? 4'ha : _GEN_19466; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19468 = 10'h79 == _T_308[9:0] ? 4'ha : _GEN_19467; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19469 = 10'h7a == _T_308[9:0] ? 4'ha : _GEN_19468; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19470 = 10'h7b == _T_308[9:0] ? 4'ha : _GEN_19469; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19471 = 10'h7c == _T_308[9:0] ? 4'ha : _GEN_19470; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19472 = 10'h7d == _T_308[9:0] ? 4'ha : _GEN_19471; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19473 = 10'h7e == _T_308[9:0] ? 4'ha : _GEN_19472; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19474 = 10'h7f == _T_308[9:0] ? 4'ha : _GEN_19473; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19475 = 10'h80 == _T_308[9:0] ? 4'ha : _GEN_19474; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19476 = 10'h81 == _T_308[9:0] ? 4'h5 : _GEN_19475; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19477 = 10'h82 == _T_308[9:0] ? 4'h5 : _GEN_19476; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19478 = 10'h83 == _T_308[9:0] ? 4'h7 : _GEN_19477; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19479 = 10'h84 == _T_308[9:0] ? 4'ha : _GEN_19478; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19480 = 10'h85 == _T_308[9:0] ? 4'ha : _GEN_19479; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19481 = 10'h86 == _T_308[9:0] ? 4'ha : _GEN_19480; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19482 = 10'h87 == _T_308[9:0] ? 4'h5 : _GEN_19481; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19483 = 10'h88 == _T_308[9:0] ? 4'h3 : _GEN_19482; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19484 = 10'h89 == _T_308[9:0] ? 4'h3 : _GEN_19483; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19485 = 10'h8a == _T_308[9:0] ? 4'h4 : _GEN_19484; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19486 = 10'h8b == _T_308[9:0] ? 4'h9 : _GEN_19485; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19487 = 10'h8c == _T_308[9:0] ? 4'ha : _GEN_19486; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19488 = 10'h8d == _T_308[9:0] ? 4'ha : _GEN_19487; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19489 = 10'h8e == _T_308[9:0] ? 4'ha : _GEN_19488; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19490 = 10'h8f == _T_308[9:0] ? 4'h6 : _GEN_19489; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19491 = 10'h90 == _T_308[9:0] ? 4'h4 : _GEN_19490; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19492 = 10'h91 == _T_308[9:0] ? 4'h3 : _GEN_19491; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19493 = 10'h92 == _T_308[9:0] ? 4'h7 : _GEN_19492; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19494 = 10'h93 == _T_308[9:0] ? 4'ha : _GEN_19493; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19495 = 10'h94 == _T_308[9:0] ? 4'ha : _GEN_19494; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19496 = 10'h95 == _T_308[9:0] ? 4'ha : _GEN_19495; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19497 = 10'h96 == _T_308[9:0] ? 4'ha : _GEN_19496; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19498 = 10'h97 == _T_308[9:0] ? 4'ha : _GEN_19497; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19499 = 10'h98 == _T_308[9:0] ? 4'ha : _GEN_19498; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19500 = 10'h99 == _T_308[9:0] ? 4'ha : _GEN_19499; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19501 = 10'h9a == _T_308[9:0] ? 4'ha : _GEN_19500; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19502 = 10'h9b == _T_308[9:0] ? 4'ha : _GEN_19501; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19503 = 10'h9c == _T_308[9:0] ? 4'ha : _GEN_19502; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19504 = 10'h9d == _T_308[9:0] ? 4'ha : _GEN_19503; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19505 = 10'h9e == _T_308[9:0] ? 4'ha : _GEN_19504; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19506 = 10'h9f == _T_308[9:0] ? 4'ha : _GEN_19505; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19507 = 10'ha0 == _T_308[9:0] ? 4'ha : _GEN_19506; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19508 = 10'ha1 == _T_308[9:0] ? 4'ha : _GEN_19507; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19509 = 10'ha2 == _T_308[9:0] ? 4'ha : _GEN_19508; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19510 = 10'ha3 == _T_308[9:0] ? 4'ha : _GEN_19509; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19511 = 10'ha4 == _T_308[9:0] ? 4'ha : _GEN_19510; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19512 = 10'ha5 == _T_308[9:0] ? 4'ha : _GEN_19511; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19513 = 10'ha6 == _T_308[9:0] ? 4'ha : _GEN_19512; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19514 = 10'ha7 == _T_308[9:0] ? 4'h9 : _GEN_19513; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19515 = 10'ha8 == _T_308[9:0] ? 4'h4 : _GEN_19514; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19516 = 10'ha9 == _T_308[9:0] ? 4'h3 : _GEN_19515; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19517 = 10'haa == _T_308[9:0] ? 4'h4 : _GEN_19516; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19518 = 10'hab == _T_308[9:0] ? 4'h7 : _GEN_19517; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19519 = 10'hac == _T_308[9:0] ? 4'h8 : _GEN_19518; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19520 = 10'had == _T_308[9:0] ? 4'h3 : _GEN_19519; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19521 = 10'hae == _T_308[9:0] ? 4'h3 : _GEN_19520; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19522 = 10'haf == _T_308[9:0] ? 4'h3 : _GEN_19521; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19523 = 10'hb0 == _T_308[9:0] ? 4'h3 : _GEN_19522; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19524 = 10'hb1 == _T_308[9:0] ? 4'h7 : _GEN_19523; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19525 = 10'hb2 == _T_308[9:0] ? 4'h9 : _GEN_19524; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19526 = 10'hb3 == _T_308[9:0] ? 4'h6 : _GEN_19525; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19527 = 10'hb4 == _T_308[9:0] ? 4'h4 : _GEN_19526; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19528 = 10'hb5 == _T_308[9:0] ? 4'h3 : _GEN_19527; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19529 = 10'hb6 == _T_308[9:0] ? 4'h3 : _GEN_19528; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19530 = 10'hb7 == _T_308[9:0] ? 4'h6 : _GEN_19529; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19531 = 10'hb8 == _T_308[9:0] ? 4'ha : _GEN_19530; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19532 = 10'hb9 == _T_308[9:0] ? 4'ha : _GEN_19531; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19533 = 10'hba == _T_308[9:0] ? 4'ha : _GEN_19532; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19534 = 10'hbb == _T_308[9:0] ? 4'ha : _GEN_19533; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19535 = 10'hbc == _T_308[9:0] ? 4'ha : _GEN_19534; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19536 = 10'hbd == _T_308[9:0] ? 4'h9 : _GEN_19535; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19537 = 10'hbe == _T_308[9:0] ? 4'ha : _GEN_19536; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19538 = 10'hbf == _T_308[9:0] ? 4'ha : _GEN_19537; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19539 = 10'hc0 == _T_308[9:0] ? 4'ha : _GEN_19538; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19540 = 10'hc1 == _T_308[9:0] ? 4'ha : _GEN_19539; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19541 = 10'hc2 == _T_308[9:0] ? 4'ha : _GEN_19540; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19542 = 10'hc3 == _T_308[9:0] ? 4'ha : _GEN_19541; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19543 = 10'hc4 == _T_308[9:0] ? 4'ha : _GEN_19542; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19544 = 10'hc5 == _T_308[9:0] ? 4'ha : _GEN_19543; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19545 = 10'hc6 == _T_308[9:0] ? 4'ha : _GEN_19544; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19546 = 10'hc7 == _T_308[9:0] ? 4'h9 : _GEN_19545; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19547 = 10'hc8 == _T_308[9:0] ? 4'h8 : _GEN_19546; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19548 = 10'hc9 == _T_308[9:0] ? 4'h8 : _GEN_19547; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19549 = 10'hca == _T_308[9:0] ? 4'h9 : _GEN_19548; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19550 = 10'hcb == _T_308[9:0] ? 4'ha : _GEN_19549; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19551 = 10'hcc == _T_308[9:0] ? 4'ha : _GEN_19550; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19552 = 10'hcd == _T_308[9:0] ? 4'ha : _GEN_19551; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19553 = 10'hce == _T_308[9:0] ? 4'h8 : _GEN_19552; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19554 = 10'hcf == _T_308[9:0] ? 4'h3 : _GEN_19553; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19555 = 10'hd0 == _T_308[9:0] ? 4'h3 : _GEN_19554; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19556 = 10'hd1 == _T_308[9:0] ? 4'h3 : _GEN_19555; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19557 = 10'hd2 == _T_308[9:0] ? 4'h4 : _GEN_19556; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19558 = 10'hd3 == _T_308[9:0] ? 4'h3 : _GEN_19557; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19559 = 10'hd4 == _T_308[9:0] ? 4'h3 : _GEN_19558; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19560 = 10'hd5 == _T_308[9:0] ? 4'h3 : _GEN_19559; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19561 = 10'hd6 == _T_308[9:0] ? 4'h3 : _GEN_19560; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19562 = 10'hd7 == _T_308[9:0] ? 4'h5 : _GEN_19561; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19563 = 10'hd8 == _T_308[9:0] ? 4'h4 : _GEN_19562; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19564 = 10'hd9 == _T_308[9:0] ? 4'h3 : _GEN_19563; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19565 = 10'hda == _T_308[9:0] ? 4'h3 : _GEN_19564; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19566 = 10'hdb == _T_308[9:0] ? 4'h3 : _GEN_19565; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19567 = 10'hdc == _T_308[9:0] ? 4'h4 : _GEN_19566; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19568 = 10'hdd == _T_308[9:0] ? 4'ha : _GEN_19567; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19569 = 10'hde == _T_308[9:0] ? 4'ha : _GEN_19568; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19570 = 10'hdf == _T_308[9:0] ? 4'ha : _GEN_19569; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19571 = 10'he0 == _T_308[9:0] ? 4'ha : _GEN_19570; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19572 = 10'he1 == _T_308[9:0] ? 4'ha : _GEN_19571; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19573 = 10'he2 == _T_308[9:0] ? 4'ha : _GEN_19572; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19574 = 10'he3 == _T_308[9:0] ? 4'h5 : _GEN_19573; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19575 = 10'he4 == _T_308[9:0] ? 4'ha : _GEN_19574; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19576 = 10'he5 == _T_308[9:0] ? 4'ha : _GEN_19575; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19577 = 10'he6 == _T_308[9:0] ? 4'ha : _GEN_19576; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19578 = 10'he7 == _T_308[9:0] ? 4'ha : _GEN_19577; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19579 = 10'he8 == _T_308[9:0] ? 4'ha : _GEN_19578; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19580 = 10'he9 == _T_308[9:0] ? 4'ha : _GEN_19579; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19581 = 10'hea == _T_308[9:0] ? 4'ha : _GEN_19580; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19582 = 10'heb == _T_308[9:0] ? 4'h9 : _GEN_19581; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19583 = 10'hec == _T_308[9:0] ? 4'h7 : _GEN_19582; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19584 = 10'hed == _T_308[9:0] ? 4'h3 : _GEN_19583; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19585 = 10'hee == _T_308[9:0] ? 4'h3 : _GEN_19584; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19586 = 10'hef == _T_308[9:0] ? 4'h3 : _GEN_19585; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19587 = 10'hf0 == _T_308[9:0] ? 4'h4 : _GEN_19586; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19588 = 10'hf1 == _T_308[9:0] ? 4'h7 : _GEN_19587; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19589 = 10'hf2 == _T_308[9:0] ? 4'ha : _GEN_19588; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19590 = 10'hf3 == _T_308[9:0] ? 4'ha : _GEN_19589; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19591 = 10'hf4 == _T_308[9:0] ? 4'ha : _GEN_19590; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19592 = 10'hf5 == _T_308[9:0] ? 4'h7 : _GEN_19591; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19593 = 10'hf6 == _T_308[9:0] ? 4'h3 : _GEN_19592; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19594 = 10'hf7 == _T_308[9:0] ? 4'h3 : _GEN_19593; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19595 = 10'hf8 == _T_308[9:0] ? 4'h3 : _GEN_19594; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19596 = 10'hf9 == _T_308[9:0] ? 4'h3 : _GEN_19595; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19597 = 10'hfa == _T_308[9:0] ? 4'h3 : _GEN_19596; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19598 = 10'hfb == _T_308[9:0] ? 4'h3 : _GEN_19597; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19599 = 10'hfc == _T_308[9:0] ? 4'h3 : _GEN_19598; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19600 = 10'hfd == _T_308[9:0] ? 4'h3 : _GEN_19599; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19601 = 10'hfe == _T_308[9:0] ? 4'h3 : _GEN_19600; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19602 = 10'hff == _T_308[9:0] ? 4'h3 : _GEN_19601; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19603 = 10'h100 == _T_308[9:0] ? 4'h3 : _GEN_19602; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19604 = 10'h101 == _T_308[9:0] ? 4'h4 : _GEN_19603; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19605 = 10'h102 == _T_308[9:0] ? 4'h6 : _GEN_19604; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19606 = 10'h103 == _T_308[9:0] ? 4'ha : _GEN_19605; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19607 = 10'h104 == _T_308[9:0] ? 4'ha : _GEN_19606; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19608 = 10'h105 == _T_308[9:0] ? 4'h9 : _GEN_19607; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19609 = 10'h106 == _T_308[9:0] ? 4'h9 : _GEN_19608; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19610 = 10'h107 == _T_308[9:0] ? 4'h9 : _GEN_19609; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19611 = 10'h108 == _T_308[9:0] ? 4'h9 : _GEN_19610; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19612 = 10'h109 == _T_308[9:0] ? 4'h3 : _GEN_19611; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19613 = 10'h10a == _T_308[9:0] ? 4'ha : _GEN_19612; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19614 = 10'h10b == _T_308[9:0] ? 4'ha : _GEN_19613; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19615 = 10'h10c == _T_308[9:0] ? 4'ha : _GEN_19614; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19616 = 10'h10d == _T_308[9:0] ? 4'ha : _GEN_19615; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19617 = 10'h10e == _T_308[9:0] ? 4'ha : _GEN_19616; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19618 = 10'h10f == _T_308[9:0] ? 4'h9 : _GEN_19617; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19619 = 10'h110 == _T_308[9:0] ? 4'h9 : _GEN_19618; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19620 = 10'h111 == _T_308[9:0] ? 4'h4 : _GEN_19619; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19621 = 10'h112 == _T_308[9:0] ? 4'h8 : _GEN_19620; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19622 = 10'h113 == _T_308[9:0] ? 4'h3 : _GEN_19621; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19623 = 10'h114 == _T_308[9:0] ? 4'h3 : _GEN_19622; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19624 = 10'h115 == _T_308[9:0] ? 4'h4 : _GEN_19623; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19625 = 10'h116 == _T_308[9:0] ? 4'h4 : _GEN_19624; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19626 = 10'h117 == _T_308[9:0] ? 4'h3 : _GEN_19625; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19627 = 10'h118 == _T_308[9:0] ? 4'h8 : _GEN_19626; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19628 = 10'h119 == _T_308[9:0] ? 4'ha : _GEN_19627; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19629 = 10'h11a == _T_308[9:0] ? 4'ha : _GEN_19628; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19630 = 10'h11b == _T_308[9:0] ? 4'ha : _GEN_19629; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19631 = 10'h11c == _T_308[9:0] ? 4'h6 : _GEN_19630; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19632 = 10'h11d == _T_308[9:0] ? 4'h3 : _GEN_19631; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19633 = 10'h11e == _T_308[9:0] ? 4'h3 : _GEN_19632; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19634 = 10'h11f == _T_308[9:0] ? 4'h3 : _GEN_19633; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19635 = 10'h120 == _T_308[9:0] ? 4'h3 : _GEN_19634; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19636 = 10'h121 == _T_308[9:0] ? 4'h3 : _GEN_19635; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19637 = 10'h122 == _T_308[9:0] ? 4'h3 : _GEN_19636; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19638 = 10'h123 == _T_308[9:0] ? 4'h3 : _GEN_19637; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19639 = 10'h124 == _T_308[9:0] ? 4'h3 : _GEN_19638; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19640 = 10'h125 == _T_308[9:0] ? 4'h3 : _GEN_19639; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19641 = 10'h126 == _T_308[9:0] ? 4'h4 : _GEN_19640; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19642 = 10'h127 == _T_308[9:0] ? 4'h6 : _GEN_19641; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19643 = 10'h128 == _T_308[9:0] ? 4'h5 : _GEN_19642; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19644 = 10'h129 == _T_308[9:0] ? 4'h8 : _GEN_19643; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19645 = 10'h12a == _T_308[9:0] ? 4'h5 : _GEN_19644; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19646 = 10'h12b == _T_308[9:0] ? 4'h3 : _GEN_19645; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19647 = 10'h12c == _T_308[9:0] ? 4'h3 : _GEN_19646; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19648 = 10'h12d == _T_308[9:0] ? 4'h3 : _GEN_19647; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19649 = 10'h12e == _T_308[9:0] ? 4'h4 : _GEN_19648; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19650 = 10'h12f == _T_308[9:0] ? 4'h4 : _GEN_19649; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19651 = 10'h130 == _T_308[9:0] ? 4'ha : _GEN_19650; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19652 = 10'h131 == _T_308[9:0] ? 4'h9 : _GEN_19651; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19653 = 10'h132 == _T_308[9:0] ? 4'h9 : _GEN_19652; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19654 = 10'h133 == _T_308[9:0] ? 4'h8 : _GEN_19653; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19655 = 10'h134 == _T_308[9:0] ? 4'h9 : _GEN_19654; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19656 = 10'h135 == _T_308[9:0] ? 4'h8 : _GEN_19655; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19657 = 10'h136 == _T_308[9:0] ? 4'h7 : _GEN_19656; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19658 = 10'h137 == _T_308[9:0] ? 4'h6 : _GEN_19657; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19659 = 10'h138 == _T_308[9:0] ? 4'h8 : _GEN_19658; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19660 = 10'h139 == _T_308[9:0] ? 4'h3 : _GEN_19659; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19661 = 10'h13a == _T_308[9:0] ? 4'h3 : _GEN_19660; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19662 = 10'h13b == _T_308[9:0] ? 4'h4 : _GEN_19661; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19663 = 10'h13c == _T_308[9:0] ? 4'h4 : _GEN_19662; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19664 = 10'h13d == _T_308[9:0] ? 4'h3 : _GEN_19663; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19665 = 10'h13e == _T_308[9:0] ? 4'h5 : _GEN_19664; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19666 = 10'h13f == _T_308[9:0] ? 4'h9 : _GEN_19665; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19667 = 10'h140 == _T_308[9:0] ? 4'ha : _GEN_19666; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19668 = 10'h141 == _T_308[9:0] ? 4'ha : _GEN_19667; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19669 = 10'h142 == _T_308[9:0] ? 4'ha : _GEN_19668; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19670 = 10'h143 == _T_308[9:0] ? 4'h5 : _GEN_19669; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19671 = 10'h144 == _T_308[9:0] ? 4'h3 : _GEN_19670; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19672 = 10'h145 == _T_308[9:0] ? 4'h3 : _GEN_19671; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19673 = 10'h146 == _T_308[9:0] ? 4'h3 : _GEN_19672; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19674 = 10'h147 == _T_308[9:0] ? 4'h4 : _GEN_19673; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19675 = 10'h148 == _T_308[9:0] ? 4'h3 : _GEN_19674; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19676 = 10'h149 == _T_308[9:0] ? 4'h3 : _GEN_19675; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19677 = 10'h14a == _T_308[9:0] ? 4'h3 : _GEN_19676; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19678 = 10'h14b == _T_308[9:0] ? 4'h6 : _GEN_19677; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19679 = 10'h14c == _T_308[9:0] ? 4'h8 : _GEN_19678; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19680 = 10'h14d == _T_308[9:0] ? 4'h5 : _GEN_19679; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19681 = 10'h14e == _T_308[9:0] ? 4'h4 : _GEN_19680; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19682 = 10'h14f == _T_308[9:0] ? 4'h3 : _GEN_19681; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19683 = 10'h150 == _T_308[9:0] ? 4'h3 : _GEN_19682; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19684 = 10'h151 == _T_308[9:0] ? 4'h3 : _GEN_19683; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19685 = 10'h152 == _T_308[9:0] ? 4'h3 : _GEN_19684; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19686 = 10'h153 == _T_308[9:0] ? 4'h3 : _GEN_19685; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19687 = 10'h154 == _T_308[9:0] ? 4'h3 : _GEN_19686; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19688 = 10'h155 == _T_308[9:0] ? 4'h4 : _GEN_19687; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19689 = 10'h156 == _T_308[9:0] ? 4'h9 : _GEN_19688; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19690 = 10'h157 == _T_308[9:0] ? 4'h8 : _GEN_19689; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19691 = 10'h158 == _T_308[9:0] ? 4'h8 : _GEN_19690; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19692 = 10'h159 == _T_308[9:0] ? 4'h8 : _GEN_19691; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19693 = 10'h15a == _T_308[9:0] ? 4'h8 : _GEN_19692; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19694 = 10'h15b == _T_308[9:0] ? 4'h8 : _GEN_19693; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19695 = 10'h15c == _T_308[9:0] ? 4'h7 : _GEN_19694; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19696 = 10'h15d == _T_308[9:0] ? 4'h7 : _GEN_19695; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19697 = 10'h15e == _T_308[9:0] ? 4'h8 : _GEN_19696; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19698 = 10'h15f == _T_308[9:0] ? 4'h3 : _GEN_19697; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19699 = 10'h160 == _T_308[9:0] ? 4'h4 : _GEN_19698; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19700 = 10'h161 == _T_308[9:0] ? 4'h4 : _GEN_19699; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19701 = 10'h162 == _T_308[9:0] ? 4'h4 : _GEN_19700; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19702 = 10'h163 == _T_308[9:0] ? 4'h4 : _GEN_19701; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19703 = 10'h164 == _T_308[9:0] ? 4'h5 : _GEN_19702; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19704 = 10'h165 == _T_308[9:0] ? 4'ha : _GEN_19703; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19705 = 10'h166 == _T_308[9:0] ? 4'h9 : _GEN_19704; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19706 = 10'h167 == _T_308[9:0] ? 4'ha : _GEN_19705; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19707 = 10'h168 == _T_308[9:0] ? 4'ha : _GEN_19706; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19708 = 10'h169 == _T_308[9:0] ? 4'h6 : _GEN_19707; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19709 = 10'h16a == _T_308[9:0] ? 4'h3 : _GEN_19708; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19710 = 10'h16b == _T_308[9:0] ? 4'h3 : _GEN_19709; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19711 = 10'h16c == _T_308[9:0] ? 4'h3 : _GEN_19710; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19712 = 10'h16d == _T_308[9:0] ? 4'h4 : _GEN_19711; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19713 = 10'h16e == _T_308[9:0] ? 4'h3 : _GEN_19712; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19714 = 10'h16f == _T_308[9:0] ? 4'h3 : _GEN_19713; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19715 = 10'h170 == _T_308[9:0] ? 4'h3 : _GEN_19714; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19716 = 10'h171 == _T_308[9:0] ? 4'h7 : _GEN_19715; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19717 = 10'h172 == _T_308[9:0] ? 4'ha : _GEN_19716; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19718 = 10'h173 == _T_308[9:0] ? 4'h5 : _GEN_19717; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19719 = 10'h174 == _T_308[9:0] ? 4'h3 : _GEN_19718; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19720 = 10'h175 == _T_308[9:0] ? 4'h4 : _GEN_19719; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19721 = 10'h176 == _T_308[9:0] ? 4'h4 : _GEN_19720; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19722 = 10'h177 == _T_308[9:0] ? 4'h4 : _GEN_19721; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19723 = 10'h178 == _T_308[9:0] ? 4'h4 : _GEN_19722; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19724 = 10'h179 == _T_308[9:0] ? 4'h3 : _GEN_19723; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19725 = 10'h17a == _T_308[9:0] ? 4'h3 : _GEN_19724; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19726 = 10'h17b == _T_308[9:0] ? 4'h3 : _GEN_19725; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19727 = 10'h17c == _T_308[9:0] ? 4'h8 : _GEN_19726; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19728 = 10'h17d == _T_308[9:0] ? 4'h8 : _GEN_19727; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19729 = 10'h17e == _T_308[9:0] ? 4'h8 : _GEN_19728; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19730 = 10'h17f == _T_308[9:0] ? 4'h8 : _GEN_19729; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19731 = 10'h180 == _T_308[9:0] ? 4'h8 : _GEN_19730; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19732 = 10'h181 == _T_308[9:0] ? 4'h8 : _GEN_19731; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19733 = 10'h182 == _T_308[9:0] ? 4'h8 : _GEN_19732; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19734 = 10'h183 == _T_308[9:0] ? 4'h8 : _GEN_19733; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19735 = 10'h184 == _T_308[9:0] ? 4'h8 : _GEN_19734; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19736 = 10'h185 == _T_308[9:0] ? 4'h5 : _GEN_19735; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19737 = 10'h186 == _T_308[9:0] ? 4'h3 : _GEN_19736; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19738 = 10'h187 == _T_308[9:0] ? 4'h4 : _GEN_19737; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19739 = 10'h188 == _T_308[9:0] ? 4'h4 : _GEN_19738; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19740 = 10'h189 == _T_308[9:0] ? 4'h4 : _GEN_19739; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19741 = 10'h18a == _T_308[9:0] ? 4'h5 : _GEN_19740; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19742 = 10'h18b == _T_308[9:0] ? 4'ha : _GEN_19741; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19743 = 10'h18c == _T_308[9:0] ? 4'ha : _GEN_19742; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19744 = 10'h18d == _T_308[9:0] ? 4'h9 : _GEN_19743; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19745 = 10'h18e == _T_308[9:0] ? 4'ha : _GEN_19744; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19746 = 10'h18f == _T_308[9:0] ? 4'h4 : _GEN_19745; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19747 = 10'h190 == _T_308[9:0] ? 4'h3 : _GEN_19746; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19748 = 10'h191 == _T_308[9:0] ? 4'h3 : _GEN_19747; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19749 = 10'h192 == _T_308[9:0] ? 4'h5 : _GEN_19748; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19750 = 10'h193 == _T_308[9:0] ? 4'h6 : _GEN_19749; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19751 = 10'h194 == _T_308[9:0] ? 4'h5 : _GEN_19750; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19752 = 10'h195 == _T_308[9:0] ? 4'h3 : _GEN_19751; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19753 = 10'h196 == _T_308[9:0] ? 4'h3 : _GEN_19752; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19754 = 10'h197 == _T_308[9:0] ? 4'h5 : _GEN_19753; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19755 = 10'h198 == _T_308[9:0] ? 4'ha : _GEN_19754; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19756 = 10'h199 == _T_308[9:0] ? 4'h3 : _GEN_19755; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19757 = 10'h19a == _T_308[9:0] ? 4'h1 : _GEN_19756; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19758 = 10'h19b == _T_308[9:0] ? 4'h2 : _GEN_19757; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19759 = 10'h19c == _T_308[9:0] ? 4'h4 : _GEN_19758; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19760 = 10'h19d == _T_308[9:0] ? 4'h3 : _GEN_19759; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19761 = 10'h19e == _T_308[9:0] ? 4'h1 : _GEN_19760; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19762 = 10'h19f == _T_308[9:0] ? 4'h2 : _GEN_19761; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19763 = 10'h1a0 == _T_308[9:0] ? 4'h3 : _GEN_19762; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19764 = 10'h1a1 == _T_308[9:0] ? 4'h4 : _GEN_19763; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19765 = 10'h1a2 == _T_308[9:0] ? 4'h8 : _GEN_19764; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19766 = 10'h1a3 == _T_308[9:0] ? 4'h8 : _GEN_19765; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19767 = 10'h1a4 == _T_308[9:0] ? 4'h8 : _GEN_19766; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19768 = 10'h1a5 == _T_308[9:0] ? 4'h8 : _GEN_19767; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19769 = 10'h1a6 == _T_308[9:0] ? 4'h7 : _GEN_19768; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19770 = 10'h1a7 == _T_308[9:0] ? 4'h8 : _GEN_19769; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19771 = 10'h1a8 == _T_308[9:0] ? 4'h8 : _GEN_19770; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19772 = 10'h1a9 == _T_308[9:0] ? 4'h8 : _GEN_19771; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19773 = 10'h1aa == _T_308[9:0] ? 4'h7 : _GEN_19772; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19774 = 10'h1ab == _T_308[9:0] ? 4'h4 : _GEN_19773; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19775 = 10'h1ac == _T_308[9:0] ? 4'h4 : _GEN_19774; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19776 = 10'h1ad == _T_308[9:0] ? 4'h3 : _GEN_19775; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19777 = 10'h1ae == _T_308[9:0] ? 4'h3 : _GEN_19776; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19778 = 10'h1af == _T_308[9:0] ? 4'h4 : _GEN_19777; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19779 = 10'h1b0 == _T_308[9:0] ? 4'h6 : _GEN_19778; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19780 = 10'h1b1 == _T_308[9:0] ? 4'ha : _GEN_19779; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19781 = 10'h1b2 == _T_308[9:0] ? 4'ha : _GEN_19780; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19782 = 10'h1b3 == _T_308[9:0] ? 4'h9 : _GEN_19781; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19783 = 10'h1b4 == _T_308[9:0] ? 4'h9 : _GEN_19782; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19784 = 10'h1b5 == _T_308[9:0] ? 4'h3 : _GEN_19783; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19785 = 10'h1b6 == _T_308[9:0] ? 4'h3 : _GEN_19784; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19786 = 10'h1b7 == _T_308[9:0] ? 4'h4 : _GEN_19785; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19787 = 10'h1b8 == _T_308[9:0] ? 4'h5 : _GEN_19786; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19788 = 10'h1b9 == _T_308[9:0] ? 4'h6 : _GEN_19787; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19789 = 10'h1ba == _T_308[9:0] ? 4'h4 : _GEN_19788; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19790 = 10'h1bb == _T_308[9:0] ? 4'h3 : _GEN_19789; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19791 = 10'h1bc == _T_308[9:0] ? 4'h3 : _GEN_19790; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19792 = 10'h1bd == _T_308[9:0] ? 4'h4 : _GEN_19791; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19793 = 10'h1be == _T_308[9:0] ? 4'ha : _GEN_19792; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19794 = 10'h1bf == _T_308[9:0] ? 4'h4 : _GEN_19793; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19795 = 10'h1c0 == _T_308[9:0] ? 4'h5 : _GEN_19794; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19796 = 10'h1c1 == _T_308[9:0] ? 4'h5 : _GEN_19795; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19797 = 10'h1c2 == _T_308[9:0] ? 4'h4 : _GEN_19796; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19798 = 10'h1c3 == _T_308[9:0] ? 4'h5 : _GEN_19797; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19799 = 10'h1c4 == _T_308[9:0] ? 4'h4 : _GEN_19798; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19800 = 10'h1c5 == _T_308[9:0] ? 4'h3 : _GEN_19799; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19801 = 10'h1c6 == _T_308[9:0] ? 4'h4 : _GEN_19800; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19802 = 10'h1c7 == _T_308[9:0] ? 4'h3 : _GEN_19801; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19803 = 10'h1c8 == _T_308[9:0] ? 4'h8 : _GEN_19802; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19804 = 10'h1c9 == _T_308[9:0] ? 4'h8 : _GEN_19803; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19805 = 10'h1ca == _T_308[9:0] ? 4'h8 : _GEN_19804; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19806 = 10'h1cb == _T_308[9:0] ? 4'h8 : _GEN_19805; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19807 = 10'h1cc == _T_308[9:0] ? 4'h8 : _GEN_19806; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19808 = 10'h1cd == _T_308[9:0] ? 4'h8 : _GEN_19807; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19809 = 10'h1ce == _T_308[9:0] ? 4'h8 : _GEN_19808; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19810 = 10'h1cf == _T_308[9:0] ? 4'h8 : _GEN_19809; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19811 = 10'h1d0 == _T_308[9:0] ? 4'h5 : _GEN_19810; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19812 = 10'h1d1 == _T_308[9:0] ? 4'h4 : _GEN_19811; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19813 = 10'h1d2 == _T_308[9:0] ? 4'h6 : _GEN_19812; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19814 = 10'h1d3 == _T_308[9:0] ? 4'h6 : _GEN_19813; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19815 = 10'h1d4 == _T_308[9:0] ? 4'h6 : _GEN_19814; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19816 = 10'h1d5 == _T_308[9:0] ? 4'h5 : _GEN_19815; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19817 = 10'h1d6 == _T_308[9:0] ? 4'h8 : _GEN_19816; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19818 = 10'h1d7 == _T_308[9:0] ? 4'ha : _GEN_19817; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19819 = 10'h1d8 == _T_308[9:0] ? 4'ha : _GEN_19818; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19820 = 10'h1d9 == _T_308[9:0] ? 4'ha : _GEN_19819; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19821 = 10'h1da == _T_308[9:0] ? 4'h6 : _GEN_19820; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19822 = 10'h1db == _T_308[9:0] ? 4'h3 : _GEN_19821; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19823 = 10'h1dc == _T_308[9:0] ? 4'h5 : _GEN_19822; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19824 = 10'h1dd == _T_308[9:0] ? 4'h2 : _GEN_19823; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19825 = 10'h1de == _T_308[9:0] ? 4'h5 : _GEN_19824; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19826 = 10'h1df == _T_308[9:0] ? 4'h5 : _GEN_19825; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19827 = 10'h1e0 == _T_308[9:0] ? 4'h5 : _GEN_19826; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19828 = 10'h1e1 == _T_308[9:0] ? 4'h3 : _GEN_19827; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19829 = 10'h1e2 == _T_308[9:0] ? 4'h3 : _GEN_19828; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19830 = 10'h1e3 == _T_308[9:0] ? 4'h3 : _GEN_19829; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19831 = 10'h1e4 == _T_308[9:0] ? 4'h9 : _GEN_19830; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19832 = 10'h1e5 == _T_308[9:0] ? 4'h4 : _GEN_19831; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19833 = 10'h1e6 == _T_308[9:0] ? 4'h4 : _GEN_19832; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19834 = 10'h1e7 == _T_308[9:0] ? 4'h4 : _GEN_19833; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19835 = 10'h1e8 == _T_308[9:0] ? 4'h4 : _GEN_19834; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19836 = 10'h1e9 == _T_308[9:0] ? 4'h4 : _GEN_19835; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19837 = 10'h1ea == _T_308[9:0] ? 4'h4 : _GEN_19836; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19838 = 10'h1eb == _T_308[9:0] ? 4'h4 : _GEN_19837; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19839 = 10'h1ec == _T_308[9:0] ? 4'h4 : _GEN_19838; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19840 = 10'h1ed == _T_308[9:0] ? 4'h4 : _GEN_19839; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19841 = 10'h1ee == _T_308[9:0] ? 4'h8 : _GEN_19840; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19842 = 10'h1ef == _T_308[9:0] ? 4'h8 : _GEN_19841; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19843 = 10'h1f0 == _T_308[9:0] ? 4'h8 : _GEN_19842; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19844 = 10'h1f1 == _T_308[9:0] ? 4'h8 : _GEN_19843; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19845 = 10'h1f2 == _T_308[9:0] ? 4'h8 : _GEN_19844; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19846 = 10'h1f3 == _T_308[9:0] ? 4'h8 : _GEN_19845; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19847 = 10'h1f4 == _T_308[9:0] ? 4'h9 : _GEN_19846; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19848 = 10'h1f5 == _T_308[9:0] ? 4'h9 : _GEN_19847; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19849 = 10'h1f6 == _T_308[9:0] ? 4'ha : _GEN_19848; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19850 = 10'h1f7 == _T_308[9:0] ? 4'h5 : _GEN_19849; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19851 = 10'h1f8 == _T_308[9:0] ? 4'h5 : _GEN_19850; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19852 = 10'h1f9 == _T_308[9:0] ? 4'h7 : _GEN_19851; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19853 = 10'h1fa == _T_308[9:0] ? 4'h7 : _GEN_19852; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19854 = 10'h1fb == _T_308[9:0] ? 4'h5 : _GEN_19853; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19855 = 10'h1fc == _T_308[9:0] ? 4'ha : _GEN_19854; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19856 = 10'h1fd == _T_308[9:0] ? 4'hb : _GEN_19855; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19857 = 10'h1fe == _T_308[9:0] ? 4'hb : _GEN_19856; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19858 = 10'h1ff == _T_308[9:0] ? 4'ha : _GEN_19857; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19859 = 10'h200 == _T_308[9:0] ? 4'h4 : _GEN_19858; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19860 = 10'h201 == _T_308[9:0] ? 4'h3 : _GEN_19859; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19861 = 10'h202 == _T_308[9:0] ? 4'h2 : _GEN_19860; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19862 = 10'h203 == _T_308[9:0] ? 4'h2 : _GEN_19861; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19863 = 10'h204 == _T_308[9:0] ? 4'h2 : _GEN_19862; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19864 = 10'h205 == _T_308[9:0] ? 4'h2 : _GEN_19863; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19865 = 10'h206 == _T_308[9:0] ? 4'h2 : _GEN_19864; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19866 = 10'h207 == _T_308[9:0] ? 4'h2 : _GEN_19865; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19867 = 10'h208 == _T_308[9:0] ? 4'h3 : _GEN_19866; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19868 = 10'h209 == _T_308[9:0] ? 4'h3 : _GEN_19867; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19869 = 10'h20a == _T_308[9:0] ? 4'h8 : _GEN_19868; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19870 = 10'h20b == _T_308[9:0] ? 4'h4 : _GEN_19869; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19871 = 10'h20c == _T_308[9:0] ? 4'h4 : _GEN_19870; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19872 = 10'h20d == _T_308[9:0] ? 4'h4 : _GEN_19871; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19873 = 10'h20e == _T_308[9:0] ? 4'h4 : _GEN_19872; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19874 = 10'h20f == _T_308[9:0] ? 4'h4 : _GEN_19873; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19875 = 10'h210 == _T_308[9:0] ? 4'h4 : _GEN_19874; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19876 = 10'h211 == _T_308[9:0] ? 4'h4 : _GEN_19875; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19877 = 10'h212 == _T_308[9:0] ? 4'h4 : _GEN_19876; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19878 = 10'h213 == _T_308[9:0] ? 4'h6 : _GEN_19877; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19879 = 10'h214 == _T_308[9:0] ? 4'h7 : _GEN_19878; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19880 = 10'h215 == _T_308[9:0] ? 4'h8 : _GEN_19879; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19881 = 10'h216 == _T_308[9:0] ? 4'h8 : _GEN_19880; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19882 = 10'h217 == _T_308[9:0] ? 4'h8 : _GEN_19881; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19883 = 10'h218 == _T_308[9:0] ? 4'h8 : _GEN_19882; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19884 = 10'h219 == _T_308[9:0] ? 4'h8 : _GEN_19883; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19885 = 10'h21a == _T_308[9:0] ? 4'h8 : _GEN_19884; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19886 = 10'h21b == _T_308[9:0] ? 4'h8 : _GEN_19885; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19887 = 10'h21c == _T_308[9:0] ? 4'ha : _GEN_19886; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19888 = 10'h21d == _T_308[9:0] ? 4'h9 : _GEN_19887; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19889 = 10'h21e == _T_308[9:0] ? 4'h6 : _GEN_19888; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19890 = 10'h21f == _T_308[9:0] ? 4'h4 : _GEN_19889; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19891 = 10'h220 == _T_308[9:0] ? 4'h4 : _GEN_19890; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19892 = 10'h221 == _T_308[9:0] ? 4'h5 : _GEN_19891; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19893 = 10'h222 == _T_308[9:0] ? 4'ha : _GEN_19892; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19894 = 10'h223 == _T_308[9:0] ? 4'ha : _GEN_19893; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19895 = 10'h224 == _T_308[9:0] ? 4'ha : _GEN_19894; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19896 = 10'h225 == _T_308[9:0] ? 4'h8 : _GEN_19895; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19897 = 10'h226 == _T_308[9:0] ? 4'h4 : _GEN_19896; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19898 = 10'h227 == _T_308[9:0] ? 4'h2 : _GEN_19897; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19899 = 10'h228 == _T_308[9:0] ? 4'h2 : _GEN_19898; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19900 = 10'h229 == _T_308[9:0] ? 4'h2 : _GEN_19899; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19901 = 10'h22a == _T_308[9:0] ? 4'h2 : _GEN_19900; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19902 = 10'h22b == _T_308[9:0] ? 4'h2 : _GEN_19901; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19903 = 10'h22c == _T_308[9:0] ? 4'h2 : _GEN_19902; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19904 = 10'h22d == _T_308[9:0] ? 4'h2 : _GEN_19903; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19905 = 10'h22e == _T_308[9:0] ? 4'h2 : _GEN_19904; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19906 = 10'h22f == _T_308[9:0] ? 4'h3 : _GEN_19905; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19907 = 10'h230 == _T_308[9:0] ? 4'h3 : _GEN_19906; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19908 = 10'h231 == _T_308[9:0] ? 4'h3 : _GEN_19907; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19909 = 10'h232 == _T_308[9:0] ? 4'h4 : _GEN_19908; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19910 = 10'h233 == _T_308[9:0] ? 4'h6 : _GEN_19909; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19911 = 10'h234 == _T_308[9:0] ? 4'h6 : _GEN_19910; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19912 = 10'h235 == _T_308[9:0] ? 4'h4 : _GEN_19911; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19913 = 10'h236 == _T_308[9:0] ? 4'h4 : _GEN_19912; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19914 = 10'h237 == _T_308[9:0] ? 4'h4 : _GEN_19913; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19915 = 10'h238 == _T_308[9:0] ? 4'h4 : _GEN_19914; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19916 = 10'h239 == _T_308[9:0] ? 4'h3 : _GEN_19915; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19917 = 10'h23a == _T_308[9:0] ? 4'h7 : _GEN_19916; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19918 = 10'h23b == _T_308[9:0] ? 4'h7 : _GEN_19917; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19919 = 10'h23c == _T_308[9:0] ? 4'h7 : _GEN_19918; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19920 = 10'h23d == _T_308[9:0] ? 4'h7 : _GEN_19919; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19921 = 10'h23e == _T_308[9:0] ? 4'h7 : _GEN_19920; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19922 = 10'h23f == _T_308[9:0] ? 4'h7 : _GEN_19921; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19923 = 10'h240 == _T_308[9:0] ? 4'h7 : _GEN_19922; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19924 = 10'h241 == _T_308[9:0] ? 4'h8 : _GEN_19923; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19925 = 10'h242 == _T_308[9:0] ? 4'ha : _GEN_19924; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19926 = 10'h243 == _T_308[9:0] ? 4'ha : _GEN_19925; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19927 = 10'h244 == _T_308[9:0] ? 4'ha : _GEN_19926; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19928 = 10'h245 == _T_308[9:0] ? 4'h8 : _GEN_19927; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19929 = 10'h246 == _T_308[9:0] ? 4'h7 : _GEN_19928; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19930 = 10'h247 == _T_308[9:0] ? 4'h8 : _GEN_19929; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19931 = 10'h248 == _T_308[9:0] ? 4'ha : _GEN_19930; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19932 = 10'h249 == _T_308[9:0] ? 4'ha : _GEN_19931; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19933 = 10'h24a == _T_308[9:0] ? 4'ha : _GEN_19932; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19934 = 10'h24b == _T_308[9:0] ? 4'h4 : _GEN_19933; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19935 = 10'h24c == _T_308[9:0] ? 4'h4 : _GEN_19934; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19936 = 10'h24d == _T_308[9:0] ? 4'h2 : _GEN_19935; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19937 = 10'h24e == _T_308[9:0] ? 4'h2 : _GEN_19936; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19938 = 10'h24f == _T_308[9:0] ? 4'h2 : _GEN_19937; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19939 = 10'h250 == _T_308[9:0] ? 4'h2 : _GEN_19938; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19940 = 10'h251 == _T_308[9:0] ? 4'h2 : _GEN_19939; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19941 = 10'h252 == _T_308[9:0] ? 4'h2 : _GEN_19940; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19942 = 10'h253 == _T_308[9:0] ? 4'h2 : _GEN_19941; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19943 = 10'h254 == _T_308[9:0] ? 4'h2 : _GEN_19942; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19944 = 10'h255 == _T_308[9:0] ? 4'h3 : _GEN_19943; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19945 = 10'h256 == _T_308[9:0] ? 4'h4 : _GEN_19944; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19946 = 10'h257 == _T_308[9:0] ? 4'h3 : _GEN_19945; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19947 = 10'h258 == _T_308[9:0] ? 4'h4 : _GEN_19946; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19948 = 10'h259 == _T_308[9:0] ? 4'h4 : _GEN_19947; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19949 = 10'h25a == _T_308[9:0] ? 4'h4 : _GEN_19948; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19950 = 10'h25b == _T_308[9:0] ? 4'h3 : _GEN_19949; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19951 = 10'h25c == _T_308[9:0] ? 4'h4 : _GEN_19950; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19952 = 10'h25d == _T_308[9:0] ? 4'h4 : _GEN_19951; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19953 = 10'h25e == _T_308[9:0] ? 4'h3 : _GEN_19952; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19954 = 10'h25f == _T_308[9:0] ? 4'h3 : _GEN_19953; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19955 = 10'h260 == _T_308[9:0] ? 4'h8 : _GEN_19954; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19956 = 10'h261 == _T_308[9:0] ? 4'h7 : _GEN_19955; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19957 = 10'h262 == _T_308[9:0] ? 4'h6 : _GEN_19956; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19958 = 10'h263 == _T_308[9:0] ? 4'h5 : _GEN_19957; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19959 = 10'h264 == _T_308[9:0] ? 4'h6 : _GEN_19958; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19960 = 10'h265 == _T_308[9:0] ? 4'h5 : _GEN_19959; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19961 = 10'h266 == _T_308[9:0] ? 4'h5 : _GEN_19960; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19962 = 10'h267 == _T_308[9:0] ? 4'h7 : _GEN_19961; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19963 = 10'h268 == _T_308[9:0] ? 4'ha : _GEN_19962; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19964 = 10'h269 == _T_308[9:0] ? 4'ha : _GEN_19963; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19965 = 10'h26a == _T_308[9:0] ? 4'ha : _GEN_19964; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19966 = 10'h26b == _T_308[9:0] ? 4'ha : _GEN_19965; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19967 = 10'h26c == _T_308[9:0] ? 4'ha : _GEN_19966; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19968 = 10'h26d == _T_308[9:0] ? 4'ha : _GEN_19967; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19969 = 10'h26e == _T_308[9:0] ? 4'ha : _GEN_19968; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19970 = 10'h26f == _T_308[9:0] ? 4'ha : _GEN_19969; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19971 = 10'h270 == _T_308[9:0] ? 4'h5 : _GEN_19970; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19972 = 10'h271 == _T_308[9:0] ? 4'h4 : _GEN_19971; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19973 = 10'h272 == _T_308[9:0] ? 4'h3 : _GEN_19972; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19974 = 10'h273 == _T_308[9:0] ? 4'h2 : _GEN_19973; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19975 = 10'h274 == _T_308[9:0] ? 4'h2 : _GEN_19974; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19976 = 10'h275 == _T_308[9:0] ? 4'h2 : _GEN_19975; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19977 = 10'h276 == _T_308[9:0] ? 4'h2 : _GEN_19976; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19978 = 10'h277 == _T_308[9:0] ? 4'h2 : _GEN_19977; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19979 = 10'h278 == _T_308[9:0] ? 4'h2 : _GEN_19978; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19980 = 10'h279 == _T_308[9:0] ? 4'h2 : _GEN_19979; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19981 = 10'h27a == _T_308[9:0] ? 4'h2 : _GEN_19980; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19982 = 10'h27b == _T_308[9:0] ? 4'h4 : _GEN_19981; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19983 = 10'h27c == _T_308[9:0] ? 4'h3 : _GEN_19982; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19984 = 10'h27d == _T_308[9:0] ? 4'h4 : _GEN_19983; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19985 = 10'h27e == _T_308[9:0] ? 4'h5 : _GEN_19984; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19986 = 10'h27f == _T_308[9:0] ? 4'h4 : _GEN_19985; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19987 = 10'h280 == _T_308[9:0] ? 4'h4 : _GEN_19986; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19988 = 10'h281 == _T_308[9:0] ? 4'h4 : _GEN_19987; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19989 = 10'h282 == _T_308[9:0] ? 4'h4 : _GEN_19988; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19990 = 10'h283 == _T_308[9:0] ? 4'h3 : _GEN_19989; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19991 = 10'h284 == _T_308[9:0] ? 4'h3 : _GEN_19990; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19992 = 10'h285 == _T_308[9:0] ? 4'h3 : _GEN_19991; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19993 = 10'h286 == _T_308[9:0] ? 4'h8 : _GEN_19992; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19994 = 10'h287 == _T_308[9:0] ? 4'h6 : _GEN_19993; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19995 = 10'h288 == _T_308[9:0] ? 4'h6 : _GEN_19994; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19996 = 10'h289 == _T_308[9:0] ? 4'h6 : _GEN_19995; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19997 = 10'h28a == _T_308[9:0] ? 4'h7 : _GEN_19996; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19998 = 10'h28b == _T_308[9:0] ? 4'h7 : _GEN_19997; // @[Filter.scala 230:62]
  wire [3:0] _GEN_19999 = 10'h28c == _T_308[9:0] ? 4'h6 : _GEN_19998; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20000 = 10'h28d == _T_308[9:0] ? 4'h6 : _GEN_19999; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20001 = 10'h28e == _T_308[9:0] ? 4'h4 : _GEN_20000; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20002 = 10'h28f == _T_308[9:0] ? 4'h7 : _GEN_20001; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20003 = 10'h290 == _T_308[9:0] ? 4'h9 : _GEN_20002; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20004 = 10'h291 == _T_308[9:0] ? 4'ha : _GEN_20003; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20005 = 10'h292 == _T_308[9:0] ? 4'ha : _GEN_20004; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20006 = 10'h293 == _T_308[9:0] ? 4'ha : _GEN_20005; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20007 = 10'h294 == _T_308[9:0] ? 4'h9 : _GEN_20006; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20008 = 10'h295 == _T_308[9:0] ? 4'h5 : _GEN_20007; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20009 = 10'h296 == _T_308[9:0] ? 4'h4 : _GEN_20008; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20010 = 10'h297 == _T_308[9:0] ? 4'h4 : _GEN_20009; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20011 = 10'h298 == _T_308[9:0] ? 4'h3 : _GEN_20010; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20012 = 10'h299 == _T_308[9:0] ? 4'h3 : _GEN_20011; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20013 = 10'h29a == _T_308[9:0] ? 4'h2 : _GEN_20012; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20014 = 10'h29b == _T_308[9:0] ? 4'h2 : _GEN_20013; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20015 = 10'h29c == _T_308[9:0] ? 4'h2 : _GEN_20014; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20016 = 10'h29d == _T_308[9:0] ? 4'h2 : _GEN_20015; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20017 = 10'h29e == _T_308[9:0] ? 4'h2 : _GEN_20016; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20018 = 10'h29f == _T_308[9:0] ? 4'h2 : _GEN_20017; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20019 = 10'h2a0 == _T_308[9:0] ? 4'h2 : _GEN_20018; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20020 = 10'h2a1 == _T_308[9:0] ? 4'h4 : _GEN_20019; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20021 = 10'h2a2 == _T_308[9:0] ? 4'h3 : _GEN_20020; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20022 = 10'h2a3 == _T_308[9:0] ? 4'h4 : _GEN_20021; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20023 = 10'h2a4 == _T_308[9:0] ? 4'h5 : _GEN_20022; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20024 = 10'h2a5 == _T_308[9:0] ? 4'h4 : _GEN_20023; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20025 = 10'h2a6 == _T_308[9:0] ? 4'h4 : _GEN_20024; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20026 = 10'h2a7 == _T_308[9:0] ? 4'h4 : _GEN_20025; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20027 = 10'h2a8 == _T_308[9:0] ? 4'h3 : _GEN_20026; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20028 = 10'h2a9 == _T_308[9:0] ? 4'h3 : _GEN_20027; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20029 = 10'h2aa == _T_308[9:0] ? 4'h3 : _GEN_20028; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20030 = 10'h2ab == _T_308[9:0] ? 4'h3 : _GEN_20029; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20031 = 10'h2ac == _T_308[9:0] ? 4'h8 : _GEN_20030; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20032 = 10'h2ad == _T_308[9:0] ? 4'h7 : _GEN_20031; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20033 = 10'h2ae == _T_308[9:0] ? 4'h5 : _GEN_20032; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20034 = 10'h2af == _T_308[9:0] ? 4'h6 : _GEN_20033; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20035 = 10'h2b0 == _T_308[9:0] ? 4'h7 : _GEN_20034; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20036 = 10'h2b1 == _T_308[9:0] ? 4'h6 : _GEN_20035; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20037 = 10'h2b2 == _T_308[9:0] ? 4'h6 : _GEN_20036; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20038 = 10'h2b3 == _T_308[9:0] ? 4'h6 : _GEN_20037; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20039 = 10'h2b4 == _T_308[9:0] ? 4'h3 : _GEN_20038; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20040 = 10'h2b5 == _T_308[9:0] ? 4'h3 : _GEN_20039; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20041 = 10'h2b6 == _T_308[9:0] ? 4'h3 : _GEN_20040; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20042 = 10'h2b7 == _T_308[9:0] ? 4'h4 : _GEN_20041; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20043 = 10'h2b8 == _T_308[9:0] ? 4'h6 : _GEN_20042; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20044 = 10'h2b9 == _T_308[9:0] ? 4'h9 : _GEN_20043; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20045 = 10'h2ba == _T_308[9:0] ? 4'h4 : _GEN_20044; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20046 = 10'h2bb == _T_308[9:0] ? 4'h3 : _GEN_20045; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20047 = 10'h2bc == _T_308[9:0] ? 4'h4 : _GEN_20046; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20048 = 10'h2bd == _T_308[9:0] ? 4'h3 : _GEN_20047; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20049 = 10'h2be == _T_308[9:0] ? 4'h3 : _GEN_20048; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20050 = 10'h2bf == _T_308[9:0] ? 4'h3 : _GEN_20049; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20051 = 10'h2c0 == _T_308[9:0] ? 4'h2 : _GEN_20050; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20052 = 10'h2c1 == _T_308[9:0] ? 4'h2 : _GEN_20051; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20053 = 10'h2c2 == _T_308[9:0] ? 4'h2 : _GEN_20052; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20054 = 10'h2c3 == _T_308[9:0] ? 4'h2 : _GEN_20053; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20055 = 10'h2c4 == _T_308[9:0] ? 4'h2 : _GEN_20054; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20056 = 10'h2c5 == _T_308[9:0] ? 4'h2 : _GEN_20055; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20057 = 10'h2c6 == _T_308[9:0] ? 4'h2 : _GEN_20056; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20058 = 10'h2c7 == _T_308[9:0] ? 4'h4 : _GEN_20057; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20059 = 10'h2c8 == _T_308[9:0] ? 4'h3 : _GEN_20058; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20060 = 10'h2c9 == _T_308[9:0] ? 4'h4 : _GEN_20059; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20061 = 10'h2ca == _T_308[9:0] ? 4'h5 : _GEN_20060; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20062 = 10'h2cb == _T_308[9:0] ? 4'h3 : _GEN_20061; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20063 = 10'h2cc == _T_308[9:0] ? 4'h3 : _GEN_20062; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20064 = 10'h2cd == _T_308[9:0] ? 4'h3 : _GEN_20063; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20065 = 10'h2ce == _T_308[9:0] ? 4'h3 : _GEN_20064; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20066 = 10'h2cf == _T_308[9:0] ? 4'h3 : _GEN_20065; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20067 = 10'h2d0 == _T_308[9:0] ? 4'h3 : _GEN_20066; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20068 = 10'h2d1 == _T_308[9:0] ? 4'h3 : _GEN_20067; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20069 = 10'h2d2 == _T_308[9:0] ? 4'h8 : _GEN_20068; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20070 = 10'h2d3 == _T_308[9:0] ? 4'h6 : _GEN_20069; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20071 = 10'h2d4 == _T_308[9:0] ? 4'h6 : _GEN_20070; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20072 = 10'h2d5 == _T_308[9:0] ? 4'h7 : _GEN_20071; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20073 = 10'h2d6 == _T_308[9:0] ? 4'h7 : _GEN_20072; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20074 = 10'h2d7 == _T_308[9:0] ? 4'h7 : _GEN_20073; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20075 = 10'h2d8 == _T_308[9:0] ? 4'h6 : _GEN_20074; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20076 = 10'h2d9 == _T_308[9:0] ? 4'h7 : _GEN_20075; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20077 = 10'h2da == _T_308[9:0] ? 4'h5 : _GEN_20076; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20078 = 10'h2db == _T_308[9:0] ? 4'h3 : _GEN_20077; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20079 = 10'h2dc == _T_308[9:0] ? 4'h3 : _GEN_20078; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20080 = 10'h2dd == _T_308[9:0] ? 4'h3 : _GEN_20079; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20081 = 10'h2de == _T_308[9:0] ? 4'h3 : _GEN_20080; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20082 = 10'h2df == _T_308[9:0] ? 4'h4 : _GEN_20081; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20083 = 10'h2e0 == _T_308[9:0] ? 4'h3 : _GEN_20082; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20084 = 10'h2e1 == _T_308[9:0] ? 4'h3 : _GEN_20083; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20085 = 10'h2e2 == _T_308[9:0] ? 4'h3 : _GEN_20084; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20086 = 10'h2e3 == _T_308[9:0] ? 4'h3 : _GEN_20085; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20087 = 10'h2e4 == _T_308[9:0] ? 4'h3 : _GEN_20086; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20088 = 10'h2e5 == _T_308[9:0] ? 4'h3 : _GEN_20087; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20089 = 10'h2e6 == _T_308[9:0] ? 4'h2 : _GEN_20088; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20090 = 10'h2e7 == _T_308[9:0] ? 4'h2 : _GEN_20089; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20091 = 10'h2e8 == _T_308[9:0] ? 4'h2 : _GEN_20090; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20092 = 10'h2e9 == _T_308[9:0] ? 4'h2 : _GEN_20091; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20093 = 10'h2ea == _T_308[9:0] ? 4'h2 : _GEN_20092; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20094 = 10'h2eb == _T_308[9:0] ? 4'h2 : _GEN_20093; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20095 = 10'h2ec == _T_308[9:0] ? 4'h3 : _GEN_20094; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20096 = 10'h2ed == _T_308[9:0] ? 4'h4 : _GEN_20095; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20097 = 10'h2ee == _T_308[9:0] ? 4'h3 : _GEN_20096; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20098 = 10'h2ef == _T_308[9:0] ? 4'h3 : _GEN_20097; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20099 = 10'h2f0 == _T_308[9:0] ? 4'h6 : _GEN_20098; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20100 = 10'h2f1 == _T_308[9:0] ? 4'h3 : _GEN_20099; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20101 = 10'h2f2 == _T_308[9:0] ? 4'h3 : _GEN_20100; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20102 = 10'h2f3 == _T_308[9:0] ? 4'h3 : _GEN_20101; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20103 = 10'h2f4 == _T_308[9:0] ? 4'h3 : _GEN_20102; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20104 = 10'h2f5 == _T_308[9:0] ? 4'h3 : _GEN_20103; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20105 = 10'h2f6 == _T_308[9:0] ? 4'h3 : _GEN_20104; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20106 = 10'h2f7 == _T_308[9:0] ? 4'h3 : _GEN_20105; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20107 = 10'h2f8 == _T_308[9:0] ? 4'h8 : _GEN_20106; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20108 = 10'h2f9 == _T_308[9:0] ? 4'h6 : _GEN_20107; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20109 = 10'h2fa == _T_308[9:0] ? 4'h7 : _GEN_20108; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20110 = 10'h2fb == _T_308[9:0] ? 4'h7 : _GEN_20109; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20111 = 10'h2fc == _T_308[9:0] ? 4'h6 : _GEN_20110; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20112 = 10'h2fd == _T_308[9:0] ? 4'h6 : _GEN_20111; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20113 = 10'h2fe == _T_308[9:0] ? 4'h6 : _GEN_20112; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20114 = 10'h2ff == _T_308[9:0] ? 4'h8 : _GEN_20113; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20115 = 10'h300 == _T_308[9:0] ? 4'h9 : _GEN_20114; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20116 = 10'h301 == _T_308[9:0] ? 4'h7 : _GEN_20115; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20117 = 10'h302 == _T_308[9:0] ? 4'h4 : _GEN_20116; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20118 = 10'h303 == _T_308[9:0] ? 4'h4 : _GEN_20117; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20119 = 10'h304 == _T_308[9:0] ? 4'h3 : _GEN_20118; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20120 = 10'h305 == _T_308[9:0] ? 4'h3 : _GEN_20119; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20121 = 10'h306 == _T_308[9:0] ? 4'h3 : _GEN_20120; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20122 = 10'h307 == _T_308[9:0] ? 4'h3 : _GEN_20121; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20123 = 10'h308 == _T_308[9:0] ? 4'h3 : _GEN_20122; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20124 = 10'h309 == _T_308[9:0] ? 4'h3 : _GEN_20123; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20125 = 10'h30a == _T_308[9:0] ? 4'h3 : _GEN_20124; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20126 = 10'h30b == _T_308[9:0] ? 4'h3 : _GEN_20125; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20127 = 10'h30c == _T_308[9:0] ? 4'h2 : _GEN_20126; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20128 = 10'h30d == _T_308[9:0] ? 4'h2 : _GEN_20127; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20129 = 10'h30e == _T_308[9:0] ? 4'h2 : _GEN_20128; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20130 = 10'h30f == _T_308[9:0] ? 4'h2 : _GEN_20129; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20131 = 10'h310 == _T_308[9:0] ? 4'h2 : _GEN_20130; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20132 = 10'h311 == _T_308[9:0] ? 4'h2 : _GEN_20131; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20133 = 10'h312 == _T_308[9:0] ? 4'h3 : _GEN_20132; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20134 = 10'h313 == _T_308[9:0] ? 4'h4 : _GEN_20133; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20135 = 10'h314 == _T_308[9:0] ? 4'h3 : _GEN_20134; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20136 = 10'h315 == _T_308[9:0] ? 4'h3 : _GEN_20135; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20137 = 10'h316 == _T_308[9:0] ? 4'h5 : _GEN_20136; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20138 = 10'h317 == _T_308[9:0] ? 4'h5 : _GEN_20137; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20139 = 10'h318 == _T_308[9:0] ? 4'h3 : _GEN_20138; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20140 = 10'h319 == _T_308[9:0] ? 4'h3 : _GEN_20139; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20141 = 10'h31a == _T_308[9:0] ? 4'h3 : _GEN_20140; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20142 = 10'h31b == _T_308[9:0] ? 4'h3 : _GEN_20141; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20143 = 10'h31c == _T_308[9:0] ? 4'h3 : _GEN_20142; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20144 = 10'h31d == _T_308[9:0] ? 4'h3 : _GEN_20143; // @[Filter.scala 230:62]
  wire [4:0] _GEN_39002 = {{1'd0}, _GEN_20144}; // @[Filter.scala 230:62]
  wire [8:0] _T_310 = _GEN_39002 * 5'h14; // @[Filter.scala 230:62]
  wire [3:0] _GEN_20168 = 10'h17 == _T_308[9:0] ? 4'hb : 4'he; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20169 = 10'h18 == _T_308[9:0] ? 4'hc : _GEN_20168; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20170 = 10'h19 == _T_308[9:0] ? 4'he : _GEN_20169; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20171 = 10'h1a == _T_308[9:0] ? 4'he : _GEN_20170; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20172 = 10'h1b == _T_308[9:0] ? 4'he : _GEN_20171; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20173 = 10'h1c == _T_308[9:0] ? 4'he : _GEN_20172; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20174 = 10'h1d == _T_308[9:0] ? 4'he : _GEN_20173; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20175 = 10'h1e == _T_308[9:0] ? 4'he : _GEN_20174; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20176 = 10'h1f == _T_308[9:0] ? 4'he : _GEN_20175; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20177 = 10'h20 == _T_308[9:0] ? 4'he : _GEN_20176; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20178 = 10'h21 == _T_308[9:0] ? 4'he : _GEN_20177; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20179 = 10'h22 == _T_308[9:0] ? 4'he : _GEN_20178; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20180 = 10'h23 == _T_308[9:0] ? 4'he : _GEN_20179; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20181 = 10'h24 == _T_308[9:0] ? 4'he : _GEN_20180; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20182 = 10'h25 == _T_308[9:0] ? 4'he : _GEN_20181; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20183 = 10'h26 == _T_308[9:0] ? 4'he : _GEN_20182; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20184 = 10'h27 == _T_308[9:0] ? 4'he : _GEN_20183; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20185 = 10'h28 == _T_308[9:0] ? 4'he : _GEN_20184; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20186 = 10'h29 == _T_308[9:0] ? 4'he : _GEN_20185; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20187 = 10'h2a == _T_308[9:0] ? 4'he : _GEN_20186; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20188 = 10'h2b == _T_308[9:0] ? 4'he : _GEN_20187; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20189 = 10'h2c == _T_308[9:0] ? 4'he : _GEN_20188; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20190 = 10'h2d == _T_308[9:0] ? 4'he : _GEN_20189; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20191 = 10'h2e == _T_308[9:0] ? 4'he : _GEN_20190; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20192 = 10'h2f == _T_308[9:0] ? 4'he : _GEN_20191; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20193 = 10'h30 == _T_308[9:0] ? 4'he : _GEN_20192; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20194 = 10'h31 == _T_308[9:0] ? 4'he : _GEN_20193; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20195 = 10'h32 == _T_308[9:0] ? 4'he : _GEN_20194; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20196 = 10'h33 == _T_308[9:0] ? 4'he : _GEN_20195; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20197 = 10'h34 == _T_308[9:0] ? 4'he : _GEN_20196; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20198 = 10'h35 == _T_308[9:0] ? 4'he : _GEN_20197; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20199 = 10'h36 == _T_308[9:0] ? 4'he : _GEN_20198; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20200 = 10'h37 == _T_308[9:0] ? 4'he : _GEN_20199; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20201 = 10'h38 == _T_308[9:0] ? 4'he : _GEN_20200; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20202 = 10'h39 == _T_308[9:0] ? 4'he : _GEN_20201; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20203 = 10'h3a == _T_308[9:0] ? 4'he : _GEN_20202; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20204 = 10'h3b == _T_308[9:0] ? 4'he : _GEN_20203; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20205 = 10'h3c == _T_308[9:0] ? 4'ha : _GEN_20204; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20206 = 10'h3d == _T_308[9:0] ? 4'hc : _GEN_20205; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20207 = 10'h3e == _T_308[9:0] ? 4'hb : _GEN_20206; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20208 = 10'h3f == _T_308[9:0] ? 4'he : _GEN_20207; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20209 = 10'h40 == _T_308[9:0] ? 4'he : _GEN_20208; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20210 = 10'h41 == _T_308[9:0] ? 4'he : _GEN_20209; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20211 = 10'h42 == _T_308[9:0] ? 4'he : _GEN_20210; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20212 = 10'h43 == _T_308[9:0] ? 4'he : _GEN_20211; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20213 = 10'h44 == _T_308[9:0] ? 4'he : _GEN_20212; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20214 = 10'h45 == _T_308[9:0] ? 4'he : _GEN_20213; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20215 = 10'h46 == _T_308[9:0] ? 4'he : _GEN_20214; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20216 = 10'h47 == _T_308[9:0] ? 4'he : _GEN_20215; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20217 = 10'h48 == _T_308[9:0] ? 4'he : _GEN_20216; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20218 = 10'h49 == _T_308[9:0] ? 4'he : _GEN_20217; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20219 = 10'h4a == _T_308[9:0] ? 4'he : _GEN_20218; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20220 = 10'h4b == _T_308[9:0] ? 4'he : _GEN_20219; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20221 = 10'h4c == _T_308[9:0] ? 4'he : _GEN_20220; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20222 = 10'h4d == _T_308[9:0] ? 4'he : _GEN_20221; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20223 = 10'h4e == _T_308[9:0] ? 4'he : _GEN_20222; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20224 = 10'h4f == _T_308[9:0] ? 4'he : _GEN_20223; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20225 = 10'h50 == _T_308[9:0] ? 4'he : _GEN_20224; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20226 = 10'h51 == _T_308[9:0] ? 4'he : _GEN_20225; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20227 = 10'h52 == _T_308[9:0] ? 4'he : _GEN_20226; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20228 = 10'h53 == _T_308[9:0] ? 4'he : _GEN_20227; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20229 = 10'h54 == _T_308[9:0] ? 4'he : _GEN_20228; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20230 = 10'h55 == _T_308[9:0] ? 4'he : _GEN_20229; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20231 = 10'h56 == _T_308[9:0] ? 4'he : _GEN_20230; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20232 = 10'h57 == _T_308[9:0] ? 4'he : _GEN_20231; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20233 = 10'h58 == _T_308[9:0] ? 4'he : _GEN_20232; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20234 = 10'h59 == _T_308[9:0] ? 4'he : _GEN_20233; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20235 = 10'h5a == _T_308[9:0] ? 4'hc : _GEN_20234; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20236 = 10'h5b == _T_308[9:0] ? 4'hd : _GEN_20235; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20237 = 10'h5c == _T_308[9:0] ? 4'he : _GEN_20236; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20238 = 10'h5d == _T_308[9:0] ? 4'he : _GEN_20237; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20239 = 10'h5e == _T_308[9:0] ? 4'he : _GEN_20238; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20240 = 10'h5f == _T_308[9:0] ? 4'he : _GEN_20239; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20241 = 10'h60 == _T_308[9:0] ? 4'he : _GEN_20240; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20242 = 10'h61 == _T_308[9:0] ? 4'hd : _GEN_20241; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20243 = 10'h62 == _T_308[9:0] ? 4'hb : _GEN_20242; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20244 = 10'h63 == _T_308[9:0] ? 4'hc : _GEN_20243; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20245 = 10'h64 == _T_308[9:0] ? 4'ha : _GEN_20244; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20246 = 10'h65 == _T_308[9:0] ? 4'hd : _GEN_20245; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20247 = 10'h66 == _T_308[9:0] ? 4'he : _GEN_20246; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20248 = 10'h67 == _T_308[9:0] ? 4'he : _GEN_20247; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20249 = 10'h68 == _T_308[9:0] ? 4'he : _GEN_20248; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20250 = 10'h69 == _T_308[9:0] ? 4'he : _GEN_20249; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20251 = 10'h6a == _T_308[9:0] ? 4'he : _GEN_20250; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20252 = 10'h6b == _T_308[9:0] ? 4'hd : _GEN_20251; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20253 = 10'h6c == _T_308[9:0] ? 4'hc : _GEN_20252; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20254 = 10'h6d == _T_308[9:0] ? 4'hc : _GEN_20253; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20255 = 10'h6e == _T_308[9:0] ? 4'he : _GEN_20254; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20256 = 10'h6f == _T_308[9:0] ? 4'he : _GEN_20255; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20257 = 10'h70 == _T_308[9:0] ? 4'he : _GEN_20256; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20258 = 10'h71 == _T_308[9:0] ? 4'he : _GEN_20257; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20259 = 10'h72 == _T_308[9:0] ? 4'he : _GEN_20258; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20260 = 10'h73 == _T_308[9:0] ? 4'he : _GEN_20259; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20261 = 10'h74 == _T_308[9:0] ? 4'he : _GEN_20260; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20262 = 10'h75 == _T_308[9:0] ? 4'he : _GEN_20261; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20263 = 10'h76 == _T_308[9:0] ? 4'he : _GEN_20262; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20264 = 10'h77 == _T_308[9:0] ? 4'he : _GEN_20263; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20265 = 10'h78 == _T_308[9:0] ? 4'he : _GEN_20264; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20266 = 10'h79 == _T_308[9:0] ? 4'he : _GEN_20265; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20267 = 10'h7a == _T_308[9:0] ? 4'he : _GEN_20266; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20268 = 10'h7b == _T_308[9:0] ? 4'he : _GEN_20267; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20269 = 10'h7c == _T_308[9:0] ? 4'he : _GEN_20268; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20270 = 10'h7d == _T_308[9:0] ? 4'he : _GEN_20269; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20271 = 10'h7e == _T_308[9:0] ? 4'he : _GEN_20270; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20272 = 10'h7f == _T_308[9:0] ? 4'he : _GEN_20271; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20273 = 10'h80 == _T_308[9:0] ? 4'he : _GEN_20272; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20274 = 10'h81 == _T_308[9:0] ? 4'hb : _GEN_20273; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20275 = 10'h82 == _T_308[9:0] ? 4'hc : _GEN_20274; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20276 = 10'h83 == _T_308[9:0] ? 4'hc : _GEN_20275; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20277 = 10'h84 == _T_308[9:0] ? 4'he : _GEN_20276; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20278 = 10'h85 == _T_308[9:0] ? 4'he : _GEN_20277; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20279 = 10'h86 == _T_308[9:0] ? 4'he : _GEN_20278; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20280 = 10'h87 == _T_308[9:0] ? 4'ha : _GEN_20279; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20281 = 10'h88 == _T_308[9:0] ? 4'hd : _GEN_20280; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20282 = 10'h89 == _T_308[9:0] ? 4'hd : _GEN_20281; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20283 = 10'h8a == _T_308[9:0] ? 4'hc : _GEN_20282; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20284 = 10'h8b == _T_308[9:0] ? 4'he : _GEN_20283; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20285 = 10'h8c == _T_308[9:0] ? 4'he : _GEN_20284; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20286 = 10'h8d == _T_308[9:0] ? 4'he : _GEN_20285; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20287 = 10'h8e == _T_308[9:0] ? 4'he : _GEN_20286; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20288 = 10'h8f == _T_308[9:0] ? 4'hb : _GEN_20287; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20289 = 10'h90 == _T_308[9:0] ? 4'hc : _GEN_20288; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20290 = 10'h91 == _T_308[9:0] ? 4'hc : _GEN_20289; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20291 = 10'h92 == _T_308[9:0] ? 4'hd : _GEN_20290; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20292 = 10'h93 == _T_308[9:0] ? 4'he : _GEN_20291; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20293 = 10'h94 == _T_308[9:0] ? 4'he : _GEN_20292; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20294 = 10'h95 == _T_308[9:0] ? 4'he : _GEN_20293; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20295 = 10'h96 == _T_308[9:0] ? 4'he : _GEN_20294; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20296 = 10'h97 == _T_308[9:0] ? 4'he : _GEN_20295; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20297 = 10'h98 == _T_308[9:0] ? 4'he : _GEN_20296; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20298 = 10'h99 == _T_308[9:0] ? 4'he : _GEN_20297; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20299 = 10'h9a == _T_308[9:0] ? 4'he : _GEN_20298; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20300 = 10'h9b == _T_308[9:0] ? 4'he : _GEN_20299; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20301 = 10'h9c == _T_308[9:0] ? 4'he : _GEN_20300; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20302 = 10'h9d == _T_308[9:0] ? 4'he : _GEN_20301; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20303 = 10'h9e == _T_308[9:0] ? 4'he : _GEN_20302; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20304 = 10'h9f == _T_308[9:0] ? 4'he : _GEN_20303; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20305 = 10'ha0 == _T_308[9:0] ? 4'he : _GEN_20304; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20306 = 10'ha1 == _T_308[9:0] ? 4'he : _GEN_20305; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20307 = 10'ha2 == _T_308[9:0] ? 4'he : _GEN_20306; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20308 = 10'ha3 == _T_308[9:0] ? 4'he : _GEN_20307; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20309 = 10'ha4 == _T_308[9:0] ? 4'he : _GEN_20308; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20310 = 10'ha5 == _T_308[9:0] ? 4'he : _GEN_20309; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20311 = 10'ha6 == _T_308[9:0] ? 4'he : _GEN_20310; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20312 = 10'ha7 == _T_308[9:0] ? 4'he : _GEN_20311; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20313 = 10'ha8 == _T_308[9:0] ? 4'hb : _GEN_20312; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20314 = 10'ha9 == _T_308[9:0] ? 4'hc : _GEN_20313; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20315 = 10'haa == _T_308[9:0] ? 4'hb : _GEN_20314; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20316 = 10'hab == _T_308[9:0] ? 4'hc : _GEN_20315; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20317 = 10'hac == _T_308[9:0] ? 4'hd : _GEN_20316; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20318 = 10'had == _T_308[9:0] ? 4'ha : _GEN_20317; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20319 = 10'hae == _T_308[9:0] ? 4'hd : _GEN_20318; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20320 = 10'haf == _T_308[9:0] ? 4'hd : _GEN_20319; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20321 = 10'hb0 == _T_308[9:0] ? 4'hb : _GEN_20320; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20322 = 10'hb1 == _T_308[9:0] ? 4'hc : _GEN_20321; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20323 = 10'hb2 == _T_308[9:0] ? 4'he : _GEN_20322; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20324 = 10'hb3 == _T_308[9:0] ? 4'hb : _GEN_20323; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20325 = 10'hb4 == _T_308[9:0] ? 4'hc : _GEN_20324; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20326 = 10'hb5 == _T_308[9:0] ? 4'hd : _GEN_20325; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20327 = 10'hb6 == _T_308[9:0] ? 4'hd : _GEN_20326; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20328 = 10'hb7 == _T_308[9:0] ? 4'hc : _GEN_20327; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20329 = 10'hb8 == _T_308[9:0] ? 4'he : _GEN_20328; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20330 = 10'hb9 == _T_308[9:0] ? 4'he : _GEN_20329; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20331 = 10'hba == _T_308[9:0] ? 4'he : _GEN_20330; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20332 = 10'hbb == _T_308[9:0] ? 4'he : _GEN_20331; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20333 = 10'hbc == _T_308[9:0] ? 4'he : _GEN_20332; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20334 = 10'hbd == _T_308[9:0] ? 4'he : _GEN_20333; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20335 = 10'hbe == _T_308[9:0] ? 4'he : _GEN_20334; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20336 = 10'hbf == _T_308[9:0] ? 4'he : _GEN_20335; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20337 = 10'hc0 == _T_308[9:0] ? 4'he : _GEN_20336; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20338 = 10'hc1 == _T_308[9:0] ? 4'he : _GEN_20337; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20339 = 10'hc2 == _T_308[9:0] ? 4'he : _GEN_20338; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20340 = 10'hc3 == _T_308[9:0] ? 4'he : _GEN_20339; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20341 = 10'hc4 == _T_308[9:0] ? 4'he : _GEN_20340; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20342 = 10'hc5 == _T_308[9:0] ? 4'he : _GEN_20341; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20343 = 10'hc6 == _T_308[9:0] ? 4'he : _GEN_20342; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20344 = 10'hc7 == _T_308[9:0] ? 4'hd : _GEN_20343; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20345 = 10'hc8 == _T_308[9:0] ? 4'hb : _GEN_20344; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20346 = 10'hc9 == _T_308[9:0] ? 4'hc : _GEN_20345; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20347 = 10'hca == _T_308[9:0] ? 4'he : _GEN_20346; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20348 = 10'hcb == _T_308[9:0] ? 4'he : _GEN_20347; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20349 = 10'hcc == _T_308[9:0] ? 4'he : _GEN_20348; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20350 = 10'hcd == _T_308[9:0] ? 4'he : _GEN_20349; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20351 = 10'hce == _T_308[9:0] ? 4'hd : _GEN_20350; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20352 = 10'hcf == _T_308[9:0] ? 4'hb : _GEN_20351; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20353 = 10'hd0 == _T_308[9:0] ? 4'hc : _GEN_20352; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20354 = 10'hd1 == _T_308[9:0] ? 4'hc : _GEN_20353; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20355 = 10'hd2 == _T_308[9:0] ? 4'hb : _GEN_20354; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20356 = 10'hd3 == _T_308[9:0] ? 4'hd : _GEN_20355; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20357 = 10'hd4 == _T_308[9:0] ? 4'hd : _GEN_20356; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20358 = 10'hd5 == _T_308[9:0] ? 4'hd : _GEN_20357; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20359 = 10'hd6 == _T_308[9:0] ? 4'hd : _GEN_20358; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20360 = 10'hd7 == _T_308[9:0] ? 4'hc : _GEN_20359; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20361 = 10'hd8 == _T_308[9:0] ? 4'hc : _GEN_20360; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20362 = 10'hd9 == _T_308[9:0] ? 4'hc : _GEN_20361; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20363 = 10'hda == _T_308[9:0] ? 4'hd : _GEN_20362; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20364 = 10'hdb == _T_308[9:0] ? 4'hc : _GEN_20363; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20365 = 10'hdc == _T_308[9:0] ? 4'h9 : _GEN_20364; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20366 = 10'hdd == _T_308[9:0] ? 4'he : _GEN_20365; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20367 = 10'hde == _T_308[9:0] ? 4'he : _GEN_20366; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20368 = 10'hdf == _T_308[9:0] ? 4'he : _GEN_20367; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20369 = 10'he0 == _T_308[9:0] ? 4'he : _GEN_20368; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20370 = 10'he1 == _T_308[9:0] ? 4'he : _GEN_20369; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20371 = 10'he2 == _T_308[9:0] ? 4'he : _GEN_20370; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20372 = 10'he3 == _T_308[9:0] ? 4'h9 : _GEN_20371; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20373 = 10'he4 == _T_308[9:0] ? 4'he : _GEN_20372; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20374 = 10'he5 == _T_308[9:0] ? 4'he : _GEN_20373; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20375 = 10'he6 == _T_308[9:0] ? 4'he : _GEN_20374; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20376 = 10'he7 == _T_308[9:0] ? 4'he : _GEN_20375; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20377 = 10'he8 == _T_308[9:0] ? 4'he : _GEN_20376; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20378 = 10'he9 == _T_308[9:0] ? 4'he : _GEN_20377; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20379 = 10'hea == _T_308[9:0] ? 4'he : _GEN_20378; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20380 = 10'heb == _T_308[9:0] ? 4'hc : _GEN_20379; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20381 = 10'hec == _T_308[9:0] ? 4'h7 : _GEN_20380; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20382 = 10'hed == _T_308[9:0] ? 4'h1 : _GEN_20381; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20383 = 10'hee == _T_308[9:0] ? 4'h0 : _GEN_20382; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20384 = 10'hef == _T_308[9:0] ? 4'h0 : _GEN_20383; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20385 = 10'hf0 == _T_308[9:0] ? 4'h2 : _GEN_20384; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20386 = 10'hf1 == _T_308[9:0] ? 4'h9 : _GEN_20385; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20387 = 10'hf2 == _T_308[9:0] ? 4'he : _GEN_20386; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20388 = 10'hf3 == _T_308[9:0] ? 4'he : _GEN_20387; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20389 = 10'hf4 == _T_308[9:0] ? 4'he : _GEN_20388; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20390 = 10'hf5 == _T_308[9:0] ? 4'hc : _GEN_20389; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20391 = 10'hf6 == _T_308[9:0] ? 4'hc : _GEN_20390; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20392 = 10'hf7 == _T_308[9:0] ? 4'hd : _GEN_20391; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20393 = 10'hf8 == _T_308[9:0] ? 4'hd : _GEN_20392; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20394 = 10'hf9 == _T_308[9:0] ? 4'hd : _GEN_20393; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20395 = 10'hfa == _T_308[9:0] ? 4'hd : _GEN_20394; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20396 = 10'hfb == _T_308[9:0] ? 4'hd : _GEN_20395; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20397 = 10'hfc == _T_308[9:0] ? 4'hd : _GEN_20396; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20398 = 10'hfd == _T_308[9:0] ? 4'hd : _GEN_20397; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20399 = 10'hfe == _T_308[9:0] ? 4'hd : _GEN_20398; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20400 = 10'hff == _T_308[9:0] ? 4'hd : _GEN_20399; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20401 = 10'h100 == _T_308[9:0] ? 4'hd : _GEN_20400; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20402 = 10'h101 == _T_308[9:0] ? 4'h9 : _GEN_20401; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20403 = 10'h102 == _T_308[9:0] ? 4'h9 : _GEN_20402; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20404 = 10'h103 == _T_308[9:0] ? 4'he : _GEN_20403; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20405 = 10'h104 == _T_308[9:0] ? 4'he : _GEN_20404; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20406 = 10'h105 == _T_308[9:0] ? 4'he : _GEN_20405; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20407 = 10'h106 == _T_308[9:0] ? 4'he : _GEN_20406; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20408 = 10'h107 == _T_308[9:0] ? 4'he : _GEN_20407; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20409 = 10'h108 == _T_308[9:0] ? 4'he : _GEN_20408; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20410 = 10'h109 == _T_308[9:0] ? 4'h6 : _GEN_20409; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20411 = 10'h10a == _T_308[9:0] ? 4'he : _GEN_20410; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20412 = 10'h10b == _T_308[9:0] ? 4'he : _GEN_20411; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20413 = 10'h10c == _T_308[9:0] ? 4'he : _GEN_20412; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20414 = 10'h10d == _T_308[9:0] ? 4'he : _GEN_20413; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20415 = 10'h10e == _T_308[9:0] ? 4'he : _GEN_20414; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20416 = 10'h10f == _T_308[9:0] ? 4'ha : _GEN_20415; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20417 = 10'h110 == _T_308[9:0] ? 4'hd : _GEN_20416; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20418 = 10'h111 == _T_308[9:0] ? 4'h4 : _GEN_20417; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20419 = 10'h112 == _T_308[9:0] ? 4'h7 : _GEN_20418; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20420 = 10'h113 == _T_308[9:0] ? 4'h0 : _GEN_20419; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20421 = 10'h114 == _T_308[9:0] ? 4'h0 : _GEN_20420; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20422 = 10'h115 == _T_308[9:0] ? 4'h0 : _GEN_20421; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20423 = 10'h116 == _T_308[9:0] ? 4'h0 : _GEN_20422; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20424 = 10'h117 == _T_308[9:0] ? 4'h0 : _GEN_20423; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20425 = 10'h118 == _T_308[9:0] ? 4'ha : _GEN_20424; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20426 = 10'h119 == _T_308[9:0] ? 4'he : _GEN_20425; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20427 = 10'h11a == _T_308[9:0] ? 4'he : _GEN_20426; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20428 = 10'h11b == _T_308[9:0] ? 4'he : _GEN_20427; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20429 = 10'h11c == _T_308[9:0] ? 4'hb : _GEN_20428; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20430 = 10'h11d == _T_308[9:0] ? 4'hc : _GEN_20429; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20431 = 10'h11e == _T_308[9:0] ? 4'hd : _GEN_20430; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20432 = 10'h11f == _T_308[9:0] ? 4'hb : _GEN_20431; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20433 = 10'h120 == _T_308[9:0] ? 4'ha : _GEN_20432; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20434 = 10'h121 == _T_308[9:0] ? 4'hc : _GEN_20433; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20435 = 10'h122 == _T_308[9:0] ? 4'ha : _GEN_20434; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20436 = 10'h123 == _T_308[9:0] ? 4'ha : _GEN_20435; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20437 = 10'h124 == _T_308[9:0] ? 4'hd : _GEN_20436; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20438 = 10'h125 == _T_308[9:0] ? 4'hd : _GEN_20437; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20439 = 10'h126 == _T_308[9:0] ? 4'hb : _GEN_20438; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20440 = 10'h127 == _T_308[9:0] ? 4'h9 : _GEN_20439; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20441 = 10'h128 == _T_308[9:0] ? 4'h7 : _GEN_20440; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20442 = 10'h129 == _T_308[9:0] ? 4'hd : _GEN_20441; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20443 = 10'h12a == _T_308[9:0] ? 4'hc : _GEN_20442; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20444 = 10'h12b == _T_308[9:0] ? 4'hb : _GEN_20443; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20445 = 10'h12c == _T_308[9:0] ? 4'hc : _GEN_20444; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20446 = 10'h12d == _T_308[9:0] ? 4'hb : _GEN_20445; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20447 = 10'h12e == _T_308[9:0] ? 4'ha : _GEN_20446; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20448 = 10'h12f == _T_308[9:0] ? 4'h6 : _GEN_20447; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20449 = 10'h130 == _T_308[9:0] ? 4'he : _GEN_20448; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20450 = 10'h131 == _T_308[9:0] ? 4'hc : _GEN_20449; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20451 = 10'h132 == _T_308[9:0] ? 4'ha : _GEN_20450; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20452 = 10'h133 == _T_308[9:0] ? 4'h9 : _GEN_20451; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20453 = 10'h134 == _T_308[9:0] ? 4'hb : _GEN_20452; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20454 = 10'h135 == _T_308[9:0] ? 4'h8 : _GEN_20453; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20455 = 10'h136 == _T_308[9:0] ? 4'h8 : _GEN_20454; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20456 = 10'h137 == _T_308[9:0] ? 4'h4 : _GEN_20455; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20457 = 10'h138 == _T_308[9:0] ? 4'h7 : _GEN_20456; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20458 = 10'h139 == _T_308[9:0] ? 4'h0 : _GEN_20457; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20459 = 10'h13a == _T_308[9:0] ? 4'h0 : _GEN_20458; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20460 = 10'h13b == _T_308[9:0] ? 4'h0 : _GEN_20459; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20461 = 10'h13c == _T_308[9:0] ? 4'h0 : _GEN_20460; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20462 = 10'h13d == _T_308[9:0] ? 4'h0 : _GEN_20461; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20463 = 10'h13e == _T_308[9:0] ? 4'h4 : _GEN_20462; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20464 = 10'h13f == _T_308[9:0] ? 4'hc : _GEN_20463; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20465 = 10'h140 == _T_308[9:0] ? 4'he : _GEN_20464; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20466 = 10'h141 == _T_308[9:0] ? 4'he : _GEN_20465; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20467 = 10'h142 == _T_308[9:0] ? 4'he : _GEN_20466; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20468 = 10'h143 == _T_308[9:0] ? 4'hc : _GEN_20467; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20469 = 10'h144 == _T_308[9:0] ? 4'hd : _GEN_20468; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20470 = 10'h145 == _T_308[9:0] ? 4'hb : _GEN_20469; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20471 = 10'h146 == _T_308[9:0] ? 4'hb : _GEN_20470; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20472 = 10'h147 == _T_308[9:0] ? 4'ha : _GEN_20471; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20473 = 10'h148 == _T_308[9:0] ? 4'ha : _GEN_20472; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20474 = 10'h149 == _T_308[9:0] ? 4'hc : _GEN_20473; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20475 = 10'h14a == _T_308[9:0] ? 4'hd : _GEN_20474; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20476 = 10'h14b == _T_308[9:0] ? 4'hc : _GEN_20475; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20477 = 10'h14c == _T_308[9:0] ? 4'hd : _GEN_20476; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20478 = 10'h14d == _T_308[9:0] ? 4'h9 : _GEN_20477; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20479 = 10'h14e == _T_308[9:0] ? 4'h7 : _GEN_20478; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20480 = 10'h14f == _T_308[9:0] ? 4'ha : _GEN_20479; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20481 = 10'h150 == _T_308[9:0] ? 4'ha : _GEN_20480; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20482 = 10'h151 == _T_308[9:0] ? 4'hb : _GEN_20481; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20483 = 10'h152 == _T_308[9:0] ? 4'hb : _GEN_20482; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20484 = 10'h153 == _T_308[9:0] ? 4'hc : _GEN_20483; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20485 = 10'h154 == _T_308[9:0] ? 4'hb : _GEN_20484; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20486 = 10'h155 == _T_308[9:0] ? 4'h6 : _GEN_20485; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20487 = 10'h156 == _T_308[9:0] ? 4'hb : _GEN_20486; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20488 = 10'h157 == _T_308[9:0] ? 4'h7 : _GEN_20487; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20489 = 10'h158 == _T_308[9:0] ? 4'h7 : _GEN_20488; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20490 = 10'h159 == _T_308[9:0] ? 4'h7 : _GEN_20489; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20491 = 10'h15a == _T_308[9:0] ? 4'h7 : _GEN_20490; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20492 = 10'h15b == _T_308[9:0] ? 4'h7 : _GEN_20491; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20493 = 10'h15c == _T_308[9:0] ? 4'h7 : _GEN_20492; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20494 = 10'h15d == _T_308[9:0] ? 4'h6 : _GEN_20493; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20495 = 10'h15e == _T_308[9:0] ? 4'h7 : _GEN_20494; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20496 = 10'h15f == _T_308[9:0] ? 4'h0 : _GEN_20495; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20497 = 10'h160 == _T_308[9:0] ? 4'h0 : _GEN_20496; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20498 = 10'h161 == _T_308[9:0] ? 4'h0 : _GEN_20497; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20499 = 10'h162 == _T_308[9:0] ? 4'h0 : _GEN_20498; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20500 = 10'h163 == _T_308[9:0] ? 4'h2 : _GEN_20499; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20501 = 10'h164 == _T_308[9:0] ? 4'h4 : _GEN_20500; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20502 = 10'h165 == _T_308[9:0] ? 4'hb : _GEN_20501; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20503 = 10'h166 == _T_308[9:0] ? 4'hb : _GEN_20502; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20504 = 10'h167 == _T_308[9:0] ? 4'he : _GEN_20503; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20505 = 10'h168 == _T_308[9:0] ? 4'he : _GEN_20504; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20506 = 10'h169 == _T_308[9:0] ? 4'hc : _GEN_20505; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20507 = 10'h16a == _T_308[9:0] ? 4'hd : _GEN_20506; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20508 = 10'h16b == _T_308[9:0] ? 4'hd : _GEN_20507; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20509 = 10'h16c == _T_308[9:0] ? 4'ha : _GEN_20508; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20510 = 10'h16d == _T_308[9:0] ? 4'ha : _GEN_20509; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20511 = 10'h16e == _T_308[9:0] ? 4'ha : _GEN_20510; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20512 = 10'h16f == _T_308[9:0] ? 4'hd : _GEN_20511; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20513 = 10'h170 == _T_308[9:0] ? 4'hd : _GEN_20512; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20514 = 10'h171 == _T_308[9:0] ? 4'hd : _GEN_20513; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20515 = 10'h172 == _T_308[9:0] ? 4'he : _GEN_20514; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20516 = 10'h173 == _T_308[9:0] ? 4'h8 : _GEN_20515; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20517 = 10'h174 == _T_308[9:0] ? 4'h5 : _GEN_20516; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20518 = 10'h175 == _T_308[9:0] ? 4'h6 : _GEN_20517; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20519 = 10'h176 == _T_308[9:0] ? 4'h6 : _GEN_20518; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20520 = 10'h177 == _T_308[9:0] ? 4'h6 : _GEN_20519; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20521 = 10'h178 == _T_308[9:0] ? 4'h7 : _GEN_20520; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20522 = 10'h179 == _T_308[9:0] ? 4'h9 : _GEN_20521; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20523 = 10'h17a == _T_308[9:0] ? 4'h9 : _GEN_20522; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20524 = 10'h17b == _T_308[9:0] ? 4'h6 : _GEN_20523; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20525 = 10'h17c == _T_308[9:0] ? 4'h7 : _GEN_20524; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20526 = 10'h17d == _T_308[9:0] ? 4'h7 : _GEN_20525; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20527 = 10'h17e == _T_308[9:0] ? 4'h7 : _GEN_20526; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20528 = 10'h17f == _T_308[9:0] ? 4'h7 : _GEN_20527; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20529 = 10'h180 == _T_308[9:0] ? 4'h7 : _GEN_20528; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20530 = 10'h181 == _T_308[9:0] ? 4'h7 : _GEN_20529; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20531 = 10'h182 == _T_308[9:0] ? 4'h8 : _GEN_20530; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20532 = 10'h183 == _T_308[9:0] ? 4'h8 : _GEN_20531; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20533 = 10'h184 == _T_308[9:0] ? 4'h8 : _GEN_20532; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20534 = 10'h185 == _T_308[9:0] ? 4'h7 : _GEN_20533; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20535 = 10'h186 == _T_308[9:0] ? 4'h1 : _GEN_20534; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20536 = 10'h187 == _T_308[9:0] ? 4'h0 : _GEN_20535; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20537 = 10'h188 == _T_308[9:0] ? 4'h0 : _GEN_20536; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20538 = 10'h189 == _T_308[9:0] ? 4'h4 : _GEN_20537; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20539 = 10'h18a == _T_308[9:0] ? 4'h4 : _GEN_20538; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20540 = 10'h18b == _T_308[9:0] ? 4'hb : _GEN_20539; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20541 = 10'h18c == _T_308[9:0] ? 4'hb : _GEN_20540; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20542 = 10'h18d == _T_308[9:0] ? 4'hc : _GEN_20541; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20543 = 10'h18e == _T_308[9:0] ? 4'he : _GEN_20542; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20544 = 10'h18f == _T_308[9:0] ? 4'hb : _GEN_20543; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20545 = 10'h190 == _T_308[9:0] ? 4'hd : _GEN_20544; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20546 = 10'h191 == _T_308[9:0] ? 4'hc : _GEN_20545; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20547 = 10'h192 == _T_308[9:0] ? 4'h9 : _GEN_20546; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20548 = 10'h193 == _T_308[9:0] ? 4'ha : _GEN_20547; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20549 = 10'h194 == _T_308[9:0] ? 4'h9 : _GEN_20548; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20550 = 10'h195 == _T_308[9:0] ? 4'hd : _GEN_20549; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20551 = 10'h196 == _T_308[9:0] ? 4'hd : _GEN_20550; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20552 = 10'h197 == _T_308[9:0] ? 4'hb : _GEN_20551; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20553 = 10'h198 == _T_308[9:0] ? 4'he : _GEN_20552; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20554 = 10'h199 == _T_308[9:0] ? 4'h5 : _GEN_20553; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20555 = 10'h19a == _T_308[9:0] ? 4'h1 : _GEN_20554; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20556 = 10'h19b == _T_308[9:0] ? 4'h3 : _GEN_20555; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20557 = 10'h19c == _T_308[9:0] ? 4'h6 : _GEN_20556; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20558 = 10'h19d == _T_308[9:0] ? 4'h4 : _GEN_20557; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20559 = 10'h19e == _T_308[9:0] ? 4'h1 : _GEN_20558; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20560 = 10'h19f == _T_308[9:0] ? 4'h3 : _GEN_20559; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20561 = 10'h1a0 == _T_308[9:0] ? 4'h6 : _GEN_20560; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20562 = 10'h1a1 == _T_308[9:0] ? 4'h6 : _GEN_20561; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20563 = 10'h1a2 == _T_308[9:0] ? 4'h7 : _GEN_20562; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20564 = 10'h1a3 == _T_308[9:0] ? 4'h7 : _GEN_20563; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20565 = 10'h1a4 == _T_308[9:0] ? 4'h7 : _GEN_20564; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20566 = 10'h1a5 == _T_308[9:0] ? 4'h7 : _GEN_20565; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20567 = 10'h1a6 == _T_308[9:0] ? 4'h7 : _GEN_20566; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20568 = 10'h1a7 == _T_308[9:0] ? 4'h7 : _GEN_20567; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20569 = 10'h1a8 == _T_308[9:0] ? 4'h8 : _GEN_20568; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20570 = 10'h1a9 == _T_308[9:0] ? 4'h8 : _GEN_20569; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20571 = 10'h1aa == _T_308[9:0] ? 4'h7 : _GEN_20570; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20572 = 10'h1ab == _T_308[9:0] ? 4'h8 : _GEN_20571; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20573 = 10'h1ac == _T_308[9:0] ? 4'h8 : _GEN_20572; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20574 = 10'h1ad == _T_308[9:0] ? 4'h3 : _GEN_20573; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20575 = 10'h1ae == _T_308[9:0] ? 4'h2 : _GEN_20574; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20576 = 10'h1af == _T_308[9:0] ? 4'h8 : _GEN_20575; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20577 = 10'h1b0 == _T_308[9:0] ? 4'h6 : _GEN_20576; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20578 = 10'h1b1 == _T_308[9:0] ? 4'hb : _GEN_20577; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20579 = 10'h1b2 == _T_308[9:0] ? 4'hb : _GEN_20578; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20580 = 10'h1b3 == _T_308[9:0] ? 4'ha : _GEN_20579; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20581 = 10'h1b4 == _T_308[9:0] ? 4'he : _GEN_20580; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20582 = 10'h1b5 == _T_308[9:0] ? 4'hb : _GEN_20581; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20583 = 10'h1b6 == _T_308[9:0] ? 4'hc : _GEN_20582; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20584 = 10'h1b7 == _T_308[9:0] ? 4'ha : _GEN_20583; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20585 = 10'h1b8 == _T_308[9:0] ? 4'h9 : _GEN_20584; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20586 = 10'h1b9 == _T_308[9:0] ? 4'h9 : _GEN_20585; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20587 = 10'h1ba == _T_308[9:0] ? 4'h9 : _GEN_20586; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20588 = 10'h1bb == _T_308[9:0] ? 4'hb : _GEN_20587; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20589 = 10'h1bc == _T_308[9:0] ? 4'hd : _GEN_20588; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20590 = 10'h1bd == _T_308[9:0] ? 4'hd : _GEN_20589; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20591 = 10'h1be == _T_308[9:0] ? 4'he : _GEN_20590; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20592 = 10'h1bf == _T_308[9:0] ? 4'h7 : _GEN_20591; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20593 = 10'h1c0 == _T_308[9:0] ? 4'h6 : _GEN_20592; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20594 = 10'h1c1 == _T_308[9:0] ? 4'h6 : _GEN_20593; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20595 = 10'h1c2 == _T_308[9:0] ? 4'h5 : _GEN_20594; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20596 = 10'h1c3 == _T_308[9:0] ? 4'h5 : _GEN_20595; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20597 = 10'h1c4 == _T_308[9:0] ? 4'h4 : _GEN_20596; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20598 = 10'h1c5 == _T_308[9:0] ? 4'h5 : _GEN_20597; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20599 = 10'h1c6 == _T_308[9:0] ? 4'h6 : _GEN_20598; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20600 = 10'h1c7 == _T_308[9:0] ? 4'h6 : _GEN_20599; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20601 = 10'h1c8 == _T_308[9:0] ? 4'h7 : _GEN_20600; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20602 = 10'h1c9 == _T_308[9:0] ? 4'h7 : _GEN_20601; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20603 = 10'h1ca == _T_308[9:0] ? 4'h7 : _GEN_20602; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20604 = 10'h1cb == _T_308[9:0] ? 4'h7 : _GEN_20603; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20605 = 10'h1cc == _T_308[9:0] ? 4'h7 : _GEN_20604; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20606 = 10'h1cd == _T_308[9:0] ? 4'h8 : _GEN_20605; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20607 = 10'h1ce == _T_308[9:0] ? 4'h8 : _GEN_20606; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20608 = 10'h1cf == _T_308[9:0] ? 4'h8 : _GEN_20607; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20609 = 10'h1d0 == _T_308[9:0] ? 4'h5 : _GEN_20608; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20610 = 10'h1d1 == _T_308[9:0] ? 4'h8 : _GEN_20609; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20611 = 10'h1d2 == _T_308[9:0] ? 4'h8 : _GEN_20610; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20612 = 10'h1d3 == _T_308[9:0] ? 4'h8 : _GEN_20611; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20613 = 10'h1d4 == _T_308[9:0] ? 4'h8 : _GEN_20612; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20614 = 10'h1d5 == _T_308[9:0] ? 4'h7 : _GEN_20613; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20615 = 10'h1d6 == _T_308[9:0] ? 4'h9 : _GEN_20614; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20616 = 10'h1d7 == _T_308[9:0] ? 4'hb : _GEN_20615; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20617 = 10'h1d8 == _T_308[9:0] ? 4'hb : _GEN_20616; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20618 = 10'h1d9 == _T_308[9:0] ? 4'hb : _GEN_20617; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20619 = 10'h1da == _T_308[9:0] ? 4'ha : _GEN_20618; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20620 = 10'h1db == _T_308[9:0] ? 4'hc : _GEN_20619; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20621 = 10'h1dc == _T_308[9:0] ? 4'hb : _GEN_20620; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20622 = 10'h1dd == _T_308[9:0] ? 4'h5 : _GEN_20621; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20623 = 10'h1de == _T_308[9:0] ? 4'h9 : _GEN_20622; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20624 = 10'h1df == _T_308[9:0] ? 4'h9 : _GEN_20623; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20625 = 10'h1e0 == _T_308[9:0] ? 4'h9 : _GEN_20624; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20626 = 10'h1e1 == _T_308[9:0] ? 4'h7 : _GEN_20625; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20627 = 10'h1e2 == _T_308[9:0] ? 4'hc : _GEN_20626; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20628 = 10'h1e3 == _T_308[9:0] ? 4'hc : _GEN_20627; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20629 = 10'h1e4 == _T_308[9:0] ? 4'hd : _GEN_20628; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20630 = 10'h1e5 == _T_308[9:0] ? 4'h7 : _GEN_20629; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20631 = 10'h1e6 == _T_308[9:0] ? 4'h6 : _GEN_20630; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20632 = 10'h1e7 == _T_308[9:0] ? 4'h6 : _GEN_20631; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20633 = 10'h1e8 == _T_308[9:0] ? 4'h6 : _GEN_20632; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20634 = 10'h1e9 == _T_308[9:0] ? 4'h6 : _GEN_20633; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20635 = 10'h1ea == _T_308[9:0] ? 4'h6 : _GEN_20634; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20636 = 10'h1eb == _T_308[9:0] ? 4'h6 : _GEN_20635; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20637 = 10'h1ec == _T_308[9:0] ? 4'h6 : _GEN_20636; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20638 = 10'h1ed == _T_308[9:0] ? 4'h8 : _GEN_20637; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20639 = 10'h1ee == _T_308[9:0] ? 4'h7 : _GEN_20638; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20640 = 10'h1ef == _T_308[9:0] ? 4'h7 : _GEN_20639; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20641 = 10'h1f0 == _T_308[9:0] ? 4'h7 : _GEN_20640; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20642 = 10'h1f1 == _T_308[9:0] ? 4'h7 : _GEN_20641; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20643 = 10'h1f2 == _T_308[9:0] ? 4'h7 : _GEN_20642; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20644 = 10'h1f3 == _T_308[9:0] ? 4'h8 : _GEN_20643; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20645 = 10'h1f4 == _T_308[9:0] ? 4'h8 : _GEN_20644; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20646 = 10'h1f5 == _T_308[9:0] ? 4'h8 : _GEN_20645; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20647 = 10'h1f6 == _T_308[9:0] ? 4'ha : _GEN_20646; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20648 = 10'h1f7 == _T_308[9:0] ? 4'h8 : _GEN_20647; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20649 = 10'h1f8 == _T_308[9:0] ? 4'h8 : _GEN_20648; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20650 = 10'h1f9 == _T_308[9:0] ? 4'h9 : _GEN_20649; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20651 = 10'h1fa == _T_308[9:0] ? 4'h9 : _GEN_20650; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20652 = 10'h1fb == _T_308[9:0] ? 4'h8 : _GEN_20651; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20653 = 10'h1fc == _T_308[9:0] ? 4'hb : _GEN_20652; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20654 = 10'h1fd == _T_308[9:0] ? 4'hb : _GEN_20653; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20655 = 10'h1fe == _T_308[9:0] ? 4'hb : _GEN_20654; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20656 = 10'h1ff == _T_308[9:0] ? 4'ha : _GEN_20655; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20657 = 10'h200 == _T_308[9:0] ? 4'h3 : _GEN_20656; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20658 = 10'h201 == _T_308[9:0] ? 4'h9 : _GEN_20657; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20659 = 10'h202 == _T_308[9:0] ? 4'h5 : _GEN_20658; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20660 = 10'h203 == _T_308[9:0] ? 4'h3 : _GEN_20659; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20661 = 10'h204 == _T_308[9:0] ? 4'h4 : _GEN_20660; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20662 = 10'h205 == _T_308[9:0] ? 4'h4 : _GEN_20661; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20663 = 10'h206 == _T_308[9:0] ? 4'h4 : _GEN_20662; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20664 = 10'h207 == _T_308[9:0] ? 4'h4 : _GEN_20663; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20665 = 10'h208 == _T_308[9:0] ? 4'h8 : _GEN_20664; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20666 = 10'h209 == _T_308[9:0] ? 4'hc : _GEN_20665; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20667 = 10'h20a == _T_308[9:0] ? 4'hd : _GEN_20666; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20668 = 10'h20b == _T_308[9:0] ? 4'h7 : _GEN_20667; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20669 = 10'h20c == _T_308[9:0] ? 4'h6 : _GEN_20668; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20670 = 10'h20d == _T_308[9:0] ? 4'h6 : _GEN_20669; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20671 = 10'h20e == _T_308[9:0] ? 4'h6 : _GEN_20670; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20672 = 10'h20f == _T_308[9:0] ? 4'h5 : _GEN_20671; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20673 = 10'h210 == _T_308[9:0] ? 4'h6 : _GEN_20672; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20674 = 10'h211 == _T_308[9:0] ? 4'h6 : _GEN_20673; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20675 = 10'h212 == _T_308[9:0] ? 4'h7 : _GEN_20674; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20676 = 10'h213 == _T_308[9:0] ? 4'ha : _GEN_20675; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20677 = 10'h214 == _T_308[9:0] ? 4'h6 : _GEN_20676; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20678 = 10'h215 == _T_308[9:0] ? 4'h7 : _GEN_20677; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20679 = 10'h216 == _T_308[9:0] ? 4'h7 : _GEN_20678; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20680 = 10'h217 == _T_308[9:0] ? 4'h7 : _GEN_20679; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20681 = 10'h218 == _T_308[9:0] ? 4'h7 : _GEN_20680; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20682 = 10'h219 == _T_308[9:0] ? 4'h8 : _GEN_20681; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20683 = 10'h21a == _T_308[9:0] ? 4'h7 : _GEN_20682; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20684 = 10'h21b == _T_308[9:0] ? 4'h8 : _GEN_20683; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20685 = 10'h21c == _T_308[9:0] ? 4'hb : _GEN_20684; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20686 = 10'h21d == _T_308[9:0] ? 4'ha : _GEN_20685; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20687 = 10'h21e == _T_308[9:0] ? 4'h9 : _GEN_20686; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20688 = 10'h21f == _T_308[9:0] ? 4'h9 : _GEN_20687; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20689 = 10'h220 == _T_308[9:0] ? 4'h8 : _GEN_20688; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20690 = 10'h221 == _T_308[9:0] ? 4'h9 : _GEN_20689; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20691 = 10'h222 == _T_308[9:0] ? 4'hb : _GEN_20690; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20692 = 10'h223 == _T_308[9:0] ? 4'hb : _GEN_20691; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20693 = 10'h224 == _T_308[9:0] ? 4'hb : _GEN_20692; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20694 = 10'h225 == _T_308[9:0] ? 4'h8 : _GEN_20693; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20695 = 10'h226 == _T_308[9:0] ? 4'h1 : _GEN_20694; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20696 = 10'h227 == _T_308[9:0] ? 4'h3 : _GEN_20695; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20697 = 10'h228 == _T_308[9:0] ? 4'h3 : _GEN_20696; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20698 = 10'h229 == _T_308[9:0] ? 4'h3 : _GEN_20697; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20699 = 10'h22a == _T_308[9:0] ? 4'h3 : _GEN_20698; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20700 = 10'h22b == _T_308[9:0] ? 4'h3 : _GEN_20699; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20701 = 10'h22c == _T_308[9:0] ? 4'h3 : _GEN_20700; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20702 = 10'h22d == _T_308[9:0] ? 4'h3 : _GEN_20701; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20703 = 10'h22e == _T_308[9:0] ? 4'h3 : _GEN_20702; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20704 = 10'h22f == _T_308[9:0] ? 4'h9 : _GEN_20703; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20705 = 10'h230 == _T_308[9:0] ? 4'h6 : _GEN_20704; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20706 = 10'h231 == _T_308[9:0] ? 4'h7 : _GEN_20705; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20707 = 10'h232 == _T_308[9:0] ? 4'h6 : _GEN_20706; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20708 = 10'h233 == _T_308[9:0] ? 4'h7 : _GEN_20707; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20709 = 10'h234 == _T_308[9:0] ? 4'h7 : _GEN_20708; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20710 = 10'h235 == _T_308[9:0] ? 4'h6 : _GEN_20709; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20711 = 10'h236 == _T_308[9:0] ? 4'h6 : _GEN_20710; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20712 = 10'h237 == _T_308[9:0] ? 4'h6 : _GEN_20711; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20713 = 10'h238 == _T_308[9:0] ? 4'h6 : _GEN_20712; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20714 = 10'h239 == _T_308[9:0] ? 4'h8 : _GEN_20713; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20715 = 10'h23a == _T_308[9:0] ? 4'h6 : _GEN_20714; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20716 = 10'h23b == _T_308[9:0] ? 4'h7 : _GEN_20715; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20717 = 10'h23c == _T_308[9:0] ? 4'h7 : _GEN_20716; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20718 = 10'h23d == _T_308[9:0] ? 4'h7 : _GEN_20717; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20719 = 10'h23e == _T_308[9:0] ? 4'h7 : _GEN_20718; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20720 = 10'h23f == _T_308[9:0] ? 4'h7 : _GEN_20719; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20721 = 10'h240 == _T_308[9:0] ? 4'h7 : _GEN_20720; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20722 = 10'h241 == _T_308[9:0] ? 4'h8 : _GEN_20721; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20723 = 10'h242 == _T_308[9:0] ? 4'hb : _GEN_20722; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20724 = 10'h243 == _T_308[9:0] ? 4'hb : _GEN_20723; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20725 = 10'h244 == _T_308[9:0] ? 4'hb : _GEN_20724; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20726 = 10'h245 == _T_308[9:0] ? 4'ha : _GEN_20725; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20727 = 10'h246 == _T_308[9:0] ? 4'h9 : _GEN_20726; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20728 = 10'h247 == _T_308[9:0] ? 4'ha : _GEN_20727; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20729 = 10'h248 == _T_308[9:0] ? 4'hb : _GEN_20728; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20730 = 10'h249 == _T_308[9:0] ? 4'hb : _GEN_20729; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20731 = 10'h24a == _T_308[9:0] ? 4'ha : _GEN_20730; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20732 = 10'h24b == _T_308[9:0] ? 4'h2 : _GEN_20731; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20733 = 10'h24c == _T_308[9:0] ? 4'h0 : _GEN_20732; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20734 = 10'h24d == _T_308[9:0] ? 4'h2 : _GEN_20733; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20735 = 10'h24e == _T_308[9:0] ? 4'h3 : _GEN_20734; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20736 = 10'h24f == _T_308[9:0] ? 4'h3 : _GEN_20735; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20737 = 10'h250 == _T_308[9:0] ? 4'h3 : _GEN_20736; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20738 = 10'h251 == _T_308[9:0] ? 4'h3 : _GEN_20737; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20739 = 10'h252 == _T_308[9:0] ? 4'h3 : _GEN_20738; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20740 = 10'h253 == _T_308[9:0] ? 4'h3 : _GEN_20739; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20741 = 10'h254 == _T_308[9:0] ? 4'h3 : _GEN_20740; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20742 = 10'h255 == _T_308[9:0] ? 4'h5 : _GEN_20741; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20743 = 10'h256 == _T_308[9:0] ? 4'h6 : _GEN_20742; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20744 = 10'h257 == _T_308[9:0] ? 4'h8 : _GEN_20743; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20745 = 10'h258 == _T_308[9:0] ? 4'h5 : _GEN_20744; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20746 = 10'h259 == _T_308[9:0] ? 4'h6 : _GEN_20745; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20747 = 10'h25a == _T_308[9:0] ? 4'h6 : _GEN_20746; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20748 = 10'h25b == _T_308[9:0] ? 4'h5 : _GEN_20747; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20749 = 10'h25c == _T_308[9:0] ? 4'h6 : _GEN_20748; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20750 = 10'h25d == _T_308[9:0] ? 4'h6 : _GEN_20749; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20751 = 10'h25e == _T_308[9:0] ? 4'h9 : _GEN_20750; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20752 = 10'h25f == _T_308[9:0] ? 4'hc : _GEN_20751; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20753 = 10'h260 == _T_308[9:0] ? 4'h7 : _GEN_20752; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20754 = 10'h261 == _T_308[9:0] ? 4'h9 : _GEN_20753; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20755 = 10'h262 == _T_308[9:0] ? 4'ha : _GEN_20754; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20756 = 10'h263 == _T_308[9:0] ? 4'h8 : _GEN_20755; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20757 = 10'h264 == _T_308[9:0] ? 4'ha : _GEN_20756; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20758 = 10'h265 == _T_308[9:0] ? 4'h9 : _GEN_20757; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20759 = 10'h266 == _T_308[9:0] ? 4'h8 : _GEN_20758; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20760 = 10'h267 == _T_308[9:0] ? 4'h8 : _GEN_20759; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20761 = 10'h268 == _T_308[9:0] ? 4'ha : _GEN_20760; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20762 = 10'h269 == _T_308[9:0] ? 4'ha : _GEN_20761; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20763 = 10'h26a == _T_308[9:0] ? 4'hb : _GEN_20762; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20764 = 10'h26b == _T_308[9:0] ? 4'hb : _GEN_20763; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20765 = 10'h26c == _T_308[9:0] ? 4'hb : _GEN_20764; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20766 = 10'h26d == _T_308[9:0] ? 4'hb : _GEN_20765; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20767 = 10'h26e == _T_308[9:0] ? 4'hb : _GEN_20766; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20768 = 10'h26f == _T_308[9:0] ? 4'ha : _GEN_20767; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20769 = 10'h270 == _T_308[9:0] ? 4'h3 : _GEN_20768; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20770 = 10'h271 == _T_308[9:0] ? 4'h0 : _GEN_20769; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20771 = 10'h272 == _T_308[9:0] ? 4'h0 : _GEN_20770; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20772 = 10'h273 == _T_308[9:0] ? 4'h2 : _GEN_20771; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20773 = 10'h274 == _T_308[9:0] ? 4'h3 : _GEN_20772; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20774 = 10'h275 == _T_308[9:0] ? 4'h3 : _GEN_20773; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20775 = 10'h276 == _T_308[9:0] ? 4'h3 : _GEN_20774; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20776 = 10'h277 == _T_308[9:0] ? 4'h3 : _GEN_20775; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20777 = 10'h278 == _T_308[9:0] ? 4'h3 : _GEN_20776; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20778 = 10'h279 == _T_308[9:0] ? 4'h3 : _GEN_20777; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20779 = 10'h27a == _T_308[9:0] ? 4'h3 : _GEN_20778; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20780 = 10'h27b == _T_308[9:0] ? 4'h6 : _GEN_20779; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20781 = 10'h27c == _T_308[9:0] ? 4'h7 : _GEN_20780; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20782 = 10'h27d == _T_308[9:0] ? 4'h7 : _GEN_20781; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20783 = 10'h27e == _T_308[9:0] ? 4'h4 : _GEN_20782; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20784 = 10'h27f == _T_308[9:0] ? 4'h6 : _GEN_20783; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20785 = 10'h280 == _T_308[9:0] ? 4'h6 : _GEN_20784; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20786 = 10'h281 == _T_308[9:0] ? 4'h6 : _GEN_20785; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20787 = 10'h282 == _T_308[9:0] ? 4'h6 : _GEN_20786; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20788 = 10'h283 == _T_308[9:0] ? 4'ha : _GEN_20787; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20789 = 10'h284 == _T_308[9:0] ? 4'hc : _GEN_20788; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20790 = 10'h285 == _T_308[9:0] ? 4'hc : _GEN_20789; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20791 = 10'h286 == _T_308[9:0] ? 4'h8 : _GEN_20790; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20792 = 10'h287 == _T_308[9:0] ? 4'ha : _GEN_20791; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20793 = 10'h288 == _T_308[9:0] ? 4'ha : _GEN_20792; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20794 = 10'h289 == _T_308[9:0] ? 4'ha : _GEN_20793; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20795 = 10'h28a == _T_308[9:0] ? 4'hc : _GEN_20794; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20796 = 10'h28b == _T_308[9:0] ? 4'hb : _GEN_20795; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20797 = 10'h28c == _T_308[9:0] ? 4'ha : _GEN_20796; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20798 = 10'h28d == _T_308[9:0] ? 4'h7 : _GEN_20797; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20799 = 10'h28e == _T_308[9:0] ? 4'h2 : _GEN_20798; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20800 = 10'h28f == _T_308[9:0] ? 4'h5 : _GEN_20799; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20801 = 10'h290 == _T_308[9:0] ? 4'h8 : _GEN_20800; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20802 = 10'h291 == _T_308[9:0] ? 4'ha : _GEN_20801; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20803 = 10'h292 == _T_308[9:0] ? 4'ha : _GEN_20802; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20804 = 10'h293 == _T_308[9:0] ? 4'ha : _GEN_20803; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20805 = 10'h294 == _T_308[9:0] ? 4'h9 : _GEN_20804; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20806 = 10'h295 == _T_308[9:0] ? 4'h3 : _GEN_20805; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20807 = 10'h296 == _T_308[9:0] ? 4'h0 : _GEN_20806; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20808 = 10'h297 == _T_308[9:0] ? 4'h0 : _GEN_20807; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20809 = 10'h298 == _T_308[9:0] ? 4'h0 : _GEN_20808; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20810 = 10'h299 == _T_308[9:0] ? 4'h1 : _GEN_20809; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20811 = 10'h29a == _T_308[9:0] ? 4'h3 : _GEN_20810; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20812 = 10'h29b == _T_308[9:0] ? 4'h3 : _GEN_20811; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20813 = 10'h29c == _T_308[9:0] ? 4'h3 : _GEN_20812; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20814 = 10'h29d == _T_308[9:0] ? 4'h3 : _GEN_20813; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20815 = 10'h29e == _T_308[9:0] ? 4'h3 : _GEN_20814; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20816 = 10'h29f == _T_308[9:0] ? 4'h3 : _GEN_20815; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20817 = 10'h2a0 == _T_308[9:0] ? 4'h4 : _GEN_20816; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20818 = 10'h2a1 == _T_308[9:0] ? 4'h6 : _GEN_20817; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20819 = 10'h2a2 == _T_308[9:0] ? 4'h7 : _GEN_20818; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20820 = 10'h2a3 == _T_308[9:0] ? 4'h6 : _GEN_20819; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20821 = 10'h2a4 == _T_308[9:0] ? 4'h4 : _GEN_20820; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20822 = 10'h2a5 == _T_308[9:0] ? 4'h6 : _GEN_20821; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20823 = 10'h2a6 == _T_308[9:0] ? 4'h6 : _GEN_20822; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20824 = 10'h2a7 == _T_308[9:0] ? 4'h7 : _GEN_20823; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20825 = 10'h2a8 == _T_308[9:0] ? 4'ha : _GEN_20824; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20826 = 10'h2a9 == _T_308[9:0] ? 4'hb : _GEN_20825; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20827 = 10'h2aa == _T_308[9:0] ? 4'hb : _GEN_20826; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20828 = 10'h2ab == _T_308[9:0] ? 4'hb : _GEN_20827; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20829 = 10'h2ac == _T_308[9:0] ? 4'h8 : _GEN_20828; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20830 = 10'h2ad == _T_308[9:0] ? 4'hb : _GEN_20829; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20831 = 10'h2ae == _T_308[9:0] ? 4'ha : _GEN_20830; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20832 = 10'h2af == _T_308[9:0] ? 4'hb : _GEN_20831; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20833 = 10'h2b0 == _T_308[9:0] ? 4'hc : _GEN_20832; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20834 = 10'h2b1 == _T_308[9:0] ? 4'hb : _GEN_20833; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20835 = 10'h2b2 == _T_308[9:0] ? 4'ha : _GEN_20834; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20836 = 10'h2b3 == _T_308[9:0] ? 4'h6 : _GEN_20835; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20837 = 10'h2b4 == _T_308[9:0] ? 4'h0 : _GEN_20836; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20838 = 10'h2b5 == _T_308[9:0] ? 4'h0 : _GEN_20837; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20839 = 10'h2b6 == _T_308[9:0] ? 4'h0 : _GEN_20838; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20840 = 10'h2b7 == _T_308[9:0] ? 4'h1 : _GEN_20839; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20841 = 10'h2b8 == _T_308[9:0] ? 4'h5 : _GEN_20840; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20842 = 10'h2b9 == _T_308[9:0] ? 4'h9 : _GEN_20841; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20843 = 10'h2ba == _T_308[9:0] ? 4'h1 : _GEN_20842; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20844 = 10'h2bb == _T_308[9:0] ? 4'h0 : _GEN_20843; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20845 = 10'h2bc == _T_308[9:0] ? 4'h0 : _GEN_20844; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20846 = 10'h2bd == _T_308[9:0] ? 4'h0 : _GEN_20845; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20847 = 10'h2be == _T_308[9:0] ? 4'h0 : _GEN_20846; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20848 = 10'h2bf == _T_308[9:0] ? 4'h0 : _GEN_20847; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20849 = 10'h2c0 == _T_308[9:0] ? 4'h3 : _GEN_20848; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20850 = 10'h2c1 == _T_308[9:0] ? 4'h3 : _GEN_20849; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20851 = 10'h2c2 == _T_308[9:0] ? 4'h3 : _GEN_20850; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20852 = 10'h2c3 == _T_308[9:0] ? 4'h3 : _GEN_20851; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20853 = 10'h2c4 == _T_308[9:0] ? 4'h3 : _GEN_20852; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20854 = 10'h2c5 == _T_308[9:0] ? 4'h3 : _GEN_20853; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20855 = 10'h2c6 == _T_308[9:0] ? 4'h4 : _GEN_20854; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20856 = 10'h2c7 == _T_308[9:0] ? 4'h5 : _GEN_20855; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20857 = 10'h2c8 == _T_308[9:0] ? 4'h7 : _GEN_20856; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20858 = 10'h2c9 == _T_308[9:0] ? 4'h7 : _GEN_20857; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20859 = 10'h2ca == _T_308[9:0] ? 4'h4 : _GEN_20858; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20860 = 10'h2cb == _T_308[9:0] ? 4'h9 : _GEN_20859; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20861 = 10'h2cc == _T_308[9:0] ? 4'h9 : _GEN_20860; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20862 = 10'h2cd == _T_308[9:0] ? 4'hb : _GEN_20861; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20863 = 10'h2ce == _T_308[9:0] ? 4'hb : _GEN_20862; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20864 = 10'h2cf == _T_308[9:0] ? 4'hb : _GEN_20863; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20865 = 10'h2d0 == _T_308[9:0] ? 4'hb : _GEN_20864; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20866 = 10'h2d1 == _T_308[9:0] ? 4'hb : _GEN_20865; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20867 = 10'h2d2 == _T_308[9:0] ? 4'h8 : _GEN_20866; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20868 = 10'h2d3 == _T_308[9:0] ? 4'ha : _GEN_20867; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20869 = 10'h2d4 == _T_308[9:0] ? 4'hb : _GEN_20868; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20870 = 10'h2d5 == _T_308[9:0] ? 4'ha : _GEN_20869; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20871 = 10'h2d6 == _T_308[9:0] ? 4'ha : _GEN_20870; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20872 = 10'h2d7 == _T_308[9:0] ? 4'ha : _GEN_20871; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20873 = 10'h2d8 == _T_308[9:0] ? 4'ha : _GEN_20872; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20874 = 10'h2d9 == _T_308[9:0] ? 4'h7 : _GEN_20873; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20875 = 10'h2da == _T_308[9:0] ? 4'h2 : _GEN_20874; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20876 = 10'h2db == _T_308[9:0] ? 4'h0 : _GEN_20875; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20877 = 10'h2dc == _T_308[9:0] ? 4'h0 : _GEN_20876; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20878 = 10'h2dd == _T_308[9:0] ? 4'h0 : _GEN_20877; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20879 = 10'h2de == _T_308[9:0] ? 4'h0 : _GEN_20878; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20880 = 10'h2df == _T_308[9:0] ? 4'h2 : _GEN_20879; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20881 = 10'h2e0 == _T_308[9:0] ? 4'h0 : _GEN_20880; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20882 = 10'h2e1 == _T_308[9:0] ? 4'h0 : _GEN_20881; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20883 = 10'h2e2 == _T_308[9:0] ? 4'h0 : _GEN_20882; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20884 = 10'h2e3 == _T_308[9:0] ? 4'h0 : _GEN_20883; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20885 = 10'h2e4 == _T_308[9:0] ? 4'h0 : _GEN_20884; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20886 = 10'h2e5 == _T_308[9:0] ? 4'h0 : _GEN_20885; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20887 = 10'h2e6 == _T_308[9:0] ? 4'h2 : _GEN_20886; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20888 = 10'h2e7 == _T_308[9:0] ? 4'h3 : _GEN_20887; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20889 = 10'h2e8 == _T_308[9:0] ? 4'h3 : _GEN_20888; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20890 = 10'h2e9 == _T_308[9:0] ? 4'h3 : _GEN_20889; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20891 = 10'h2ea == _T_308[9:0] ? 4'h3 : _GEN_20890; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20892 = 10'h2eb == _T_308[9:0] ? 4'h3 : _GEN_20891; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20893 = 10'h2ec == _T_308[9:0] ? 4'h4 : _GEN_20892; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20894 = 10'h2ed == _T_308[9:0] ? 4'h5 : _GEN_20893; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20895 = 10'h2ee == _T_308[9:0] ? 4'h6 : _GEN_20894; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20896 = 10'h2ef == _T_308[9:0] ? 4'h8 : _GEN_20895; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20897 = 10'h2f0 == _T_308[9:0] ? 4'h4 : _GEN_20896; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20898 = 10'h2f1 == _T_308[9:0] ? 4'h9 : _GEN_20897; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20899 = 10'h2f2 == _T_308[9:0] ? 4'hb : _GEN_20898; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20900 = 10'h2f3 == _T_308[9:0] ? 4'hb : _GEN_20899; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20901 = 10'h2f4 == _T_308[9:0] ? 4'hb : _GEN_20900; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20902 = 10'h2f5 == _T_308[9:0] ? 4'hb : _GEN_20901; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20903 = 10'h2f6 == _T_308[9:0] ? 4'hb : _GEN_20902; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20904 = 10'h2f7 == _T_308[9:0] ? 4'hb : _GEN_20903; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20905 = 10'h2f8 == _T_308[9:0] ? 4'h8 : _GEN_20904; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20906 = 10'h2f9 == _T_308[9:0] ? 4'h9 : _GEN_20905; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20907 = 10'h2fa == _T_308[9:0] ? 4'hb : _GEN_20906; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20908 = 10'h2fb == _T_308[9:0] ? 4'hb : _GEN_20907; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20909 = 10'h2fc == _T_308[9:0] ? 4'ha : _GEN_20908; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20910 = 10'h2fd == _T_308[9:0] ? 4'ha : _GEN_20909; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20911 = 10'h2fe == _T_308[9:0] ? 4'h9 : _GEN_20910; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20912 = 10'h2ff == _T_308[9:0] ? 4'h8 : _GEN_20911; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20913 = 10'h300 == _T_308[9:0] ? 4'h8 : _GEN_20912; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20914 = 10'h301 == _T_308[9:0] ? 4'h6 : _GEN_20913; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20915 = 10'h302 == _T_308[9:0] ? 4'h1 : _GEN_20914; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20916 = 10'h303 == _T_308[9:0] ? 4'h0 : _GEN_20915; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20917 = 10'h304 == _T_308[9:0] ? 4'h0 : _GEN_20916; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20918 = 10'h305 == _T_308[9:0] ? 4'h0 : _GEN_20917; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20919 = 10'h306 == _T_308[9:0] ? 4'h0 : _GEN_20918; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20920 = 10'h307 == _T_308[9:0] ? 4'h0 : _GEN_20919; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20921 = 10'h308 == _T_308[9:0] ? 4'h0 : _GEN_20920; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20922 = 10'h309 == _T_308[9:0] ? 4'h0 : _GEN_20921; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20923 = 10'h30a == _T_308[9:0] ? 4'h0 : _GEN_20922; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20924 = 10'h30b == _T_308[9:0] ? 4'h0 : _GEN_20923; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20925 = 10'h30c == _T_308[9:0] ? 4'h2 : _GEN_20924; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20926 = 10'h30d == _T_308[9:0] ? 4'h3 : _GEN_20925; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20927 = 10'h30e == _T_308[9:0] ? 4'h3 : _GEN_20926; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20928 = 10'h30f == _T_308[9:0] ? 4'h3 : _GEN_20927; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20929 = 10'h310 == _T_308[9:0] ? 4'h3 : _GEN_20928; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20930 = 10'h311 == _T_308[9:0] ? 4'h3 : _GEN_20929; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20931 = 10'h312 == _T_308[9:0] ? 4'h4 : _GEN_20930; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20932 = 10'h313 == _T_308[9:0] ? 4'h5 : _GEN_20931; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20933 = 10'h314 == _T_308[9:0] ? 4'h5 : _GEN_20932; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20934 = 10'h315 == _T_308[9:0] ? 4'h8 : _GEN_20933; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20935 = 10'h316 == _T_308[9:0] ? 4'h4 : _GEN_20934; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20936 = 10'h317 == _T_308[9:0] ? 4'h6 : _GEN_20935; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20937 = 10'h318 == _T_308[9:0] ? 4'hb : _GEN_20936; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20938 = 10'h319 == _T_308[9:0] ? 4'hb : _GEN_20937; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20939 = 10'h31a == _T_308[9:0] ? 4'hb : _GEN_20938; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20940 = 10'h31b == _T_308[9:0] ? 4'hb : _GEN_20939; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20941 = 10'h31c == _T_308[9:0] ? 4'hb : _GEN_20940; // @[Filter.scala 230:102]
  wire [3:0] _GEN_20942 = 10'h31d == _T_308[9:0] ? 4'hb : _GEN_20941; // @[Filter.scala 230:102]
  wire [6:0] _GEN_39004 = {{3'd0}, _GEN_20942}; // @[Filter.scala 230:102]
  wire [10:0] _T_315 = _GEN_39004 * 7'h46; // @[Filter.scala 230:102]
  wire [10:0] _GEN_39005 = {{2'd0}, _T_310}; // @[Filter.scala 230:69]
  wire [10:0] _T_317 = _GEN_39005 + _T_315; // @[Filter.scala 230:69]
  wire [3:0] _GEN_20965 = 10'h16 == _T_308[9:0] ? 4'hb : 4'hc; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20966 = 10'h17 == _T_308[9:0] ? 4'h8 : _GEN_20965; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20967 = 10'h18 == _T_308[9:0] ? 4'ha : _GEN_20966; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20968 = 10'h19 == _T_308[9:0] ? 4'hc : _GEN_20967; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20969 = 10'h1a == _T_308[9:0] ? 4'hc : _GEN_20968; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20970 = 10'h1b == _T_308[9:0] ? 4'hc : _GEN_20969; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20971 = 10'h1c == _T_308[9:0] ? 4'hc : _GEN_20970; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20972 = 10'h1d == _T_308[9:0] ? 4'hc : _GEN_20971; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20973 = 10'h1e == _T_308[9:0] ? 4'hc : _GEN_20972; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20974 = 10'h1f == _T_308[9:0] ? 4'hc : _GEN_20973; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20975 = 10'h20 == _T_308[9:0] ? 4'hc : _GEN_20974; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20976 = 10'h21 == _T_308[9:0] ? 4'hc : _GEN_20975; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20977 = 10'h22 == _T_308[9:0] ? 4'hc : _GEN_20976; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20978 = 10'h23 == _T_308[9:0] ? 4'hc : _GEN_20977; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20979 = 10'h24 == _T_308[9:0] ? 4'hc : _GEN_20978; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20980 = 10'h25 == _T_308[9:0] ? 4'hc : _GEN_20979; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20981 = 10'h26 == _T_308[9:0] ? 4'hc : _GEN_20980; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20982 = 10'h27 == _T_308[9:0] ? 4'hc : _GEN_20981; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20983 = 10'h28 == _T_308[9:0] ? 4'hc : _GEN_20982; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20984 = 10'h29 == _T_308[9:0] ? 4'hc : _GEN_20983; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20985 = 10'h2a == _T_308[9:0] ? 4'hc : _GEN_20984; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20986 = 10'h2b == _T_308[9:0] ? 4'hc : _GEN_20985; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20987 = 10'h2c == _T_308[9:0] ? 4'hc : _GEN_20986; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20988 = 10'h2d == _T_308[9:0] ? 4'hc : _GEN_20987; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20989 = 10'h2e == _T_308[9:0] ? 4'hc : _GEN_20988; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20990 = 10'h2f == _T_308[9:0] ? 4'hc : _GEN_20989; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20991 = 10'h30 == _T_308[9:0] ? 4'hc : _GEN_20990; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20992 = 10'h31 == _T_308[9:0] ? 4'hc : _GEN_20991; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20993 = 10'h32 == _T_308[9:0] ? 4'hc : _GEN_20992; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20994 = 10'h33 == _T_308[9:0] ? 4'hc : _GEN_20993; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20995 = 10'h34 == _T_308[9:0] ? 4'hc : _GEN_20994; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20996 = 10'h35 == _T_308[9:0] ? 4'hc : _GEN_20995; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20997 = 10'h36 == _T_308[9:0] ? 4'hc : _GEN_20996; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20998 = 10'h37 == _T_308[9:0] ? 4'hc : _GEN_20997; // @[Filter.scala 230:142]
  wire [3:0] _GEN_20999 = 10'h38 == _T_308[9:0] ? 4'hc : _GEN_20998; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21000 = 10'h39 == _T_308[9:0] ? 4'hc : _GEN_20999; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21001 = 10'h3a == _T_308[9:0] ? 4'hc : _GEN_21000; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21002 = 10'h3b == _T_308[9:0] ? 4'hc : _GEN_21001; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21003 = 10'h3c == _T_308[9:0] ? 4'h7 : _GEN_21002; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21004 = 10'h3d == _T_308[9:0] ? 4'h9 : _GEN_21003; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21005 = 10'h3e == _T_308[9:0] ? 4'h8 : _GEN_21004; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21006 = 10'h3f == _T_308[9:0] ? 4'hc : _GEN_21005; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21007 = 10'h40 == _T_308[9:0] ? 4'hc : _GEN_21006; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21008 = 10'h41 == _T_308[9:0] ? 4'hc : _GEN_21007; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21009 = 10'h42 == _T_308[9:0] ? 4'hc : _GEN_21008; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21010 = 10'h43 == _T_308[9:0] ? 4'hc : _GEN_21009; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21011 = 10'h44 == _T_308[9:0] ? 4'hc : _GEN_21010; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21012 = 10'h45 == _T_308[9:0] ? 4'hc : _GEN_21011; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21013 = 10'h46 == _T_308[9:0] ? 4'hc : _GEN_21012; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21014 = 10'h47 == _T_308[9:0] ? 4'hc : _GEN_21013; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21015 = 10'h48 == _T_308[9:0] ? 4'hc : _GEN_21014; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21016 = 10'h49 == _T_308[9:0] ? 4'hc : _GEN_21015; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21017 = 10'h4a == _T_308[9:0] ? 4'hc : _GEN_21016; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21018 = 10'h4b == _T_308[9:0] ? 4'hc : _GEN_21017; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21019 = 10'h4c == _T_308[9:0] ? 4'hc : _GEN_21018; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21020 = 10'h4d == _T_308[9:0] ? 4'hc : _GEN_21019; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21021 = 10'h4e == _T_308[9:0] ? 4'hc : _GEN_21020; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21022 = 10'h4f == _T_308[9:0] ? 4'hc : _GEN_21021; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21023 = 10'h50 == _T_308[9:0] ? 4'hc : _GEN_21022; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21024 = 10'h51 == _T_308[9:0] ? 4'hc : _GEN_21023; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21025 = 10'h52 == _T_308[9:0] ? 4'hc : _GEN_21024; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21026 = 10'h53 == _T_308[9:0] ? 4'hc : _GEN_21025; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21027 = 10'h54 == _T_308[9:0] ? 4'hc : _GEN_21026; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21028 = 10'h55 == _T_308[9:0] ? 4'hc : _GEN_21027; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21029 = 10'h56 == _T_308[9:0] ? 4'hc : _GEN_21028; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21030 = 10'h57 == _T_308[9:0] ? 4'hc : _GEN_21029; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21031 = 10'h58 == _T_308[9:0] ? 4'hc : _GEN_21030; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21032 = 10'h59 == _T_308[9:0] ? 4'hc : _GEN_21031; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21033 = 10'h5a == _T_308[9:0] ? 4'h9 : _GEN_21032; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21034 = 10'h5b == _T_308[9:0] ? 4'ha : _GEN_21033; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21035 = 10'h5c == _T_308[9:0] ? 4'hc : _GEN_21034; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21036 = 10'h5d == _T_308[9:0] ? 4'hc : _GEN_21035; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21037 = 10'h5e == _T_308[9:0] ? 4'hc : _GEN_21036; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21038 = 10'h5f == _T_308[9:0] ? 4'hc : _GEN_21037; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21039 = 10'h60 == _T_308[9:0] ? 4'hc : _GEN_21038; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21040 = 10'h61 == _T_308[9:0] ? 4'hb : _GEN_21039; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21041 = 10'h62 == _T_308[9:0] ? 4'h8 : _GEN_21040; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21042 = 10'h63 == _T_308[9:0] ? 4'h9 : _GEN_21041; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21043 = 10'h64 == _T_308[9:0] ? 4'h7 : _GEN_21042; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21044 = 10'h65 == _T_308[9:0] ? 4'hb : _GEN_21043; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21045 = 10'h66 == _T_308[9:0] ? 4'hc : _GEN_21044; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21046 = 10'h67 == _T_308[9:0] ? 4'hc : _GEN_21045; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21047 = 10'h68 == _T_308[9:0] ? 4'hc : _GEN_21046; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21048 = 10'h69 == _T_308[9:0] ? 4'hc : _GEN_21047; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21049 = 10'h6a == _T_308[9:0] ? 4'hc : _GEN_21048; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21050 = 10'h6b == _T_308[9:0] ? 4'hb : _GEN_21049; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21051 = 10'h6c == _T_308[9:0] ? 4'h9 : _GEN_21050; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21052 = 10'h6d == _T_308[9:0] ? 4'ha : _GEN_21051; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21053 = 10'h6e == _T_308[9:0] ? 4'hc : _GEN_21052; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21054 = 10'h6f == _T_308[9:0] ? 4'hc : _GEN_21053; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21055 = 10'h70 == _T_308[9:0] ? 4'hc : _GEN_21054; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21056 = 10'h71 == _T_308[9:0] ? 4'hc : _GEN_21055; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21057 = 10'h72 == _T_308[9:0] ? 4'hc : _GEN_21056; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21058 = 10'h73 == _T_308[9:0] ? 4'hc : _GEN_21057; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21059 = 10'h74 == _T_308[9:0] ? 4'hc : _GEN_21058; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21060 = 10'h75 == _T_308[9:0] ? 4'hc : _GEN_21059; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21061 = 10'h76 == _T_308[9:0] ? 4'hc : _GEN_21060; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21062 = 10'h77 == _T_308[9:0] ? 4'hc : _GEN_21061; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21063 = 10'h78 == _T_308[9:0] ? 4'hc : _GEN_21062; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21064 = 10'h79 == _T_308[9:0] ? 4'hc : _GEN_21063; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21065 = 10'h7a == _T_308[9:0] ? 4'hc : _GEN_21064; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21066 = 10'h7b == _T_308[9:0] ? 4'hc : _GEN_21065; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21067 = 10'h7c == _T_308[9:0] ? 4'hc : _GEN_21066; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21068 = 10'h7d == _T_308[9:0] ? 4'hc : _GEN_21067; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21069 = 10'h7e == _T_308[9:0] ? 4'hc : _GEN_21068; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21070 = 10'h7f == _T_308[9:0] ? 4'hc : _GEN_21069; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21071 = 10'h80 == _T_308[9:0] ? 4'hc : _GEN_21070; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21072 = 10'h81 == _T_308[9:0] ? 4'h9 : _GEN_21071; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21073 = 10'h82 == _T_308[9:0] ? 4'h9 : _GEN_21072; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21074 = 10'h83 == _T_308[9:0] ? 4'h9 : _GEN_21073; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21075 = 10'h84 == _T_308[9:0] ? 4'hc : _GEN_21074; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21076 = 10'h85 == _T_308[9:0] ? 4'hc : _GEN_21075; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21077 = 10'h86 == _T_308[9:0] ? 4'hc : _GEN_21076; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21078 = 10'h87 == _T_308[9:0] ? 4'h8 : _GEN_21077; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21079 = 10'h88 == _T_308[9:0] ? 4'h9 : _GEN_21078; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21080 = 10'h89 == _T_308[9:0] ? 4'h9 : _GEN_21079; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21081 = 10'h8a == _T_308[9:0] ? 4'h9 : _GEN_21080; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21082 = 10'h8b == _T_308[9:0] ? 4'hc : _GEN_21081; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21083 = 10'h8c == _T_308[9:0] ? 4'hc : _GEN_21082; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21084 = 10'h8d == _T_308[9:0] ? 4'hc : _GEN_21083; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21085 = 10'h8e == _T_308[9:0] ? 4'hc : _GEN_21084; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21086 = 10'h8f == _T_308[9:0] ? 4'h9 : _GEN_21085; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21087 = 10'h90 == _T_308[9:0] ? 4'h9 : _GEN_21086; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21088 = 10'h91 == _T_308[9:0] ? 4'h9 : _GEN_21087; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21089 = 10'h92 == _T_308[9:0] ? 4'ha : _GEN_21088; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21090 = 10'h93 == _T_308[9:0] ? 4'hc : _GEN_21089; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21091 = 10'h94 == _T_308[9:0] ? 4'hc : _GEN_21090; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21092 = 10'h95 == _T_308[9:0] ? 4'hc : _GEN_21091; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21093 = 10'h96 == _T_308[9:0] ? 4'hc : _GEN_21092; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21094 = 10'h97 == _T_308[9:0] ? 4'hc : _GEN_21093; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21095 = 10'h98 == _T_308[9:0] ? 4'hc : _GEN_21094; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21096 = 10'h99 == _T_308[9:0] ? 4'hc : _GEN_21095; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21097 = 10'h9a == _T_308[9:0] ? 4'hc : _GEN_21096; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21098 = 10'h9b == _T_308[9:0] ? 4'hc : _GEN_21097; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21099 = 10'h9c == _T_308[9:0] ? 4'hc : _GEN_21098; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21100 = 10'h9d == _T_308[9:0] ? 4'hc : _GEN_21099; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21101 = 10'h9e == _T_308[9:0] ? 4'hc : _GEN_21100; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21102 = 10'h9f == _T_308[9:0] ? 4'hc : _GEN_21101; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21103 = 10'ha0 == _T_308[9:0] ? 4'hc : _GEN_21102; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21104 = 10'ha1 == _T_308[9:0] ? 4'hc : _GEN_21103; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21105 = 10'ha2 == _T_308[9:0] ? 4'hc : _GEN_21104; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21106 = 10'ha3 == _T_308[9:0] ? 4'hc : _GEN_21105; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21107 = 10'ha4 == _T_308[9:0] ? 4'hc : _GEN_21106; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21108 = 10'ha5 == _T_308[9:0] ? 4'hc : _GEN_21107; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21109 = 10'ha6 == _T_308[9:0] ? 4'hc : _GEN_21108; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21110 = 10'ha7 == _T_308[9:0] ? 4'hc : _GEN_21109; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21111 = 10'ha8 == _T_308[9:0] ? 4'h9 : _GEN_21110; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21112 = 10'ha9 == _T_308[9:0] ? 4'h8 : _GEN_21111; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21113 = 10'haa == _T_308[9:0] ? 4'h8 : _GEN_21112; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21114 = 10'hab == _T_308[9:0] ? 4'ha : _GEN_21113; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21115 = 10'hac == _T_308[9:0] ? 4'hb : _GEN_21114; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21116 = 10'had == _T_308[9:0] ? 4'h7 : _GEN_21115; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21117 = 10'hae == _T_308[9:0] ? 4'h9 : _GEN_21116; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21118 = 10'haf == _T_308[9:0] ? 4'h9 : _GEN_21117; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21119 = 10'hb0 == _T_308[9:0] ? 4'h8 : _GEN_21118; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21120 = 10'hb1 == _T_308[9:0] ? 4'h9 : _GEN_21119; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21121 = 10'hb2 == _T_308[9:0] ? 4'hc : _GEN_21120; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21122 = 10'hb3 == _T_308[9:0] ? 4'h9 : _GEN_21121; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21123 = 10'hb4 == _T_308[9:0] ? 4'h9 : _GEN_21122; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21124 = 10'hb5 == _T_308[9:0] ? 4'h9 : _GEN_21123; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21125 = 10'hb6 == _T_308[9:0] ? 4'h9 : _GEN_21124; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21126 = 10'hb7 == _T_308[9:0] ? 4'ha : _GEN_21125; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21127 = 10'hb8 == _T_308[9:0] ? 4'hc : _GEN_21126; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21128 = 10'hb9 == _T_308[9:0] ? 4'hc : _GEN_21127; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21129 = 10'hba == _T_308[9:0] ? 4'hc : _GEN_21128; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21130 = 10'hbb == _T_308[9:0] ? 4'hc : _GEN_21129; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21131 = 10'hbc == _T_308[9:0] ? 4'hc : _GEN_21130; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21132 = 10'hbd == _T_308[9:0] ? 4'hb : _GEN_21131; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21133 = 10'hbe == _T_308[9:0] ? 4'hc : _GEN_21132; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21134 = 10'hbf == _T_308[9:0] ? 4'hc : _GEN_21133; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21135 = 10'hc0 == _T_308[9:0] ? 4'hc : _GEN_21134; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21136 = 10'hc1 == _T_308[9:0] ? 4'hc : _GEN_21135; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21137 = 10'hc2 == _T_308[9:0] ? 4'hc : _GEN_21136; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21138 = 10'hc3 == _T_308[9:0] ? 4'hc : _GEN_21137; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21139 = 10'hc4 == _T_308[9:0] ? 4'hc : _GEN_21138; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21140 = 10'hc5 == _T_308[9:0] ? 4'hc : _GEN_21139; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21141 = 10'hc6 == _T_308[9:0] ? 4'hb : _GEN_21140; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21142 = 10'hc7 == _T_308[9:0] ? 4'hb : _GEN_21141; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21143 = 10'hc8 == _T_308[9:0] ? 4'ha : _GEN_21142; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21144 = 10'hc9 == _T_308[9:0] ? 4'ha : _GEN_21143; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21145 = 10'hca == _T_308[9:0] ? 4'hb : _GEN_21144; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21146 = 10'hcb == _T_308[9:0] ? 4'hc : _GEN_21145; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21147 = 10'hcc == _T_308[9:0] ? 4'hc : _GEN_21146; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21148 = 10'hcd == _T_308[9:0] ? 4'hc : _GEN_21147; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21149 = 10'hce == _T_308[9:0] ? 4'ha : _GEN_21148; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21150 = 10'hcf == _T_308[9:0] ? 4'h8 : _GEN_21149; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21151 = 10'hd0 == _T_308[9:0] ? 4'h9 : _GEN_21150; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21152 = 10'hd1 == _T_308[9:0] ? 4'h8 : _GEN_21151; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21153 = 10'hd2 == _T_308[9:0] ? 4'h9 : _GEN_21152; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21154 = 10'hd3 == _T_308[9:0] ? 4'h9 : _GEN_21153; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21155 = 10'hd4 == _T_308[9:0] ? 4'h9 : _GEN_21154; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21156 = 10'hd5 == _T_308[9:0] ? 4'h9 : _GEN_21155; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21157 = 10'hd6 == _T_308[9:0] ? 4'ha : _GEN_21156; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21158 = 10'hd7 == _T_308[9:0] ? 4'h9 : _GEN_21157; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21159 = 10'hd8 == _T_308[9:0] ? 4'h9 : _GEN_21158; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21160 = 10'hd9 == _T_308[9:0] ? 4'h9 : _GEN_21159; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21161 = 10'hda == _T_308[9:0] ? 4'ha : _GEN_21160; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21162 = 10'hdb == _T_308[9:0] ? 4'h9 : _GEN_21161; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21163 = 10'hdc == _T_308[9:0] ? 4'h7 : _GEN_21162; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21164 = 10'hdd == _T_308[9:0] ? 4'hc : _GEN_21163; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21165 = 10'hde == _T_308[9:0] ? 4'hc : _GEN_21164; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21166 = 10'hdf == _T_308[9:0] ? 4'hc : _GEN_21165; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21167 = 10'he0 == _T_308[9:0] ? 4'hc : _GEN_21166; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21168 = 10'he1 == _T_308[9:0] ? 4'hc : _GEN_21167; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21169 = 10'he2 == _T_308[9:0] ? 4'hc : _GEN_21168; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21170 = 10'he3 == _T_308[9:0] ? 4'h8 : _GEN_21169; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21171 = 10'he4 == _T_308[9:0] ? 4'hc : _GEN_21170; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21172 = 10'he5 == _T_308[9:0] ? 4'hc : _GEN_21171; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21173 = 10'he6 == _T_308[9:0] ? 4'hc : _GEN_21172; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21174 = 10'he7 == _T_308[9:0] ? 4'hc : _GEN_21173; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21175 = 10'he8 == _T_308[9:0] ? 4'hc : _GEN_21174; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21176 = 10'he9 == _T_308[9:0] ? 4'hc : _GEN_21175; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21177 = 10'hea == _T_308[9:0] ? 4'hc : _GEN_21176; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21178 = 10'heb == _T_308[9:0] ? 4'ha : _GEN_21177; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21179 = 10'hec == _T_308[9:0] ? 4'h7 : _GEN_21178; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21180 = 10'hed == _T_308[9:0] ? 4'h3 : _GEN_21179; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21181 = 10'hee == _T_308[9:0] ? 4'h3 : _GEN_21180; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21182 = 10'hef == _T_308[9:0] ? 4'h3 : _GEN_21181; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21183 = 10'hf0 == _T_308[9:0] ? 4'h3 : _GEN_21182; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21184 = 10'hf1 == _T_308[9:0] ? 4'h8 : _GEN_21183; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21185 = 10'hf2 == _T_308[9:0] ? 4'hc : _GEN_21184; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21186 = 10'hf3 == _T_308[9:0] ? 4'hc : _GEN_21185; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21187 = 10'hf4 == _T_308[9:0] ? 4'hc : _GEN_21186; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21188 = 10'hf5 == _T_308[9:0] ? 4'h9 : _GEN_21187; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21189 = 10'hf6 == _T_308[9:0] ? 4'h9 : _GEN_21188; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21190 = 10'hf7 == _T_308[9:0] ? 4'h9 : _GEN_21189; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21191 = 10'hf8 == _T_308[9:0] ? 4'h9 : _GEN_21190; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21192 = 10'hf9 == _T_308[9:0] ? 4'ha : _GEN_21191; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21193 = 10'hfa == _T_308[9:0] ? 4'h9 : _GEN_21192; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21194 = 10'hfb == _T_308[9:0] ? 4'h9 : _GEN_21193; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21195 = 10'hfc == _T_308[9:0] ? 4'h9 : _GEN_21194; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21196 = 10'hfd == _T_308[9:0] ? 4'h9 : _GEN_21195; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21197 = 10'hfe == _T_308[9:0] ? 4'h9 : _GEN_21196; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21198 = 10'hff == _T_308[9:0] ? 4'ha : _GEN_21197; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21199 = 10'h100 == _T_308[9:0] ? 4'ha : _GEN_21198; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21200 = 10'h101 == _T_308[9:0] ? 4'h7 : _GEN_21199; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21201 = 10'h102 == _T_308[9:0] ? 4'h9 : _GEN_21200; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21202 = 10'h103 == _T_308[9:0] ? 4'hc : _GEN_21201; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21203 = 10'h104 == _T_308[9:0] ? 4'hc : _GEN_21202; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21204 = 10'h105 == _T_308[9:0] ? 4'hb : _GEN_21203; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21205 = 10'h106 == _T_308[9:0] ? 4'hb : _GEN_21204; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21206 = 10'h107 == _T_308[9:0] ? 4'hb : _GEN_21205; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21207 = 10'h108 == _T_308[9:0] ? 4'hb : _GEN_21206; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21208 = 10'h109 == _T_308[9:0] ? 4'h7 : _GEN_21207; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21209 = 10'h10a == _T_308[9:0] ? 4'hc : _GEN_21208; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21210 = 10'h10b == _T_308[9:0] ? 4'hc : _GEN_21209; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21211 = 10'h10c == _T_308[9:0] ? 4'hc : _GEN_21210; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21212 = 10'h10d == _T_308[9:0] ? 4'hc : _GEN_21211; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21213 = 10'h10e == _T_308[9:0] ? 4'hc : _GEN_21212; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21214 = 10'h10f == _T_308[9:0] ? 4'h9 : _GEN_21213; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21215 = 10'h110 == _T_308[9:0] ? 4'hb : _GEN_21214; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21216 = 10'h111 == _T_308[9:0] ? 4'h4 : _GEN_21215; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21217 = 10'h112 == _T_308[9:0] ? 4'h7 : _GEN_21216; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21218 = 10'h113 == _T_308[9:0] ? 4'h3 : _GEN_21217; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21219 = 10'h114 == _T_308[9:0] ? 4'h3 : _GEN_21218; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21220 = 10'h115 == _T_308[9:0] ? 4'h3 : _GEN_21219; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21221 = 10'h116 == _T_308[9:0] ? 4'h3 : _GEN_21220; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21222 = 10'h117 == _T_308[9:0] ? 4'h2 : _GEN_21221; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21223 = 10'h118 == _T_308[9:0] ? 4'h9 : _GEN_21222; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21224 = 10'h119 == _T_308[9:0] ? 4'hc : _GEN_21223; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21225 = 10'h11a == _T_308[9:0] ? 4'hc : _GEN_21224; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21226 = 10'h11b == _T_308[9:0] ? 4'hc : _GEN_21225; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21227 = 10'h11c == _T_308[9:0] ? 4'h9 : _GEN_21226; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21228 = 10'h11d == _T_308[9:0] ? 4'h9 : _GEN_21227; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21229 = 10'h11e == _T_308[9:0] ? 4'h9 : _GEN_21228; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21230 = 10'h11f == _T_308[9:0] ? 4'h8 : _GEN_21229; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21231 = 10'h120 == _T_308[9:0] ? 4'h7 : _GEN_21230; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21232 = 10'h121 == _T_308[9:0] ? 4'h9 : _GEN_21231; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21233 = 10'h122 == _T_308[9:0] ? 4'h7 : _GEN_21232; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21234 = 10'h123 == _T_308[9:0] ? 4'h7 : _GEN_21233; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21235 = 10'h124 == _T_308[9:0] ? 4'h9 : _GEN_21234; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21236 = 10'h125 == _T_308[9:0] ? 4'h9 : _GEN_21235; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21237 = 10'h126 == _T_308[9:0] ? 4'h8 : _GEN_21236; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21238 = 10'h127 == _T_308[9:0] ? 4'h9 : _GEN_21237; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21239 = 10'h128 == _T_308[9:0] ? 4'h8 : _GEN_21238; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21240 = 10'h129 == _T_308[9:0] ? 4'ha : _GEN_21239; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21241 = 10'h12a == _T_308[9:0] ? 4'h5 : _GEN_21240; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21242 = 10'h12b == _T_308[9:0] ? 4'h3 : _GEN_21241; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21243 = 10'h12c == _T_308[9:0] ? 4'h3 : _GEN_21242; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21244 = 10'h12d == _T_308[9:0] ? 4'h3 : _GEN_21243; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21245 = 10'h12e == _T_308[9:0] ? 4'h5 : _GEN_21244; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21246 = 10'h12f == _T_308[9:0] ? 4'h8 : _GEN_21245; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21247 = 10'h130 == _T_308[9:0] ? 4'hc : _GEN_21246; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21248 = 10'h131 == _T_308[9:0] ? 4'hb : _GEN_21247; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21249 = 10'h132 == _T_308[9:0] ? 4'h9 : _GEN_21248; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21250 = 10'h133 == _T_308[9:0] ? 4'h8 : _GEN_21249; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21251 = 10'h134 == _T_308[9:0] ? 4'h9 : _GEN_21250; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21252 = 10'h135 == _T_308[9:0] ? 4'h7 : _GEN_21251; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21253 = 10'h136 == _T_308[9:0] ? 4'h7 : _GEN_21252; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21254 = 10'h137 == _T_308[9:0] ? 4'h5 : _GEN_21253; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21255 = 10'h138 == _T_308[9:0] ? 4'h7 : _GEN_21254; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21256 = 10'h139 == _T_308[9:0] ? 4'h3 : _GEN_21255; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21257 = 10'h13a == _T_308[9:0] ? 4'h3 : _GEN_21256; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21258 = 10'h13b == _T_308[9:0] ? 4'h3 : _GEN_21257; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21259 = 10'h13c == _T_308[9:0] ? 4'h3 : _GEN_21258; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21260 = 10'h13d == _T_308[9:0] ? 4'h3 : _GEN_21259; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21261 = 10'h13e == _T_308[9:0] ? 4'h5 : _GEN_21260; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21262 = 10'h13f == _T_308[9:0] ? 4'ha : _GEN_21261; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21263 = 10'h140 == _T_308[9:0] ? 4'hc : _GEN_21262; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21264 = 10'h141 == _T_308[9:0] ? 4'hc : _GEN_21263; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21265 = 10'h142 == _T_308[9:0] ? 4'hc : _GEN_21264; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21266 = 10'h143 == _T_308[9:0] ? 4'h9 : _GEN_21265; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21267 = 10'h144 == _T_308[9:0] ? 4'h9 : _GEN_21266; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21268 = 10'h145 == _T_308[9:0] ? 4'h8 : _GEN_21267; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21269 = 10'h146 == _T_308[9:0] ? 4'h8 : _GEN_21268; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21270 = 10'h147 == _T_308[9:0] ? 4'h7 : _GEN_21269; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21271 = 10'h148 == _T_308[9:0] ? 4'h8 : _GEN_21270; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21272 = 10'h149 == _T_308[9:0] ? 4'h9 : _GEN_21271; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21273 = 10'h14a == _T_308[9:0] ? 4'ha : _GEN_21272; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21274 = 10'h14b == _T_308[9:0] ? 4'h9 : _GEN_21273; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21275 = 10'h14c == _T_308[9:0] ? 4'ha : _GEN_21274; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21276 = 10'h14d == _T_308[9:0] ? 4'h9 : _GEN_21275; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21277 = 10'h14e == _T_308[9:0] ? 4'h7 : _GEN_21276; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21278 = 10'h14f == _T_308[9:0] ? 4'h3 : _GEN_21277; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21279 = 10'h150 == _T_308[9:0] ? 4'h3 : _GEN_21278; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21280 = 10'h151 == _T_308[9:0] ? 4'h3 : _GEN_21279; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21281 = 10'h152 == _T_308[9:0] ? 4'h3 : _GEN_21280; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21282 = 10'h153 == _T_308[9:0] ? 4'h3 : _GEN_21281; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21283 = 10'h154 == _T_308[9:0] ? 4'h3 : _GEN_21282; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21284 = 10'h155 == _T_308[9:0] ? 4'h8 : _GEN_21283; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21285 = 10'h156 == _T_308[9:0] ? 4'ha : _GEN_21284; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21286 = 10'h157 == _T_308[9:0] ? 4'h7 : _GEN_21285; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21287 = 10'h158 == _T_308[9:0] ? 4'h7 : _GEN_21286; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21288 = 10'h159 == _T_308[9:0] ? 4'h7 : _GEN_21287; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21289 = 10'h15a == _T_308[9:0] ? 4'h7 : _GEN_21288; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21290 = 10'h15b == _T_308[9:0] ? 4'h7 : _GEN_21289; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21291 = 10'h15c == _T_308[9:0] ? 4'h7 : _GEN_21290; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21292 = 10'h15d == _T_308[9:0] ? 4'h7 : _GEN_21291; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21293 = 10'h15e == _T_308[9:0] ? 4'h7 : _GEN_21292; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21294 = 10'h15f == _T_308[9:0] ? 4'h3 : _GEN_21293; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21295 = 10'h160 == _T_308[9:0] ? 4'h3 : _GEN_21294; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21296 = 10'h161 == _T_308[9:0] ? 4'h3 : _GEN_21295; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21297 = 10'h162 == _T_308[9:0] ? 4'h3 : _GEN_21296; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21298 = 10'h163 == _T_308[9:0] ? 4'h3 : _GEN_21297; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21299 = 10'h164 == _T_308[9:0] ? 4'h4 : _GEN_21298; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21300 = 10'h165 == _T_308[9:0] ? 4'ha : _GEN_21299; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21301 = 10'h166 == _T_308[9:0] ? 4'ha : _GEN_21300; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21302 = 10'h167 == _T_308[9:0] ? 4'hc : _GEN_21301; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21303 = 10'h168 == _T_308[9:0] ? 4'hc : _GEN_21302; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21304 = 10'h169 == _T_308[9:0] ? 4'h9 : _GEN_21303; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21305 = 10'h16a == _T_308[9:0] ? 4'h9 : _GEN_21304; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21306 = 10'h16b == _T_308[9:0] ? 4'ha : _GEN_21305; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21307 = 10'h16c == _T_308[9:0] ? 4'h7 : _GEN_21306; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21308 = 10'h16d == _T_308[9:0] ? 4'h7 : _GEN_21307; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21309 = 10'h16e == _T_308[9:0] ? 4'h7 : _GEN_21308; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21310 = 10'h16f == _T_308[9:0] ? 4'ha : _GEN_21309; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21311 = 10'h170 == _T_308[9:0] ? 4'ha : _GEN_21310; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21312 = 10'h171 == _T_308[9:0] ? 4'ha : _GEN_21311; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21313 = 10'h172 == _T_308[9:0] ? 4'hc : _GEN_21312; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21314 = 10'h173 == _T_308[9:0] ? 4'h8 : _GEN_21313; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21315 = 10'h174 == _T_308[9:0] ? 4'h5 : _GEN_21314; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21316 = 10'h175 == _T_308[9:0] ? 4'h8 : _GEN_21315; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21317 = 10'h176 == _T_308[9:0] ? 4'h7 : _GEN_21316; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21318 = 10'h177 == _T_308[9:0] ? 4'h8 : _GEN_21317; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21319 = 10'h178 == _T_308[9:0] ? 4'h7 : _GEN_21318; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21320 = 10'h179 == _T_308[9:0] ? 4'h5 : _GEN_21319; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21321 = 10'h17a == _T_308[9:0] ? 4'h5 : _GEN_21320; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21322 = 10'h17b == _T_308[9:0] ? 4'h7 : _GEN_21321; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21323 = 10'h17c == _T_308[9:0] ? 4'h7 : _GEN_21322; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21324 = 10'h17d == _T_308[9:0] ? 4'h7 : _GEN_21323; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21325 = 10'h17e == _T_308[9:0] ? 4'h7 : _GEN_21324; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21326 = 10'h17f == _T_308[9:0] ? 4'h7 : _GEN_21325; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21327 = 10'h180 == _T_308[9:0] ? 4'h7 : _GEN_21326; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21328 = 10'h181 == _T_308[9:0] ? 4'h7 : _GEN_21327; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21329 = 10'h182 == _T_308[9:0] ? 4'h7 : _GEN_21328; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21330 = 10'h183 == _T_308[9:0] ? 4'h7 : _GEN_21329; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21331 = 10'h184 == _T_308[9:0] ? 4'h7 : _GEN_21330; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21332 = 10'h185 == _T_308[9:0] ? 4'h5 : _GEN_21331; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21333 = 10'h186 == _T_308[9:0] ? 4'h3 : _GEN_21332; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21334 = 10'h187 == _T_308[9:0] ? 4'h3 : _GEN_21333; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21335 = 10'h188 == _T_308[9:0] ? 4'h3 : _GEN_21334; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21336 = 10'h189 == _T_308[9:0] ? 4'h4 : _GEN_21335; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21337 = 10'h18a == _T_308[9:0] ? 4'h5 : _GEN_21336; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21338 = 10'h18b == _T_308[9:0] ? 4'ha : _GEN_21337; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21339 = 10'h18c == _T_308[9:0] ? 4'ha : _GEN_21338; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21340 = 10'h18d == _T_308[9:0] ? 4'ha : _GEN_21339; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21341 = 10'h18e == _T_308[9:0] ? 4'hc : _GEN_21340; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21342 = 10'h18f == _T_308[9:0] ? 4'h8 : _GEN_21341; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21343 = 10'h190 == _T_308[9:0] ? 4'h9 : _GEN_21342; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21344 = 10'h191 == _T_308[9:0] ? 4'h8 : _GEN_21343; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21345 = 10'h192 == _T_308[9:0] ? 4'h7 : _GEN_21344; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21346 = 10'h193 == _T_308[9:0] ? 4'h7 : _GEN_21345; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21347 = 10'h194 == _T_308[9:0] ? 4'h7 : _GEN_21346; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21348 = 10'h195 == _T_308[9:0] ? 4'h9 : _GEN_21347; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21349 = 10'h196 == _T_308[9:0] ? 4'ha : _GEN_21348; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21350 = 10'h197 == _T_308[9:0] ? 4'h8 : _GEN_21349; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21351 = 10'h198 == _T_308[9:0] ? 4'hc : _GEN_21350; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21352 = 10'h199 == _T_308[9:0] ? 4'h5 : _GEN_21351; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21353 = 10'h19a == _T_308[9:0] ? 4'h1 : _GEN_21352; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21354 = 10'h19b == _T_308[9:0] ? 4'h4 : _GEN_21353; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21355 = 10'h19c == _T_308[9:0] ? 4'h7 : _GEN_21354; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21356 = 10'h19d == _T_308[9:0] ? 4'h5 : _GEN_21355; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21357 = 10'h19e == _T_308[9:0] ? 4'h2 : _GEN_21356; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21358 = 10'h19f == _T_308[9:0] ? 4'h3 : _GEN_21357; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21359 = 10'h1a0 == _T_308[9:0] ? 4'h7 : _GEN_21358; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21360 = 10'h1a1 == _T_308[9:0] ? 4'h7 : _GEN_21359; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21361 = 10'h1a2 == _T_308[9:0] ? 4'h7 : _GEN_21360; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21362 = 10'h1a3 == _T_308[9:0] ? 4'h7 : _GEN_21361; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21363 = 10'h1a4 == _T_308[9:0] ? 4'h7 : _GEN_21362; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21364 = 10'h1a5 == _T_308[9:0] ? 4'h7 : _GEN_21363; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21365 = 10'h1a6 == _T_308[9:0] ? 4'h7 : _GEN_21364; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21366 = 10'h1a7 == _T_308[9:0] ? 4'h7 : _GEN_21365; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21367 = 10'h1a8 == _T_308[9:0] ? 4'h8 : _GEN_21366; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21368 = 10'h1a9 == _T_308[9:0] ? 4'h8 : _GEN_21367; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21369 = 10'h1aa == _T_308[9:0] ? 4'h6 : _GEN_21368; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21370 = 10'h1ab == _T_308[9:0] ? 4'h6 : _GEN_21369; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21371 = 10'h1ac == _T_308[9:0] ? 4'h5 : _GEN_21370; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21372 = 10'h1ad == _T_308[9:0] ? 4'h4 : _GEN_21371; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21373 = 10'h1ae == _T_308[9:0] ? 4'h3 : _GEN_21372; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21374 = 10'h1af == _T_308[9:0] ? 4'h6 : _GEN_21373; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21375 = 10'h1b0 == _T_308[9:0] ? 4'h6 : _GEN_21374; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21376 = 10'h1b1 == _T_308[9:0] ? 4'ha : _GEN_21375; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21377 = 10'h1b2 == _T_308[9:0] ? 4'ha : _GEN_21376; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21378 = 10'h1b3 == _T_308[9:0] ? 4'h9 : _GEN_21377; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21379 = 10'h1b4 == _T_308[9:0] ? 4'hb : _GEN_21378; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21380 = 10'h1b5 == _T_308[9:0] ? 4'h8 : _GEN_21379; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21381 = 10'h1b6 == _T_308[9:0] ? 4'h8 : _GEN_21380; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21382 = 10'h1b7 == _T_308[9:0] ? 4'h7 : _GEN_21381; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21383 = 10'h1b8 == _T_308[9:0] ? 4'h6 : _GEN_21382; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21384 = 10'h1b9 == _T_308[9:0] ? 4'h7 : _GEN_21383; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21385 = 10'h1ba == _T_308[9:0] ? 4'h6 : _GEN_21384; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21386 = 10'h1bb == _T_308[9:0] ? 4'h8 : _GEN_21385; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21387 = 10'h1bc == _T_308[9:0] ? 4'ha : _GEN_21386; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21388 = 10'h1bd == _T_308[9:0] ? 4'h9 : _GEN_21387; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21389 = 10'h1be == _T_308[9:0] ? 4'hc : _GEN_21388; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21390 = 10'h1bf == _T_308[9:0] ? 4'h7 : _GEN_21389; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21391 = 10'h1c0 == _T_308[9:0] ? 4'h6 : _GEN_21390; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21392 = 10'h1c1 == _T_308[9:0] ? 4'h7 : _GEN_21391; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21393 = 10'h1c2 == _T_308[9:0] ? 4'h7 : _GEN_21392; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21394 = 10'h1c3 == _T_308[9:0] ? 4'h6 : _GEN_21393; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21395 = 10'h1c4 == _T_308[9:0] ? 4'h5 : _GEN_21394; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21396 = 10'h1c5 == _T_308[9:0] ? 4'h6 : _GEN_21395; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21397 = 10'h1c6 == _T_308[9:0] ? 4'h8 : _GEN_21396; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21398 = 10'h1c7 == _T_308[9:0] ? 4'h7 : _GEN_21397; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21399 = 10'h1c8 == _T_308[9:0] ? 4'h7 : _GEN_21398; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21400 = 10'h1c9 == _T_308[9:0] ? 4'h7 : _GEN_21399; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21401 = 10'h1ca == _T_308[9:0] ? 4'h7 : _GEN_21400; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21402 = 10'h1cb == _T_308[9:0] ? 4'h7 : _GEN_21401; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21403 = 10'h1cc == _T_308[9:0] ? 4'h7 : _GEN_21402; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21404 = 10'h1cd == _T_308[9:0] ? 4'h8 : _GEN_21403; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21405 = 10'h1ce == _T_308[9:0] ? 4'h8 : _GEN_21404; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21406 = 10'h1cf == _T_308[9:0] ? 4'h8 : _GEN_21405; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21407 = 10'h1d0 == _T_308[9:0] ? 4'h5 : _GEN_21406; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21408 = 10'h1d1 == _T_308[9:0] ? 4'h6 : _GEN_21407; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21409 = 10'h1d2 == _T_308[9:0] ? 4'h7 : _GEN_21408; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21410 = 10'h1d3 == _T_308[9:0] ? 4'h7 : _GEN_21409; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21411 = 10'h1d4 == _T_308[9:0] ? 4'h7 : _GEN_21410; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21412 = 10'h1d5 == _T_308[9:0] ? 4'h6 : _GEN_21411; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21413 = 10'h1d6 == _T_308[9:0] ? 4'h8 : _GEN_21412; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21414 = 10'h1d7 == _T_308[9:0] ? 4'ha : _GEN_21413; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21415 = 10'h1d8 == _T_308[9:0] ? 4'ha : _GEN_21414; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21416 = 10'h1d9 == _T_308[9:0] ? 4'ha : _GEN_21415; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21417 = 10'h1da == _T_308[9:0] ? 4'h8 : _GEN_21416; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21418 = 10'h1db == _T_308[9:0] ? 4'h9 : _GEN_21417; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21419 = 10'h1dc == _T_308[9:0] ? 4'h9 : _GEN_21418; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21420 = 10'h1dd == _T_308[9:0] ? 4'h5 : _GEN_21419; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21421 = 10'h1de == _T_308[9:0] ? 4'h7 : _GEN_21420; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21422 = 10'h1df == _T_308[9:0] ? 4'h7 : _GEN_21421; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21423 = 10'h1e0 == _T_308[9:0] ? 4'h7 : _GEN_21422; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21424 = 10'h1e1 == _T_308[9:0] ? 4'h6 : _GEN_21423; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21425 = 10'h1e2 == _T_308[9:0] ? 4'h9 : _GEN_21424; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21426 = 10'h1e3 == _T_308[9:0] ? 4'h9 : _GEN_21425; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21427 = 10'h1e4 == _T_308[9:0] ? 4'hb : _GEN_21426; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21428 = 10'h1e5 == _T_308[9:0] ? 4'h8 : _GEN_21427; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21429 = 10'h1e6 == _T_308[9:0] ? 4'h7 : _GEN_21428; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21430 = 10'h1e7 == _T_308[9:0] ? 4'h8 : _GEN_21429; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21431 = 10'h1e8 == _T_308[9:0] ? 4'h8 : _GEN_21430; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21432 = 10'h1e9 == _T_308[9:0] ? 4'h8 : _GEN_21431; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21433 = 10'h1ea == _T_308[9:0] ? 4'h8 : _GEN_21432; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21434 = 10'h1eb == _T_308[9:0] ? 4'h8 : _GEN_21433; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21435 = 10'h1ec == _T_308[9:0] ? 4'h8 : _GEN_21434; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21436 = 10'h1ed == _T_308[9:0] ? 4'h6 : _GEN_21435; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21437 = 10'h1ee == _T_308[9:0] ? 4'h7 : _GEN_21436; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21438 = 10'h1ef == _T_308[9:0] ? 4'h7 : _GEN_21437; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21439 = 10'h1f0 == _T_308[9:0] ? 4'h7 : _GEN_21438; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21440 = 10'h1f1 == _T_308[9:0] ? 4'h7 : _GEN_21439; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21441 = 10'h1f2 == _T_308[9:0] ? 4'h7 : _GEN_21440; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21442 = 10'h1f3 == _T_308[9:0] ? 4'h8 : _GEN_21441; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21443 = 10'h1f4 == _T_308[9:0] ? 4'h8 : _GEN_21442; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21444 = 10'h1f5 == _T_308[9:0] ? 4'h8 : _GEN_21443; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21445 = 10'h1f6 == _T_308[9:0] ? 4'ha : _GEN_21444; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21446 = 10'h1f7 == _T_308[9:0] ? 4'h6 : _GEN_21445; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21447 = 10'h1f8 == _T_308[9:0] ? 4'h6 : _GEN_21446; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21448 = 10'h1f9 == _T_308[9:0] ? 4'h8 : _GEN_21447; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21449 = 10'h1fa == _T_308[9:0] ? 4'h8 : _GEN_21448; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21450 = 10'h1fb == _T_308[9:0] ? 4'h6 : _GEN_21449; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21451 = 10'h1fc == _T_308[9:0] ? 4'ha : _GEN_21450; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21452 = 10'h1fd == _T_308[9:0] ? 4'hb : _GEN_21451; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21453 = 10'h1fe == _T_308[9:0] ? 4'ha : _GEN_21452; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21454 = 10'h1ff == _T_308[9:0] ? 4'ha : _GEN_21453; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21455 = 10'h200 == _T_308[9:0] ? 4'h4 : _GEN_21454; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21456 = 10'h201 == _T_308[9:0] ? 4'h7 : _GEN_21455; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21457 = 10'h202 == _T_308[9:0] ? 4'h6 : _GEN_21456; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21458 = 10'h203 == _T_308[9:0] ? 4'h6 : _GEN_21457; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21459 = 10'h204 == _T_308[9:0] ? 4'h5 : _GEN_21458; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21460 = 10'h205 == _T_308[9:0] ? 4'h6 : _GEN_21459; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21461 = 10'h206 == _T_308[9:0] ? 4'h6 : _GEN_21460; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21462 = 10'h207 == _T_308[9:0] ? 4'h5 : _GEN_21461; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21463 = 10'h208 == _T_308[9:0] ? 4'h7 : _GEN_21462; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21464 = 10'h209 == _T_308[9:0] ? 4'h9 : _GEN_21463; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21465 = 10'h20a == _T_308[9:0] ? 4'hb : _GEN_21464; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21466 = 10'h20b == _T_308[9:0] ? 4'h7 : _GEN_21465; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21467 = 10'h20c == _T_308[9:0] ? 4'h7 : _GEN_21466; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21468 = 10'h20d == _T_308[9:0] ? 4'h7 : _GEN_21467; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21469 = 10'h20e == _T_308[9:0] ? 4'h7 : _GEN_21468; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21470 = 10'h20f == _T_308[9:0] ? 4'h7 : _GEN_21469; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21471 = 10'h210 == _T_308[9:0] ? 4'h7 : _GEN_21470; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21472 = 10'h211 == _T_308[9:0] ? 4'h8 : _GEN_21471; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21473 = 10'h212 == _T_308[9:0] ? 4'h8 : _GEN_21472; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21474 = 10'h213 == _T_308[9:0] ? 4'h9 : _GEN_21473; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21475 = 10'h214 == _T_308[9:0] ? 4'h6 : _GEN_21474; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21476 = 10'h215 == _T_308[9:0] ? 4'h7 : _GEN_21475; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21477 = 10'h216 == _T_308[9:0] ? 4'h7 : _GEN_21476; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21478 = 10'h217 == _T_308[9:0] ? 4'h7 : _GEN_21477; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21479 = 10'h218 == _T_308[9:0] ? 4'h7 : _GEN_21478; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21480 = 10'h219 == _T_308[9:0] ? 4'h8 : _GEN_21479; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21481 = 10'h21a == _T_308[9:0] ? 4'h7 : _GEN_21480; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21482 = 10'h21b == _T_308[9:0] ? 4'h8 : _GEN_21481; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21483 = 10'h21c == _T_308[9:0] ? 4'ha : _GEN_21482; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21484 = 10'h21d == _T_308[9:0] ? 4'ha : _GEN_21483; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21485 = 10'h21e == _T_308[9:0] ? 4'h7 : _GEN_21484; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21486 = 10'h21f == _T_308[9:0] ? 4'h6 : _GEN_21485; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21487 = 10'h220 == _T_308[9:0] ? 4'h6 : _GEN_21486; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21488 = 10'h221 == _T_308[9:0] ? 4'h7 : _GEN_21487; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21489 = 10'h222 == _T_308[9:0] ? 4'ha : _GEN_21488; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21490 = 10'h223 == _T_308[9:0] ? 4'ha : _GEN_21489; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21491 = 10'h224 == _T_308[9:0] ? 4'ha : _GEN_21490; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21492 = 10'h225 == _T_308[9:0] ? 4'h8 : _GEN_21491; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21493 = 10'h226 == _T_308[9:0] ? 4'h3 : _GEN_21492; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21494 = 10'h227 == _T_308[9:0] ? 4'h4 : _GEN_21493; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21495 = 10'h228 == _T_308[9:0] ? 4'h6 : _GEN_21494; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21496 = 10'h229 == _T_308[9:0] ? 4'h6 : _GEN_21495; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21497 = 10'h22a == _T_308[9:0] ? 4'h6 : _GEN_21496; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21498 = 10'h22b == _T_308[9:0] ? 4'h6 : _GEN_21497; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21499 = 10'h22c == _T_308[9:0] ? 4'h5 : _GEN_21498; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21500 = 10'h22d == _T_308[9:0] ? 4'h6 : _GEN_21499; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21501 = 10'h22e == _T_308[9:0] ? 4'h6 : _GEN_21500; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21502 = 10'h22f == _T_308[9:0] ? 4'h8 : _GEN_21501; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21503 = 10'h230 == _T_308[9:0] ? 4'h7 : _GEN_21502; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21504 = 10'h231 == _T_308[9:0] ? 4'h5 : _GEN_21503; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21505 = 10'h232 == _T_308[9:0] ? 4'h6 : _GEN_21504; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21506 = 10'h233 == _T_308[9:0] ? 4'h8 : _GEN_21505; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21507 = 10'h234 == _T_308[9:0] ? 4'h8 : _GEN_21506; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21508 = 10'h235 == _T_308[9:0] ? 4'h8 : _GEN_21507; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21509 = 10'h236 == _T_308[9:0] ? 4'h8 : _GEN_21508; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21510 = 10'h237 == _T_308[9:0] ? 4'h8 : _GEN_21509; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21511 = 10'h238 == _T_308[9:0] ? 4'h8 : _GEN_21510; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21512 = 10'h239 == _T_308[9:0] ? 4'h6 : _GEN_21511; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21513 = 10'h23a == _T_308[9:0] ? 4'h6 : _GEN_21512; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21514 = 10'h23b == _T_308[9:0] ? 4'h7 : _GEN_21513; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21515 = 10'h23c == _T_308[9:0] ? 4'h6 : _GEN_21514; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21516 = 10'h23d == _T_308[9:0] ? 4'h7 : _GEN_21515; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21517 = 10'h23e == _T_308[9:0] ? 4'h7 : _GEN_21516; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21518 = 10'h23f == _T_308[9:0] ? 4'h6 : _GEN_21517; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21519 = 10'h240 == _T_308[9:0] ? 4'h6 : _GEN_21518; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21520 = 10'h241 == _T_308[9:0] ? 4'h8 : _GEN_21519; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21521 = 10'h242 == _T_308[9:0] ? 4'ha : _GEN_21520; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21522 = 10'h243 == _T_308[9:0] ? 4'ha : _GEN_21521; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21523 = 10'h244 == _T_308[9:0] ? 4'ha : _GEN_21522; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21524 = 10'h245 == _T_308[9:0] ? 4'h8 : _GEN_21523; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21525 = 10'h246 == _T_308[9:0] ? 4'h8 : _GEN_21524; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21526 = 10'h247 == _T_308[9:0] ? 4'h9 : _GEN_21525; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21527 = 10'h248 == _T_308[9:0] ? 4'ha : _GEN_21526; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21528 = 10'h249 == _T_308[9:0] ? 4'ha : _GEN_21527; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21529 = 10'h24a == _T_308[9:0] ? 4'ha : _GEN_21528; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21530 = 10'h24b == _T_308[9:0] ? 4'h4 : _GEN_21529; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21531 = 10'h24c == _T_308[9:0] ? 4'h3 : _GEN_21530; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21532 = 10'h24d == _T_308[9:0] ? 4'h4 : _GEN_21531; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21533 = 10'h24e == _T_308[9:0] ? 4'h5 : _GEN_21532; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21534 = 10'h24f == _T_308[9:0] ? 4'h5 : _GEN_21533; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21535 = 10'h250 == _T_308[9:0] ? 4'h5 : _GEN_21534; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21536 = 10'h251 == _T_308[9:0] ? 4'h5 : _GEN_21535; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21537 = 10'h252 == _T_308[9:0] ? 4'h5 : _GEN_21536; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21538 = 10'h253 == _T_308[9:0] ? 4'h5 : _GEN_21537; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21539 = 10'h254 == _T_308[9:0] ? 4'h5 : _GEN_21538; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21540 = 10'h255 == _T_308[9:0] ? 4'h6 : _GEN_21539; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21541 = 10'h256 == _T_308[9:0] ? 4'h7 : _GEN_21540; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21542 = 10'h257 == _T_308[9:0] ? 4'h3 : _GEN_21541; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21543 = 10'h258 == _T_308[9:0] ? 4'h6 : _GEN_21542; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21544 = 10'h259 == _T_308[9:0] ? 4'h7 : _GEN_21543; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21545 = 10'h25a == _T_308[9:0] ? 4'h7 : _GEN_21544; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21546 = 10'h25b == _T_308[9:0] ? 4'h7 : _GEN_21545; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21547 = 10'h25c == _T_308[9:0] ? 4'h8 : _GEN_21546; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21548 = 10'h25d == _T_308[9:0] ? 4'h8 : _GEN_21547; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21549 = 10'h25e == _T_308[9:0] ? 4'h4 : _GEN_21548; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21550 = 10'h25f == _T_308[9:0] ? 4'h3 : _GEN_21549; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21551 = 10'h260 == _T_308[9:0] ? 4'h7 : _GEN_21550; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21552 = 10'h261 == _T_308[9:0] ? 4'h7 : _GEN_21551; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21553 = 10'h262 == _T_308[9:0] ? 4'h7 : _GEN_21552; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21554 = 10'h263 == _T_308[9:0] ? 4'h6 : _GEN_21553; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21555 = 10'h264 == _T_308[9:0] ? 4'h7 : _GEN_21554; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21556 = 10'h265 == _T_308[9:0] ? 4'h6 : _GEN_21555; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21557 = 10'h266 == _T_308[9:0] ? 4'h5 : _GEN_21556; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21558 = 10'h267 == _T_308[9:0] ? 4'h7 : _GEN_21557; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21559 = 10'h268 == _T_308[9:0] ? 4'ha : _GEN_21558; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21560 = 10'h269 == _T_308[9:0] ? 4'ha : _GEN_21559; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21561 = 10'h26a == _T_308[9:0] ? 4'ha : _GEN_21560; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21562 = 10'h26b == _T_308[9:0] ? 4'ha : _GEN_21561; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21563 = 10'h26c == _T_308[9:0] ? 4'ha : _GEN_21562; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21564 = 10'h26d == _T_308[9:0] ? 4'ha : _GEN_21563; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21565 = 10'h26e == _T_308[9:0] ? 4'ha : _GEN_21564; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21566 = 10'h26f == _T_308[9:0] ? 4'ha : _GEN_21565; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21567 = 10'h270 == _T_308[9:0] ? 4'h5 : _GEN_21566; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21568 = 10'h271 == _T_308[9:0] ? 4'h3 : _GEN_21567; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21569 = 10'h272 == _T_308[9:0] ? 4'h3 : _GEN_21568; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21570 = 10'h273 == _T_308[9:0] ? 4'h4 : _GEN_21569; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21571 = 10'h274 == _T_308[9:0] ? 4'h6 : _GEN_21570; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21572 = 10'h275 == _T_308[9:0] ? 4'h5 : _GEN_21571; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21573 = 10'h276 == _T_308[9:0] ? 4'h6 : _GEN_21572; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21574 = 10'h277 == _T_308[9:0] ? 4'h5 : _GEN_21573; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21575 = 10'h278 == _T_308[9:0] ? 4'h6 : _GEN_21574; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21576 = 10'h279 == _T_308[9:0] ? 4'h6 : _GEN_21575; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21577 = 10'h27a == _T_308[9:0] ? 4'h6 : _GEN_21576; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21578 = 10'h27b == _T_308[9:0] ? 4'h8 : _GEN_21577; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21579 = 10'h27c == _T_308[9:0] ? 4'h6 : _GEN_21578; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21580 = 10'h27d == _T_308[9:0] ? 4'h2 : _GEN_21579; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21581 = 10'h27e == _T_308[9:0] ? 4'h5 : _GEN_21580; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21582 = 10'h27f == _T_308[9:0] ? 4'h7 : _GEN_21581; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21583 = 10'h280 == _T_308[9:0] ? 4'h7 : _GEN_21582; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21584 = 10'h281 == _T_308[9:0] ? 4'h8 : _GEN_21583; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21585 = 10'h282 == _T_308[9:0] ? 4'h7 : _GEN_21584; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21586 = 10'h283 == _T_308[9:0] ? 4'h3 : _GEN_21585; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21587 = 10'h284 == _T_308[9:0] ? 4'h3 : _GEN_21586; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21588 = 10'h285 == _T_308[9:0] ? 4'h3 : _GEN_21587; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21589 = 10'h286 == _T_308[9:0] ? 4'h7 : _GEN_21588; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21590 = 10'h287 == _T_308[9:0] ? 4'h7 : _GEN_21589; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21591 = 10'h288 == _T_308[9:0] ? 4'h7 : _GEN_21590; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21592 = 10'h289 == _T_308[9:0] ? 4'h7 : _GEN_21591; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21593 = 10'h28a == _T_308[9:0] ? 4'h8 : _GEN_21592; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21594 = 10'h28b == _T_308[9:0] ? 4'h8 : _GEN_21593; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21595 = 10'h28c == _T_308[9:0] ? 4'h7 : _GEN_21594; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21596 = 10'h28d == _T_308[9:0] ? 4'h6 : _GEN_21595; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21597 = 10'h28e == _T_308[9:0] ? 4'h3 : _GEN_21596; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21598 = 10'h28f == _T_308[9:0] ? 4'h6 : _GEN_21597; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21599 = 10'h290 == _T_308[9:0] ? 4'h8 : _GEN_21598; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21600 = 10'h291 == _T_308[9:0] ? 4'ha : _GEN_21599; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21601 = 10'h292 == _T_308[9:0] ? 4'ha : _GEN_21600; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21602 = 10'h293 == _T_308[9:0] ? 4'ha : _GEN_21601; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21603 = 10'h294 == _T_308[9:0] ? 4'h9 : _GEN_21602; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21604 = 10'h295 == _T_308[9:0] ? 4'h4 : _GEN_21603; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21605 = 10'h296 == _T_308[9:0] ? 4'h3 : _GEN_21604; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21606 = 10'h297 == _T_308[9:0] ? 4'h3 : _GEN_21605; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21607 = 10'h298 == _T_308[9:0] ? 4'h3 : _GEN_21606; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21608 = 10'h299 == _T_308[9:0] ? 4'h4 : _GEN_21607; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21609 = 10'h29a == _T_308[9:0] ? 4'h5 : _GEN_21608; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21610 = 10'h29b == _T_308[9:0] ? 4'h5 : _GEN_21609; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21611 = 10'h29c == _T_308[9:0] ? 4'h5 : _GEN_21610; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21612 = 10'h29d == _T_308[9:0] ? 4'h5 : _GEN_21611; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21613 = 10'h29e == _T_308[9:0] ? 4'h5 : _GEN_21612; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21614 = 10'h29f == _T_308[9:0] ? 4'h5 : _GEN_21613; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21615 = 10'h2a0 == _T_308[9:0] ? 4'h6 : _GEN_21614; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21616 = 10'h2a1 == _T_308[9:0] ? 4'h7 : _GEN_21615; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21617 = 10'h2a2 == _T_308[9:0] ? 4'h5 : _GEN_21616; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21618 = 10'h2a3 == _T_308[9:0] ? 4'h2 : _GEN_21617; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21619 = 10'h2a4 == _T_308[9:0] ? 4'h3 : _GEN_21618; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21620 = 10'h2a5 == _T_308[9:0] ? 4'h7 : _GEN_21619; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21621 = 10'h2a6 == _T_308[9:0] ? 4'h8 : _GEN_21620; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21622 = 10'h2a7 == _T_308[9:0] ? 4'h7 : _GEN_21621; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21623 = 10'h2a8 == _T_308[9:0] ? 4'h3 : _GEN_21622; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21624 = 10'h2a9 == _T_308[9:0] ? 4'h2 : _GEN_21623; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21625 = 10'h2aa == _T_308[9:0] ? 4'h3 : _GEN_21624; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21626 = 10'h2ab == _T_308[9:0] ? 4'h3 : _GEN_21625; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21627 = 10'h2ac == _T_308[9:0] ? 4'h7 : _GEN_21626; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21628 = 10'h2ad == _T_308[9:0] ? 4'h8 : _GEN_21627; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21629 = 10'h2ae == _T_308[9:0] ? 4'h7 : _GEN_21628; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21630 = 10'h2af == _T_308[9:0] ? 4'h8 : _GEN_21629; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21631 = 10'h2b0 == _T_308[9:0] ? 4'h8 : _GEN_21630; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21632 = 10'h2b1 == _T_308[9:0] ? 4'h8 : _GEN_21631; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21633 = 10'h2b2 == _T_308[9:0] ? 4'h7 : _GEN_21632; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21634 = 10'h2b3 == _T_308[9:0] ? 4'h6 : _GEN_21633; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21635 = 10'h2b4 == _T_308[9:0] ? 4'h2 : _GEN_21634; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21636 = 10'h2b5 == _T_308[9:0] ? 4'h2 : _GEN_21635; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21637 = 10'h2b6 == _T_308[9:0] ? 4'h3 : _GEN_21636; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21638 = 10'h2b7 == _T_308[9:0] ? 4'h3 : _GEN_21637; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21639 = 10'h2b8 == _T_308[9:0] ? 4'h6 : _GEN_21638; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21640 = 10'h2b9 == _T_308[9:0] ? 4'h9 : _GEN_21639; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21641 = 10'h2ba == _T_308[9:0] ? 4'h3 : _GEN_21640; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21642 = 10'h2bb == _T_308[9:0] ? 4'h3 : _GEN_21641; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21643 = 10'h2bc == _T_308[9:0] ? 4'h3 : _GEN_21642; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21644 = 10'h2bd == _T_308[9:0] ? 4'h2 : _GEN_21643; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21645 = 10'h2be == _T_308[9:0] ? 4'h3 : _GEN_21644; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21646 = 10'h2bf == _T_308[9:0] ? 4'h3 : _GEN_21645; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21647 = 10'h2c0 == _T_308[9:0] ? 4'h5 : _GEN_21646; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21648 = 10'h2c1 == _T_308[9:0] ? 4'h5 : _GEN_21647; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21649 = 10'h2c2 == _T_308[9:0] ? 4'h5 : _GEN_21648; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21650 = 10'h2c3 == _T_308[9:0] ? 4'h5 : _GEN_21649; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21651 = 10'h2c4 == _T_308[9:0] ? 4'h5 : _GEN_21650; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21652 = 10'h2c5 == _T_308[9:0] ? 4'h5 : _GEN_21651; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21653 = 10'h2c6 == _T_308[9:0] ? 4'h6 : _GEN_21652; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21654 = 10'h2c7 == _T_308[9:0] ? 4'h7 : _GEN_21653; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21655 = 10'h2c8 == _T_308[9:0] ? 4'h5 : _GEN_21654; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21656 = 10'h2c9 == _T_308[9:0] ? 4'h2 : _GEN_21655; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21657 = 10'h2ca == _T_308[9:0] ? 4'h2 : _GEN_21656; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21658 = 10'h2cb == _T_308[9:0] ? 4'h3 : _GEN_21657; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21659 = 10'h2cc == _T_308[9:0] ? 4'h3 : _GEN_21658; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21660 = 10'h2cd == _T_308[9:0] ? 4'h2 : _GEN_21659; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21661 = 10'h2ce == _T_308[9:0] ? 4'h2 : _GEN_21660; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21662 = 10'h2cf == _T_308[9:0] ? 4'h2 : _GEN_21661; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21663 = 10'h2d0 == _T_308[9:0] ? 4'h2 : _GEN_21662; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21664 = 10'h2d1 == _T_308[9:0] ? 4'h2 : _GEN_21663; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21665 = 10'h2d2 == _T_308[9:0] ? 4'h7 : _GEN_21664; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21666 = 10'h2d3 == _T_308[9:0] ? 4'h7 : _GEN_21665; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21667 = 10'h2d4 == _T_308[9:0] ? 4'h8 : _GEN_21666; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21668 = 10'h2d5 == _T_308[9:0] ? 4'h8 : _GEN_21667; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21669 = 10'h2d6 == _T_308[9:0] ? 4'h8 : _GEN_21668; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21670 = 10'h2d7 == _T_308[9:0] ? 4'h8 : _GEN_21669; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21671 = 10'h2d8 == _T_308[9:0] ? 4'h7 : _GEN_21670; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21672 = 10'h2d9 == _T_308[9:0] ? 4'h6 : _GEN_21671; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21673 = 10'h2da == _T_308[9:0] ? 4'h4 : _GEN_21672; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21674 = 10'h2db == _T_308[9:0] ? 4'h2 : _GEN_21673; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21675 = 10'h2dc == _T_308[9:0] ? 4'h2 : _GEN_21674; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21676 = 10'h2dd == _T_308[9:0] ? 4'h3 : _GEN_21675; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21677 = 10'h2de == _T_308[9:0] ? 4'h3 : _GEN_21676; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21678 = 10'h2df == _T_308[9:0] ? 4'h3 : _GEN_21677; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21679 = 10'h2e0 == _T_308[9:0] ? 4'h3 : _GEN_21678; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21680 = 10'h2e1 == _T_308[9:0] ? 4'h3 : _GEN_21679; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21681 = 10'h2e2 == _T_308[9:0] ? 4'h3 : _GEN_21680; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21682 = 10'h2e3 == _T_308[9:0] ? 4'h2 : _GEN_21681; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21683 = 10'h2e4 == _T_308[9:0] ? 4'h3 : _GEN_21682; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21684 = 10'h2e5 == _T_308[9:0] ? 4'h2 : _GEN_21683; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21685 = 10'h2e6 == _T_308[9:0] ? 4'h5 : _GEN_21684; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21686 = 10'h2e7 == _T_308[9:0] ? 4'h5 : _GEN_21685; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21687 = 10'h2e8 == _T_308[9:0] ? 4'h5 : _GEN_21686; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21688 = 10'h2e9 == _T_308[9:0] ? 4'h5 : _GEN_21687; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21689 = 10'h2ea == _T_308[9:0] ? 4'h5 : _GEN_21688; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21690 = 10'h2eb == _T_308[9:0] ? 4'h5 : _GEN_21689; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21691 = 10'h2ec == _T_308[9:0] ? 4'h6 : _GEN_21690; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21692 = 10'h2ed == _T_308[9:0] ? 4'h7 : _GEN_21691; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21693 = 10'h2ee == _T_308[9:0] ? 4'h6 : _GEN_21692; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21694 = 10'h2ef == _T_308[9:0] ? 4'h2 : _GEN_21693; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21695 = 10'h2f0 == _T_308[9:0] ? 4'h2 : _GEN_21694; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21696 = 10'h2f1 == _T_308[9:0] ? 4'h2 : _GEN_21695; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21697 = 10'h2f2 == _T_308[9:0] ? 4'h2 : _GEN_21696; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21698 = 10'h2f3 == _T_308[9:0] ? 4'h2 : _GEN_21697; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21699 = 10'h2f4 == _T_308[9:0] ? 4'h2 : _GEN_21698; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21700 = 10'h2f5 == _T_308[9:0] ? 4'h2 : _GEN_21699; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21701 = 10'h2f6 == _T_308[9:0] ? 4'h2 : _GEN_21700; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21702 = 10'h2f7 == _T_308[9:0] ? 4'h2 : _GEN_21701; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21703 = 10'h2f8 == _T_308[9:0] ? 4'h7 : _GEN_21702; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21704 = 10'h2f9 == _T_308[9:0] ? 4'h7 : _GEN_21703; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21705 = 10'h2fa == _T_308[9:0] ? 4'h8 : _GEN_21704; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21706 = 10'h2fb == _T_308[9:0] ? 4'h8 : _GEN_21705; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21707 = 10'h2fc == _T_308[9:0] ? 4'h7 : _GEN_21706; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21708 = 10'h2fd == _T_308[9:0] ? 4'h7 : _GEN_21707; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21709 = 10'h2fe == _T_308[9:0] ? 4'h7 : _GEN_21708; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21710 = 10'h2ff == _T_308[9:0] ? 4'h7 : _GEN_21709; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21711 = 10'h300 == _T_308[9:0] ? 4'h8 : _GEN_21710; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21712 = 10'h301 == _T_308[9:0] ? 4'h7 : _GEN_21711; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21713 = 10'h302 == _T_308[9:0] ? 4'h3 : _GEN_21712; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21714 = 10'h303 == _T_308[9:0] ? 4'h3 : _GEN_21713; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21715 = 10'h304 == _T_308[9:0] ? 4'h2 : _GEN_21714; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21716 = 10'h305 == _T_308[9:0] ? 4'h2 : _GEN_21715; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21717 = 10'h306 == _T_308[9:0] ? 4'h2 : _GEN_21716; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21718 = 10'h307 == _T_308[9:0] ? 4'h2 : _GEN_21717; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21719 = 10'h308 == _T_308[9:0] ? 4'h2 : _GEN_21718; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21720 = 10'h309 == _T_308[9:0] ? 4'h2 : _GEN_21719; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21721 = 10'h30a == _T_308[9:0] ? 4'h2 : _GEN_21720; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21722 = 10'h30b == _T_308[9:0] ? 4'h3 : _GEN_21721; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21723 = 10'h30c == _T_308[9:0] ? 4'h4 : _GEN_21722; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21724 = 10'h30d == _T_308[9:0] ? 4'h5 : _GEN_21723; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21725 = 10'h30e == _T_308[9:0] ? 4'h5 : _GEN_21724; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21726 = 10'h30f == _T_308[9:0] ? 4'h5 : _GEN_21725; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21727 = 10'h310 == _T_308[9:0] ? 4'h5 : _GEN_21726; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21728 = 10'h311 == _T_308[9:0] ? 4'h5 : _GEN_21727; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21729 = 10'h312 == _T_308[9:0] ? 4'h6 : _GEN_21728; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21730 = 10'h313 == _T_308[9:0] ? 4'h7 : _GEN_21729; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21731 = 10'h314 == _T_308[9:0] ? 4'h7 : _GEN_21730; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21732 = 10'h315 == _T_308[9:0] ? 4'h3 : _GEN_21731; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21733 = 10'h316 == _T_308[9:0] ? 4'h2 : _GEN_21732; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21734 = 10'h317 == _T_308[9:0] ? 4'h2 : _GEN_21733; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21735 = 10'h318 == _T_308[9:0] ? 4'h2 : _GEN_21734; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21736 = 10'h319 == _T_308[9:0] ? 4'h2 : _GEN_21735; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21737 = 10'h31a == _T_308[9:0] ? 4'h2 : _GEN_21736; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21738 = 10'h31b == _T_308[9:0] ? 4'h2 : _GEN_21737; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21739 = 10'h31c == _T_308[9:0] ? 4'h2 : _GEN_21738; // @[Filter.scala 230:142]
  wire [3:0] _GEN_21740 = 10'h31d == _T_308[9:0] ? 4'h2 : _GEN_21739; // @[Filter.scala 230:142]
  wire [7:0] _T_322 = _GEN_21740 * 4'ha; // @[Filter.scala 230:142]
  wire [10:0] _GEN_39007 = {{3'd0}, _T_322}; // @[Filter.scala 230:109]
  wire [10:0] _T_324 = _T_317 + _GEN_39007; // @[Filter.scala 230:109]
  wire [10:0] _T_325 = _T_324 / 11'h64; // @[Filter.scala 230:150]
  wire  _T_327 = _T_298 >= 6'h20; // @[Filter.scala 233:31]
  wire  _T_331 = _T_305 >= 32'h12; // @[Filter.scala 233:63]
  wire  _T_332 = _T_327 | _T_331; // @[Filter.scala 233:58]
  wire [10:0] _GEN_22539 = io_SPI_distort ? _T_325 : {{7'd0}, _GEN_20144}; // @[Filter.scala 235:35]
  wire [10:0] _GEN_22540 = _T_332 ? 11'h0 : _GEN_22539; // @[Filter.scala 233:80]
  wire [10:0] _GEN_23339 = io_SPI_distort ? _T_325 : {{7'd0}, _GEN_20942}; // @[Filter.scala 235:35]
  wire [10:0] _GEN_23340 = _T_332 ? 11'h0 : _GEN_23339; // @[Filter.scala 233:80]
  wire [10:0] _GEN_24139 = io_SPI_distort ? _T_325 : {{7'd0}, _GEN_21740}; // @[Filter.scala 235:35]
  wire [10:0] _GEN_24140 = _T_332 ? 11'h0 : _GEN_24139; // @[Filter.scala 233:80]
  wire [31:0] _T_360 = pixelIndex + 32'h5; // @[Filter.scala 228:31]
  wire [31:0] _GEN_5 = _T_360 % 32'h20; // @[Filter.scala 228:38]
  wire [5:0] _T_361 = _GEN_5[5:0]; // @[Filter.scala 228:38]
  wire [5:0] _T_363 = _T_361 + _GEN_38951; // @[Filter.scala 228:53]
  wire [5:0] _T_365 = _T_363 - 6'h1; // @[Filter.scala 228:69]
  wire [31:0] _T_368 = _T_360 / 32'h20; // @[Filter.scala 229:38]
  wire [31:0] _T_370 = _T_368 + _GEN_38952; // @[Filter.scala 229:53]
  wire [31:0] _T_372 = _T_370 - 32'h1; // @[Filter.scala 229:69]
  wire [37:0] _T_373 = _T_372 * 32'h20; // @[Filter.scala 230:42]
  wire [37:0] _GEN_39013 = {{32'd0}, _T_365}; // @[Filter.scala 230:57]
  wire [37:0] _T_375 = _T_373 + _GEN_39013; // @[Filter.scala 230:57]
  wire [3:0] _GEN_24163 = 10'h16 == _T_375[9:0] ? 4'h9 : 4'ha; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24164 = 10'h17 == _T_375[9:0] ? 4'h3 : _GEN_24163; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24165 = 10'h18 == _T_375[9:0] ? 4'h6 : _GEN_24164; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24166 = 10'h19 == _T_375[9:0] ? 4'ha : _GEN_24165; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24167 = 10'h1a == _T_375[9:0] ? 4'ha : _GEN_24166; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24168 = 10'h1b == _T_375[9:0] ? 4'ha : _GEN_24167; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24169 = 10'h1c == _T_375[9:0] ? 4'ha : _GEN_24168; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24170 = 10'h1d == _T_375[9:0] ? 4'ha : _GEN_24169; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24171 = 10'h1e == _T_375[9:0] ? 4'ha : _GEN_24170; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24172 = 10'h1f == _T_375[9:0] ? 4'ha : _GEN_24171; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24173 = 10'h20 == _T_375[9:0] ? 4'ha : _GEN_24172; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24174 = 10'h21 == _T_375[9:0] ? 4'ha : _GEN_24173; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24175 = 10'h22 == _T_375[9:0] ? 4'ha : _GEN_24174; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24176 = 10'h23 == _T_375[9:0] ? 4'ha : _GEN_24175; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24177 = 10'h24 == _T_375[9:0] ? 4'ha : _GEN_24176; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24178 = 10'h25 == _T_375[9:0] ? 4'ha : _GEN_24177; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24179 = 10'h26 == _T_375[9:0] ? 4'ha : _GEN_24178; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24180 = 10'h27 == _T_375[9:0] ? 4'ha : _GEN_24179; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24181 = 10'h28 == _T_375[9:0] ? 4'ha : _GEN_24180; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24182 = 10'h29 == _T_375[9:0] ? 4'ha : _GEN_24181; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24183 = 10'h2a == _T_375[9:0] ? 4'ha : _GEN_24182; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24184 = 10'h2b == _T_375[9:0] ? 4'ha : _GEN_24183; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24185 = 10'h2c == _T_375[9:0] ? 4'ha : _GEN_24184; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24186 = 10'h2d == _T_375[9:0] ? 4'ha : _GEN_24185; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24187 = 10'h2e == _T_375[9:0] ? 4'ha : _GEN_24186; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24188 = 10'h2f == _T_375[9:0] ? 4'ha : _GEN_24187; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24189 = 10'h30 == _T_375[9:0] ? 4'ha : _GEN_24188; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24190 = 10'h31 == _T_375[9:0] ? 4'ha : _GEN_24189; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24191 = 10'h32 == _T_375[9:0] ? 4'ha : _GEN_24190; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24192 = 10'h33 == _T_375[9:0] ? 4'ha : _GEN_24191; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24193 = 10'h34 == _T_375[9:0] ? 4'ha : _GEN_24192; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24194 = 10'h35 == _T_375[9:0] ? 4'ha : _GEN_24193; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24195 = 10'h36 == _T_375[9:0] ? 4'ha : _GEN_24194; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24196 = 10'h37 == _T_375[9:0] ? 4'ha : _GEN_24195; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24197 = 10'h38 == _T_375[9:0] ? 4'ha : _GEN_24196; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24198 = 10'h39 == _T_375[9:0] ? 4'ha : _GEN_24197; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24199 = 10'h3a == _T_375[9:0] ? 4'ha : _GEN_24198; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24200 = 10'h3b == _T_375[9:0] ? 4'h9 : _GEN_24199; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24201 = 10'h3c == _T_375[9:0] ? 4'h4 : _GEN_24200; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24202 = 10'h3d == _T_375[9:0] ? 4'h3 : _GEN_24201; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24203 = 10'h3e == _T_375[9:0] ? 4'h4 : _GEN_24202; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24204 = 10'h3f == _T_375[9:0] ? 4'ha : _GEN_24203; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24205 = 10'h40 == _T_375[9:0] ? 4'ha : _GEN_24204; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24206 = 10'h41 == _T_375[9:0] ? 4'ha : _GEN_24205; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24207 = 10'h42 == _T_375[9:0] ? 4'ha : _GEN_24206; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24208 = 10'h43 == _T_375[9:0] ? 4'ha : _GEN_24207; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24209 = 10'h44 == _T_375[9:0] ? 4'ha : _GEN_24208; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24210 = 10'h45 == _T_375[9:0] ? 4'ha : _GEN_24209; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24211 = 10'h46 == _T_375[9:0] ? 4'ha : _GEN_24210; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24212 = 10'h47 == _T_375[9:0] ? 4'ha : _GEN_24211; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24213 = 10'h48 == _T_375[9:0] ? 4'ha : _GEN_24212; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24214 = 10'h49 == _T_375[9:0] ? 4'ha : _GEN_24213; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24215 = 10'h4a == _T_375[9:0] ? 4'ha : _GEN_24214; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24216 = 10'h4b == _T_375[9:0] ? 4'ha : _GEN_24215; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24217 = 10'h4c == _T_375[9:0] ? 4'ha : _GEN_24216; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24218 = 10'h4d == _T_375[9:0] ? 4'ha : _GEN_24217; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24219 = 10'h4e == _T_375[9:0] ? 4'ha : _GEN_24218; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24220 = 10'h4f == _T_375[9:0] ? 4'ha : _GEN_24219; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24221 = 10'h50 == _T_375[9:0] ? 4'ha : _GEN_24220; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24222 = 10'h51 == _T_375[9:0] ? 4'ha : _GEN_24221; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24223 = 10'h52 == _T_375[9:0] ? 4'ha : _GEN_24222; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24224 = 10'h53 == _T_375[9:0] ? 4'ha : _GEN_24223; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24225 = 10'h54 == _T_375[9:0] ? 4'ha : _GEN_24224; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24226 = 10'h55 == _T_375[9:0] ? 4'ha : _GEN_24225; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24227 = 10'h56 == _T_375[9:0] ? 4'ha : _GEN_24226; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24228 = 10'h57 == _T_375[9:0] ? 4'ha : _GEN_24227; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24229 = 10'h58 == _T_375[9:0] ? 4'ha : _GEN_24228; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24230 = 10'h59 == _T_375[9:0] ? 4'ha : _GEN_24229; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24231 = 10'h5a == _T_375[9:0] ? 4'h7 : _GEN_24230; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24232 = 10'h5b == _T_375[9:0] ? 4'h7 : _GEN_24231; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24233 = 10'h5c == _T_375[9:0] ? 4'ha : _GEN_24232; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24234 = 10'h5d == _T_375[9:0] ? 4'ha : _GEN_24233; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24235 = 10'h5e == _T_375[9:0] ? 4'ha : _GEN_24234; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24236 = 10'h5f == _T_375[9:0] ? 4'ha : _GEN_24235; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24237 = 10'h60 == _T_375[9:0] ? 4'ha : _GEN_24236; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24238 = 10'h61 == _T_375[9:0] ? 4'h8 : _GEN_24237; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24239 = 10'h62 == _T_375[9:0] ? 4'h3 : _GEN_24238; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24240 = 10'h63 == _T_375[9:0] ? 4'h3 : _GEN_24239; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24241 = 10'h64 == _T_375[9:0] ? 4'h3 : _GEN_24240; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24242 = 10'h65 == _T_375[9:0] ? 4'h9 : _GEN_24241; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24243 = 10'h66 == _T_375[9:0] ? 4'ha : _GEN_24242; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24244 = 10'h67 == _T_375[9:0] ? 4'ha : _GEN_24243; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24245 = 10'h68 == _T_375[9:0] ? 4'ha : _GEN_24244; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24246 = 10'h69 == _T_375[9:0] ? 4'ha : _GEN_24245; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24247 = 10'h6a == _T_375[9:0] ? 4'ha : _GEN_24246; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24248 = 10'h6b == _T_375[9:0] ? 4'h8 : _GEN_24247; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24249 = 10'h6c == _T_375[9:0] ? 4'h5 : _GEN_24248; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24250 = 10'h6d == _T_375[9:0] ? 4'h8 : _GEN_24249; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24251 = 10'h6e == _T_375[9:0] ? 4'ha : _GEN_24250; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24252 = 10'h6f == _T_375[9:0] ? 4'ha : _GEN_24251; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24253 = 10'h70 == _T_375[9:0] ? 4'ha : _GEN_24252; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24254 = 10'h71 == _T_375[9:0] ? 4'ha : _GEN_24253; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24255 = 10'h72 == _T_375[9:0] ? 4'ha : _GEN_24254; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24256 = 10'h73 == _T_375[9:0] ? 4'ha : _GEN_24255; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24257 = 10'h74 == _T_375[9:0] ? 4'ha : _GEN_24256; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24258 = 10'h75 == _T_375[9:0] ? 4'ha : _GEN_24257; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24259 = 10'h76 == _T_375[9:0] ? 4'ha : _GEN_24258; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24260 = 10'h77 == _T_375[9:0] ? 4'ha : _GEN_24259; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24261 = 10'h78 == _T_375[9:0] ? 4'ha : _GEN_24260; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24262 = 10'h79 == _T_375[9:0] ? 4'ha : _GEN_24261; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24263 = 10'h7a == _T_375[9:0] ? 4'ha : _GEN_24262; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24264 = 10'h7b == _T_375[9:0] ? 4'ha : _GEN_24263; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24265 = 10'h7c == _T_375[9:0] ? 4'ha : _GEN_24264; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24266 = 10'h7d == _T_375[9:0] ? 4'ha : _GEN_24265; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24267 = 10'h7e == _T_375[9:0] ? 4'ha : _GEN_24266; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24268 = 10'h7f == _T_375[9:0] ? 4'ha : _GEN_24267; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24269 = 10'h80 == _T_375[9:0] ? 4'ha : _GEN_24268; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24270 = 10'h81 == _T_375[9:0] ? 4'h5 : _GEN_24269; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24271 = 10'h82 == _T_375[9:0] ? 4'h5 : _GEN_24270; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24272 = 10'h83 == _T_375[9:0] ? 4'h7 : _GEN_24271; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24273 = 10'h84 == _T_375[9:0] ? 4'ha : _GEN_24272; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24274 = 10'h85 == _T_375[9:0] ? 4'ha : _GEN_24273; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24275 = 10'h86 == _T_375[9:0] ? 4'ha : _GEN_24274; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24276 = 10'h87 == _T_375[9:0] ? 4'h5 : _GEN_24275; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24277 = 10'h88 == _T_375[9:0] ? 4'h3 : _GEN_24276; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24278 = 10'h89 == _T_375[9:0] ? 4'h3 : _GEN_24277; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24279 = 10'h8a == _T_375[9:0] ? 4'h4 : _GEN_24278; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24280 = 10'h8b == _T_375[9:0] ? 4'h9 : _GEN_24279; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24281 = 10'h8c == _T_375[9:0] ? 4'ha : _GEN_24280; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24282 = 10'h8d == _T_375[9:0] ? 4'ha : _GEN_24281; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24283 = 10'h8e == _T_375[9:0] ? 4'ha : _GEN_24282; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24284 = 10'h8f == _T_375[9:0] ? 4'h6 : _GEN_24283; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24285 = 10'h90 == _T_375[9:0] ? 4'h4 : _GEN_24284; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24286 = 10'h91 == _T_375[9:0] ? 4'h3 : _GEN_24285; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24287 = 10'h92 == _T_375[9:0] ? 4'h7 : _GEN_24286; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24288 = 10'h93 == _T_375[9:0] ? 4'ha : _GEN_24287; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24289 = 10'h94 == _T_375[9:0] ? 4'ha : _GEN_24288; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24290 = 10'h95 == _T_375[9:0] ? 4'ha : _GEN_24289; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24291 = 10'h96 == _T_375[9:0] ? 4'ha : _GEN_24290; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24292 = 10'h97 == _T_375[9:0] ? 4'ha : _GEN_24291; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24293 = 10'h98 == _T_375[9:0] ? 4'ha : _GEN_24292; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24294 = 10'h99 == _T_375[9:0] ? 4'ha : _GEN_24293; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24295 = 10'h9a == _T_375[9:0] ? 4'ha : _GEN_24294; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24296 = 10'h9b == _T_375[9:0] ? 4'ha : _GEN_24295; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24297 = 10'h9c == _T_375[9:0] ? 4'ha : _GEN_24296; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24298 = 10'h9d == _T_375[9:0] ? 4'ha : _GEN_24297; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24299 = 10'h9e == _T_375[9:0] ? 4'ha : _GEN_24298; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24300 = 10'h9f == _T_375[9:0] ? 4'ha : _GEN_24299; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24301 = 10'ha0 == _T_375[9:0] ? 4'ha : _GEN_24300; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24302 = 10'ha1 == _T_375[9:0] ? 4'ha : _GEN_24301; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24303 = 10'ha2 == _T_375[9:0] ? 4'ha : _GEN_24302; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24304 = 10'ha3 == _T_375[9:0] ? 4'ha : _GEN_24303; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24305 = 10'ha4 == _T_375[9:0] ? 4'ha : _GEN_24304; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24306 = 10'ha5 == _T_375[9:0] ? 4'ha : _GEN_24305; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24307 = 10'ha6 == _T_375[9:0] ? 4'ha : _GEN_24306; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24308 = 10'ha7 == _T_375[9:0] ? 4'h9 : _GEN_24307; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24309 = 10'ha8 == _T_375[9:0] ? 4'h4 : _GEN_24308; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24310 = 10'ha9 == _T_375[9:0] ? 4'h3 : _GEN_24309; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24311 = 10'haa == _T_375[9:0] ? 4'h4 : _GEN_24310; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24312 = 10'hab == _T_375[9:0] ? 4'h7 : _GEN_24311; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24313 = 10'hac == _T_375[9:0] ? 4'h8 : _GEN_24312; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24314 = 10'had == _T_375[9:0] ? 4'h3 : _GEN_24313; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24315 = 10'hae == _T_375[9:0] ? 4'h3 : _GEN_24314; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24316 = 10'haf == _T_375[9:0] ? 4'h3 : _GEN_24315; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24317 = 10'hb0 == _T_375[9:0] ? 4'h3 : _GEN_24316; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24318 = 10'hb1 == _T_375[9:0] ? 4'h7 : _GEN_24317; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24319 = 10'hb2 == _T_375[9:0] ? 4'h9 : _GEN_24318; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24320 = 10'hb3 == _T_375[9:0] ? 4'h6 : _GEN_24319; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24321 = 10'hb4 == _T_375[9:0] ? 4'h4 : _GEN_24320; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24322 = 10'hb5 == _T_375[9:0] ? 4'h3 : _GEN_24321; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24323 = 10'hb6 == _T_375[9:0] ? 4'h3 : _GEN_24322; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24324 = 10'hb7 == _T_375[9:0] ? 4'h6 : _GEN_24323; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24325 = 10'hb8 == _T_375[9:0] ? 4'ha : _GEN_24324; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24326 = 10'hb9 == _T_375[9:0] ? 4'ha : _GEN_24325; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24327 = 10'hba == _T_375[9:0] ? 4'ha : _GEN_24326; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24328 = 10'hbb == _T_375[9:0] ? 4'ha : _GEN_24327; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24329 = 10'hbc == _T_375[9:0] ? 4'ha : _GEN_24328; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24330 = 10'hbd == _T_375[9:0] ? 4'h9 : _GEN_24329; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24331 = 10'hbe == _T_375[9:0] ? 4'ha : _GEN_24330; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24332 = 10'hbf == _T_375[9:0] ? 4'ha : _GEN_24331; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24333 = 10'hc0 == _T_375[9:0] ? 4'ha : _GEN_24332; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24334 = 10'hc1 == _T_375[9:0] ? 4'ha : _GEN_24333; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24335 = 10'hc2 == _T_375[9:0] ? 4'ha : _GEN_24334; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24336 = 10'hc3 == _T_375[9:0] ? 4'ha : _GEN_24335; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24337 = 10'hc4 == _T_375[9:0] ? 4'ha : _GEN_24336; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24338 = 10'hc5 == _T_375[9:0] ? 4'ha : _GEN_24337; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24339 = 10'hc6 == _T_375[9:0] ? 4'ha : _GEN_24338; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24340 = 10'hc7 == _T_375[9:0] ? 4'h9 : _GEN_24339; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24341 = 10'hc8 == _T_375[9:0] ? 4'h8 : _GEN_24340; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24342 = 10'hc9 == _T_375[9:0] ? 4'h8 : _GEN_24341; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24343 = 10'hca == _T_375[9:0] ? 4'h9 : _GEN_24342; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24344 = 10'hcb == _T_375[9:0] ? 4'ha : _GEN_24343; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24345 = 10'hcc == _T_375[9:0] ? 4'ha : _GEN_24344; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24346 = 10'hcd == _T_375[9:0] ? 4'ha : _GEN_24345; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24347 = 10'hce == _T_375[9:0] ? 4'h8 : _GEN_24346; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24348 = 10'hcf == _T_375[9:0] ? 4'h3 : _GEN_24347; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24349 = 10'hd0 == _T_375[9:0] ? 4'h3 : _GEN_24348; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24350 = 10'hd1 == _T_375[9:0] ? 4'h3 : _GEN_24349; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24351 = 10'hd2 == _T_375[9:0] ? 4'h4 : _GEN_24350; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24352 = 10'hd3 == _T_375[9:0] ? 4'h3 : _GEN_24351; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24353 = 10'hd4 == _T_375[9:0] ? 4'h3 : _GEN_24352; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24354 = 10'hd5 == _T_375[9:0] ? 4'h3 : _GEN_24353; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24355 = 10'hd6 == _T_375[9:0] ? 4'h3 : _GEN_24354; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24356 = 10'hd7 == _T_375[9:0] ? 4'h5 : _GEN_24355; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24357 = 10'hd8 == _T_375[9:0] ? 4'h4 : _GEN_24356; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24358 = 10'hd9 == _T_375[9:0] ? 4'h3 : _GEN_24357; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24359 = 10'hda == _T_375[9:0] ? 4'h3 : _GEN_24358; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24360 = 10'hdb == _T_375[9:0] ? 4'h3 : _GEN_24359; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24361 = 10'hdc == _T_375[9:0] ? 4'h4 : _GEN_24360; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24362 = 10'hdd == _T_375[9:0] ? 4'ha : _GEN_24361; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24363 = 10'hde == _T_375[9:0] ? 4'ha : _GEN_24362; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24364 = 10'hdf == _T_375[9:0] ? 4'ha : _GEN_24363; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24365 = 10'he0 == _T_375[9:0] ? 4'ha : _GEN_24364; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24366 = 10'he1 == _T_375[9:0] ? 4'ha : _GEN_24365; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24367 = 10'he2 == _T_375[9:0] ? 4'ha : _GEN_24366; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24368 = 10'he3 == _T_375[9:0] ? 4'h5 : _GEN_24367; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24369 = 10'he4 == _T_375[9:0] ? 4'ha : _GEN_24368; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24370 = 10'he5 == _T_375[9:0] ? 4'ha : _GEN_24369; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24371 = 10'he6 == _T_375[9:0] ? 4'ha : _GEN_24370; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24372 = 10'he7 == _T_375[9:0] ? 4'ha : _GEN_24371; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24373 = 10'he8 == _T_375[9:0] ? 4'ha : _GEN_24372; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24374 = 10'he9 == _T_375[9:0] ? 4'ha : _GEN_24373; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24375 = 10'hea == _T_375[9:0] ? 4'ha : _GEN_24374; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24376 = 10'heb == _T_375[9:0] ? 4'h9 : _GEN_24375; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24377 = 10'hec == _T_375[9:0] ? 4'h7 : _GEN_24376; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24378 = 10'hed == _T_375[9:0] ? 4'h3 : _GEN_24377; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24379 = 10'hee == _T_375[9:0] ? 4'h3 : _GEN_24378; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24380 = 10'hef == _T_375[9:0] ? 4'h3 : _GEN_24379; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24381 = 10'hf0 == _T_375[9:0] ? 4'h4 : _GEN_24380; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24382 = 10'hf1 == _T_375[9:0] ? 4'h7 : _GEN_24381; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24383 = 10'hf2 == _T_375[9:0] ? 4'ha : _GEN_24382; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24384 = 10'hf3 == _T_375[9:0] ? 4'ha : _GEN_24383; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24385 = 10'hf4 == _T_375[9:0] ? 4'ha : _GEN_24384; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24386 = 10'hf5 == _T_375[9:0] ? 4'h7 : _GEN_24385; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24387 = 10'hf6 == _T_375[9:0] ? 4'h3 : _GEN_24386; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24388 = 10'hf7 == _T_375[9:0] ? 4'h3 : _GEN_24387; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24389 = 10'hf8 == _T_375[9:0] ? 4'h3 : _GEN_24388; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24390 = 10'hf9 == _T_375[9:0] ? 4'h3 : _GEN_24389; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24391 = 10'hfa == _T_375[9:0] ? 4'h3 : _GEN_24390; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24392 = 10'hfb == _T_375[9:0] ? 4'h3 : _GEN_24391; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24393 = 10'hfc == _T_375[9:0] ? 4'h3 : _GEN_24392; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24394 = 10'hfd == _T_375[9:0] ? 4'h3 : _GEN_24393; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24395 = 10'hfe == _T_375[9:0] ? 4'h3 : _GEN_24394; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24396 = 10'hff == _T_375[9:0] ? 4'h3 : _GEN_24395; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24397 = 10'h100 == _T_375[9:0] ? 4'h3 : _GEN_24396; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24398 = 10'h101 == _T_375[9:0] ? 4'h4 : _GEN_24397; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24399 = 10'h102 == _T_375[9:0] ? 4'h6 : _GEN_24398; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24400 = 10'h103 == _T_375[9:0] ? 4'ha : _GEN_24399; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24401 = 10'h104 == _T_375[9:0] ? 4'ha : _GEN_24400; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24402 = 10'h105 == _T_375[9:0] ? 4'h9 : _GEN_24401; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24403 = 10'h106 == _T_375[9:0] ? 4'h9 : _GEN_24402; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24404 = 10'h107 == _T_375[9:0] ? 4'h9 : _GEN_24403; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24405 = 10'h108 == _T_375[9:0] ? 4'h9 : _GEN_24404; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24406 = 10'h109 == _T_375[9:0] ? 4'h3 : _GEN_24405; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24407 = 10'h10a == _T_375[9:0] ? 4'ha : _GEN_24406; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24408 = 10'h10b == _T_375[9:0] ? 4'ha : _GEN_24407; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24409 = 10'h10c == _T_375[9:0] ? 4'ha : _GEN_24408; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24410 = 10'h10d == _T_375[9:0] ? 4'ha : _GEN_24409; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24411 = 10'h10e == _T_375[9:0] ? 4'ha : _GEN_24410; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24412 = 10'h10f == _T_375[9:0] ? 4'h9 : _GEN_24411; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24413 = 10'h110 == _T_375[9:0] ? 4'h9 : _GEN_24412; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24414 = 10'h111 == _T_375[9:0] ? 4'h4 : _GEN_24413; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24415 = 10'h112 == _T_375[9:0] ? 4'h8 : _GEN_24414; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24416 = 10'h113 == _T_375[9:0] ? 4'h3 : _GEN_24415; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24417 = 10'h114 == _T_375[9:0] ? 4'h3 : _GEN_24416; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24418 = 10'h115 == _T_375[9:0] ? 4'h4 : _GEN_24417; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24419 = 10'h116 == _T_375[9:0] ? 4'h4 : _GEN_24418; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24420 = 10'h117 == _T_375[9:0] ? 4'h3 : _GEN_24419; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24421 = 10'h118 == _T_375[9:0] ? 4'h8 : _GEN_24420; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24422 = 10'h119 == _T_375[9:0] ? 4'ha : _GEN_24421; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24423 = 10'h11a == _T_375[9:0] ? 4'ha : _GEN_24422; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24424 = 10'h11b == _T_375[9:0] ? 4'ha : _GEN_24423; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24425 = 10'h11c == _T_375[9:0] ? 4'h6 : _GEN_24424; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24426 = 10'h11d == _T_375[9:0] ? 4'h3 : _GEN_24425; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24427 = 10'h11e == _T_375[9:0] ? 4'h3 : _GEN_24426; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24428 = 10'h11f == _T_375[9:0] ? 4'h3 : _GEN_24427; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24429 = 10'h120 == _T_375[9:0] ? 4'h3 : _GEN_24428; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24430 = 10'h121 == _T_375[9:0] ? 4'h3 : _GEN_24429; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24431 = 10'h122 == _T_375[9:0] ? 4'h3 : _GEN_24430; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24432 = 10'h123 == _T_375[9:0] ? 4'h3 : _GEN_24431; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24433 = 10'h124 == _T_375[9:0] ? 4'h3 : _GEN_24432; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24434 = 10'h125 == _T_375[9:0] ? 4'h3 : _GEN_24433; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24435 = 10'h126 == _T_375[9:0] ? 4'h4 : _GEN_24434; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24436 = 10'h127 == _T_375[9:0] ? 4'h6 : _GEN_24435; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24437 = 10'h128 == _T_375[9:0] ? 4'h5 : _GEN_24436; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24438 = 10'h129 == _T_375[9:0] ? 4'h8 : _GEN_24437; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24439 = 10'h12a == _T_375[9:0] ? 4'h5 : _GEN_24438; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24440 = 10'h12b == _T_375[9:0] ? 4'h3 : _GEN_24439; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24441 = 10'h12c == _T_375[9:0] ? 4'h3 : _GEN_24440; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24442 = 10'h12d == _T_375[9:0] ? 4'h3 : _GEN_24441; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24443 = 10'h12e == _T_375[9:0] ? 4'h4 : _GEN_24442; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24444 = 10'h12f == _T_375[9:0] ? 4'h4 : _GEN_24443; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24445 = 10'h130 == _T_375[9:0] ? 4'ha : _GEN_24444; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24446 = 10'h131 == _T_375[9:0] ? 4'h9 : _GEN_24445; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24447 = 10'h132 == _T_375[9:0] ? 4'h9 : _GEN_24446; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24448 = 10'h133 == _T_375[9:0] ? 4'h8 : _GEN_24447; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24449 = 10'h134 == _T_375[9:0] ? 4'h9 : _GEN_24448; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24450 = 10'h135 == _T_375[9:0] ? 4'h8 : _GEN_24449; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24451 = 10'h136 == _T_375[9:0] ? 4'h7 : _GEN_24450; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24452 = 10'h137 == _T_375[9:0] ? 4'h6 : _GEN_24451; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24453 = 10'h138 == _T_375[9:0] ? 4'h8 : _GEN_24452; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24454 = 10'h139 == _T_375[9:0] ? 4'h3 : _GEN_24453; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24455 = 10'h13a == _T_375[9:0] ? 4'h3 : _GEN_24454; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24456 = 10'h13b == _T_375[9:0] ? 4'h4 : _GEN_24455; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24457 = 10'h13c == _T_375[9:0] ? 4'h4 : _GEN_24456; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24458 = 10'h13d == _T_375[9:0] ? 4'h3 : _GEN_24457; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24459 = 10'h13e == _T_375[9:0] ? 4'h5 : _GEN_24458; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24460 = 10'h13f == _T_375[9:0] ? 4'h9 : _GEN_24459; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24461 = 10'h140 == _T_375[9:0] ? 4'ha : _GEN_24460; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24462 = 10'h141 == _T_375[9:0] ? 4'ha : _GEN_24461; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24463 = 10'h142 == _T_375[9:0] ? 4'ha : _GEN_24462; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24464 = 10'h143 == _T_375[9:0] ? 4'h5 : _GEN_24463; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24465 = 10'h144 == _T_375[9:0] ? 4'h3 : _GEN_24464; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24466 = 10'h145 == _T_375[9:0] ? 4'h3 : _GEN_24465; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24467 = 10'h146 == _T_375[9:0] ? 4'h3 : _GEN_24466; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24468 = 10'h147 == _T_375[9:0] ? 4'h4 : _GEN_24467; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24469 = 10'h148 == _T_375[9:0] ? 4'h3 : _GEN_24468; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24470 = 10'h149 == _T_375[9:0] ? 4'h3 : _GEN_24469; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24471 = 10'h14a == _T_375[9:0] ? 4'h3 : _GEN_24470; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24472 = 10'h14b == _T_375[9:0] ? 4'h6 : _GEN_24471; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24473 = 10'h14c == _T_375[9:0] ? 4'h8 : _GEN_24472; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24474 = 10'h14d == _T_375[9:0] ? 4'h5 : _GEN_24473; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24475 = 10'h14e == _T_375[9:0] ? 4'h4 : _GEN_24474; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24476 = 10'h14f == _T_375[9:0] ? 4'h3 : _GEN_24475; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24477 = 10'h150 == _T_375[9:0] ? 4'h3 : _GEN_24476; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24478 = 10'h151 == _T_375[9:0] ? 4'h3 : _GEN_24477; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24479 = 10'h152 == _T_375[9:0] ? 4'h3 : _GEN_24478; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24480 = 10'h153 == _T_375[9:0] ? 4'h3 : _GEN_24479; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24481 = 10'h154 == _T_375[9:0] ? 4'h3 : _GEN_24480; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24482 = 10'h155 == _T_375[9:0] ? 4'h4 : _GEN_24481; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24483 = 10'h156 == _T_375[9:0] ? 4'h9 : _GEN_24482; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24484 = 10'h157 == _T_375[9:0] ? 4'h8 : _GEN_24483; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24485 = 10'h158 == _T_375[9:0] ? 4'h8 : _GEN_24484; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24486 = 10'h159 == _T_375[9:0] ? 4'h8 : _GEN_24485; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24487 = 10'h15a == _T_375[9:0] ? 4'h8 : _GEN_24486; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24488 = 10'h15b == _T_375[9:0] ? 4'h8 : _GEN_24487; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24489 = 10'h15c == _T_375[9:0] ? 4'h7 : _GEN_24488; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24490 = 10'h15d == _T_375[9:0] ? 4'h7 : _GEN_24489; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24491 = 10'h15e == _T_375[9:0] ? 4'h8 : _GEN_24490; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24492 = 10'h15f == _T_375[9:0] ? 4'h3 : _GEN_24491; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24493 = 10'h160 == _T_375[9:0] ? 4'h4 : _GEN_24492; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24494 = 10'h161 == _T_375[9:0] ? 4'h4 : _GEN_24493; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24495 = 10'h162 == _T_375[9:0] ? 4'h4 : _GEN_24494; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24496 = 10'h163 == _T_375[9:0] ? 4'h4 : _GEN_24495; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24497 = 10'h164 == _T_375[9:0] ? 4'h5 : _GEN_24496; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24498 = 10'h165 == _T_375[9:0] ? 4'ha : _GEN_24497; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24499 = 10'h166 == _T_375[9:0] ? 4'h9 : _GEN_24498; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24500 = 10'h167 == _T_375[9:0] ? 4'ha : _GEN_24499; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24501 = 10'h168 == _T_375[9:0] ? 4'ha : _GEN_24500; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24502 = 10'h169 == _T_375[9:0] ? 4'h6 : _GEN_24501; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24503 = 10'h16a == _T_375[9:0] ? 4'h3 : _GEN_24502; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24504 = 10'h16b == _T_375[9:0] ? 4'h3 : _GEN_24503; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24505 = 10'h16c == _T_375[9:0] ? 4'h3 : _GEN_24504; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24506 = 10'h16d == _T_375[9:0] ? 4'h4 : _GEN_24505; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24507 = 10'h16e == _T_375[9:0] ? 4'h3 : _GEN_24506; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24508 = 10'h16f == _T_375[9:0] ? 4'h3 : _GEN_24507; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24509 = 10'h170 == _T_375[9:0] ? 4'h3 : _GEN_24508; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24510 = 10'h171 == _T_375[9:0] ? 4'h7 : _GEN_24509; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24511 = 10'h172 == _T_375[9:0] ? 4'ha : _GEN_24510; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24512 = 10'h173 == _T_375[9:0] ? 4'h5 : _GEN_24511; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24513 = 10'h174 == _T_375[9:0] ? 4'h3 : _GEN_24512; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24514 = 10'h175 == _T_375[9:0] ? 4'h4 : _GEN_24513; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24515 = 10'h176 == _T_375[9:0] ? 4'h4 : _GEN_24514; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24516 = 10'h177 == _T_375[9:0] ? 4'h4 : _GEN_24515; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24517 = 10'h178 == _T_375[9:0] ? 4'h4 : _GEN_24516; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24518 = 10'h179 == _T_375[9:0] ? 4'h3 : _GEN_24517; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24519 = 10'h17a == _T_375[9:0] ? 4'h3 : _GEN_24518; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24520 = 10'h17b == _T_375[9:0] ? 4'h3 : _GEN_24519; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24521 = 10'h17c == _T_375[9:0] ? 4'h8 : _GEN_24520; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24522 = 10'h17d == _T_375[9:0] ? 4'h8 : _GEN_24521; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24523 = 10'h17e == _T_375[9:0] ? 4'h8 : _GEN_24522; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24524 = 10'h17f == _T_375[9:0] ? 4'h8 : _GEN_24523; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24525 = 10'h180 == _T_375[9:0] ? 4'h8 : _GEN_24524; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24526 = 10'h181 == _T_375[9:0] ? 4'h8 : _GEN_24525; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24527 = 10'h182 == _T_375[9:0] ? 4'h8 : _GEN_24526; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24528 = 10'h183 == _T_375[9:0] ? 4'h8 : _GEN_24527; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24529 = 10'h184 == _T_375[9:0] ? 4'h8 : _GEN_24528; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24530 = 10'h185 == _T_375[9:0] ? 4'h5 : _GEN_24529; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24531 = 10'h186 == _T_375[9:0] ? 4'h3 : _GEN_24530; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24532 = 10'h187 == _T_375[9:0] ? 4'h4 : _GEN_24531; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24533 = 10'h188 == _T_375[9:0] ? 4'h4 : _GEN_24532; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24534 = 10'h189 == _T_375[9:0] ? 4'h4 : _GEN_24533; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24535 = 10'h18a == _T_375[9:0] ? 4'h5 : _GEN_24534; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24536 = 10'h18b == _T_375[9:0] ? 4'ha : _GEN_24535; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24537 = 10'h18c == _T_375[9:0] ? 4'ha : _GEN_24536; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24538 = 10'h18d == _T_375[9:0] ? 4'h9 : _GEN_24537; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24539 = 10'h18e == _T_375[9:0] ? 4'ha : _GEN_24538; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24540 = 10'h18f == _T_375[9:0] ? 4'h4 : _GEN_24539; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24541 = 10'h190 == _T_375[9:0] ? 4'h3 : _GEN_24540; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24542 = 10'h191 == _T_375[9:0] ? 4'h3 : _GEN_24541; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24543 = 10'h192 == _T_375[9:0] ? 4'h5 : _GEN_24542; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24544 = 10'h193 == _T_375[9:0] ? 4'h6 : _GEN_24543; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24545 = 10'h194 == _T_375[9:0] ? 4'h5 : _GEN_24544; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24546 = 10'h195 == _T_375[9:0] ? 4'h3 : _GEN_24545; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24547 = 10'h196 == _T_375[9:0] ? 4'h3 : _GEN_24546; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24548 = 10'h197 == _T_375[9:0] ? 4'h5 : _GEN_24547; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24549 = 10'h198 == _T_375[9:0] ? 4'ha : _GEN_24548; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24550 = 10'h199 == _T_375[9:0] ? 4'h3 : _GEN_24549; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24551 = 10'h19a == _T_375[9:0] ? 4'h1 : _GEN_24550; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24552 = 10'h19b == _T_375[9:0] ? 4'h2 : _GEN_24551; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24553 = 10'h19c == _T_375[9:0] ? 4'h4 : _GEN_24552; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24554 = 10'h19d == _T_375[9:0] ? 4'h3 : _GEN_24553; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24555 = 10'h19e == _T_375[9:0] ? 4'h1 : _GEN_24554; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24556 = 10'h19f == _T_375[9:0] ? 4'h2 : _GEN_24555; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24557 = 10'h1a0 == _T_375[9:0] ? 4'h3 : _GEN_24556; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24558 = 10'h1a1 == _T_375[9:0] ? 4'h4 : _GEN_24557; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24559 = 10'h1a2 == _T_375[9:0] ? 4'h8 : _GEN_24558; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24560 = 10'h1a3 == _T_375[9:0] ? 4'h8 : _GEN_24559; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24561 = 10'h1a4 == _T_375[9:0] ? 4'h8 : _GEN_24560; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24562 = 10'h1a5 == _T_375[9:0] ? 4'h8 : _GEN_24561; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24563 = 10'h1a6 == _T_375[9:0] ? 4'h7 : _GEN_24562; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24564 = 10'h1a7 == _T_375[9:0] ? 4'h8 : _GEN_24563; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24565 = 10'h1a8 == _T_375[9:0] ? 4'h8 : _GEN_24564; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24566 = 10'h1a9 == _T_375[9:0] ? 4'h8 : _GEN_24565; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24567 = 10'h1aa == _T_375[9:0] ? 4'h7 : _GEN_24566; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24568 = 10'h1ab == _T_375[9:0] ? 4'h4 : _GEN_24567; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24569 = 10'h1ac == _T_375[9:0] ? 4'h4 : _GEN_24568; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24570 = 10'h1ad == _T_375[9:0] ? 4'h3 : _GEN_24569; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24571 = 10'h1ae == _T_375[9:0] ? 4'h3 : _GEN_24570; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24572 = 10'h1af == _T_375[9:0] ? 4'h4 : _GEN_24571; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24573 = 10'h1b0 == _T_375[9:0] ? 4'h6 : _GEN_24572; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24574 = 10'h1b1 == _T_375[9:0] ? 4'ha : _GEN_24573; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24575 = 10'h1b2 == _T_375[9:0] ? 4'ha : _GEN_24574; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24576 = 10'h1b3 == _T_375[9:0] ? 4'h9 : _GEN_24575; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24577 = 10'h1b4 == _T_375[9:0] ? 4'h9 : _GEN_24576; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24578 = 10'h1b5 == _T_375[9:0] ? 4'h3 : _GEN_24577; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24579 = 10'h1b6 == _T_375[9:0] ? 4'h3 : _GEN_24578; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24580 = 10'h1b7 == _T_375[9:0] ? 4'h4 : _GEN_24579; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24581 = 10'h1b8 == _T_375[9:0] ? 4'h5 : _GEN_24580; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24582 = 10'h1b9 == _T_375[9:0] ? 4'h6 : _GEN_24581; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24583 = 10'h1ba == _T_375[9:0] ? 4'h4 : _GEN_24582; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24584 = 10'h1bb == _T_375[9:0] ? 4'h3 : _GEN_24583; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24585 = 10'h1bc == _T_375[9:0] ? 4'h3 : _GEN_24584; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24586 = 10'h1bd == _T_375[9:0] ? 4'h4 : _GEN_24585; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24587 = 10'h1be == _T_375[9:0] ? 4'ha : _GEN_24586; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24588 = 10'h1bf == _T_375[9:0] ? 4'h4 : _GEN_24587; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24589 = 10'h1c0 == _T_375[9:0] ? 4'h5 : _GEN_24588; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24590 = 10'h1c1 == _T_375[9:0] ? 4'h5 : _GEN_24589; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24591 = 10'h1c2 == _T_375[9:0] ? 4'h4 : _GEN_24590; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24592 = 10'h1c3 == _T_375[9:0] ? 4'h5 : _GEN_24591; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24593 = 10'h1c4 == _T_375[9:0] ? 4'h4 : _GEN_24592; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24594 = 10'h1c5 == _T_375[9:0] ? 4'h3 : _GEN_24593; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24595 = 10'h1c6 == _T_375[9:0] ? 4'h4 : _GEN_24594; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24596 = 10'h1c7 == _T_375[9:0] ? 4'h3 : _GEN_24595; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24597 = 10'h1c8 == _T_375[9:0] ? 4'h8 : _GEN_24596; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24598 = 10'h1c9 == _T_375[9:0] ? 4'h8 : _GEN_24597; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24599 = 10'h1ca == _T_375[9:0] ? 4'h8 : _GEN_24598; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24600 = 10'h1cb == _T_375[9:0] ? 4'h8 : _GEN_24599; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24601 = 10'h1cc == _T_375[9:0] ? 4'h8 : _GEN_24600; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24602 = 10'h1cd == _T_375[9:0] ? 4'h8 : _GEN_24601; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24603 = 10'h1ce == _T_375[9:0] ? 4'h8 : _GEN_24602; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24604 = 10'h1cf == _T_375[9:0] ? 4'h8 : _GEN_24603; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24605 = 10'h1d0 == _T_375[9:0] ? 4'h5 : _GEN_24604; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24606 = 10'h1d1 == _T_375[9:0] ? 4'h4 : _GEN_24605; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24607 = 10'h1d2 == _T_375[9:0] ? 4'h6 : _GEN_24606; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24608 = 10'h1d3 == _T_375[9:0] ? 4'h6 : _GEN_24607; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24609 = 10'h1d4 == _T_375[9:0] ? 4'h6 : _GEN_24608; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24610 = 10'h1d5 == _T_375[9:0] ? 4'h5 : _GEN_24609; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24611 = 10'h1d6 == _T_375[9:0] ? 4'h8 : _GEN_24610; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24612 = 10'h1d7 == _T_375[9:0] ? 4'ha : _GEN_24611; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24613 = 10'h1d8 == _T_375[9:0] ? 4'ha : _GEN_24612; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24614 = 10'h1d9 == _T_375[9:0] ? 4'ha : _GEN_24613; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24615 = 10'h1da == _T_375[9:0] ? 4'h6 : _GEN_24614; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24616 = 10'h1db == _T_375[9:0] ? 4'h3 : _GEN_24615; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24617 = 10'h1dc == _T_375[9:0] ? 4'h5 : _GEN_24616; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24618 = 10'h1dd == _T_375[9:0] ? 4'h2 : _GEN_24617; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24619 = 10'h1de == _T_375[9:0] ? 4'h5 : _GEN_24618; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24620 = 10'h1df == _T_375[9:0] ? 4'h5 : _GEN_24619; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24621 = 10'h1e0 == _T_375[9:0] ? 4'h5 : _GEN_24620; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24622 = 10'h1e1 == _T_375[9:0] ? 4'h3 : _GEN_24621; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24623 = 10'h1e2 == _T_375[9:0] ? 4'h3 : _GEN_24622; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24624 = 10'h1e3 == _T_375[9:0] ? 4'h3 : _GEN_24623; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24625 = 10'h1e4 == _T_375[9:0] ? 4'h9 : _GEN_24624; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24626 = 10'h1e5 == _T_375[9:0] ? 4'h4 : _GEN_24625; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24627 = 10'h1e6 == _T_375[9:0] ? 4'h4 : _GEN_24626; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24628 = 10'h1e7 == _T_375[9:0] ? 4'h4 : _GEN_24627; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24629 = 10'h1e8 == _T_375[9:0] ? 4'h4 : _GEN_24628; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24630 = 10'h1e9 == _T_375[9:0] ? 4'h4 : _GEN_24629; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24631 = 10'h1ea == _T_375[9:0] ? 4'h4 : _GEN_24630; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24632 = 10'h1eb == _T_375[9:0] ? 4'h4 : _GEN_24631; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24633 = 10'h1ec == _T_375[9:0] ? 4'h4 : _GEN_24632; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24634 = 10'h1ed == _T_375[9:0] ? 4'h4 : _GEN_24633; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24635 = 10'h1ee == _T_375[9:0] ? 4'h8 : _GEN_24634; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24636 = 10'h1ef == _T_375[9:0] ? 4'h8 : _GEN_24635; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24637 = 10'h1f0 == _T_375[9:0] ? 4'h8 : _GEN_24636; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24638 = 10'h1f1 == _T_375[9:0] ? 4'h8 : _GEN_24637; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24639 = 10'h1f2 == _T_375[9:0] ? 4'h8 : _GEN_24638; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24640 = 10'h1f3 == _T_375[9:0] ? 4'h8 : _GEN_24639; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24641 = 10'h1f4 == _T_375[9:0] ? 4'h9 : _GEN_24640; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24642 = 10'h1f5 == _T_375[9:0] ? 4'h9 : _GEN_24641; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24643 = 10'h1f6 == _T_375[9:0] ? 4'ha : _GEN_24642; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24644 = 10'h1f7 == _T_375[9:0] ? 4'h5 : _GEN_24643; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24645 = 10'h1f8 == _T_375[9:0] ? 4'h5 : _GEN_24644; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24646 = 10'h1f9 == _T_375[9:0] ? 4'h7 : _GEN_24645; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24647 = 10'h1fa == _T_375[9:0] ? 4'h7 : _GEN_24646; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24648 = 10'h1fb == _T_375[9:0] ? 4'h5 : _GEN_24647; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24649 = 10'h1fc == _T_375[9:0] ? 4'ha : _GEN_24648; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24650 = 10'h1fd == _T_375[9:0] ? 4'hb : _GEN_24649; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24651 = 10'h1fe == _T_375[9:0] ? 4'hb : _GEN_24650; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24652 = 10'h1ff == _T_375[9:0] ? 4'ha : _GEN_24651; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24653 = 10'h200 == _T_375[9:0] ? 4'h4 : _GEN_24652; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24654 = 10'h201 == _T_375[9:0] ? 4'h3 : _GEN_24653; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24655 = 10'h202 == _T_375[9:0] ? 4'h2 : _GEN_24654; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24656 = 10'h203 == _T_375[9:0] ? 4'h2 : _GEN_24655; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24657 = 10'h204 == _T_375[9:0] ? 4'h2 : _GEN_24656; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24658 = 10'h205 == _T_375[9:0] ? 4'h2 : _GEN_24657; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24659 = 10'h206 == _T_375[9:0] ? 4'h2 : _GEN_24658; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24660 = 10'h207 == _T_375[9:0] ? 4'h2 : _GEN_24659; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24661 = 10'h208 == _T_375[9:0] ? 4'h3 : _GEN_24660; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24662 = 10'h209 == _T_375[9:0] ? 4'h3 : _GEN_24661; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24663 = 10'h20a == _T_375[9:0] ? 4'h8 : _GEN_24662; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24664 = 10'h20b == _T_375[9:0] ? 4'h4 : _GEN_24663; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24665 = 10'h20c == _T_375[9:0] ? 4'h4 : _GEN_24664; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24666 = 10'h20d == _T_375[9:0] ? 4'h4 : _GEN_24665; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24667 = 10'h20e == _T_375[9:0] ? 4'h4 : _GEN_24666; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24668 = 10'h20f == _T_375[9:0] ? 4'h4 : _GEN_24667; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24669 = 10'h210 == _T_375[9:0] ? 4'h4 : _GEN_24668; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24670 = 10'h211 == _T_375[9:0] ? 4'h4 : _GEN_24669; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24671 = 10'h212 == _T_375[9:0] ? 4'h4 : _GEN_24670; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24672 = 10'h213 == _T_375[9:0] ? 4'h6 : _GEN_24671; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24673 = 10'h214 == _T_375[9:0] ? 4'h7 : _GEN_24672; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24674 = 10'h215 == _T_375[9:0] ? 4'h8 : _GEN_24673; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24675 = 10'h216 == _T_375[9:0] ? 4'h8 : _GEN_24674; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24676 = 10'h217 == _T_375[9:0] ? 4'h8 : _GEN_24675; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24677 = 10'h218 == _T_375[9:0] ? 4'h8 : _GEN_24676; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24678 = 10'h219 == _T_375[9:0] ? 4'h8 : _GEN_24677; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24679 = 10'h21a == _T_375[9:0] ? 4'h8 : _GEN_24678; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24680 = 10'h21b == _T_375[9:0] ? 4'h8 : _GEN_24679; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24681 = 10'h21c == _T_375[9:0] ? 4'ha : _GEN_24680; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24682 = 10'h21d == _T_375[9:0] ? 4'h9 : _GEN_24681; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24683 = 10'h21e == _T_375[9:0] ? 4'h6 : _GEN_24682; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24684 = 10'h21f == _T_375[9:0] ? 4'h4 : _GEN_24683; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24685 = 10'h220 == _T_375[9:0] ? 4'h4 : _GEN_24684; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24686 = 10'h221 == _T_375[9:0] ? 4'h5 : _GEN_24685; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24687 = 10'h222 == _T_375[9:0] ? 4'ha : _GEN_24686; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24688 = 10'h223 == _T_375[9:0] ? 4'ha : _GEN_24687; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24689 = 10'h224 == _T_375[9:0] ? 4'ha : _GEN_24688; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24690 = 10'h225 == _T_375[9:0] ? 4'h8 : _GEN_24689; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24691 = 10'h226 == _T_375[9:0] ? 4'h4 : _GEN_24690; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24692 = 10'h227 == _T_375[9:0] ? 4'h2 : _GEN_24691; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24693 = 10'h228 == _T_375[9:0] ? 4'h2 : _GEN_24692; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24694 = 10'h229 == _T_375[9:0] ? 4'h2 : _GEN_24693; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24695 = 10'h22a == _T_375[9:0] ? 4'h2 : _GEN_24694; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24696 = 10'h22b == _T_375[9:0] ? 4'h2 : _GEN_24695; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24697 = 10'h22c == _T_375[9:0] ? 4'h2 : _GEN_24696; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24698 = 10'h22d == _T_375[9:0] ? 4'h2 : _GEN_24697; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24699 = 10'h22e == _T_375[9:0] ? 4'h2 : _GEN_24698; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24700 = 10'h22f == _T_375[9:0] ? 4'h3 : _GEN_24699; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24701 = 10'h230 == _T_375[9:0] ? 4'h3 : _GEN_24700; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24702 = 10'h231 == _T_375[9:0] ? 4'h3 : _GEN_24701; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24703 = 10'h232 == _T_375[9:0] ? 4'h4 : _GEN_24702; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24704 = 10'h233 == _T_375[9:0] ? 4'h6 : _GEN_24703; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24705 = 10'h234 == _T_375[9:0] ? 4'h6 : _GEN_24704; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24706 = 10'h235 == _T_375[9:0] ? 4'h4 : _GEN_24705; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24707 = 10'h236 == _T_375[9:0] ? 4'h4 : _GEN_24706; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24708 = 10'h237 == _T_375[9:0] ? 4'h4 : _GEN_24707; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24709 = 10'h238 == _T_375[9:0] ? 4'h4 : _GEN_24708; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24710 = 10'h239 == _T_375[9:0] ? 4'h3 : _GEN_24709; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24711 = 10'h23a == _T_375[9:0] ? 4'h7 : _GEN_24710; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24712 = 10'h23b == _T_375[9:0] ? 4'h7 : _GEN_24711; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24713 = 10'h23c == _T_375[9:0] ? 4'h7 : _GEN_24712; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24714 = 10'h23d == _T_375[9:0] ? 4'h7 : _GEN_24713; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24715 = 10'h23e == _T_375[9:0] ? 4'h7 : _GEN_24714; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24716 = 10'h23f == _T_375[9:0] ? 4'h7 : _GEN_24715; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24717 = 10'h240 == _T_375[9:0] ? 4'h7 : _GEN_24716; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24718 = 10'h241 == _T_375[9:0] ? 4'h8 : _GEN_24717; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24719 = 10'h242 == _T_375[9:0] ? 4'ha : _GEN_24718; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24720 = 10'h243 == _T_375[9:0] ? 4'ha : _GEN_24719; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24721 = 10'h244 == _T_375[9:0] ? 4'ha : _GEN_24720; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24722 = 10'h245 == _T_375[9:0] ? 4'h8 : _GEN_24721; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24723 = 10'h246 == _T_375[9:0] ? 4'h7 : _GEN_24722; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24724 = 10'h247 == _T_375[9:0] ? 4'h8 : _GEN_24723; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24725 = 10'h248 == _T_375[9:0] ? 4'ha : _GEN_24724; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24726 = 10'h249 == _T_375[9:0] ? 4'ha : _GEN_24725; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24727 = 10'h24a == _T_375[9:0] ? 4'ha : _GEN_24726; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24728 = 10'h24b == _T_375[9:0] ? 4'h4 : _GEN_24727; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24729 = 10'h24c == _T_375[9:0] ? 4'h4 : _GEN_24728; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24730 = 10'h24d == _T_375[9:0] ? 4'h2 : _GEN_24729; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24731 = 10'h24e == _T_375[9:0] ? 4'h2 : _GEN_24730; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24732 = 10'h24f == _T_375[9:0] ? 4'h2 : _GEN_24731; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24733 = 10'h250 == _T_375[9:0] ? 4'h2 : _GEN_24732; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24734 = 10'h251 == _T_375[9:0] ? 4'h2 : _GEN_24733; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24735 = 10'h252 == _T_375[9:0] ? 4'h2 : _GEN_24734; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24736 = 10'h253 == _T_375[9:0] ? 4'h2 : _GEN_24735; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24737 = 10'h254 == _T_375[9:0] ? 4'h2 : _GEN_24736; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24738 = 10'h255 == _T_375[9:0] ? 4'h3 : _GEN_24737; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24739 = 10'h256 == _T_375[9:0] ? 4'h4 : _GEN_24738; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24740 = 10'h257 == _T_375[9:0] ? 4'h3 : _GEN_24739; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24741 = 10'h258 == _T_375[9:0] ? 4'h4 : _GEN_24740; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24742 = 10'h259 == _T_375[9:0] ? 4'h4 : _GEN_24741; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24743 = 10'h25a == _T_375[9:0] ? 4'h4 : _GEN_24742; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24744 = 10'h25b == _T_375[9:0] ? 4'h3 : _GEN_24743; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24745 = 10'h25c == _T_375[9:0] ? 4'h4 : _GEN_24744; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24746 = 10'h25d == _T_375[9:0] ? 4'h4 : _GEN_24745; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24747 = 10'h25e == _T_375[9:0] ? 4'h3 : _GEN_24746; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24748 = 10'h25f == _T_375[9:0] ? 4'h3 : _GEN_24747; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24749 = 10'h260 == _T_375[9:0] ? 4'h8 : _GEN_24748; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24750 = 10'h261 == _T_375[9:0] ? 4'h7 : _GEN_24749; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24751 = 10'h262 == _T_375[9:0] ? 4'h6 : _GEN_24750; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24752 = 10'h263 == _T_375[9:0] ? 4'h5 : _GEN_24751; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24753 = 10'h264 == _T_375[9:0] ? 4'h6 : _GEN_24752; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24754 = 10'h265 == _T_375[9:0] ? 4'h5 : _GEN_24753; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24755 = 10'h266 == _T_375[9:0] ? 4'h5 : _GEN_24754; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24756 = 10'h267 == _T_375[9:0] ? 4'h7 : _GEN_24755; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24757 = 10'h268 == _T_375[9:0] ? 4'ha : _GEN_24756; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24758 = 10'h269 == _T_375[9:0] ? 4'ha : _GEN_24757; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24759 = 10'h26a == _T_375[9:0] ? 4'ha : _GEN_24758; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24760 = 10'h26b == _T_375[9:0] ? 4'ha : _GEN_24759; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24761 = 10'h26c == _T_375[9:0] ? 4'ha : _GEN_24760; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24762 = 10'h26d == _T_375[9:0] ? 4'ha : _GEN_24761; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24763 = 10'h26e == _T_375[9:0] ? 4'ha : _GEN_24762; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24764 = 10'h26f == _T_375[9:0] ? 4'ha : _GEN_24763; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24765 = 10'h270 == _T_375[9:0] ? 4'h5 : _GEN_24764; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24766 = 10'h271 == _T_375[9:0] ? 4'h4 : _GEN_24765; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24767 = 10'h272 == _T_375[9:0] ? 4'h3 : _GEN_24766; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24768 = 10'h273 == _T_375[9:0] ? 4'h2 : _GEN_24767; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24769 = 10'h274 == _T_375[9:0] ? 4'h2 : _GEN_24768; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24770 = 10'h275 == _T_375[9:0] ? 4'h2 : _GEN_24769; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24771 = 10'h276 == _T_375[9:0] ? 4'h2 : _GEN_24770; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24772 = 10'h277 == _T_375[9:0] ? 4'h2 : _GEN_24771; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24773 = 10'h278 == _T_375[9:0] ? 4'h2 : _GEN_24772; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24774 = 10'h279 == _T_375[9:0] ? 4'h2 : _GEN_24773; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24775 = 10'h27a == _T_375[9:0] ? 4'h2 : _GEN_24774; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24776 = 10'h27b == _T_375[9:0] ? 4'h4 : _GEN_24775; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24777 = 10'h27c == _T_375[9:0] ? 4'h3 : _GEN_24776; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24778 = 10'h27d == _T_375[9:0] ? 4'h4 : _GEN_24777; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24779 = 10'h27e == _T_375[9:0] ? 4'h5 : _GEN_24778; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24780 = 10'h27f == _T_375[9:0] ? 4'h4 : _GEN_24779; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24781 = 10'h280 == _T_375[9:0] ? 4'h4 : _GEN_24780; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24782 = 10'h281 == _T_375[9:0] ? 4'h4 : _GEN_24781; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24783 = 10'h282 == _T_375[9:0] ? 4'h4 : _GEN_24782; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24784 = 10'h283 == _T_375[9:0] ? 4'h3 : _GEN_24783; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24785 = 10'h284 == _T_375[9:0] ? 4'h3 : _GEN_24784; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24786 = 10'h285 == _T_375[9:0] ? 4'h3 : _GEN_24785; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24787 = 10'h286 == _T_375[9:0] ? 4'h8 : _GEN_24786; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24788 = 10'h287 == _T_375[9:0] ? 4'h6 : _GEN_24787; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24789 = 10'h288 == _T_375[9:0] ? 4'h6 : _GEN_24788; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24790 = 10'h289 == _T_375[9:0] ? 4'h6 : _GEN_24789; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24791 = 10'h28a == _T_375[9:0] ? 4'h7 : _GEN_24790; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24792 = 10'h28b == _T_375[9:0] ? 4'h7 : _GEN_24791; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24793 = 10'h28c == _T_375[9:0] ? 4'h6 : _GEN_24792; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24794 = 10'h28d == _T_375[9:0] ? 4'h6 : _GEN_24793; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24795 = 10'h28e == _T_375[9:0] ? 4'h4 : _GEN_24794; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24796 = 10'h28f == _T_375[9:0] ? 4'h7 : _GEN_24795; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24797 = 10'h290 == _T_375[9:0] ? 4'h9 : _GEN_24796; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24798 = 10'h291 == _T_375[9:0] ? 4'ha : _GEN_24797; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24799 = 10'h292 == _T_375[9:0] ? 4'ha : _GEN_24798; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24800 = 10'h293 == _T_375[9:0] ? 4'ha : _GEN_24799; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24801 = 10'h294 == _T_375[9:0] ? 4'h9 : _GEN_24800; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24802 = 10'h295 == _T_375[9:0] ? 4'h5 : _GEN_24801; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24803 = 10'h296 == _T_375[9:0] ? 4'h4 : _GEN_24802; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24804 = 10'h297 == _T_375[9:0] ? 4'h4 : _GEN_24803; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24805 = 10'h298 == _T_375[9:0] ? 4'h3 : _GEN_24804; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24806 = 10'h299 == _T_375[9:0] ? 4'h3 : _GEN_24805; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24807 = 10'h29a == _T_375[9:0] ? 4'h2 : _GEN_24806; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24808 = 10'h29b == _T_375[9:0] ? 4'h2 : _GEN_24807; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24809 = 10'h29c == _T_375[9:0] ? 4'h2 : _GEN_24808; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24810 = 10'h29d == _T_375[9:0] ? 4'h2 : _GEN_24809; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24811 = 10'h29e == _T_375[9:0] ? 4'h2 : _GEN_24810; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24812 = 10'h29f == _T_375[9:0] ? 4'h2 : _GEN_24811; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24813 = 10'h2a0 == _T_375[9:0] ? 4'h2 : _GEN_24812; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24814 = 10'h2a1 == _T_375[9:0] ? 4'h4 : _GEN_24813; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24815 = 10'h2a2 == _T_375[9:0] ? 4'h3 : _GEN_24814; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24816 = 10'h2a3 == _T_375[9:0] ? 4'h4 : _GEN_24815; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24817 = 10'h2a4 == _T_375[9:0] ? 4'h5 : _GEN_24816; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24818 = 10'h2a5 == _T_375[9:0] ? 4'h4 : _GEN_24817; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24819 = 10'h2a6 == _T_375[9:0] ? 4'h4 : _GEN_24818; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24820 = 10'h2a7 == _T_375[9:0] ? 4'h4 : _GEN_24819; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24821 = 10'h2a8 == _T_375[9:0] ? 4'h3 : _GEN_24820; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24822 = 10'h2a9 == _T_375[9:0] ? 4'h3 : _GEN_24821; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24823 = 10'h2aa == _T_375[9:0] ? 4'h3 : _GEN_24822; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24824 = 10'h2ab == _T_375[9:0] ? 4'h3 : _GEN_24823; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24825 = 10'h2ac == _T_375[9:0] ? 4'h8 : _GEN_24824; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24826 = 10'h2ad == _T_375[9:0] ? 4'h7 : _GEN_24825; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24827 = 10'h2ae == _T_375[9:0] ? 4'h5 : _GEN_24826; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24828 = 10'h2af == _T_375[9:0] ? 4'h6 : _GEN_24827; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24829 = 10'h2b0 == _T_375[9:0] ? 4'h7 : _GEN_24828; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24830 = 10'h2b1 == _T_375[9:0] ? 4'h6 : _GEN_24829; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24831 = 10'h2b2 == _T_375[9:0] ? 4'h6 : _GEN_24830; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24832 = 10'h2b3 == _T_375[9:0] ? 4'h6 : _GEN_24831; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24833 = 10'h2b4 == _T_375[9:0] ? 4'h3 : _GEN_24832; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24834 = 10'h2b5 == _T_375[9:0] ? 4'h3 : _GEN_24833; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24835 = 10'h2b6 == _T_375[9:0] ? 4'h3 : _GEN_24834; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24836 = 10'h2b7 == _T_375[9:0] ? 4'h4 : _GEN_24835; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24837 = 10'h2b8 == _T_375[9:0] ? 4'h6 : _GEN_24836; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24838 = 10'h2b9 == _T_375[9:0] ? 4'h9 : _GEN_24837; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24839 = 10'h2ba == _T_375[9:0] ? 4'h4 : _GEN_24838; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24840 = 10'h2bb == _T_375[9:0] ? 4'h3 : _GEN_24839; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24841 = 10'h2bc == _T_375[9:0] ? 4'h4 : _GEN_24840; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24842 = 10'h2bd == _T_375[9:0] ? 4'h3 : _GEN_24841; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24843 = 10'h2be == _T_375[9:0] ? 4'h3 : _GEN_24842; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24844 = 10'h2bf == _T_375[9:0] ? 4'h3 : _GEN_24843; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24845 = 10'h2c0 == _T_375[9:0] ? 4'h2 : _GEN_24844; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24846 = 10'h2c1 == _T_375[9:0] ? 4'h2 : _GEN_24845; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24847 = 10'h2c2 == _T_375[9:0] ? 4'h2 : _GEN_24846; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24848 = 10'h2c3 == _T_375[9:0] ? 4'h2 : _GEN_24847; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24849 = 10'h2c4 == _T_375[9:0] ? 4'h2 : _GEN_24848; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24850 = 10'h2c5 == _T_375[9:0] ? 4'h2 : _GEN_24849; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24851 = 10'h2c6 == _T_375[9:0] ? 4'h2 : _GEN_24850; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24852 = 10'h2c7 == _T_375[9:0] ? 4'h4 : _GEN_24851; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24853 = 10'h2c8 == _T_375[9:0] ? 4'h3 : _GEN_24852; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24854 = 10'h2c9 == _T_375[9:0] ? 4'h4 : _GEN_24853; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24855 = 10'h2ca == _T_375[9:0] ? 4'h5 : _GEN_24854; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24856 = 10'h2cb == _T_375[9:0] ? 4'h3 : _GEN_24855; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24857 = 10'h2cc == _T_375[9:0] ? 4'h3 : _GEN_24856; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24858 = 10'h2cd == _T_375[9:0] ? 4'h3 : _GEN_24857; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24859 = 10'h2ce == _T_375[9:0] ? 4'h3 : _GEN_24858; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24860 = 10'h2cf == _T_375[9:0] ? 4'h3 : _GEN_24859; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24861 = 10'h2d0 == _T_375[9:0] ? 4'h3 : _GEN_24860; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24862 = 10'h2d1 == _T_375[9:0] ? 4'h3 : _GEN_24861; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24863 = 10'h2d2 == _T_375[9:0] ? 4'h8 : _GEN_24862; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24864 = 10'h2d3 == _T_375[9:0] ? 4'h6 : _GEN_24863; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24865 = 10'h2d4 == _T_375[9:0] ? 4'h6 : _GEN_24864; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24866 = 10'h2d5 == _T_375[9:0] ? 4'h7 : _GEN_24865; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24867 = 10'h2d6 == _T_375[9:0] ? 4'h7 : _GEN_24866; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24868 = 10'h2d7 == _T_375[9:0] ? 4'h7 : _GEN_24867; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24869 = 10'h2d8 == _T_375[9:0] ? 4'h6 : _GEN_24868; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24870 = 10'h2d9 == _T_375[9:0] ? 4'h7 : _GEN_24869; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24871 = 10'h2da == _T_375[9:0] ? 4'h5 : _GEN_24870; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24872 = 10'h2db == _T_375[9:0] ? 4'h3 : _GEN_24871; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24873 = 10'h2dc == _T_375[9:0] ? 4'h3 : _GEN_24872; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24874 = 10'h2dd == _T_375[9:0] ? 4'h3 : _GEN_24873; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24875 = 10'h2de == _T_375[9:0] ? 4'h3 : _GEN_24874; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24876 = 10'h2df == _T_375[9:0] ? 4'h4 : _GEN_24875; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24877 = 10'h2e0 == _T_375[9:0] ? 4'h3 : _GEN_24876; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24878 = 10'h2e1 == _T_375[9:0] ? 4'h3 : _GEN_24877; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24879 = 10'h2e2 == _T_375[9:0] ? 4'h3 : _GEN_24878; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24880 = 10'h2e3 == _T_375[9:0] ? 4'h3 : _GEN_24879; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24881 = 10'h2e4 == _T_375[9:0] ? 4'h3 : _GEN_24880; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24882 = 10'h2e5 == _T_375[9:0] ? 4'h3 : _GEN_24881; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24883 = 10'h2e6 == _T_375[9:0] ? 4'h2 : _GEN_24882; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24884 = 10'h2e7 == _T_375[9:0] ? 4'h2 : _GEN_24883; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24885 = 10'h2e8 == _T_375[9:0] ? 4'h2 : _GEN_24884; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24886 = 10'h2e9 == _T_375[9:0] ? 4'h2 : _GEN_24885; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24887 = 10'h2ea == _T_375[9:0] ? 4'h2 : _GEN_24886; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24888 = 10'h2eb == _T_375[9:0] ? 4'h2 : _GEN_24887; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24889 = 10'h2ec == _T_375[9:0] ? 4'h3 : _GEN_24888; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24890 = 10'h2ed == _T_375[9:0] ? 4'h4 : _GEN_24889; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24891 = 10'h2ee == _T_375[9:0] ? 4'h3 : _GEN_24890; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24892 = 10'h2ef == _T_375[9:0] ? 4'h3 : _GEN_24891; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24893 = 10'h2f0 == _T_375[9:0] ? 4'h6 : _GEN_24892; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24894 = 10'h2f1 == _T_375[9:0] ? 4'h3 : _GEN_24893; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24895 = 10'h2f2 == _T_375[9:0] ? 4'h3 : _GEN_24894; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24896 = 10'h2f3 == _T_375[9:0] ? 4'h3 : _GEN_24895; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24897 = 10'h2f4 == _T_375[9:0] ? 4'h3 : _GEN_24896; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24898 = 10'h2f5 == _T_375[9:0] ? 4'h3 : _GEN_24897; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24899 = 10'h2f6 == _T_375[9:0] ? 4'h3 : _GEN_24898; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24900 = 10'h2f7 == _T_375[9:0] ? 4'h3 : _GEN_24899; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24901 = 10'h2f8 == _T_375[9:0] ? 4'h8 : _GEN_24900; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24902 = 10'h2f9 == _T_375[9:0] ? 4'h6 : _GEN_24901; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24903 = 10'h2fa == _T_375[9:0] ? 4'h7 : _GEN_24902; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24904 = 10'h2fb == _T_375[9:0] ? 4'h7 : _GEN_24903; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24905 = 10'h2fc == _T_375[9:0] ? 4'h6 : _GEN_24904; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24906 = 10'h2fd == _T_375[9:0] ? 4'h6 : _GEN_24905; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24907 = 10'h2fe == _T_375[9:0] ? 4'h6 : _GEN_24906; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24908 = 10'h2ff == _T_375[9:0] ? 4'h8 : _GEN_24907; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24909 = 10'h300 == _T_375[9:0] ? 4'h9 : _GEN_24908; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24910 = 10'h301 == _T_375[9:0] ? 4'h7 : _GEN_24909; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24911 = 10'h302 == _T_375[9:0] ? 4'h4 : _GEN_24910; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24912 = 10'h303 == _T_375[9:0] ? 4'h4 : _GEN_24911; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24913 = 10'h304 == _T_375[9:0] ? 4'h3 : _GEN_24912; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24914 = 10'h305 == _T_375[9:0] ? 4'h3 : _GEN_24913; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24915 = 10'h306 == _T_375[9:0] ? 4'h3 : _GEN_24914; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24916 = 10'h307 == _T_375[9:0] ? 4'h3 : _GEN_24915; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24917 = 10'h308 == _T_375[9:0] ? 4'h3 : _GEN_24916; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24918 = 10'h309 == _T_375[9:0] ? 4'h3 : _GEN_24917; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24919 = 10'h30a == _T_375[9:0] ? 4'h3 : _GEN_24918; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24920 = 10'h30b == _T_375[9:0] ? 4'h3 : _GEN_24919; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24921 = 10'h30c == _T_375[9:0] ? 4'h2 : _GEN_24920; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24922 = 10'h30d == _T_375[9:0] ? 4'h2 : _GEN_24921; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24923 = 10'h30e == _T_375[9:0] ? 4'h2 : _GEN_24922; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24924 = 10'h30f == _T_375[9:0] ? 4'h2 : _GEN_24923; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24925 = 10'h310 == _T_375[9:0] ? 4'h2 : _GEN_24924; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24926 = 10'h311 == _T_375[9:0] ? 4'h2 : _GEN_24925; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24927 = 10'h312 == _T_375[9:0] ? 4'h3 : _GEN_24926; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24928 = 10'h313 == _T_375[9:0] ? 4'h4 : _GEN_24927; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24929 = 10'h314 == _T_375[9:0] ? 4'h3 : _GEN_24928; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24930 = 10'h315 == _T_375[9:0] ? 4'h3 : _GEN_24929; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24931 = 10'h316 == _T_375[9:0] ? 4'h5 : _GEN_24930; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24932 = 10'h317 == _T_375[9:0] ? 4'h5 : _GEN_24931; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24933 = 10'h318 == _T_375[9:0] ? 4'h3 : _GEN_24932; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24934 = 10'h319 == _T_375[9:0] ? 4'h3 : _GEN_24933; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24935 = 10'h31a == _T_375[9:0] ? 4'h3 : _GEN_24934; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24936 = 10'h31b == _T_375[9:0] ? 4'h3 : _GEN_24935; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24937 = 10'h31c == _T_375[9:0] ? 4'h3 : _GEN_24936; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24938 = 10'h31d == _T_375[9:0] ? 4'h3 : _GEN_24937; // @[Filter.scala 230:62]
  wire [4:0] _GEN_39014 = {{1'd0}, _GEN_24938}; // @[Filter.scala 230:62]
  wire [8:0] _T_377 = _GEN_39014 * 5'h14; // @[Filter.scala 230:62]
  wire [3:0] _GEN_24962 = 10'h17 == _T_375[9:0] ? 4'hb : 4'he; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24963 = 10'h18 == _T_375[9:0] ? 4'hc : _GEN_24962; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24964 = 10'h19 == _T_375[9:0] ? 4'he : _GEN_24963; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24965 = 10'h1a == _T_375[9:0] ? 4'he : _GEN_24964; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24966 = 10'h1b == _T_375[9:0] ? 4'he : _GEN_24965; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24967 = 10'h1c == _T_375[9:0] ? 4'he : _GEN_24966; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24968 = 10'h1d == _T_375[9:0] ? 4'he : _GEN_24967; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24969 = 10'h1e == _T_375[9:0] ? 4'he : _GEN_24968; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24970 = 10'h1f == _T_375[9:0] ? 4'he : _GEN_24969; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24971 = 10'h20 == _T_375[9:0] ? 4'he : _GEN_24970; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24972 = 10'h21 == _T_375[9:0] ? 4'he : _GEN_24971; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24973 = 10'h22 == _T_375[9:0] ? 4'he : _GEN_24972; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24974 = 10'h23 == _T_375[9:0] ? 4'he : _GEN_24973; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24975 = 10'h24 == _T_375[9:0] ? 4'he : _GEN_24974; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24976 = 10'h25 == _T_375[9:0] ? 4'he : _GEN_24975; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24977 = 10'h26 == _T_375[9:0] ? 4'he : _GEN_24976; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24978 = 10'h27 == _T_375[9:0] ? 4'he : _GEN_24977; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24979 = 10'h28 == _T_375[9:0] ? 4'he : _GEN_24978; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24980 = 10'h29 == _T_375[9:0] ? 4'he : _GEN_24979; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24981 = 10'h2a == _T_375[9:0] ? 4'he : _GEN_24980; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24982 = 10'h2b == _T_375[9:0] ? 4'he : _GEN_24981; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24983 = 10'h2c == _T_375[9:0] ? 4'he : _GEN_24982; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24984 = 10'h2d == _T_375[9:0] ? 4'he : _GEN_24983; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24985 = 10'h2e == _T_375[9:0] ? 4'he : _GEN_24984; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24986 = 10'h2f == _T_375[9:0] ? 4'he : _GEN_24985; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24987 = 10'h30 == _T_375[9:0] ? 4'he : _GEN_24986; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24988 = 10'h31 == _T_375[9:0] ? 4'he : _GEN_24987; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24989 = 10'h32 == _T_375[9:0] ? 4'he : _GEN_24988; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24990 = 10'h33 == _T_375[9:0] ? 4'he : _GEN_24989; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24991 = 10'h34 == _T_375[9:0] ? 4'he : _GEN_24990; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24992 = 10'h35 == _T_375[9:0] ? 4'he : _GEN_24991; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24993 = 10'h36 == _T_375[9:0] ? 4'he : _GEN_24992; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24994 = 10'h37 == _T_375[9:0] ? 4'he : _GEN_24993; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24995 = 10'h38 == _T_375[9:0] ? 4'he : _GEN_24994; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24996 = 10'h39 == _T_375[9:0] ? 4'he : _GEN_24995; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24997 = 10'h3a == _T_375[9:0] ? 4'he : _GEN_24996; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24998 = 10'h3b == _T_375[9:0] ? 4'he : _GEN_24997; // @[Filter.scala 230:102]
  wire [3:0] _GEN_24999 = 10'h3c == _T_375[9:0] ? 4'ha : _GEN_24998; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25000 = 10'h3d == _T_375[9:0] ? 4'hc : _GEN_24999; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25001 = 10'h3e == _T_375[9:0] ? 4'hb : _GEN_25000; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25002 = 10'h3f == _T_375[9:0] ? 4'he : _GEN_25001; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25003 = 10'h40 == _T_375[9:0] ? 4'he : _GEN_25002; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25004 = 10'h41 == _T_375[9:0] ? 4'he : _GEN_25003; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25005 = 10'h42 == _T_375[9:0] ? 4'he : _GEN_25004; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25006 = 10'h43 == _T_375[9:0] ? 4'he : _GEN_25005; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25007 = 10'h44 == _T_375[9:0] ? 4'he : _GEN_25006; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25008 = 10'h45 == _T_375[9:0] ? 4'he : _GEN_25007; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25009 = 10'h46 == _T_375[9:0] ? 4'he : _GEN_25008; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25010 = 10'h47 == _T_375[9:0] ? 4'he : _GEN_25009; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25011 = 10'h48 == _T_375[9:0] ? 4'he : _GEN_25010; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25012 = 10'h49 == _T_375[9:0] ? 4'he : _GEN_25011; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25013 = 10'h4a == _T_375[9:0] ? 4'he : _GEN_25012; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25014 = 10'h4b == _T_375[9:0] ? 4'he : _GEN_25013; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25015 = 10'h4c == _T_375[9:0] ? 4'he : _GEN_25014; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25016 = 10'h4d == _T_375[9:0] ? 4'he : _GEN_25015; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25017 = 10'h4e == _T_375[9:0] ? 4'he : _GEN_25016; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25018 = 10'h4f == _T_375[9:0] ? 4'he : _GEN_25017; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25019 = 10'h50 == _T_375[9:0] ? 4'he : _GEN_25018; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25020 = 10'h51 == _T_375[9:0] ? 4'he : _GEN_25019; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25021 = 10'h52 == _T_375[9:0] ? 4'he : _GEN_25020; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25022 = 10'h53 == _T_375[9:0] ? 4'he : _GEN_25021; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25023 = 10'h54 == _T_375[9:0] ? 4'he : _GEN_25022; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25024 = 10'h55 == _T_375[9:0] ? 4'he : _GEN_25023; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25025 = 10'h56 == _T_375[9:0] ? 4'he : _GEN_25024; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25026 = 10'h57 == _T_375[9:0] ? 4'he : _GEN_25025; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25027 = 10'h58 == _T_375[9:0] ? 4'he : _GEN_25026; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25028 = 10'h59 == _T_375[9:0] ? 4'he : _GEN_25027; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25029 = 10'h5a == _T_375[9:0] ? 4'hc : _GEN_25028; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25030 = 10'h5b == _T_375[9:0] ? 4'hd : _GEN_25029; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25031 = 10'h5c == _T_375[9:0] ? 4'he : _GEN_25030; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25032 = 10'h5d == _T_375[9:0] ? 4'he : _GEN_25031; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25033 = 10'h5e == _T_375[9:0] ? 4'he : _GEN_25032; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25034 = 10'h5f == _T_375[9:0] ? 4'he : _GEN_25033; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25035 = 10'h60 == _T_375[9:0] ? 4'he : _GEN_25034; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25036 = 10'h61 == _T_375[9:0] ? 4'hd : _GEN_25035; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25037 = 10'h62 == _T_375[9:0] ? 4'hb : _GEN_25036; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25038 = 10'h63 == _T_375[9:0] ? 4'hc : _GEN_25037; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25039 = 10'h64 == _T_375[9:0] ? 4'ha : _GEN_25038; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25040 = 10'h65 == _T_375[9:0] ? 4'hd : _GEN_25039; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25041 = 10'h66 == _T_375[9:0] ? 4'he : _GEN_25040; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25042 = 10'h67 == _T_375[9:0] ? 4'he : _GEN_25041; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25043 = 10'h68 == _T_375[9:0] ? 4'he : _GEN_25042; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25044 = 10'h69 == _T_375[9:0] ? 4'he : _GEN_25043; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25045 = 10'h6a == _T_375[9:0] ? 4'he : _GEN_25044; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25046 = 10'h6b == _T_375[9:0] ? 4'hd : _GEN_25045; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25047 = 10'h6c == _T_375[9:0] ? 4'hc : _GEN_25046; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25048 = 10'h6d == _T_375[9:0] ? 4'hc : _GEN_25047; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25049 = 10'h6e == _T_375[9:0] ? 4'he : _GEN_25048; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25050 = 10'h6f == _T_375[9:0] ? 4'he : _GEN_25049; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25051 = 10'h70 == _T_375[9:0] ? 4'he : _GEN_25050; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25052 = 10'h71 == _T_375[9:0] ? 4'he : _GEN_25051; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25053 = 10'h72 == _T_375[9:0] ? 4'he : _GEN_25052; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25054 = 10'h73 == _T_375[9:0] ? 4'he : _GEN_25053; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25055 = 10'h74 == _T_375[9:0] ? 4'he : _GEN_25054; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25056 = 10'h75 == _T_375[9:0] ? 4'he : _GEN_25055; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25057 = 10'h76 == _T_375[9:0] ? 4'he : _GEN_25056; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25058 = 10'h77 == _T_375[9:0] ? 4'he : _GEN_25057; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25059 = 10'h78 == _T_375[9:0] ? 4'he : _GEN_25058; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25060 = 10'h79 == _T_375[9:0] ? 4'he : _GEN_25059; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25061 = 10'h7a == _T_375[9:0] ? 4'he : _GEN_25060; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25062 = 10'h7b == _T_375[9:0] ? 4'he : _GEN_25061; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25063 = 10'h7c == _T_375[9:0] ? 4'he : _GEN_25062; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25064 = 10'h7d == _T_375[9:0] ? 4'he : _GEN_25063; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25065 = 10'h7e == _T_375[9:0] ? 4'he : _GEN_25064; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25066 = 10'h7f == _T_375[9:0] ? 4'he : _GEN_25065; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25067 = 10'h80 == _T_375[9:0] ? 4'he : _GEN_25066; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25068 = 10'h81 == _T_375[9:0] ? 4'hb : _GEN_25067; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25069 = 10'h82 == _T_375[9:0] ? 4'hc : _GEN_25068; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25070 = 10'h83 == _T_375[9:0] ? 4'hc : _GEN_25069; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25071 = 10'h84 == _T_375[9:0] ? 4'he : _GEN_25070; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25072 = 10'h85 == _T_375[9:0] ? 4'he : _GEN_25071; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25073 = 10'h86 == _T_375[9:0] ? 4'he : _GEN_25072; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25074 = 10'h87 == _T_375[9:0] ? 4'ha : _GEN_25073; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25075 = 10'h88 == _T_375[9:0] ? 4'hd : _GEN_25074; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25076 = 10'h89 == _T_375[9:0] ? 4'hd : _GEN_25075; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25077 = 10'h8a == _T_375[9:0] ? 4'hc : _GEN_25076; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25078 = 10'h8b == _T_375[9:0] ? 4'he : _GEN_25077; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25079 = 10'h8c == _T_375[9:0] ? 4'he : _GEN_25078; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25080 = 10'h8d == _T_375[9:0] ? 4'he : _GEN_25079; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25081 = 10'h8e == _T_375[9:0] ? 4'he : _GEN_25080; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25082 = 10'h8f == _T_375[9:0] ? 4'hb : _GEN_25081; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25083 = 10'h90 == _T_375[9:0] ? 4'hc : _GEN_25082; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25084 = 10'h91 == _T_375[9:0] ? 4'hc : _GEN_25083; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25085 = 10'h92 == _T_375[9:0] ? 4'hd : _GEN_25084; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25086 = 10'h93 == _T_375[9:0] ? 4'he : _GEN_25085; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25087 = 10'h94 == _T_375[9:0] ? 4'he : _GEN_25086; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25088 = 10'h95 == _T_375[9:0] ? 4'he : _GEN_25087; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25089 = 10'h96 == _T_375[9:0] ? 4'he : _GEN_25088; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25090 = 10'h97 == _T_375[9:0] ? 4'he : _GEN_25089; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25091 = 10'h98 == _T_375[9:0] ? 4'he : _GEN_25090; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25092 = 10'h99 == _T_375[9:0] ? 4'he : _GEN_25091; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25093 = 10'h9a == _T_375[9:0] ? 4'he : _GEN_25092; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25094 = 10'h9b == _T_375[9:0] ? 4'he : _GEN_25093; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25095 = 10'h9c == _T_375[9:0] ? 4'he : _GEN_25094; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25096 = 10'h9d == _T_375[9:0] ? 4'he : _GEN_25095; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25097 = 10'h9e == _T_375[9:0] ? 4'he : _GEN_25096; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25098 = 10'h9f == _T_375[9:0] ? 4'he : _GEN_25097; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25099 = 10'ha0 == _T_375[9:0] ? 4'he : _GEN_25098; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25100 = 10'ha1 == _T_375[9:0] ? 4'he : _GEN_25099; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25101 = 10'ha2 == _T_375[9:0] ? 4'he : _GEN_25100; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25102 = 10'ha3 == _T_375[9:0] ? 4'he : _GEN_25101; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25103 = 10'ha4 == _T_375[9:0] ? 4'he : _GEN_25102; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25104 = 10'ha5 == _T_375[9:0] ? 4'he : _GEN_25103; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25105 = 10'ha6 == _T_375[9:0] ? 4'he : _GEN_25104; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25106 = 10'ha7 == _T_375[9:0] ? 4'he : _GEN_25105; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25107 = 10'ha8 == _T_375[9:0] ? 4'hb : _GEN_25106; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25108 = 10'ha9 == _T_375[9:0] ? 4'hc : _GEN_25107; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25109 = 10'haa == _T_375[9:0] ? 4'hb : _GEN_25108; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25110 = 10'hab == _T_375[9:0] ? 4'hc : _GEN_25109; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25111 = 10'hac == _T_375[9:0] ? 4'hd : _GEN_25110; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25112 = 10'had == _T_375[9:0] ? 4'ha : _GEN_25111; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25113 = 10'hae == _T_375[9:0] ? 4'hd : _GEN_25112; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25114 = 10'haf == _T_375[9:0] ? 4'hd : _GEN_25113; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25115 = 10'hb0 == _T_375[9:0] ? 4'hb : _GEN_25114; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25116 = 10'hb1 == _T_375[9:0] ? 4'hc : _GEN_25115; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25117 = 10'hb2 == _T_375[9:0] ? 4'he : _GEN_25116; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25118 = 10'hb3 == _T_375[9:0] ? 4'hb : _GEN_25117; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25119 = 10'hb4 == _T_375[9:0] ? 4'hc : _GEN_25118; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25120 = 10'hb5 == _T_375[9:0] ? 4'hd : _GEN_25119; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25121 = 10'hb6 == _T_375[9:0] ? 4'hd : _GEN_25120; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25122 = 10'hb7 == _T_375[9:0] ? 4'hc : _GEN_25121; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25123 = 10'hb8 == _T_375[9:0] ? 4'he : _GEN_25122; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25124 = 10'hb9 == _T_375[9:0] ? 4'he : _GEN_25123; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25125 = 10'hba == _T_375[9:0] ? 4'he : _GEN_25124; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25126 = 10'hbb == _T_375[9:0] ? 4'he : _GEN_25125; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25127 = 10'hbc == _T_375[9:0] ? 4'he : _GEN_25126; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25128 = 10'hbd == _T_375[9:0] ? 4'he : _GEN_25127; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25129 = 10'hbe == _T_375[9:0] ? 4'he : _GEN_25128; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25130 = 10'hbf == _T_375[9:0] ? 4'he : _GEN_25129; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25131 = 10'hc0 == _T_375[9:0] ? 4'he : _GEN_25130; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25132 = 10'hc1 == _T_375[9:0] ? 4'he : _GEN_25131; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25133 = 10'hc2 == _T_375[9:0] ? 4'he : _GEN_25132; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25134 = 10'hc3 == _T_375[9:0] ? 4'he : _GEN_25133; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25135 = 10'hc4 == _T_375[9:0] ? 4'he : _GEN_25134; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25136 = 10'hc5 == _T_375[9:0] ? 4'he : _GEN_25135; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25137 = 10'hc6 == _T_375[9:0] ? 4'he : _GEN_25136; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25138 = 10'hc7 == _T_375[9:0] ? 4'hd : _GEN_25137; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25139 = 10'hc8 == _T_375[9:0] ? 4'hb : _GEN_25138; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25140 = 10'hc9 == _T_375[9:0] ? 4'hc : _GEN_25139; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25141 = 10'hca == _T_375[9:0] ? 4'he : _GEN_25140; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25142 = 10'hcb == _T_375[9:0] ? 4'he : _GEN_25141; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25143 = 10'hcc == _T_375[9:0] ? 4'he : _GEN_25142; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25144 = 10'hcd == _T_375[9:0] ? 4'he : _GEN_25143; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25145 = 10'hce == _T_375[9:0] ? 4'hd : _GEN_25144; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25146 = 10'hcf == _T_375[9:0] ? 4'hb : _GEN_25145; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25147 = 10'hd0 == _T_375[9:0] ? 4'hc : _GEN_25146; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25148 = 10'hd1 == _T_375[9:0] ? 4'hc : _GEN_25147; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25149 = 10'hd2 == _T_375[9:0] ? 4'hb : _GEN_25148; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25150 = 10'hd3 == _T_375[9:0] ? 4'hd : _GEN_25149; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25151 = 10'hd4 == _T_375[9:0] ? 4'hd : _GEN_25150; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25152 = 10'hd5 == _T_375[9:0] ? 4'hd : _GEN_25151; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25153 = 10'hd6 == _T_375[9:0] ? 4'hd : _GEN_25152; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25154 = 10'hd7 == _T_375[9:0] ? 4'hc : _GEN_25153; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25155 = 10'hd8 == _T_375[9:0] ? 4'hc : _GEN_25154; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25156 = 10'hd9 == _T_375[9:0] ? 4'hc : _GEN_25155; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25157 = 10'hda == _T_375[9:0] ? 4'hd : _GEN_25156; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25158 = 10'hdb == _T_375[9:0] ? 4'hc : _GEN_25157; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25159 = 10'hdc == _T_375[9:0] ? 4'h9 : _GEN_25158; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25160 = 10'hdd == _T_375[9:0] ? 4'he : _GEN_25159; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25161 = 10'hde == _T_375[9:0] ? 4'he : _GEN_25160; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25162 = 10'hdf == _T_375[9:0] ? 4'he : _GEN_25161; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25163 = 10'he0 == _T_375[9:0] ? 4'he : _GEN_25162; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25164 = 10'he1 == _T_375[9:0] ? 4'he : _GEN_25163; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25165 = 10'he2 == _T_375[9:0] ? 4'he : _GEN_25164; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25166 = 10'he3 == _T_375[9:0] ? 4'h9 : _GEN_25165; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25167 = 10'he4 == _T_375[9:0] ? 4'he : _GEN_25166; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25168 = 10'he5 == _T_375[9:0] ? 4'he : _GEN_25167; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25169 = 10'he6 == _T_375[9:0] ? 4'he : _GEN_25168; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25170 = 10'he7 == _T_375[9:0] ? 4'he : _GEN_25169; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25171 = 10'he8 == _T_375[9:0] ? 4'he : _GEN_25170; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25172 = 10'he9 == _T_375[9:0] ? 4'he : _GEN_25171; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25173 = 10'hea == _T_375[9:0] ? 4'he : _GEN_25172; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25174 = 10'heb == _T_375[9:0] ? 4'hc : _GEN_25173; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25175 = 10'hec == _T_375[9:0] ? 4'h7 : _GEN_25174; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25176 = 10'hed == _T_375[9:0] ? 4'h1 : _GEN_25175; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25177 = 10'hee == _T_375[9:0] ? 4'h0 : _GEN_25176; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25178 = 10'hef == _T_375[9:0] ? 4'h0 : _GEN_25177; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25179 = 10'hf0 == _T_375[9:0] ? 4'h2 : _GEN_25178; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25180 = 10'hf1 == _T_375[9:0] ? 4'h9 : _GEN_25179; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25181 = 10'hf2 == _T_375[9:0] ? 4'he : _GEN_25180; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25182 = 10'hf3 == _T_375[9:0] ? 4'he : _GEN_25181; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25183 = 10'hf4 == _T_375[9:0] ? 4'he : _GEN_25182; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25184 = 10'hf5 == _T_375[9:0] ? 4'hc : _GEN_25183; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25185 = 10'hf6 == _T_375[9:0] ? 4'hc : _GEN_25184; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25186 = 10'hf7 == _T_375[9:0] ? 4'hd : _GEN_25185; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25187 = 10'hf8 == _T_375[9:0] ? 4'hd : _GEN_25186; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25188 = 10'hf9 == _T_375[9:0] ? 4'hd : _GEN_25187; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25189 = 10'hfa == _T_375[9:0] ? 4'hd : _GEN_25188; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25190 = 10'hfb == _T_375[9:0] ? 4'hd : _GEN_25189; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25191 = 10'hfc == _T_375[9:0] ? 4'hd : _GEN_25190; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25192 = 10'hfd == _T_375[9:0] ? 4'hd : _GEN_25191; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25193 = 10'hfe == _T_375[9:0] ? 4'hd : _GEN_25192; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25194 = 10'hff == _T_375[9:0] ? 4'hd : _GEN_25193; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25195 = 10'h100 == _T_375[9:0] ? 4'hd : _GEN_25194; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25196 = 10'h101 == _T_375[9:0] ? 4'h9 : _GEN_25195; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25197 = 10'h102 == _T_375[9:0] ? 4'h9 : _GEN_25196; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25198 = 10'h103 == _T_375[9:0] ? 4'he : _GEN_25197; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25199 = 10'h104 == _T_375[9:0] ? 4'he : _GEN_25198; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25200 = 10'h105 == _T_375[9:0] ? 4'he : _GEN_25199; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25201 = 10'h106 == _T_375[9:0] ? 4'he : _GEN_25200; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25202 = 10'h107 == _T_375[9:0] ? 4'he : _GEN_25201; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25203 = 10'h108 == _T_375[9:0] ? 4'he : _GEN_25202; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25204 = 10'h109 == _T_375[9:0] ? 4'h6 : _GEN_25203; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25205 = 10'h10a == _T_375[9:0] ? 4'he : _GEN_25204; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25206 = 10'h10b == _T_375[9:0] ? 4'he : _GEN_25205; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25207 = 10'h10c == _T_375[9:0] ? 4'he : _GEN_25206; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25208 = 10'h10d == _T_375[9:0] ? 4'he : _GEN_25207; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25209 = 10'h10e == _T_375[9:0] ? 4'he : _GEN_25208; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25210 = 10'h10f == _T_375[9:0] ? 4'ha : _GEN_25209; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25211 = 10'h110 == _T_375[9:0] ? 4'hd : _GEN_25210; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25212 = 10'h111 == _T_375[9:0] ? 4'h4 : _GEN_25211; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25213 = 10'h112 == _T_375[9:0] ? 4'h7 : _GEN_25212; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25214 = 10'h113 == _T_375[9:0] ? 4'h0 : _GEN_25213; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25215 = 10'h114 == _T_375[9:0] ? 4'h0 : _GEN_25214; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25216 = 10'h115 == _T_375[9:0] ? 4'h0 : _GEN_25215; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25217 = 10'h116 == _T_375[9:0] ? 4'h0 : _GEN_25216; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25218 = 10'h117 == _T_375[9:0] ? 4'h0 : _GEN_25217; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25219 = 10'h118 == _T_375[9:0] ? 4'ha : _GEN_25218; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25220 = 10'h119 == _T_375[9:0] ? 4'he : _GEN_25219; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25221 = 10'h11a == _T_375[9:0] ? 4'he : _GEN_25220; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25222 = 10'h11b == _T_375[9:0] ? 4'he : _GEN_25221; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25223 = 10'h11c == _T_375[9:0] ? 4'hb : _GEN_25222; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25224 = 10'h11d == _T_375[9:0] ? 4'hc : _GEN_25223; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25225 = 10'h11e == _T_375[9:0] ? 4'hd : _GEN_25224; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25226 = 10'h11f == _T_375[9:0] ? 4'hb : _GEN_25225; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25227 = 10'h120 == _T_375[9:0] ? 4'ha : _GEN_25226; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25228 = 10'h121 == _T_375[9:0] ? 4'hc : _GEN_25227; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25229 = 10'h122 == _T_375[9:0] ? 4'ha : _GEN_25228; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25230 = 10'h123 == _T_375[9:0] ? 4'ha : _GEN_25229; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25231 = 10'h124 == _T_375[9:0] ? 4'hd : _GEN_25230; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25232 = 10'h125 == _T_375[9:0] ? 4'hd : _GEN_25231; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25233 = 10'h126 == _T_375[9:0] ? 4'hb : _GEN_25232; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25234 = 10'h127 == _T_375[9:0] ? 4'h9 : _GEN_25233; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25235 = 10'h128 == _T_375[9:0] ? 4'h7 : _GEN_25234; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25236 = 10'h129 == _T_375[9:0] ? 4'hd : _GEN_25235; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25237 = 10'h12a == _T_375[9:0] ? 4'hc : _GEN_25236; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25238 = 10'h12b == _T_375[9:0] ? 4'hb : _GEN_25237; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25239 = 10'h12c == _T_375[9:0] ? 4'hc : _GEN_25238; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25240 = 10'h12d == _T_375[9:0] ? 4'hb : _GEN_25239; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25241 = 10'h12e == _T_375[9:0] ? 4'ha : _GEN_25240; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25242 = 10'h12f == _T_375[9:0] ? 4'h6 : _GEN_25241; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25243 = 10'h130 == _T_375[9:0] ? 4'he : _GEN_25242; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25244 = 10'h131 == _T_375[9:0] ? 4'hc : _GEN_25243; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25245 = 10'h132 == _T_375[9:0] ? 4'ha : _GEN_25244; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25246 = 10'h133 == _T_375[9:0] ? 4'h9 : _GEN_25245; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25247 = 10'h134 == _T_375[9:0] ? 4'hb : _GEN_25246; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25248 = 10'h135 == _T_375[9:0] ? 4'h8 : _GEN_25247; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25249 = 10'h136 == _T_375[9:0] ? 4'h8 : _GEN_25248; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25250 = 10'h137 == _T_375[9:0] ? 4'h4 : _GEN_25249; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25251 = 10'h138 == _T_375[9:0] ? 4'h7 : _GEN_25250; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25252 = 10'h139 == _T_375[9:0] ? 4'h0 : _GEN_25251; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25253 = 10'h13a == _T_375[9:0] ? 4'h0 : _GEN_25252; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25254 = 10'h13b == _T_375[9:0] ? 4'h0 : _GEN_25253; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25255 = 10'h13c == _T_375[9:0] ? 4'h0 : _GEN_25254; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25256 = 10'h13d == _T_375[9:0] ? 4'h0 : _GEN_25255; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25257 = 10'h13e == _T_375[9:0] ? 4'h4 : _GEN_25256; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25258 = 10'h13f == _T_375[9:0] ? 4'hc : _GEN_25257; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25259 = 10'h140 == _T_375[9:0] ? 4'he : _GEN_25258; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25260 = 10'h141 == _T_375[9:0] ? 4'he : _GEN_25259; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25261 = 10'h142 == _T_375[9:0] ? 4'he : _GEN_25260; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25262 = 10'h143 == _T_375[9:0] ? 4'hc : _GEN_25261; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25263 = 10'h144 == _T_375[9:0] ? 4'hd : _GEN_25262; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25264 = 10'h145 == _T_375[9:0] ? 4'hb : _GEN_25263; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25265 = 10'h146 == _T_375[9:0] ? 4'hb : _GEN_25264; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25266 = 10'h147 == _T_375[9:0] ? 4'ha : _GEN_25265; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25267 = 10'h148 == _T_375[9:0] ? 4'ha : _GEN_25266; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25268 = 10'h149 == _T_375[9:0] ? 4'hc : _GEN_25267; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25269 = 10'h14a == _T_375[9:0] ? 4'hd : _GEN_25268; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25270 = 10'h14b == _T_375[9:0] ? 4'hc : _GEN_25269; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25271 = 10'h14c == _T_375[9:0] ? 4'hd : _GEN_25270; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25272 = 10'h14d == _T_375[9:0] ? 4'h9 : _GEN_25271; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25273 = 10'h14e == _T_375[9:0] ? 4'h7 : _GEN_25272; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25274 = 10'h14f == _T_375[9:0] ? 4'ha : _GEN_25273; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25275 = 10'h150 == _T_375[9:0] ? 4'ha : _GEN_25274; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25276 = 10'h151 == _T_375[9:0] ? 4'hb : _GEN_25275; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25277 = 10'h152 == _T_375[9:0] ? 4'hb : _GEN_25276; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25278 = 10'h153 == _T_375[9:0] ? 4'hc : _GEN_25277; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25279 = 10'h154 == _T_375[9:0] ? 4'hb : _GEN_25278; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25280 = 10'h155 == _T_375[9:0] ? 4'h6 : _GEN_25279; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25281 = 10'h156 == _T_375[9:0] ? 4'hb : _GEN_25280; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25282 = 10'h157 == _T_375[9:0] ? 4'h7 : _GEN_25281; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25283 = 10'h158 == _T_375[9:0] ? 4'h7 : _GEN_25282; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25284 = 10'h159 == _T_375[9:0] ? 4'h7 : _GEN_25283; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25285 = 10'h15a == _T_375[9:0] ? 4'h7 : _GEN_25284; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25286 = 10'h15b == _T_375[9:0] ? 4'h7 : _GEN_25285; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25287 = 10'h15c == _T_375[9:0] ? 4'h7 : _GEN_25286; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25288 = 10'h15d == _T_375[9:0] ? 4'h6 : _GEN_25287; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25289 = 10'h15e == _T_375[9:0] ? 4'h7 : _GEN_25288; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25290 = 10'h15f == _T_375[9:0] ? 4'h0 : _GEN_25289; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25291 = 10'h160 == _T_375[9:0] ? 4'h0 : _GEN_25290; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25292 = 10'h161 == _T_375[9:0] ? 4'h0 : _GEN_25291; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25293 = 10'h162 == _T_375[9:0] ? 4'h0 : _GEN_25292; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25294 = 10'h163 == _T_375[9:0] ? 4'h2 : _GEN_25293; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25295 = 10'h164 == _T_375[9:0] ? 4'h4 : _GEN_25294; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25296 = 10'h165 == _T_375[9:0] ? 4'hb : _GEN_25295; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25297 = 10'h166 == _T_375[9:0] ? 4'hb : _GEN_25296; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25298 = 10'h167 == _T_375[9:0] ? 4'he : _GEN_25297; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25299 = 10'h168 == _T_375[9:0] ? 4'he : _GEN_25298; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25300 = 10'h169 == _T_375[9:0] ? 4'hc : _GEN_25299; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25301 = 10'h16a == _T_375[9:0] ? 4'hd : _GEN_25300; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25302 = 10'h16b == _T_375[9:0] ? 4'hd : _GEN_25301; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25303 = 10'h16c == _T_375[9:0] ? 4'ha : _GEN_25302; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25304 = 10'h16d == _T_375[9:0] ? 4'ha : _GEN_25303; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25305 = 10'h16e == _T_375[9:0] ? 4'ha : _GEN_25304; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25306 = 10'h16f == _T_375[9:0] ? 4'hd : _GEN_25305; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25307 = 10'h170 == _T_375[9:0] ? 4'hd : _GEN_25306; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25308 = 10'h171 == _T_375[9:0] ? 4'hd : _GEN_25307; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25309 = 10'h172 == _T_375[9:0] ? 4'he : _GEN_25308; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25310 = 10'h173 == _T_375[9:0] ? 4'h8 : _GEN_25309; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25311 = 10'h174 == _T_375[9:0] ? 4'h5 : _GEN_25310; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25312 = 10'h175 == _T_375[9:0] ? 4'h6 : _GEN_25311; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25313 = 10'h176 == _T_375[9:0] ? 4'h6 : _GEN_25312; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25314 = 10'h177 == _T_375[9:0] ? 4'h6 : _GEN_25313; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25315 = 10'h178 == _T_375[9:0] ? 4'h7 : _GEN_25314; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25316 = 10'h179 == _T_375[9:0] ? 4'h9 : _GEN_25315; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25317 = 10'h17a == _T_375[9:0] ? 4'h9 : _GEN_25316; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25318 = 10'h17b == _T_375[9:0] ? 4'h6 : _GEN_25317; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25319 = 10'h17c == _T_375[9:0] ? 4'h7 : _GEN_25318; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25320 = 10'h17d == _T_375[9:0] ? 4'h7 : _GEN_25319; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25321 = 10'h17e == _T_375[9:0] ? 4'h7 : _GEN_25320; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25322 = 10'h17f == _T_375[9:0] ? 4'h7 : _GEN_25321; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25323 = 10'h180 == _T_375[9:0] ? 4'h7 : _GEN_25322; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25324 = 10'h181 == _T_375[9:0] ? 4'h7 : _GEN_25323; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25325 = 10'h182 == _T_375[9:0] ? 4'h8 : _GEN_25324; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25326 = 10'h183 == _T_375[9:0] ? 4'h8 : _GEN_25325; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25327 = 10'h184 == _T_375[9:0] ? 4'h8 : _GEN_25326; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25328 = 10'h185 == _T_375[9:0] ? 4'h7 : _GEN_25327; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25329 = 10'h186 == _T_375[9:0] ? 4'h1 : _GEN_25328; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25330 = 10'h187 == _T_375[9:0] ? 4'h0 : _GEN_25329; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25331 = 10'h188 == _T_375[9:0] ? 4'h0 : _GEN_25330; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25332 = 10'h189 == _T_375[9:0] ? 4'h4 : _GEN_25331; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25333 = 10'h18a == _T_375[9:0] ? 4'h4 : _GEN_25332; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25334 = 10'h18b == _T_375[9:0] ? 4'hb : _GEN_25333; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25335 = 10'h18c == _T_375[9:0] ? 4'hb : _GEN_25334; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25336 = 10'h18d == _T_375[9:0] ? 4'hc : _GEN_25335; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25337 = 10'h18e == _T_375[9:0] ? 4'he : _GEN_25336; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25338 = 10'h18f == _T_375[9:0] ? 4'hb : _GEN_25337; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25339 = 10'h190 == _T_375[9:0] ? 4'hd : _GEN_25338; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25340 = 10'h191 == _T_375[9:0] ? 4'hc : _GEN_25339; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25341 = 10'h192 == _T_375[9:0] ? 4'h9 : _GEN_25340; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25342 = 10'h193 == _T_375[9:0] ? 4'ha : _GEN_25341; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25343 = 10'h194 == _T_375[9:0] ? 4'h9 : _GEN_25342; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25344 = 10'h195 == _T_375[9:0] ? 4'hd : _GEN_25343; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25345 = 10'h196 == _T_375[9:0] ? 4'hd : _GEN_25344; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25346 = 10'h197 == _T_375[9:0] ? 4'hb : _GEN_25345; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25347 = 10'h198 == _T_375[9:0] ? 4'he : _GEN_25346; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25348 = 10'h199 == _T_375[9:0] ? 4'h5 : _GEN_25347; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25349 = 10'h19a == _T_375[9:0] ? 4'h1 : _GEN_25348; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25350 = 10'h19b == _T_375[9:0] ? 4'h3 : _GEN_25349; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25351 = 10'h19c == _T_375[9:0] ? 4'h6 : _GEN_25350; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25352 = 10'h19d == _T_375[9:0] ? 4'h4 : _GEN_25351; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25353 = 10'h19e == _T_375[9:0] ? 4'h1 : _GEN_25352; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25354 = 10'h19f == _T_375[9:0] ? 4'h3 : _GEN_25353; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25355 = 10'h1a0 == _T_375[9:0] ? 4'h6 : _GEN_25354; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25356 = 10'h1a1 == _T_375[9:0] ? 4'h6 : _GEN_25355; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25357 = 10'h1a2 == _T_375[9:0] ? 4'h7 : _GEN_25356; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25358 = 10'h1a3 == _T_375[9:0] ? 4'h7 : _GEN_25357; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25359 = 10'h1a4 == _T_375[9:0] ? 4'h7 : _GEN_25358; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25360 = 10'h1a5 == _T_375[9:0] ? 4'h7 : _GEN_25359; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25361 = 10'h1a6 == _T_375[9:0] ? 4'h7 : _GEN_25360; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25362 = 10'h1a7 == _T_375[9:0] ? 4'h7 : _GEN_25361; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25363 = 10'h1a8 == _T_375[9:0] ? 4'h8 : _GEN_25362; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25364 = 10'h1a9 == _T_375[9:0] ? 4'h8 : _GEN_25363; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25365 = 10'h1aa == _T_375[9:0] ? 4'h7 : _GEN_25364; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25366 = 10'h1ab == _T_375[9:0] ? 4'h8 : _GEN_25365; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25367 = 10'h1ac == _T_375[9:0] ? 4'h8 : _GEN_25366; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25368 = 10'h1ad == _T_375[9:0] ? 4'h3 : _GEN_25367; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25369 = 10'h1ae == _T_375[9:0] ? 4'h2 : _GEN_25368; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25370 = 10'h1af == _T_375[9:0] ? 4'h8 : _GEN_25369; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25371 = 10'h1b0 == _T_375[9:0] ? 4'h6 : _GEN_25370; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25372 = 10'h1b1 == _T_375[9:0] ? 4'hb : _GEN_25371; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25373 = 10'h1b2 == _T_375[9:0] ? 4'hb : _GEN_25372; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25374 = 10'h1b3 == _T_375[9:0] ? 4'ha : _GEN_25373; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25375 = 10'h1b4 == _T_375[9:0] ? 4'he : _GEN_25374; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25376 = 10'h1b5 == _T_375[9:0] ? 4'hb : _GEN_25375; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25377 = 10'h1b6 == _T_375[9:0] ? 4'hc : _GEN_25376; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25378 = 10'h1b7 == _T_375[9:0] ? 4'ha : _GEN_25377; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25379 = 10'h1b8 == _T_375[9:0] ? 4'h9 : _GEN_25378; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25380 = 10'h1b9 == _T_375[9:0] ? 4'h9 : _GEN_25379; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25381 = 10'h1ba == _T_375[9:0] ? 4'h9 : _GEN_25380; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25382 = 10'h1bb == _T_375[9:0] ? 4'hb : _GEN_25381; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25383 = 10'h1bc == _T_375[9:0] ? 4'hd : _GEN_25382; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25384 = 10'h1bd == _T_375[9:0] ? 4'hd : _GEN_25383; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25385 = 10'h1be == _T_375[9:0] ? 4'he : _GEN_25384; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25386 = 10'h1bf == _T_375[9:0] ? 4'h7 : _GEN_25385; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25387 = 10'h1c0 == _T_375[9:0] ? 4'h6 : _GEN_25386; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25388 = 10'h1c1 == _T_375[9:0] ? 4'h6 : _GEN_25387; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25389 = 10'h1c2 == _T_375[9:0] ? 4'h5 : _GEN_25388; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25390 = 10'h1c3 == _T_375[9:0] ? 4'h5 : _GEN_25389; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25391 = 10'h1c4 == _T_375[9:0] ? 4'h4 : _GEN_25390; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25392 = 10'h1c5 == _T_375[9:0] ? 4'h5 : _GEN_25391; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25393 = 10'h1c6 == _T_375[9:0] ? 4'h6 : _GEN_25392; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25394 = 10'h1c7 == _T_375[9:0] ? 4'h6 : _GEN_25393; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25395 = 10'h1c8 == _T_375[9:0] ? 4'h7 : _GEN_25394; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25396 = 10'h1c9 == _T_375[9:0] ? 4'h7 : _GEN_25395; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25397 = 10'h1ca == _T_375[9:0] ? 4'h7 : _GEN_25396; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25398 = 10'h1cb == _T_375[9:0] ? 4'h7 : _GEN_25397; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25399 = 10'h1cc == _T_375[9:0] ? 4'h7 : _GEN_25398; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25400 = 10'h1cd == _T_375[9:0] ? 4'h8 : _GEN_25399; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25401 = 10'h1ce == _T_375[9:0] ? 4'h8 : _GEN_25400; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25402 = 10'h1cf == _T_375[9:0] ? 4'h8 : _GEN_25401; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25403 = 10'h1d0 == _T_375[9:0] ? 4'h5 : _GEN_25402; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25404 = 10'h1d1 == _T_375[9:0] ? 4'h8 : _GEN_25403; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25405 = 10'h1d2 == _T_375[9:0] ? 4'h8 : _GEN_25404; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25406 = 10'h1d3 == _T_375[9:0] ? 4'h8 : _GEN_25405; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25407 = 10'h1d4 == _T_375[9:0] ? 4'h8 : _GEN_25406; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25408 = 10'h1d5 == _T_375[9:0] ? 4'h7 : _GEN_25407; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25409 = 10'h1d6 == _T_375[9:0] ? 4'h9 : _GEN_25408; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25410 = 10'h1d7 == _T_375[9:0] ? 4'hb : _GEN_25409; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25411 = 10'h1d8 == _T_375[9:0] ? 4'hb : _GEN_25410; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25412 = 10'h1d9 == _T_375[9:0] ? 4'hb : _GEN_25411; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25413 = 10'h1da == _T_375[9:0] ? 4'ha : _GEN_25412; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25414 = 10'h1db == _T_375[9:0] ? 4'hc : _GEN_25413; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25415 = 10'h1dc == _T_375[9:0] ? 4'hb : _GEN_25414; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25416 = 10'h1dd == _T_375[9:0] ? 4'h5 : _GEN_25415; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25417 = 10'h1de == _T_375[9:0] ? 4'h9 : _GEN_25416; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25418 = 10'h1df == _T_375[9:0] ? 4'h9 : _GEN_25417; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25419 = 10'h1e0 == _T_375[9:0] ? 4'h9 : _GEN_25418; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25420 = 10'h1e1 == _T_375[9:0] ? 4'h7 : _GEN_25419; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25421 = 10'h1e2 == _T_375[9:0] ? 4'hc : _GEN_25420; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25422 = 10'h1e3 == _T_375[9:0] ? 4'hc : _GEN_25421; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25423 = 10'h1e4 == _T_375[9:0] ? 4'hd : _GEN_25422; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25424 = 10'h1e5 == _T_375[9:0] ? 4'h7 : _GEN_25423; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25425 = 10'h1e6 == _T_375[9:0] ? 4'h6 : _GEN_25424; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25426 = 10'h1e7 == _T_375[9:0] ? 4'h6 : _GEN_25425; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25427 = 10'h1e8 == _T_375[9:0] ? 4'h6 : _GEN_25426; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25428 = 10'h1e9 == _T_375[9:0] ? 4'h6 : _GEN_25427; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25429 = 10'h1ea == _T_375[9:0] ? 4'h6 : _GEN_25428; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25430 = 10'h1eb == _T_375[9:0] ? 4'h6 : _GEN_25429; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25431 = 10'h1ec == _T_375[9:0] ? 4'h6 : _GEN_25430; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25432 = 10'h1ed == _T_375[9:0] ? 4'h8 : _GEN_25431; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25433 = 10'h1ee == _T_375[9:0] ? 4'h7 : _GEN_25432; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25434 = 10'h1ef == _T_375[9:0] ? 4'h7 : _GEN_25433; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25435 = 10'h1f0 == _T_375[9:0] ? 4'h7 : _GEN_25434; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25436 = 10'h1f1 == _T_375[9:0] ? 4'h7 : _GEN_25435; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25437 = 10'h1f2 == _T_375[9:0] ? 4'h7 : _GEN_25436; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25438 = 10'h1f3 == _T_375[9:0] ? 4'h8 : _GEN_25437; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25439 = 10'h1f4 == _T_375[9:0] ? 4'h8 : _GEN_25438; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25440 = 10'h1f5 == _T_375[9:0] ? 4'h8 : _GEN_25439; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25441 = 10'h1f6 == _T_375[9:0] ? 4'ha : _GEN_25440; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25442 = 10'h1f7 == _T_375[9:0] ? 4'h8 : _GEN_25441; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25443 = 10'h1f8 == _T_375[9:0] ? 4'h8 : _GEN_25442; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25444 = 10'h1f9 == _T_375[9:0] ? 4'h9 : _GEN_25443; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25445 = 10'h1fa == _T_375[9:0] ? 4'h9 : _GEN_25444; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25446 = 10'h1fb == _T_375[9:0] ? 4'h8 : _GEN_25445; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25447 = 10'h1fc == _T_375[9:0] ? 4'hb : _GEN_25446; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25448 = 10'h1fd == _T_375[9:0] ? 4'hb : _GEN_25447; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25449 = 10'h1fe == _T_375[9:0] ? 4'hb : _GEN_25448; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25450 = 10'h1ff == _T_375[9:0] ? 4'ha : _GEN_25449; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25451 = 10'h200 == _T_375[9:0] ? 4'h3 : _GEN_25450; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25452 = 10'h201 == _T_375[9:0] ? 4'h9 : _GEN_25451; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25453 = 10'h202 == _T_375[9:0] ? 4'h5 : _GEN_25452; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25454 = 10'h203 == _T_375[9:0] ? 4'h3 : _GEN_25453; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25455 = 10'h204 == _T_375[9:0] ? 4'h4 : _GEN_25454; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25456 = 10'h205 == _T_375[9:0] ? 4'h4 : _GEN_25455; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25457 = 10'h206 == _T_375[9:0] ? 4'h4 : _GEN_25456; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25458 = 10'h207 == _T_375[9:0] ? 4'h4 : _GEN_25457; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25459 = 10'h208 == _T_375[9:0] ? 4'h8 : _GEN_25458; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25460 = 10'h209 == _T_375[9:0] ? 4'hc : _GEN_25459; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25461 = 10'h20a == _T_375[9:0] ? 4'hd : _GEN_25460; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25462 = 10'h20b == _T_375[9:0] ? 4'h7 : _GEN_25461; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25463 = 10'h20c == _T_375[9:0] ? 4'h6 : _GEN_25462; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25464 = 10'h20d == _T_375[9:0] ? 4'h6 : _GEN_25463; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25465 = 10'h20e == _T_375[9:0] ? 4'h6 : _GEN_25464; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25466 = 10'h20f == _T_375[9:0] ? 4'h5 : _GEN_25465; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25467 = 10'h210 == _T_375[9:0] ? 4'h6 : _GEN_25466; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25468 = 10'h211 == _T_375[9:0] ? 4'h6 : _GEN_25467; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25469 = 10'h212 == _T_375[9:0] ? 4'h7 : _GEN_25468; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25470 = 10'h213 == _T_375[9:0] ? 4'ha : _GEN_25469; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25471 = 10'h214 == _T_375[9:0] ? 4'h6 : _GEN_25470; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25472 = 10'h215 == _T_375[9:0] ? 4'h7 : _GEN_25471; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25473 = 10'h216 == _T_375[9:0] ? 4'h7 : _GEN_25472; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25474 = 10'h217 == _T_375[9:0] ? 4'h7 : _GEN_25473; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25475 = 10'h218 == _T_375[9:0] ? 4'h7 : _GEN_25474; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25476 = 10'h219 == _T_375[9:0] ? 4'h8 : _GEN_25475; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25477 = 10'h21a == _T_375[9:0] ? 4'h7 : _GEN_25476; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25478 = 10'h21b == _T_375[9:0] ? 4'h8 : _GEN_25477; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25479 = 10'h21c == _T_375[9:0] ? 4'hb : _GEN_25478; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25480 = 10'h21d == _T_375[9:0] ? 4'ha : _GEN_25479; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25481 = 10'h21e == _T_375[9:0] ? 4'h9 : _GEN_25480; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25482 = 10'h21f == _T_375[9:0] ? 4'h9 : _GEN_25481; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25483 = 10'h220 == _T_375[9:0] ? 4'h8 : _GEN_25482; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25484 = 10'h221 == _T_375[9:0] ? 4'h9 : _GEN_25483; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25485 = 10'h222 == _T_375[9:0] ? 4'hb : _GEN_25484; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25486 = 10'h223 == _T_375[9:0] ? 4'hb : _GEN_25485; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25487 = 10'h224 == _T_375[9:0] ? 4'hb : _GEN_25486; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25488 = 10'h225 == _T_375[9:0] ? 4'h8 : _GEN_25487; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25489 = 10'h226 == _T_375[9:0] ? 4'h1 : _GEN_25488; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25490 = 10'h227 == _T_375[9:0] ? 4'h3 : _GEN_25489; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25491 = 10'h228 == _T_375[9:0] ? 4'h3 : _GEN_25490; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25492 = 10'h229 == _T_375[9:0] ? 4'h3 : _GEN_25491; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25493 = 10'h22a == _T_375[9:0] ? 4'h3 : _GEN_25492; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25494 = 10'h22b == _T_375[9:0] ? 4'h3 : _GEN_25493; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25495 = 10'h22c == _T_375[9:0] ? 4'h3 : _GEN_25494; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25496 = 10'h22d == _T_375[9:0] ? 4'h3 : _GEN_25495; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25497 = 10'h22e == _T_375[9:0] ? 4'h3 : _GEN_25496; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25498 = 10'h22f == _T_375[9:0] ? 4'h9 : _GEN_25497; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25499 = 10'h230 == _T_375[9:0] ? 4'h6 : _GEN_25498; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25500 = 10'h231 == _T_375[9:0] ? 4'h7 : _GEN_25499; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25501 = 10'h232 == _T_375[9:0] ? 4'h6 : _GEN_25500; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25502 = 10'h233 == _T_375[9:0] ? 4'h7 : _GEN_25501; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25503 = 10'h234 == _T_375[9:0] ? 4'h7 : _GEN_25502; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25504 = 10'h235 == _T_375[9:0] ? 4'h6 : _GEN_25503; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25505 = 10'h236 == _T_375[9:0] ? 4'h6 : _GEN_25504; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25506 = 10'h237 == _T_375[9:0] ? 4'h6 : _GEN_25505; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25507 = 10'h238 == _T_375[9:0] ? 4'h6 : _GEN_25506; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25508 = 10'h239 == _T_375[9:0] ? 4'h8 : _GEN_25507; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25509 = 10'h23a == _T_375[9:0] ? 4'h6 : _GEN_25508; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25510 = 10'h23b == _T_375[9:0] ? 4'h7 : _GEN_25509; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25511 = 10'h23c == _T_375[9:0] ? 4'h7 : _GEN_25510; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25512 = 10'h23d == _T_375[9:0] ? 4'h7 : _GEN_25511; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25513 = 10'h23e == _T_375[9:0] ? 4'h7 : _GEN_25512; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25514 = 10'h23f == _T_375[9:0] ? 4'h7 : _GEN_25513; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25515 = 10'h240 == _T_375[9:0] ? 4'h7 : _GEN_25514; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25516 = 10'h241 == _T_375[9:0] ? 4'h8 : _GEN_25515; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25517 = 10'h242 == _T_375[9:0] ? 4'hb : _GEN_25516; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25518 = 10'h243 == _T_375[9:0] ? 4'hb : _GEN_25517; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25519 = 10'h244 == _T_375[9:0] ? 4'hb : _GEN_25518; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25520 = 10'h245 == _T_375[9:0] ? 4'ha : _GEN_25519; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25521 = 10'h246 == _T_375[9:0] ? 4'h9 : _GEN_25520; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25522 = 10'h247 == _T_375[9:0] ? 4'ha : _GEN_25521; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25523 = 10'h248 == _T_375[9:0] ? 4'hb : _GEN_25522; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25524 = 10'h249 == _T_375[9:0] ? 4'hb : _GEN_25523; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25525 = 10'h24a == _T_375[9:0] ? 4'ha : _GEN_25524; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25526 = 10'h24b == _T_375[9:0] ? 4'h2 : _GEN_25525; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25527 = 10'h24c == _T_375[9:0] ? 4'h0 : _GEN_25526; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25528 = 10'h24d == _T_375[9:0] ? 4'h2 : _GEN_25527; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25529 = 10'h24e == _T_375[9:0] ? 4'h3 : _GEN_25528; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25530 = 10'h24f == _T_375[9:0] ? 4'h3 : _GEN_25529; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25531 = 10'h250 == _T_375[9:0] ? 4'h3 : _GEN_25530; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25532 = 10'h251 == _T_375[9:0] ? 4'h3 : _GEN_25531; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25533 = 10'h252 == _T_375[9:0] ? 4'h3 : _GEN_25532; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25534 = 10'h253 == _T_375[9:0] ? 4'h3 : _GEN_25533; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25535 = 10'h254 == _T_375[9:0] ? 4'h3 : _GEN_25534; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25536 = 10'h255 == _T_375[9:0] ? 4'h5 : _GEN_25535; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25537 = 10'h256 == _T_375[9:0] ? 4'h6 : _GEN_25536; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25538 = 10'h257 == _T_375[9:0] ? 4'h8 : _GEN_25537; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25539 = 10'h258 == _T_375[9:0] ? 4'h5 : _GEN_25538; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25540 = 10'h259 == _T_375[9:0] ? 4'h6 : _GEN_25539; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25541 = 10'h25a == _T_375[9:0] ? 4'h6 : _GEN_25540; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25542 = 10'h25b == _T_375[9:0] ? 4'h5 : _GEN_25541; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25543 = 10'h25c == _T_375[9:0] ? 4'h6 : _GEN_25542; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25544 = 10'h25d == _T_375[9:0] ? 4'h6 : _GEN_25543; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25545 = 10'h25e == _T_375[9:0] ? 4'h9 : _GEN_25544; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25546 = 10'h25f == _T_375[9:0] ? 4'hc : _GEN_25545; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25547 = 10'h260 == _T_375[9:0] ? 4'h7 : _GEN_25546; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25548 = 10'h261 == _T_375[9:0] ? 4'h9 : _GEN_25547; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25549 = 10'h262 == _T_375[9:0] ? 4'ha : _GEN_25548; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25550 = 10'h263 == _T_375[9:0] ? 4'h8 : _GEN_25549; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25551 = 10'h264 == _T_375[9:0] ? 4'ha : _GEN_25550; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25552 = 10'h265 == _T_375[9:0] ? 4'h9 : _GEN_25551; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25553 = 10'h266 == _T_375[9:0] ? 4'h8 : _GEN_25552; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25554 = 10'h267 == _T_375[9:0] ? 4'h8 : _GEN_25553; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25555 = 10'h268 == _T_375[9:0] ? 4'ha : _GEN_25554; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25556 = 10'h269 == _T_375[9:0] ? 4'ha : _GEN_25555; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25557 = 10'h26a == _T_375[9:0] ? 4'hb : _GEN_25556; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25558 = 10'h26b == _T_375[9:0] ? 4'hb : _GEN_25557; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25559 = 10'h26c == _T_375[9:0] ? 4'hb : _GEN_25558; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25560 = 10'h26d == _T_375[9:0] ? 4'hb : _GEN_25559; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25561 = 10'h26e == _T_375[9:0] ? 4'hb : _GEN_25560; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25562 = 10'h26f == _T_375[9:0] ? 4'ha : _GEN_25561; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25563 = 10'h270 == _T_375[9:0] ? 4'h3 : _GEN_25562; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25564 = 10'h271 == _T_375[9:0] ? 4'h0 : _GEN_25563; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25565 = 10'h272 == _T_375[9:0] ? 4'h0 : _GEN_25564; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25566 = 10'h273 == _T_375[9:0] ? 4'h2 : _GEN_25565; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25567 = 10'h274 == _T_375[9:0] ? 4'h3 : _GEN_25566; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25568 = 10'h275 == _T_375[9:0] ? 4'h3 : _GEN_25567; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25569 = 10'h276 == _T_375[9:0] ? 4'h3 : _GEN_25568; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25570 = 10'h277 == _T_375[9:0] ? 4'h3 : _GEN_25569; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25571 = 10'h278 == _T_375[9:0] ? 4'h3 : _GEN_25570; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25572 = 10'h279 == _T_375[9:0] ? 4'h3 : _GEN_25571; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25573 = 10'h27a == _T_375[9:0] ? 4'h3 : _GEN_25572; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25574 = 10'h27b == _T_375[9:0] ? 4'h6 : _GEN_25573; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25575 = 10'h27c == _T_375[9:0] ? 4'h7 : _GEN_25574; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25576 = 10'h27d == _T_375[9:0] ? 4'h7 : _GEN_25575; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25577 = 10'h27e == _T_375[9:0] ? 4'h4 : _GEN_25576; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25578 = 10'h27f == _T_375[9:0] ? 4'h6 : _GEN_25577; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25579 = 10'h280 == _T_375[9:0] ? 4'h6 : _GEN_25578; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25580 = 10'h281 == _T_375[9:0] ? 4'h6 : _GEN_25579; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25581 = 10'h282 == _T_375[9:0] ? 4'h6 : _GEN_25580; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25582 = 10'h283 == _T_375[9:0] ? 4'ha : _GEN_25581; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25583 = 10'h284 == _T_375[9:0] ? 4'hc : _GEN_25582; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25584 = 10'h285 == _T_375[9:0] ? 4'hc : _GEN_25583; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25585 = 10'h286 == _T_375[9:0] ? 4'h8 : _GEN_25584; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25586 = 10'h287 == _T_375[9:0] ? 4'ha : _GEN_25585; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25587 = 10'h288 == _T_375[9:0] ? 4'ha : _GEN_25586; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25588 = 10'h289 == _T_375[9:0] ? 4'ha : _GEN_25587; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25589 = 10'h28a == _T_375[9:0] ? 4'hc : _GEN_25588; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25590 = 10'h28b == _T_375[9:0] ? 4'hb : _GEN_25589; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25591 = 10'h28c == _T_375[9:0] ? 4'ha : _GEN_25590; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25592 = 10'h28d == _T_375[9:0] ? 4'h7 : _GEN_25591; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25593 = 10'h28e == _T_375[9:0] ? 4'h2 : _GEN_25592; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25594 = 10'h28f == _T_375[9:0] ? 4'h5 : _GEN_25593; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25595 = 10'h290 == _T_375[9:0] ? 4'h8 : _GEN_25594; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25596 = 10'h291 == _T_375[9:0] ? 4'ha : _GEN_25595; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25597 = 10'h292 == _T_375[9:0] ? 4'ha : _GEN_25596; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25598 = 10'h293 == _T_375[9:0] ? 4'ha : _GEN_25597; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25599 = 10'h294 == _T_375[9:0] ? 4'h9 : _GEN_25598; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25600 = 10'h295 == _T_375[9:0] ? 4'h3 : _GEN_25599; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25601 = 10'h296 == _T_375[9:0] ? 4'h0 : _GEN_25600; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25602 = 10'h297 == _T_375[9:0] ? 4'h0 : _GEN_25601; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25603 = 10'h298 == _T_375[9:0] ? 4'h0 : _GEN_25602; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25604 = 10'h299 == _T_375[9:0] ? 4'h1 : _GEN_25603; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25605 = 10'h29a == _T_375[9:0] ? 4'h3 : _GEN_25604; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25606 = 10'h29b == _T_375[9:0] ? 4'h3 : _GEN_25605; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25607 = 10'h29c == _T_375[9:0] ? 4'h3 : _GEN_25606; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25608 = 10'h29d == _T_375[9:0] ? 4'h3 : _GEN_25607; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25609 = 10'h29e == _T_375[9:0] ? 4'h3 : _GEN_25608; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25610 = 10'h29f == _T_375[9:0] ? 4'h3 : _GEN_25609; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25611 = 10'h2a0 == _T_375[9:0] ? 4'h4 : _GEN_25610; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25612 = 10'h2a1 == _T_375[9:0] ? 4'h6 : _GEN_25611; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25613 = 10'h2a2 == _T_375[9:0] ? 4'h7 : _GEN_25612; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25614 = 10'h2a3 == _T_375[9:0] ? 4'h6 : _GEN_25613; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25615 = 10'h2a4 == _T_375[9:0] ? 4'h4 : _GEN_25614; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25616 = 10'h2a5 == _T_375[9:0] ? 4'h6 : _GEN_25615; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25617 = 10'h2a6 == _T_375[9:0] ? 4'h6 : _GEN_25616; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25618 = 10'h2a7 == _T_375[9:0] ? 4'h7 : _GEN_25617; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25619 = 10'h2a8 == _T_375[9:0] ? 4'ha : _GEN_25618; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25620 = 10'h2a9 == _T_375[9:0] ? 4'hb : _GEN_25619; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25621 = 10'h2aa == _T_375[9:0] ? 4'hb : _GEN_25620; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25622 = 10'h2ab == _T_375[9:0] ? 4'hb : _GEN_25621; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25623 = 10'h2ac == _T_375[9:0] ? 4'h8 : _GEN_25622; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25624 = 10'h2ad == _T_375[9:0] ? 4'hb : _GEN_25623; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25625 = 10'h2ae == _T_375[9:0] ? 4'ha : _GEN_25624; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25626 = 10'h2af == _T_375[9:0] ? 4'hb : _GEN_25625; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25627 = 10'h2b0 == _T_375[9:0] ? 4'hc : _GEN_25626; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25628 = 10'h2b1 == _T_375[9:0] ? 4'hb : _GEN_25627; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25629 = 10'h2b2 == _T_375[9:0] ? 4'ha : _GEN_25628; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25630 = 10'h2b3 == _T_375[9:0] ? 4'h6 : _GEN_25629; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25631 = 10'h2b4 == _T_375[9:0] ? 4'h0 : _GEN_25630; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25632 = 10'h2b5 == _T_375[9:0] ? 4'h0 : _GEN_25631; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25633 = 10'h2b6 == _T_375[9:0] ? 4'h0 : _GEN_25632; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25634 = 10'h2b7 == _T_375[9:0] ? 4'h1 : _GEN_25633; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25635 = 10'h2b8 == _T_375[9:0] ? 4'h5 : _GEN_25634; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25636 = 10'h2b9 == _T_375[9:0] ? 4'h9 : _GEN_25635; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25637 = 10'h2ba == _T_375[9:0] ? 4'h1 : _GEN_25636; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25638 = 10'h2bb == _T_375[9:0] ? 4'h0 : _GEN_25637; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25639 = 10'h2bc == _T_375[9:0] ? 4'h0 : _GEN_25638; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25640 = 10'h2bd == _T_375[9:0] ? 4'h0 : _GEN_25639; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25641 = 10'h2be == _T_375[9:0] ? 4'h0 : _GEN_25640; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25642 = 10'h2bf == _T_375[9:0] ? 4'h0 : _GEN_25641; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25643 = 10'h2c0 == _T_375[9:0] ? 4'h3 : _GEN_25642; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25644 = 10'h2c1 == _T_375[9:0] ? 4'h3 : _GEN_25643; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25645 = 10'h2c2 == _T_375[9:0] ? 4'h3 : _GEN_25644; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25646 = 10'h2c3 == _T_375[9:0] ? 4'h3 : _GEN_25645; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25647 = 10'h2c4 == _T_375[9:0] ? 4'h3 : _GEN_25646; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25648 = 10'h2c5 == _T_375[9:0] ? 4'h3 : _GEN_25647; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25649 = 10'h2c6 == _T_375[9:0] ? 4'h4 : _GEN_25648; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25650 = 10'h2c7 == _T_375[9:0] ? 4'h5 : _GEN_25649; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25651 = 10'h2c8 == _T_375[9:0] ? 4'h7 : _GEN_25650; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25652 = 10'h2c9 == _T_375[9:0] ? 4'h7 : _GEN_25651; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25653 = 10'h2ca == _T_375[9:0] ? 4'h4 : _GEN_25652; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25654 = 10'h2cb == _T_375[9:0] ? 4'h9 : _GEN_25653; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25655 = 10'h2cc == _T_375[9:0] ? 4'h9 : _GEN_25654; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25656 = 10'h2cd == _T_375[9:0] ? 4'hb : _GEN_25655; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25657 = 10'h2ce == _T_375[9:0] ? 4'hb : _GEN_25656; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25658 = 10'h2cf == _T_375[9:0] ? 4'hb : _GEN_25657; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25659 = 10'h2d0 == _T_375[9:0] ? 4'hb : _GEN_25658; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25660 = 10'h2d1 == _T_375[9:0] ? 4'hb : _GEN_25659; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25661 = 10'h2d2 == _T_375[9:0] ? 4'h8 : _GEN_25660; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25662 = 10'h2d3 == _T_375[9:0] ? 4'ha : _GEN_25661; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25663 = 10'h2d4 == _T_375[9:0] ? 4'hb : _GEN_25662; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25664 = 10'h2d5 == _T_375[9:0] ? 4'ha : _GEN_25663; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25665 = 10'h2d6 == _T_375[9:0] ? 4'ha : _GEN_25664; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25666 = 10'h2d7 == _T_375[9:0] ? 4'ha : _GEN_25665; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25667 = 10'h2d8 == _T_375[9:0] ? 4'ha : _GEN_25666; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25668 = 10'h2d9 == _T_375[9:0] ? 4'h7 : _GEN_25667; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25669 = 10'h2da == _T_375[9:0] ? 4'h2 : _GEN_25668; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25670 = 10'h2db == _T_375[9:0] ? 4'h0 : _GEN_25669; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25671 = 10'h2dc == _T_375[9:0] ? 4'h0 : _GEN_25670; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25672 = 10'h2dd == _T_375[9:0] ? 4'h0 : _GEN_25671; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25673 = 10'h2de == _T_375[9:0] ? 4'h0 : _GEN_25672; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25674 = 10'h2df == _T_375[9:0] ? 4'h2 : _GEN_25673; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25675 = 10'h2e0 == _T_375[9:0] ? 4'h0 : _GEN_25674; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25676 = 10'h2e1 == _T_375[9:0] ? 4'h0 : _GEN_25675; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25677 = 10'h2e2 == _T_375[9:0] ? 4'h0 : _GEN_25676; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25678 = 10'h2e3 == _T_375[9:0] ? 4'h0 : _GEN_25677; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25679 = 10'h2e4 == _T_375[9:0] ? 4'h0 : _GEN_25678; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25680 = 10'h2e5 == _T_375[9:0] ? 4'h0 : _GEN_25679; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25681 = 10'h2e6 == _T_375[9:0] ? 4'h2 : _GEN_25680; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25682 = 10'h2e7 == _T_375[9:0] ? 4'h3 : _GEN_25681; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25683 = 10'h2e8 == _T_375[9:0] ? 4'h3 : _GEN_25682; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25684 = 10'h2e9 == _T_375[9:0] ? 4'h3 : _GEN_25683; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25685 = 10'h2ea == _T_375[9:0] ? 4'h3 : _GEN_25684; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25686 = 10'h2eb == _T_375[9:0] ? 4'h3 : _GEN_25685; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25687 = 10'h2ec == _T_375[9:0] ? 4'h4 : _GEN_25686; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25688 = 10'h2ed == _T_375[9:0] ? 4'h5 : _GEN_25687; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25689 = 10'h2ee == _T_375[9:0] ? 4'h6 : _GEN_25688; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25690 = 10'h2ef == _T_375[9:0] ? 4'h8 : _GEN_25689; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25691 = 10'h2f0 == _T_375[9:0] ? 4'h4 : _GEN_25690; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25692 = 10'h2f1 == _T_375[9:0] ? 4'h9 : _GEN_25691; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25693 = 10'h2f2 == _T_375[9:0] ? 4'hb : _GEN_25692; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25694 = 10'h2f3 == _T_375[9:0] ? 4'hb : _GEN_25693; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25695 = 10'h2f4 == _T_375[9:0] ? 4'hb : _GEN_25694; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25696 = 10'h2f5 == _T_375[9:0] ? 4'hb : _GEN_25695; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25697 = 10'h2f6 == _T_375[9:0] ? 4'hb : _GEN_25696; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25698 = 10'h2f7 == _T_375[9:0] ? 4'hb : _GEN_25697; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25699 = 10'h2f8 == _T_375[9:0] ? 4'h8 : _GEN_25698; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25700 = 10'h2f9 == _T_375[9:0] ? 4'h9 : _GEN_25699; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25701 = 10'h2fa == _T_375[9:0] ? 4'hb : _GEN_25700; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25702 = 10'h2fb == _T_375[9:0] ? 4'hb : _GEN_25701; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25703 = 10'h2fc == _T_375[9:0] ? 4'ha : _GEN_25702; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25704 = 10'h2fd == _T_375[9:0] ? 4'ha : _GEN_25703; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25705 = 10'h2fe == _T_375[9:0] ? 4'h9 : _GEN_25704; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25706 = 10'h2ff == _T_375[9:0] ? 4'h8 : _GEN_25705; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25707 = 10'h300 == _T_375[9:0] ? 4'h8 : _GEN_25706; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25708 = 10'h301 == _T_375[9:0] ? 4'h6 : _GEN_25707; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25709 = 10'h302 == _T_375[9:0] ? 4'h1 : _GEN_25708; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25710 = 10'h303 == _T_375[9:0] ? 4'h0 : _GEN_25709; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25711 = 10'h304 == _T_375[9:0] ? 4'h0 : _GEN_25710; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25712 = 10'h305 == _T_375[9:0] ? 4'h0 : _GEN_25711; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25713 = 10'h306 == _T_375[9:0] ? 4'h0 : _GEN_25712; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25714 = 10'h307 == _T_375[9:0] ? 4'h0 : _GEN_25713; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25715 = 10'h308 == _T_375[9:0] ? 4'h0 : _GEN_25714; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25716 = 10'h309 == _T_375[9:0] ? 4'h0 : _GEN_25715; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25717 = 10'h30a == _T_375[9:0] ? 4'h0 : _GEN_25716; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25718 = 10'h30b == _T_375[9:0] ? 4'h0 : _GEN_25717; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25719 = 10'h30c == _T_375[9:0] ? 4'h2 : _GEN_25718; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25720 = 10'h30d == _T_375[9:0] ? 4'h3 : _GEN_25719; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25721 = 10'h30e == _T_375[9:0] ? 4'h3 : _GEN_25720; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25722 = 10'h30f == _T_375[9:0] ? 4'h3 : _GEN_25721; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25723 = 10'h310 == _T_375[9:0] ? 4'h3 : _GEN_25722; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25724 = 10'h311 == _T_375[9:0] ? 4'h3 : _GEN_25723; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25725 = 10'h312 == _T_375[9:0] ? 4'h4 : _GEN_25724; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25726 = 10'h313 == _T_375[9:0] ? 4'h5 : _GEN_25725; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25727 = 10'h314 == _T_375[9:0] ? 4'h5 : _GEN_25726; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25728 = 10'h315 == _T_375[9:0] ? 4'h8 : _GEN_25727; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25729 = 10'h316 == _T_375[9:0] ? 4'h4 : _GEN_25728; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25730 = 10'h317 == _T_375[9:0] ? 4'h6 : _GEN_25729; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25731 = 10'h318 == _T_375[9:0] ? 4'hb : _GEN_25730; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25732 = 10'h319 == _T_375[9:0] ? 4'hb : _GEN_25731; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25733 = 10'h31a == _T_375[9:0] ? 4'hb : _GEN_25732; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25734 = 10'h31b == _T_375[9:0] ? 4'hb : _GEN_25733; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25735 = 10'h31c == _T_375[9:0] ? 4'hb : _GEN_25734; // @[Filter.scala 230:102]
  wire [3:0] _GEN_25736 = 10'h31d == _T_375[9:0] ? 4'hb : _GEN_25735; // @[Filter.scala 230:102]
  wire [6:0] _GEN_39016 = {{3'd0}, _GEN_25736}; // @[Filter.scala 230:102]
  wire [10:0] _T_382 = _GEN_39016 * 7'h46; // @[Filter.scala 230:102]
  wire [10:0] _GEN_39017 = {{2'd0}, _T_377}; // @[Filter.scala 230:69]
  wire [10:0] _T_384 = _GEN_39017 + _T_382; // @[Filter.scala 230:69]
  wire [3:0] _GEN_25759 = 10'h16 == _T_375[9:0] ? 4'hb : 4'hc; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25760 = 10'h17 == _T_375[9:0] ? 4'h8 : _GEN_25759; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25761 = 10'h18 == _T_375[9:0] ? 4'ha : _GEN_25760; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25762 = 10'h19 == _T_375[9:0] ? 4'hc : _GEN_25761; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25763 = 10'h1a == _T_375[9:0] ? 4'hc : _GEN_25762; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25764 = 10'h1b == _T_375[9:0] ? 4'hc : _GEN_25763; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25765 = 10'h1c == _T_375[9:0] ? 4'hc : _GEN_25764; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25766 = 10'h1d == _T_375[9:0] ? 4'hc : _GEN_25765; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25767 = 10'h1e == _T_375[9:0] ? 4'hc : _GEN_25766; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25768 = 10'h1f == _T_375[9:0] ? 4'hc : _GEN_25767; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25769 = 10'h20 == _T_375[9:0] ? 4'hc : _GEN_25768; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25770 = 10'h21 == _T_375[9:0] ? 4'hc : _GEN_25769; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25771 = 10'h22 == _T_375[9:0] ? 4'hc : _GEN_25770; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25772 = 10'h23 == _T_375[9:0] ? 4'hc : _GEN_25771; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25773 = 10'h24 == _T_375[9:0] ? 4'hc : _GEN_25772; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25774 = 10'h25 == _T_375[9:0] ? 4'hc : _GEN_25773; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25775 = 10'h26 == _T_375[9:0] ? 4'hc : _GEN_25774; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25776 = 10'h27 == _T_375[9:0] ? 4'hc : _GEN_25775; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25777 = 10'h28 == _T_375[9:0] ? 4'hc : _GEN_25776; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25778 = 10'h29 == _T_375[9:0] ? 4'hc : _GEN_25777; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25779 = 10'h2a == _T_375[9:0] ? 4'hc : _GEN_25778; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25780 = 10'h2b == _T_375[9:0] ? 4'hc : _GEN_25779; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25781 = 10'h2c == _T_375[9:0] ? 4'hc : _GEN_25780; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25782 = 10'h2d == _T_375[9:0] ? 4'hc : _GEN_25781; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25783 = 10'h2e == _T_375[9:0] ? 4'hc : _GEN_25782; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25784 = 10'h2f == _T_375[9:0] ? 4'hc : _GEN_25783; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25785 = 10'h30 == _T_375[9:0] ? 4'hc : _GEN_25784; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25786 = 10'h31 == _T_375[9:0] ? 4'hc : _GEN_25785; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25787 = 10'h32 == _T_375[9:0] ? 4'hc : _GEN_25786; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25788 = 10'h33 == _T_375[9:0] ? 4'hc : _GEN_25787; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25789 = 10'h34 == _T_375[9:0] ? 4'hc : _GEN_25788; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25790 = 10'h35 == _T_375[9:0] ? 4'hc : _GEN_25789; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25791 = 10'h36 == _T_375[9:0] ? 4'hc : _GEN_25790; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25792 = 10'h37 == _T_375[9:0] ? 4'hc : _GEN_25791; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25793 = 10'h38 == _T_375[9:0] ? 4'hc : _GEN_25792; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25794 = 10'h39 == _T_375[9:0] ? 4'hc : _GEN_25793; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25795 = 10'h3a == _T_375[9:0] ? 4'hc : _GEN_25794; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25796 = 10'h3b == _T_375[9:0] ? 4'hc : _GEN_25795; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25797 = 10'h3c == _T_375[9:0] ? 4'h7 : _GEN_25796; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25798 = 10'h3d == _T_375[9:0] ? 4'h9 : _GEN_25797; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25799 = 10'h3e == _T_375[9:0] ? 4'h8 : _GEN_25798; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25800 = 10'h3f == _T_375[9:0] ? 4'hc : _GEN_25799; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25801 = 10'h40 == _T_375[9:0] ? 4'hc : _GEN_25800; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25802 = 10'h41 == _T_375[9:0] ? 4'hc : _GEN_25801; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25803 = 10'h42 == _T_375[9:0] ? 4'hc : _GEN_25802; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25804 = 10'h43 == _T_375[9:0] ? 4'hc : _GEN_25803; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25805 = 10'h44 == _T_375[9:0] ? 4'hc : _GEN_25804; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25806 = 10'h45 == _T_375[9:0] ? 4'hc : _GEN_25805; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25807 = 10'h46 == _T_375[9:0] ? 4'hc : _GEN_25806; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25808 = 10'h47 == _T_375[9:0] ? 4'hc : _GEN_25807; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25809 = 10'h48 == _T_375[9:0] ? 4'hc : _GEN_25808; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25810 = 10'h49 == _T_375[9:0] ? 4'hc : _GEN_25809; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25811 = 10'h4a == _T_375[9:0] ? 4'hc : _GEN_25810; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25812 = 10'h4b == _T_375[9:0] ? 4'hc : _GEN_25811; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25813 = 10'h4c == _T_375[9:0] ? 4'hc : _GEN_25812; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25814 = 10'h4d == _T_375[9:0] ? 4'hc : _GEN_25813; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25815 = 10'h4e == _T_375[9:0] ? 4'hc : _GEN_25814; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25816 = 10'h4f == _T_375[9:0] ? 4'hc : _GEN_25815; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25817 = 10'h50 == _T_375[9:0] ? 4'hc : _GEN_25816; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25818 = 10'h51 == _T_375[9:0] ? 4'hc : _GEN_25817; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25819 = 10'h52 == _T_375[9:0] ? 4'hc : _GEN_25818; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25820 = 10'h53 == _T_375[9:0] ? 4'hc : _GEN_25819; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25821 = 10'h54 == _T_375[9:0] ? 4'hc : _GEN_25820; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25822 = 10'h55 == _T_375[9:0] ? 4'hc : _GEN_25821; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25823 = 10'h56 == _T_375[9:0] ? 4'hc : _GEN_25822; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25824 = 10'h57 == _T_375[9:0] ? 4'hc : _GEN_25823; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25825 = 10'h58 == _T_375[9:0] ? 4'hc : _GEN_25824; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25826 = 10'h59 == _T_375[9:0] ? 4'hc : _GEN_25825; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25827 = 10'h5a == _T_375[9:0] ? 4'h9 : _GEN_25826; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25828 = 10'h5b == _T_375[9:0] ? 4'ha : _GEN_25827; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25829 = 10'h5c == _T_375[9:0] ? 4'hc : _GEN_25828; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25830 = 10'h5d == _T_375[9:0] ? 4'hc : _GEN_25829; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25831 = 10'h5e == _T_375[9:0] ? 4'hc : _GEN_25830; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25832 = 10'h5f == _T_375[9:0] ? 4'hc : _GEN_25831; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25833 = 10'h60 == _T_375[9:0] ? 4'hc : _GEN_25832; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25834 = 10'h61 == _T_375[9:0] ? 4'hb : _GEN_25833; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25835 = 10'h62 == _T_375[9:0] ? 4'h8 : _GEN_25834; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25836 = 10'h63 == _T_375[9:0] ? 4'h9 : _GEN_25835; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25837 = 10'h64 == _T_375[9:0] ? 4'h7 : _GEN_25836; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25838 = 10'h65 == _T_375[9:0] ? 4'hb : _GEN_25837; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25839 = 10'h66 == _T_375[9:0] ? 4'hc : _GEN_25838; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25840 = 10'h67 == _T_375[9:0] ? 4'hc : _GEN_25839; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25841 = 10'h68 == _T_375[9:0] ? 4'hc : _GEN_25840; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25842 = 10'h69 == _T_375[9:0] ? 4'hc : _GEN_25841; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25843 = 10'h6a == _T_375[9:0] ? 4'hc : _GEN_25842; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25844 = 10'h6b == _T_375[9:0] ? 4'hb : _GEN_25843; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25845 = 10'h6c == _T_375[9:0] ? 4'h9 : _GEN_25844; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25846 = 10'h6d == _T_375[9:0] ? 4'ha : _GEN_25845; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25847 = 10'h6e == _T_375[9:0] ? 4'hc : _GEN_25846; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25848 = 10'h6f == _T_375[9:0] ? 4'hc : _GEN_25847; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25849 = 10'h70 == _T_375[9:0] ? 4'hc : _GEN_25848; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25850 = 10'h71 == _T_375[9:0] ? 4'hc : _GEN_25849; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25851 = 10'h72 == _T_375[9:0] ? 4'hc : _GEN_25850; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25852 = 10'h73 == _T_375[9:0] ? 4'hc : _GEN_25851; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25853 = 10'h74 == _T_375[9:0] ? 4'hc : _GEN_25852; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25854 = 10'h75 == _T_375[9:0] ? 4'hc : _GEN_25853; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25855 = 10'h76 == _T_375[9:0] ? 4'hc : _GEN_25854; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25856 = 10'h77 == _T_375[9:0] ? 4'hc : _GEN_25855; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25857 = 10'h78 == _T_375[9:0] ? 4'hc : _GEN_25856; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25858 = 10'h79 == _T_375[9:0] ? 4'hc : _GEN_25857; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25859 = 10'h7a == _T_375[9:0] ? 4'hc : _GEN_25858; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25860 = 10'h7b == _T_375[9:0] ? 4'hc : _GEN_25859; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25861 = 10'h7c == _T_375[9:0] ? 4'hc : _GEN_25860; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25862 = 10'h7d == _T_375[9:0] ? 4'hc : _GEN_25861; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25863 = 10'h7e == _T_375[9:0] ? 4'hc : _GEN_25862; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25864 = 10'h7f == _T_375[9:0] ? 4'hc : _GEN_25863; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25865 = 10'h80 == _T_375[9:0] ? 4'hc : _GEN_25864; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25866 = 10'h81 == _T_375[9:0] ? 4'h9 : _GEN_25865; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25867 = 10'h82 == _T_375[9:0] ? 4'h9 : _GEN_25866; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25868 = 10'h83 == _T_375[9:0] ? 4'h9 : _GEN_25867; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25869 = 10'h84 == _T_375[9:0] ? 4'hc : _GEN_25868; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25870 = 10'h85 == _T_375[9:0] ? 4'hc : _GEN_25869; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25871 = 10'h86 == _T_375[9:0] ? 4'hc : _GEN_25870; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25872 = 10'h87 == _T_375[9:0] ? 4'h8 : _GEN_25871; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25873 = 10'h88 == _T_375[9:0] ? 4'h9 : _GEN_25872; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25874 = 10'h89 == _T_375[9:0] ? 4'h9 : _GEN_25873; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25875 = 10'h8a == _T_375[9:0] ? 4'h9 : _GEN_25874; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25876 = 10'h8b == _T_375[9:0] ? 4'hc : _GEN_25875; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25877 = 10'h8c == _T_375[9:0] ? 4'hc : _GEN_25876; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25878 = 10'h8d == _T_375[9:0] ? 4'hc : _GEN_25877; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25879 = 10'h8e == _T_375[9:0] ? 4'hc : _GEN_25878; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25880 = 10'h8f == _T_375[9:0] ? 4'h9 : _GEN_25879; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25881 = 10'h90 == _T_375[9:0] ? 4'h9 : _GEN_25880; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25882 = 10'h91 == _T_375[9:0] ? 4'h9 : _GEN_25881; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25883 = 10'h92 == _T_375[9:0] ? 4'ha : _GEN_25882; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25884 = 10'h93 == _T_375[9:0] ? 4'hc : _GEN_25883; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25885 = 10'h94 == _T_375[9:0] ? 4'hc : _GEN_25884; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25886 = 10'h95 == _T_375[9:0] ? 4'hc : _GEN_25885; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25887 = 10'h96 == _T_375[9:0] ? 4'hc : _GEN_25886; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25888 = 10'h97 == _T_375[9:0] ? 4'hc : _GEN_25887; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25889 = 10'h98 == _T_375[9:0] ? 4'hc : _GEN_25888; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25890 = 10'h99 == _T_375[9:0] ? 4'hc : _GEN_25889; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25891 = 10'h9a == _T_375[9:0] ? 4'hc : _GEN_25890; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25892 = 10'h9b == _T_375[9:0] ? 4'hc : _GEN_25891; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25893 = 10'h9c == _T_375[9:0] ? 4'hc : _GEN_25892; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25894 = 10'h9d == _T_375[9:0] ? 4'hc : _GEN_25893; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25895 = 10'h9e == _T_375[9:0] ? 4'hc : _GEN_25894; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25896 = 10'h9f == _T_375[9:0] ? 4'hc : _GEN_25895; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25897 = 10'ha0 == _T_375[9:0] ? 4'hc : _GEN_25896; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25898 = 10'ha1 == _T_375[9:0] ? 4'hc : _GEN_25897; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25899 = 10'ha2 == _T_375[9:0] ? 4'hc : _GEN_25898; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25900 = 10'ha3 == _T_375[9:0] ? 4'hc : _GEN_25899; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25901 = 10'ha4 == _T_375[9:0] ? 4'hc : _GEN_25900; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25902 = 10'ha5 == _T_375[9:0] ? 4'hc : _GEN_25901; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25903 = 10'ha6 == _T_375[9:0] ? 4'hc : _GEN_25902; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25904 = 10'ha7 == _T_375[9:0] ? 4'hc : _GEN_25903; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25905 = 10'ha8 == _T_375[9:0] ? 4'h9 : _GEN_25904; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25906 = 10'ha9 == _T_375[9:0] ? 4'h8 : _GEN_25905; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25907 = 10'haa == _T_375[9:0] ? 4'h8 : _GEN_25906; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25908 = 10'hab == _T_375[9:0] ? 4'ha : _GEN_25907; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25909 = 10'hac == _T_375[9:0] ? 4'hb : _GEN_25908; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25910 = 10'had == _T_375[9:0] ? 4'h7 : _GEN_25909; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25911 = 10'hae == _T_375[9:0] ? 4'h9 : _GEN_25910; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25912 = 10'haf == _T_375[9:0] ? 4'h9 : _GEN_25911; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25913 = 10'hb0 == _T_375[9:0] ? 4'h8 : _GEN_25912; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25914 = 10'hb1 == _T_375[9:0] ? 4'h9 : _GEN_25913; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25915 = 10'hb2 == _T_375[9:0] ? 4'hc : _GEN_25914; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25916 = 10'hb3 == _T_375[9:0] ? 4'h9 : _GEN_25915; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25917 = 10'hb4 == _T_375[9:0] ? 4'h9 : _GEN_25916; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25918 = 10'hb5 == _T_375[9:0] ? 4'h9 : _GEN_25917; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25919 = 10'hb6 == _T_375[9:0] ? 4'h9 : _GEN_25918; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25920 = 10'hb7 == _T_375[9:0] ? 4'ha : _GEN_25919; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25921 = 10'hb8 == _T_375[9:0] ? 4'hc : _GEN_25920; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25922 = 10'hb9 == _T_375[9:0] ? 4'hc : _GEN_25921; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25923 = 10'hba == _T_375[9:0] ? 4'hc : _GEN_25922; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25924 = 10'hbb == _T_375[9:0] ? 4'hc : _GEN_25923; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25925 = 10'hbc == _T_375[9:0] ? 4'hc : _GEN_25924; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25926 = 10'hbd == _T_375[9:0] ? 4'hb : _GEN_25925; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25927 = 10'hbe == _T_375[9:0] ? 4'hc : _GEN_25926; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25928 = 10'hbf == _T_375[9:0] ? 4'hc : _GEN_25927; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25929 = 10'hc0 == _T_375[9:0] ? 4'hc : _GEN_25928; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25930 = 10'hc1 == _T_375[9:0] ? 4'hc : _GEN_25929; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25931 = 10'hc2 == _T_375[9:0] ? 4'hc : _GEN_25930; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25932 = 10'hc3 == _T_375[9:0] ? 4'hc : _GEN_25931; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25933 = 10'hc4 == _T_375[9:0] ? 4'hc : _GEN_25932; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25934 = 10'hc5 == _T_375[9:0] ? 4'hc : _GEN_25933; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25935 = 10'hc6 == _T_375[9:0] ? 4'hb : _GEN_25934; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25936 = 10'hc7 == _T_375[9:0] ? 4'hb : _GEN_25935; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25937 = 10'hc8 == _T_375[9:0] ? 4'ha : _GEN_25936; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25938 = 10'hc9 == _T_375[9:0] ? 4'ha : _GEN_25937; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25939 = 10'hca == _T_375[9:0] ? 4'hb : _GEN_25938; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25940 = 10'hcb == _T_375[9:0] ? 4'hc : _GEN_25939; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25941 = 10'hcc == _T_375[9:0] ? 4'hc : _GEN_25940; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25942 = 10'hcd == _T_375[9:0] ? 4'hc : _GEN_25941; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25943 = 10'hce == _T_375[9:0] ? 4'ha : _GEN_25942; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25944 = 10'hcf == _T_375[9:0] ? 4'h8 : _GEN_25943; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25945 = 10'hd0 == _T_375[9:0] ? 4'h9 : _GEN_25944; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25946 = 10'hd1 == _T_375[9:0] ? 4'h8 : _GEN_25945; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25947 = 10'hd2 == _T_375[9:0] ? 4'h9 : _GEN_25946; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25948 = 10'hd3 == _T_375[9:0] ? 4'h9 : _GEN_25947; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25949 = 10'hd4 == _T_375[9:0] ? 4'h9 : _GEN_25948; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25950 = 10'hd5 == _T_375[9:0] ? 4'h9 : _GEN_25949; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25951 = 10'hd6 == _T_375[9:0] ? 4'ha : _GEN_25950; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25952 = 10'hd7 == _T_375[9:0] ? 4'h9 : _GEN_25951; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25953 = 10'hd8 == _T_375[9:0] ? 4'h9 : _GEN_25952; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25954 = 10'hd9 == _T_375[9:0] ? 4'h9 : _GEN_25953; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25955 = 10'hda == _T_375[9:0] ? 4'ha : _GEN_25954; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25956 = 10'hdb == _T_375[9:0] ? 4'h9 : _GEN_25955; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25957 = 10'hdc == _T_375[9:0] ? 4'h7 : _GEN_25956; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25958 = 10'hdd == _T_375[9:0] ? 4'hc : _GEN_25957; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25959 = 10'hde == _T_375[9:0] ? 4'hc : _GEN_25958; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25960 = 10'hdf == _T_375[9:0] ? 4'hc : _GEN_25959; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25961 = 10'he0 == _T_375[9:0] ? 4'hc : _GEN_25960; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25962 = 10'he1 == _T_375[9:0] ? 4'hc : _GEN_25961; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25963 = 10'he2 == _T_375[9:0] ? 4'hc : _GEN_25962; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25964 = 10'he3 == _T_375[9:0] ? 4'h8 : _GEN_25963; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25965 = 10'he4 == _T_375[9:0] ? 4'hc : _GEN_25964; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25966 = 10'he5 == _T_375[9:0] ? 4'hc : _GEN_25965; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25967 = 10'he6 == _T_375[9:0] ? 4'hc : _GEN_25966; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25968 = 10'he7 == _T_375[9:0] ? 4'hc : _GEN_25967; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25969 = 10'he8 == _T_375[9:0] ? 4'hc : _GEN_25968; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25970 = 10'he9 == _T_375[9:0] ? 4'hc : _GEN_25969; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25971 = 10'hea == _T_375[9:0] ? 4'hc : _GEN_25970; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25972 = 10'heb == _T_375[9:0] ? 4'ha : _GEN_25971; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25973 = 10'hec == _T_375[9:0] ? 4'h7 : _GEN_25972; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25974 = 10'hed == _T_375[9:0] ? 4'h3 : _GEN_25973; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25975 = 10'hee == _T_375[9:0] ? 4'h3 : _GEN_25974; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25976 = 10'hef == _T_375[9:0] ? 4'h3 : _GEN_25975; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25977 = 10'hf0 == _T_375[9:0] ? 4'h3 : _GEN_25976; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25978 = 10'hf1 == _T_375[9:0] ? 4'h8 : _GEN_25977; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25979 = 10'hf2 == _T_375[9:0] ? 4'hc : _GEN_25978; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25980 = 10'hf3 == _T_375[9:0] ? 4'hc : _GEN_25979; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25981 = 10'hf4 == _T_375[9:0] ? 4'hc : _GEN_25980; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25982 = 10'hf5 == _T_375[9:0] ? 4'h9 : _GEN_25981; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25983 = 10'hf6 == _T_375[9:0] ? 4'h9 : _GEN_25982; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25984 = 10'hf7 == _T_375[9:0] ? 4'h9 : _GEN_25983; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25985 = 10'hf8 == _T_375[9:0] ? 4'h9 : _GEN_25984; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25986 = 10'hf9 == _T_375[9:0] ? 4'ha : _GEN_25985; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25987 = 10'hfa == _T_375[9:0] ? 4'h9 : _GEN_25986; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25988 = 10'hfb == _T_375[9:0] ? 4'h9 : _GEN_25987; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25989 = 10'hfc == _T_375[9:0] ? 4'h9 : _GEN_25988; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25990 = 10'hfd == _T_375[9:0] ? 4'h9 : _GEN_25989; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25991 = 10'hfe == _T_375[9:0] ? 4'h9 : _GEN_25990; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25992 = 10'hff == _T_375[9:0] ? 4'ha : _GEN_25991; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25993 = 10'h100 == _T_375[9:0] ? 4'ha : _GEN_25992; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25994 = 10'h101 == _T_375[9:0] ? 4'h7 : _GEN_25993; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25995 = 10'h102 == _T_375[9:0] ? 4'h9 : _GEN_25994; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25996 = 10'h103 == _T_375[9:0] ? 4'hc : _GEN_25995; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25997 = 10'h104 == _T_375[9:0] ? 4'hc : _GEN_25996; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25998 = 10'h105 == _T_375[9:0] ? 4'hb : _GEN_25997; // @[Filter.scala 230:142]
  wire [3:0] _GEN_25999 = 10'h106 == _T_375[9:0] ? 4'hb : _GEN_25998; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26000 = 10'h107 == _T_375[9:0] ? 4'hb : _GEN_25999; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26001 = 10'h108 == _T_375[9:0] ? 4'hb : _GEN_26000; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26002 = 10'h109 == _T_375[9:0] ? 4'h7 : _GEN_26001; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26003 = 10'h10a == _T_375[9:0] ? 4'hc : _GEN_26002; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26004 = 10'h10b == _T_375[9:0] ? 4'hc : _GEN_26003; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26005 = 10'h10c == _T_375[9:0] ? 4'hc : _GEN_26004; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26006 = 10'h10d == _T_375[9:0] ? 4'hc : _GEN_26005; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26007 = 10'h10e == _T_375[9:0] ? 4'hc : _GEN_26006; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26008 = 10'h10f == _T_375[9:0] ? 4'h9 : _GEN_26007; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26009 = 10'h110 == _T_375[9:0] ? 4'hb : _GEN_26008; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26010 = 10'h111 == _T_375[9:0] ? 4'h4 : _GEN_26009; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26011 = 10'h112 == _T_375[9:0] ? 4'h7 : _GEN_26010; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26012 = 10'h113 == _T_375[9:0] ? 4'h3 : _GEN_26011; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26013 = 10'h114 == _T_375[9:0] ? 4'h3 : _GEN_26012; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26014 = 10'h115 == _T_375[9:0] ? 4'h3 : _GEN_26013; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26015 = 10'h116 == _T_375[9:0] ? 4'h3 : _GEN_26014; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26016 = 10'h117 == _T_375[9:0] ? 4'h2 : _GEN_26015; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26017 = 10'h118 == _T_375[9:0] ? 4'h9 : _GEN_26016; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26018 = 10'h119 == _T_375[9:0] ? 4'hc : _GEN_26017; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26019 = 10'h11a == _T_375[9:0] ? 4'hc : _GEN_26018; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26020 = 10'h11b == _T_375[9:0] ? 4'hc : _GEN_26019; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26021 = 10'h11c == _T_375[9:0] ? 4'h9 : _GEN_26020; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26022 = 10'h11d == _T_375[9:0] ? 4'h9 : _GEN_26021; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26023 = 10'h11e == _T_375[9:0] ? 4'h9 : _GEN_26022; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26024 = 10'h11f == _T_375[9:0] ? 4'h8 : _GEN_26023; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26025 = 10'h120 == _T_375[9:0] ? 4'h7 : _GEN_26024; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26026 = 10'h121 == _T_375[9:0] ? 4'h9 : _GEN_26025; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26027 = 10'h122 == _T_375[9:0] ? 4'h7 : _GEN_26026; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26028 = 10'h123 == _T_375[9:0] ? 4'h7 : _GEN_26027; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26029 = 10'h124 == _T_375[9:0] ? 4'h9 : _GEN_26028; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26030 = 10'h125 == _T_375[9:0] ? 4'h9 : _GEN_26029; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26031 = 10'h126 == _T_375[9:0] ? 4'h8 : _GEN_26030; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26032 = 10'h127 == _T_375[9:0] ? 4'h9 : _GEN_26031; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26033 = 10'h128 == _T_375[9:0] ? 4'h8 : _GEN_26032; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26034 = 10'h129 == _T_375[9:0] ? 4'ha : _GEN_26033; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26035 = 10'h12a == _T_375[9:0] ? 4'h5 : _GEN_26034; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26036 = 10'h12b == _T_375[9:0] ? 4'h3 : _GEN_26035; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26037 = 10'h12c == _T_375[9:0] ? 4'h3 : _GEN_26036; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26038 = 10'h12d == _T_375[9:0] ? 4'h3 : _GEN_26037; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26039 = 10'h12e == _T_375[9:0] ? 4'h5 : _GEN_26038; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26040 = 10'h12f == _T_375[9:0] ? 4'h8 : _GEN_26039; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26041 = 10'h130 == _T_375[9:0] ? 4'hc : _GEN_26040; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26042 = 10'h131 == _T_375[9:0] ? 4'hb : _GEN_26041; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26043 = 10'h132 == _T_375[9:0] ? 4'h9 : _GEN_26042; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26044 = 10'h133 == _T_375[9:0] ? 4'h8 : _GEN_26043; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26045 = 10'h134 == _T_375[9:0] ? 4'h9 : _GEN_26044; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26046 = 10'h135 == _T_375[9:0] ? 4'h7 : _GEN_26045; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26047 = 10'h136 == _T_375[9:0] ? 4'h7 : _GEN_26046; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26048 = 10'h137 == _T_375[9:0] ? 4'h5 : _GEN_26047; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26049 = 10'h138 == _T_375[9:0] ? 4'h7 : _GEN_26048; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26050 = 10'h139 == _T_375[9:0] ? 4'h3 : _GEN_26049; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26051 = 10'h13a == _T_375[9:0] ? 4'h3 : _GEN_26050; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26052 = 10'h13b == _T_375[9:0] ? 4'h3 : _GEN_26051; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26053 = 10'h13c == _T_375[9:0] ? 4'h3 : _GEN_26052; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26054 = 10'h13d == _T_375[9:0] ? 4'h3 : _GEN_26053; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26055 = 10'h13e == _T_375[9:0] ? 4'h5 : _GEN_26054; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26056 = 10'h13f == _T_375[9:0] ? 4'ha : _GEN_26055; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26057 = 10'h140 == _T_375[9:0] ? 4'hc : _GEN_26056; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26058 = 10'h141 == _T_375[9:0] ? 4'hc : _GEN_26057; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26059 = 10'h142 == _T_375[9:0] ? 4'hc : _GEN_26058; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26060 = 10'h143 == _T_375[9:0] ? 4'h9 : _GEN_26059; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26061 = 10'h144 == _T_375[9:0] ? 4'h9 : _GEN_26060; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26062 = 10'h145 == _T_375[9:0] ? 4'h8 : _GEN_26061; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26063 = 10'h146 == _T_375[9:0] ? 4'h8 : _GEN_26062; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26064 = 10'h147 == _T_375[9:0] ? 4'h7 : _GEN_26063; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26065 = 10'h148 == _T_375[9:0] ? 4'h8 : _GEN_26064; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26066 = 10'h149 == _T_375[9:0] ? 4'h9 : _GEN_26065; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26067 = 10'h14a == _T_375[9:0] ? 4'ha : _GEN_26066; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26068 = 10'h14b == _T_375[9:0] ? 4'h9 : _GEN_26067; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26069 = 10'h14c == _T_375[9:0] ? 4'ha : _GEN_26068; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26070 = 10'h14d == _T_375[9:0] ? 4'h9 : _GEN_26069; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26071 = 10'h14e == _T_375[9:0] ? 4'h7 : _GEN_26070; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26072 = 10'h14f == _T_375[9:0] ? 4'h3 : _GEN_26071; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26073 = 10'h150 == _T_375[9:0] ? 4'h3 : _GEN_26072; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26074 = 10'h151 == _T_375[9:0] ? 4'h3 : _GEN_26073; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26075 = 10'h152 == _T_375[9:0] ? 4'h3 : _GEN_26074; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26076 = 10'h153 == _T_375[9:0] ? 4'h3 : _GEN_26075; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26077 = 10'h154 == _T_375[9:0] ? 4'h3 : _GEN_26076; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26078 = 10'h155 == _T_375[9:0] ? 4'h8 : _GEN_26077; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26079 = 10'h156 == _T_375[9:0] ? 4'ha : _GEN_26078; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26080 = 10'h157 == _T_375[9:0] ? 4'h7 : _GEN_26079; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26081 = 10'h158 == _T_375[9:0] ? 4'h7 : _GEN_26080; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26082 = 10'h159 == _T_375[9:0] ? 4'h7 : _GEN_26081; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26083 = 10'h15a == _T_375[9:0] ? 4'h7 : _GEN_26082; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26084 = 10'h15b == _T_375[9:0] ? 4'h7 : _GEN_26083; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26085 = 10'h15c == _T_375[9:0] ? 4'h7 : _GEN_26084; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26086 = 10'h15d == _T_375[9:0] ? 4'h7 : _GEN_26085; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26087 = 10'h15e == _T_375[9:0] ? 4'h7 : _GEN_26086; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26088 = 10'h15f == _T_375[9:0] ? 4'h3 : _GEN_26087; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26089 = 10'h160 == _T_375[9:0] ? 4'h3 : _GEN_26088; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26090 = 10'h161 == _T_375[9:0] ? 4'h3 : _GEN_26089; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26091 = 10'h162 == _T_375[9:0] ? 4'h3 : _GEN_26090; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26092 = 10'h163 == _T_375[9:0] ? 4'h3 : _GEN_26091; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26093 = 10'h164 == _T_375[9:0] ? 4'h4 : _GEN_26092; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26094 = 10'h165 == _T_375[9:0] ? 4'ha : _GEN_26093; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26095 = 10'h166 == _T_375[9:0] ? 4'ha : _GEN_26094; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26096 = 10'h167 == _T_375[9:0] ? 4'hc : _GEN_26095; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26097 = 10'h168 == _T_375[9:0] ? 4'hc : _GEN_26096; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26098 = 10'h169 == _T_375[9:0] ? 4'h9 : _GEN_26097; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26099 = 10'h16a == _T_375[9:0] ? 4'h9 : _GEN_26098; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26100 = 10'h16b == _T_375[9:0] ? 4'ha : _GEN_26099; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26101 = 10'h16c == _T_375[9:0] ? 4'h7 : _GEN_26100; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26102 = 10'h16d == _T_375[9:0] ? 4'h7 : _GEN_26101; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26103 = 10'h16e == _T_375[9:0] ? 4'h7 : _GEN_26102; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26104 = 10'h16f == _T_375[9:0] ? 4'ha : _GEN_26103; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26105 = 10'h170 == _T_375[9:0] ? 4'ha : _GEN_26104; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26106 = 10'h171 == _T_375[9:0] ? 4'ha : _GEN_26105; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26107 = 10'h172 == _T_375[9:0] ? 4'hc : _GEN_26106; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26108 = 10'h173 == _T_375[9:0] ? 4'h8 : _GEN_26107; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26109 = 10'h174 == _T_375[9:0] ? 4'h5 : _GEN_26108; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26110 = 10'h175 == _T_375[9:0] ? 4'h8 : _GEN_26109; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26111 = 10'h176 == _T_375[9:0] ? 4'h7 : _GEN_26110; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26112 = 10'h177 == _T_375[9:0] ? 4'h8 : _GEN_26111; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26113 = 10'h178 == _T_375[9:0] ? 4'h7 : _GEN_26112; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26114 = 10'h179 == _T_375[9:0] ? 4'h5 : _GEN_26113; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26115 = 10'h17a == _T_375[9:0] ? 4'h5 : _GEN_26114; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26116 = 10'h17b == _T_375[9:0] ? 4'h7 : _GEN_26115; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26117 = 10'h17c == _T_375[9:0] ? 4'h7 : _GEN_26116; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26118 = 10'h17d == _T_375[9:0] ? 4'h7 : _GEN_26117; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26119 = 10'h17e == _T_375[9:0] ? 4'h7 : _GEN_26118; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26120 = 10'h17f == _T_375[9:0] ? 4'h7 : _GEN_26119; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26121 = 10'h180 == _T_375[9:0] ? 4'h7 : _GEN_26120; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26122 = 10'h181 == _T_375[9:0] ? 4'h7 : _GEN_26121; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26123 = 10'h182 == _T_375[9:0] ? 4'h7 : _GEN_26122; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26124 = 10'h183 == _T_375[9:0] ? 4'h7 : _GEN_26123; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26125 = 10'h184 == _T_375[9:0] ? 4'h7 : _GEN_26124; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26126 = 10'h185 == _T_375[9:0] ? 4'h5 : _GEN_26125; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26127 = 10'h186 == _T_375[9:0] ? 4'h3 : _GEN_26126; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26128 = 10'h187 == _T_375[9:0] ? 4'h3 : _GEN_26127; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26129 = 10'h188 == _T_375[9:0] ? 4'h3 : _GEN_26128; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26130 = 10'h189 == _T_375[9:0] ? 4'h4 : _GEN_26129; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26131 = 10'h18a == _T_375[9:0] ? 4'h5 : _GEN_26130; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26132 = 10'h18b == _T_375[9:0] ? 4'ha : _GEN_26131; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26133 = 10'h18c == _T_375[9:0] ? 4'ha : _GEN_26132; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26134 = 10'h18d == _T_375[9:0] ? 4'ha : _GEN_26133; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26135 = 10'h18e == _T_375[9:0] ? 4'hc : _GEN_26134; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26136 = 10'h18f == _T_375[9:0] ? 4'h8 : _GEN_26135; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26137 = 10'h190 == _T_375[9:0] ? 4'h9 : _GEN_26136; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26138 = 10'h191 == _T_375[9:0] ? 4'h8 : _GEN_26137; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26139 = 10'h192 == _T_375[9:0] ? 4'h7 : _GEN_26138; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26140 = 10'h193 == _T_375[9:0] ? 4'h7 : _GEN_26139; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26141 = 10'h194 == _T_375[9:0] ? 4'h7 : _GEN_26140; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26142 = 10'h195 == _T_375[9:0] ? 4'h9 : _GEN_26141; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26143 = 10'h196 == _T_375[9:0] ? 4'ha : _GEN_26142; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26144 = 10'h197 == _T_375[9:0] ? 4'h8 : _GEN_26143; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26145 = 10'h198 == _T_375[9:0] ? 4'hc : _GEN_26144; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26146 = 10'h199 == _T_375[9:0] ? 4'h5 : _GEN_26145; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26147 = 10'h19a == _T_375[9:0] ? 4'h1 : _GEN_26146; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26148 = 10'h19b == _T_375[9:0] ? 4'h4 : _GEN_26147; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26149 = 10'h19c == _T_375[9:0] ? 4'h7 : _GEN_26148; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26150 = 10'h19d == _T_375[9:0] ? 4'h5 : _GEN_26149; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26151 = 10'h19e == _T_375[9:0] ? 4'h2 : _GEN_26150; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26152 = 10'h19f == _T_375[9:0] ? 4'h3 : _GEN_26151; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26153 = 10'h1a0 == _T_375[9:0] ? 4'h7 : _GEN_26152; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26154 = 10'h1a1 == _T_375[9:0] ? 4'h7 : _GEN_26153; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26155 = 10'h1a2 == _T_375[9:0] ? 4'h7 : _GEN_26154; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26156 = 10'h1a3 == _T_375[9:0] ? 4'h7 : _GEN_26155; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26157 = 10'h1a4 == _T_375[9:0] ? 4'h7 : _GEN_26156; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26158 = 10'h1a5 == _T_375[9:0] ? 4'h7 : _GEN_26157; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26159 = 10'h1a6 == _T_375[9:0] ? 4'h7 : _GEN_26158; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26160 = 10'h1a7 == _T_375[9:0] ? 4'h7 : _GEN_26159; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26161 = 10'h1a8 == _T_375[9:0] ? 4'h8 : _GEN_26160; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26162 = 10'h1a9 == _T_375[9:0] ? 4'h8 : _GEN_26161; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26163 = 10'h1aa == _T_375[9:0] ? 4'h6 : _GEN_26162; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26164 = 10'h1ab == _T_375[9:0] ? 4'h6 : _GEN_26163; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26165 = 10'h1ac == _T_375[9:0] ? 4'h5 : _GEN_26164; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26166 = 10'h1ad == _T_375[9:0] ? 4'h4 : _GEN_26165; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26167 = 10'h1ae == _T_375[9:0] ? 4'h3 : _GEN_26166; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26168 = 10'h1af == _T_375[9:0] ? 4'h6 : _GEN_26167; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26169 = 10'h1b0 == _T_375[9:0] ? 4'h6 : _GEN_26168; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26170 = 10'h1b1 == _T_375[9:0] ? 4'ha : _GEN_26169; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26171 = 10'h1b2 == _T_375[9:0] ? 4'ha : _GEN_26170; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26172 = 10'h1b3 == _T_375[9:0] ? 4'h9 : _GEN_26171; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26173 = 10'h1b4 == _T_375[9:0] ? 4'hb : _GEN_26172; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26174 = 10'h1b5 == _T_375[9:0] ? 4'h8 : _GEN_26173; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26175 = 10'h1b6 == _T_375[9:0] ? 4'h8 : _GEN_26174; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26176 = 10'h1b7 == _T_375[9:0] ? 4'h7 : _GEN_26175; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26177 = 10'h1b8 == _T_375[9:0] ? 4'h6 : _GEN_26176; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26178 = 10'h1b9 == _T_375[9:0] ? 4'h7 : _GEN_26177; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26179 = 10'h1ba == _T_375[9:0] ? 4'h6 : _GEN_26178; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26180 = 10'h1bb == _T_375[9:0] ? 4'h8 : _GEN_26179; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26181 = 10'h1bc == _T_375[9:0] ? 4'ha : _GEN_26180; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26182 = 10'h1bd == _T_375[9:0] ? 4'h9 : _GEN_26181; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26183 = 10'h1be == _T_375[9:0] ? 4'hc : _GEN_26182; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26184 = 10'h1bf == _T_375[9:0] ? 4'h7 : _GEN_26183; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26185 = 10'h1c0 == _T_375[9:0] ? 4'h6 : _GEN_26184; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26186 = 10'h1c1 == _T_375[9:0] ? 4'h7 : _GEN_26185; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26187 = 10'h1c2 == _T_375[9:0] ? 4'h7 : _GEN_26186; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26188 = 10'h1c3 == _T_375[9:0] ? 4'h6 : _GEN_26187; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26189 = 10'h1c4 == _T_375[9:0] ? 4'h5 : _GEN_26188; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26190 = 10'h1c5 == _T_375[9:0] ? 4'h6 : _GEN_26189; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26191 = 10'h1c6 == _T_375[9:0] ? 4'h8 : _GEN_26190; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26192 = 10'h1c7 == _T_375[9:0] ? 4'h7 : _GEN_26191; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26193 = 10'h1c8 == _T_375[9:0] ? 4'h7 : _GEN_26192; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26194 = 10'h1c9 == _T_375[9:0] ? 4'h7 : _GEN_26193; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26195 = 10'h1ca == _T_375[9:0] ? 4'h7 : _GEN_26194; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26196 = 10'h1cb == _T_375[9:0] ? 4'h7 : _GEN_26195; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26197 = 10'h1cc == _T_375[9:0] ? 4'h7 : _GEN_26196; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26198 = 10'h1cd == _T_375[9:0] ? 4'h8 : _GEN_26197; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26199 = 10'h1ce == _T_375[9:0] ? 4'h8 : _GEN_26198; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26200 = 10'h1cf == _T_375[9:0] ? 4'h8 : _GEN_26199; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26201 = 10'h1d0 == _T_375[9:0] ? 4'h5 : _GEN_26200; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26202 = 10'h1d1 == _T_375[9:0] ? 4'h6 : _GEN_26201; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26203 = 10'h1d2 == _T_375[9:0] ? 4'h7 : _GEN_26202; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26204 = 10'h1d3 == _T_375[9:0] ? 4'h7 : _GEN_26203; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26205 = 10'h1d4 == _T_375[9:0] ? 4'h7 : _GEN_26204; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26206 = 10'h1d5 == _T_375[9:0] ? 4'h6 : _GEN_26205; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26207 = 10'h1d6 == _T_375[9:0] ? 4'h8 : _GEN_26206; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26208 = 10'h1d7 == _T_375[9:0] ? 4'ha : _GEN_26207; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26209 = 10'h1d8 == _T_375[9:0] ? 4'ha : _GEN_26208; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26210 = 10'h1d9 == _T_375[9:0] ? 4'ha : _GEN_26209; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26211 = 10'h1da == _T_375[9:0] ? 4'h8 : _GEN_26210; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26212 = 10'h1db == _T_375[9:0] ? 4'h9 : _GEN_26211; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26213 = 10'h1dc == _T_375[9:0] ? 4'h9 : _GEN_26212; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26214 = 10'h1dd == _T_375[9:0] ? 4'h5 : _GEN_26213; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26215 = 10'h1de == _T_375[9:0] ? 4'h7 : _GEN_26214; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26216 = 10'h1df == _T_375[9:0] ? 4'h7 : _GEN_26215; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26217 = 10'h1e0 == _T_375[9:0] ? 4'h7 : _GEN_26216; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26218 = 10'h1e1 == _T_375[9:0] ? 4'h6 : _GEN_26217; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26219 = 10'h1e2 == _T_375[9:0] ? 4'h9 : _GEN_26218; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26220 = 10'h1e3 == _T_375[9:0] ? 4'h9 : _GEN_26219; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26221 = 10'h1e4 == _T_375[9:0] ? 4'hb : _GEN_26220; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26222 = 10'h1e5 == _T_375[9:0] ? 4'h8 : _GEN_26221; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26223 = 10'h1e6 == _T_375[9:0] ? 4'h7 : _GEN_26222; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26224 = 10'h1e7 == _T_375[9:0] ? 4'h8 : _GEN_26223; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26225 = 10'h1e8 == _T_375[9:0] ? 4'h8 : _GEN_26224; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26226 = 10'h1e9 == _T_375[9:0] ? 4'h8 : _GEN_26225; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26227 = 10'h1ea == _T_375[9:0] ? 4'h8 : _GEN_26226; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26228 = 10'h1eb == _T_375[9:0] ? 4'h8 : _GEN_26227; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26229 = 10'h1ec == _T_375[9:0] ? 4'h8 : _GEN_26228; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26230 = 10'h1ed == _T_375[9:0] ? 4'h6 : _GEN_26229; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26231 = 10'h1ee == _T_375[9:0] ? 4'h7 : _GEN_26230; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26232 = 10'h1ef == _T_375[9:0] ? 4'h7 : _GEN_26231; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26233 = 10'h1f0 == _T_375[9:0] ? 4'h7 : _GEN_26232; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26234 = 10'h1f1 == _T_375[9:0] ? 4'h7 : _GEN_26233; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26235 = 10'h1f2 == _T_375[9:0] ? 4'h7 : _GEN_26234; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26236 = 10'h1f3 == _T_375[9:0] ? 4'h8 : _GEN_26235; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26237 = 10'h1f4 == _T_375[9:0] ? 4'h8 : _GEN_26236; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26238 = 10'h1f5 == _T_375[9:0] ? 4'h8 : _GEN_26237; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26239 = 10'h1f6 == _T_375[9:0] ? 4'ha : _GEN_26238; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26240 = 10'h1f7 == _T_375[9:0] ? 4'h6 : _GEN_26239; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26241 = 10'h1f8 == _T_375[9:0] ? 4'h6 : _GEN_26240; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26242 = 10'h1f9 == _T_375[9:0] ? 4'h8 : _GEN_26241; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26243 = 10'h1fa == _T_375[9:0] ? 4'h8 : _GEN_26242; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26244 = 10'h1fb == _T_375[9:0] ? 4'h6 : _GEN_26243; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26245 = 10'h1fc == _T_375[9:0] ? 4'ha : _GEN_26244; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26246 = 10'h1fd == _T_375[9:0] ? 4'hb : _GEN_26245; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26247 = 10'h1fe == _T_375[9:0] ? 4'ha : _GEN_26246; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26248 = 10'h1ff == _T_375[9:0] ? 4'ha : _GEN_26247; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26249 = 10'h200 == _T_375[9:0] ? 4'h4 : _GEN_26248; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26250 = 10'h201 == _T_375[9:0] ? 4'h7 : _GEN_26249; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26251 = 10'h202 == _T_375[9:0] ? 4'h6 : _GEN_26250; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26252 = 10'h203 == _T_375[9:0] ? 4'h6 : _GEN_26251; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26253 = 10'h204 == _T_375[9:0] ? 4'h5 : _GEN_26252; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26254 = 10'h205 == _T_375[9:0] ? 4'h6 : _GEN_26253; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26255 = 10'h206 == _T_375[9:0] ? 4'h6 : _GEN_26254; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26256 = 10'h207 == _T_375[9:0] ? 4'h5 : _GEN_26255; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26257 = 10'h208 == _T_375[9:0] ? 4'h7 : _GEN_26256; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26258 = 10'h209 == _T_375[9:0] ? 4'h9 : _GEN_26257; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26259 = 10'h20a == _T_375[9:0] ? 4'hb : _GEN_26258; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26260 = 10'h20b == _T_375[9:0] ? 4'h7 : _GEN_26259; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26261 = 10'h20c == _T_375[9:0] ? 4'h7 : _GEN_26260; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26262 = 10'h20d == _T_375[9:0] ? 4'h7 : _GEN_26261; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26263 = 10'h20e == _T_375[9:0] ? 4'h7 : _GEN_26262; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26264 = 10'h20f == _T_375[9:0] ? 4'h7 : _GEN_26263; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26265 = 10'h210 == _T_375[9:0] ? 4'h7 : _GEN_26264; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26266 = 10'h211 == _T_375[9:0] ? 4'h8 : _GEN_26265; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26267 = 10'h212 == _T_375[9:0] ? 4'h8 : _GEN_26266; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26268 = 10'h213 == _T_375[9:0] ? 4'h9 : _GEN_26267; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26269 = 10'h214 == _T_375[9:0] ? 4'h6 : _GEN_26268; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26270 = 10'h215 == _T_375[9:0] ? 4'h7 : _GEN_26269; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26271 = 10'h216 == _T_375[9:0] ? 4'h7 : _GEN_26270; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26272 = 10'h217 == _T_375[9:0] ? 4'h7 : _GEN_26271; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26273 = 10'h218 == _T_375[9:0] ? 4'h7 : _GEN_26272; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26274 = 10'h219 == _T_375[9:0] ? 4'h8 : _GEN_26273; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26275 = 10'h21a == _T_375[9:0] ? 4'h7 : _GEN_26274; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26276 = 10'h21b == _T_375[9:0] ? 4'h8 : _GEN_26275; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26277 = 10'h21c == _T_375[9:0] ? 4'ha : _GEN_26276; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26278 = 10'h21d == _T_375[9:0] ? 4'ha : _GEN_26277; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26279 = 10'h21e == _T_375[9:0] ? 4'h7 : _GEN_26278; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26280 = 10'h21f == _T_375[9:0] ? 4'h6 : _GEN_26279; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26281 = 10'h220 == _T_375[9:0] ? 4'h6 : _GEN_26280; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26282 = 10'h221 == _T_375[9:0] ? 4'h7 : _GEN_26281; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26283 = 10'h222 == _T_375[9:0] ? 4'ha : _GEN_26282; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26284 = 10'h223 == _T_375[9:0] ? 4'ha : _GEN_26283; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26285 = 10'h224 == _T_375[9:0] ? 4'ha : _GEN_26284; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26286 = 10'h225 == _T_375[9:0] ? 4'h8 : _GEN_26285; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26287 = 10'h226 == _T_375[9:0] ? 4'h3 : _GEN_26286; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26288 = 10'h227 == _T_375[9:0] ? 4'h4 : _GEN_26287; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26289 = 10'h228 == _T_375[9:0] ? 4'h6 : _GEN_26288; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26290 = 10'h229 == _T_375[9:0] ? 4'h6 : _GEN_26289; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26291 = 10'h22a == _T_375[9:0] ? 4'h6 : _GEN_26290; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26292 = 10'h22b == _T_375[9:0] ? 4'h6 : _GEN_26291; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26293 = 10'h22c == _T_375[9:0] ? 4'h5 : _GEN_26292; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26294 = 10'h22d == _T_375[9:0] ? 4'h6 : _GEN_26293; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26295 = 10'h22e == _T_375[9:0] ? 4'h6 : _GEN_26294; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26296 = 10'h22f == _T_375[9:0] ? 4'h8 : _GEN_26295; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26297 = 10'h230 == _T_375[9:0] ? 4'h7 : _GEN_26296; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26298 = 10'h231 == _T_375[9:0] ? 4'h5 : _GEN_26297; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26299 = 10'h232 == _T_375[9:0] ? 4'h6 : _GEN_26298; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26300 = 10'h233 == _T_375[9:0] ? 4'h8 : _GEN_26299; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26301 = 10'h234 == _T_375[9:0] ? 4'h8 : _GEN_26300; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26302 = 10'h235 == _T_375[9:0] ? 4'h8 : _GEN_26301; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26303 = 10'h236 == _T_375[9:0] ? 4'h8 : _GEN_26302; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26304 = 10'h237 == _T_375[9:0] ? 4'h8 : _GEN_26303; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26305 = 10'h238 == _T_375[9:0] ? 4'h8 : _GEN_26304; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26306 = 10'h239 == _T_375[9:0] ? 4'h6 : _GEN_26305; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26307 = 10'h23a == _T_375[9:0] ? 4'h6 : _GEN_26306; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26308 = 10'h23b == _T_375[9:0] ? 4'h7 : _GEN_26307; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26309 = 10'h23c == _T_375[9:0] ? 4'h6 : _GEN_26308; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26310 = 10'h23d == _T_375[9:0] ? 4'h7 : _GEN_26309; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26311 = 10'h23e == _T_375[9:0] ? 4'h7 : _GEN_26310; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26312 = 10'h23f == _T_375[9:0] ? 4'h6 : _GEN_26311; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26313 = 10'h240 == _T_375[9:0] ? 4'h6 : _GEN_26312; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26314 = 10'h241 == _T_375[9:0] ? 4'h8 : _GEN_26313; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26315 = 10'h242 == _T_375[9:0] ? 4'ha : _GEN_26314; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26316 = 10'h243 == _T_375[9:0] ? 4'ha : _GEN_26315; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26317 = 10'h244 == _T_375[9:0] ? 4'ha : _GEN_26316; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26318 = 10'h245 == _T_375[9:0] ? 4'h8 : _GEN_26317; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26319 = 10'h246 == _T_375[9:0] ? 4'h8 : _GEN_26318; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26320 = 10'h247 == _T_375[9:0] ? 4'h9 : _GEN_26319; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26321 = 10'h248 == _T_375[9:0] ? 4'ha : _GEN_26320; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26322 = 10'h249 == _T_375[9:0] ? 4'ha : _GEN_26321; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26323 = 10'h24a == _T_375[9:0] ? 4'ha : _GEN_26322; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26324 = 10'h24b == _T_375[9:0] ? 4'h4 : _GEN_26323; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26325 = 10'h24c == _T_375[9:0] ? 4'h3 : _GEN_26324; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26326 = 10'h24d == _T_375[9:0] ? 4'h4 : _GEN_26325; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26327 = 10'h24e == _T_375[9:0] ? 4'h5 : _GEN_26326; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26328 = 10'h24f == _T_375[9:0] ? 4'h5 : _GEN_26327; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26329 = 10'h250 == _T_375[9:0] ? 4'h5 : _GEN_26328; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26330 = 10'h251 == _T_375[9:0] ? 4'h5 : _GEN_26329; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26331 = 10'h252 == _T_375[9:0] ? 4'h5 : _GEN_26330; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26332 = 10'h253 == _T_375[9:0] ? 4'h5 : _GEN_26331; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26333 = 10'h254 == _T_375[9:0] ? 4'h5 : _GEN_26332; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26334 = 10'h255 == _T_375[9:0] ? 4'h6 : _GEN_26333; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26335 = 10'h256 == _T_375[9:0] ? 4'h7 : _GEN_26334; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26336 = 10'h257 == _T_375[9:0] ? 4'h3 : _GEN_26335; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26337 = 10'h258 == _T_375[9:0] ? 4'h6 : _GEN_26336; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26338 = 10'h259 == _T_375[9:0] ? 4'h7 : _GEN_26337; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26339 = 10'h25a == _T_375[9:0] ? 4'h7 : _GEN_26338; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26340 = 10'h25b == _T_375[9:0] ? 4'h7 : _GEN_26339; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26341 = 10'h25c == _T_375[9:0] ? 4'h8 : _GEN_26340; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26342 = 10'h25d == _T_375[9:0] ? 4'h8 : _GEN_26341; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26343 = 10'h25e == _T_375[9:0] ? 4'h4 : _GEN_26342; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26344 = 10'h25f == _T_375[9:0] ? 4'h3 : _GEN_26343; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26345 = 10'h260 == _T_375[9:0] ? 4'h7 : _GEN_26344; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26346 = 10'h261 == _T_375[9:0] ? 4'h7 : _GEN_26345; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26347 = 10'h262 == _T_375[9:0] ? 4'h7 : _GEN_26346; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26348 = 10'h263 == _T_375[9:0] ? 4'h6 : _GEN_26347; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26349 = 10'h264 == _T_375[9:0] ? 4'h7 : _GEN_26348; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26350 = 10'h265 == _T_375[9:0] ? 4'h6 : _GEN_26349; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26351 = 10'h266 == _T_375[9:0] ? 4'h5 : _GEN_26350; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26352 = 10'h267 == _T_375[9:0] ? 4'h7 : _GEN_26351; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26353 = 10'h268 == _T_375[9:0] ? 4'ha : _GEN_26352; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26354 = 10'h269 == _T_375[9:0] ? 4'ha : _GEN_26353; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26355 = 10'h26a == _T_375[9:0] ? 4'ha : _GEN_26354; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26356 = 10'h26b == _T_375[9:0] ? 4'ha : _GEN_26355; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26357 = 10'h26c == _T_375[9:0] ? 4'ha : _GEN_26356; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26358 = 10'h26d == _T_375[9:0] ? 4'ha : _GEN_26357; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26359 = 10'h26e == _T_375[9:0] ? 4'ha : _GEN_26358; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26360 = 10'h26f == _T_375[9:0] ? 4'ha : _GEN_26359; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26361 = 10'h270 == _T_375[9:0] ? 4'h5 : _GEN_26360; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26362 = 10'h271 == _T_375[9:0] ? 4'h3 : _GEN_26361; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26363 = 10'h272 == _T_375[9:0] ? 4'h3 : _GEN_26362; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26364 = 10'h273 == _T_375[9:0] ? 4'h4 : _GEN_26363; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26365 = 10'h274 == _T_375[9:0] ? 4'h6 : _GEN_26364; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26366 = 10'h275 == _T_375[9:0] ? 4'h5 : _GEN_26365; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26367 = 10'h276 == _T_375[9:0] ? 4'h6 : _GEN_26366; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26368 = 10'h277 == _T_375[9:0] ? 4'h5 : _GEN_26367; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26369 = 10'h278 == _T_375[9:0] ? 4'h6 : _GEN_26368; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26370 = 10'h279 == _T_375[9:0] ? 4'h6 : _GEN_26369; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26371 = 10'h27a == _T_375[9:0] ? 4'h6 : _GEN_26370; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26372 = 10'h27b == _T_375[9:0] ? 4'h8 : _GEN_26371; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26373 = 10'h27c == _T_375[9:0] ? 4'h6 : _GEN_26372; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26374 = 10'h27d == _T_375[9:0] ? 4'h2 : _GEN_26373; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26375 = 10'h27e == _T_375[9:0] ? 4'h5 : _GEN_26374; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26376 = 10'h27f == _T_375[9:0] ? 4'h7 : _GEN_26375; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26377 = 10'h280 == _T_375[9:0] ? 4'h7 : _GEN_26376; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26378 = 10'h281 == _T_375[9:0] ? 4'h8 : _GEN_26377; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26379 = 10'h282 == _T_375[9:0] ? 4'h7 : _GEN_26378; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26380 = 10'h283 == _T_375[9:0] ? 4'h3 : _GEN_26379; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26381 = 10'h284 == _T_375[9:0] ? 4'h3 : _GEN_26380; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26382 = 10'h285 == _T_375[9:0] ? 4'h3 : _GEN_26381; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26383 = 10'h286 == _T_375[9:0] ? 4'h7 : _GEN_26382; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26384 = 10'h287 == _T_375[9:0] ? 4'h7 : _GEN_26383; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26385 = 10'h288 == _T_375[9:0] ? 4'h7 : _GEN_26384; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26386 = 10'h289 == _T_375[9:0] ? 4'h7 : _GEN_26385; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26387 = 10'h28a == _T_375[9:0] ? 4'h8 : _GEN_26386; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26388 = 10'h28b == _T_375[9:0] ? 4'h8 : _GEN_26387; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26389 = 10'h28c == _T_375[9:0] ? 4'h7 : _GEN_26388; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26390 = 10'h28d == _T_375[9:0] ? 4'h6 : _GEN_26389; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26391 = 10'h28e == _T_375[9:0] ? 4'h3 : _GEN_26390; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26392 = 10'h28f == _T_375[9:0] ? 4'h6 : _GEN_26391; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26393 = 10'h290 == _T_375[9:0] ? 4'h8 : _GEN_26392; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26394 = 10'h291 == _T_375[9:0] ? 4'ha : _GEN_26393; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26395 = 10'h292 == _T_375[9:0] ? 4'ha : _GEN_26394; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26396 = 10'h293 == _T_375[9:0] ? 4'ha : _GEN_26395; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26397 = 10'h294 == _T_375[9:0] ? 4'h9 : _GEN_26396; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26398 = 10'h295 == _T_375[9:0] ? 4'h4 : _GEN_26397; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26399 = 10'h296 == _T_375[9:0] ? 4'h3 : _GEN_26398; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26400 = 10'h297 == _T_375[9:0] ? 4'h3 : _GEN_26399; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26401 = 10'h298 == _T_375[9:0] ? 4'h3 : _GEN_26400; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26402 = 10'h299 == _T_375[9:0] ? 4'h4 : _GEN_26401; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26403 = 10'h29a == _T_375[9:0] ? 4'h5 : _GEN_26402; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26404 = 10'h29b == _T_375[9:0] ? 4'h5 : _GEN_26403; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26405 = 10'h29c == _T_375[9:0] ? 4'h5 : _GEN_26404; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26406 = 10'h29d == _T_375[9:0] ? 4'h5 : _GEN_26405; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26407 = 10'h29e == _T_375[9:0] ? 4'h5 : _GEN_26406; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26408 = 10'h29f == _T_375[9:0] ? 4'h5 : _GEN_26407; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26409 = 10'h2a0 == _T_375[9:0] ? 4'h6 : _GEN_26408; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26410 = 10'h2a1 == _T_375[9:0] ? 4'h7 : _GEN_26409; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26411 = 10'h2a2 == _T_375[9:0] ? 4'h5 : _GEN_26410; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26412 = 10'h2a3 == _T_375[9:0] ? 4'h2 : _GEN_26411; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26413 = 10'h2a4 == _T_375[9:0] ? 4'h3 : _GEN_26412; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26414 = 10'h2a5 == _T_375[9:0] ? 4'h7 : _GEN_26413; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26415 = 10'h2a6 == _T_375[9:0] ? 4'h8 : _GEN_26414; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26416 = 10'h2a7 == _T_375[9:0] ? 4'h7 : _GEN_26415; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26417 = 10'h2a8 == _T_375[9:0] ? 4'h3 : _GEN_26416; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26418 = 10'h2a9 == _T_375[9:0] ? 4'h2 : _GEN_26417; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26419 = 10'h2aa == _T_375[9:0] ? 4'h3 : _GEN_26418; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26420 = 10'h2ab == _T_375[9:0] ? 4'h3 : _GEN_26419; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26421 = 10'h2ac == _T_375[9:0] ? 4'h7 : _GEN_26420; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26422 = 10'h2ad == _T_375[9:0] ? 4'h8 : _GEN_26421; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26423 = 10'h2ae == _T_375[9:0] ? 4'h7 : _GEN_26422; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26424 = 10'h2af == _T_375[9:0] ? 4'h8 : _GEN_26423; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26425 = 10'h2b0 == _T_375[9:0] ? 4'h8 : _GEN_26424; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26426 = 10'h2b1 == _T_375[9:0] ? 4'h8 : _GEN_26425; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26427 = 10'h2b2 == _T_375[9:0] ? 4'h7 : _GEN_26426; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26428 = 10'h2b3 == _T_375[9:0] ? 4'h6 : _GEN_26427; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26429 = 10'h2b4 == _T_375[9:0] ? 4'h2 : _GEN_26428; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26430 = 10'h2b5 == _T_375[9:0] ? 4'h2 : _GEN_26429; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26431 = 10'h2b6 == _T_375[9:0] ? 4'h3 : _GEN_26430; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26432 = 10'h2b7 == _T_375[9:0] ? 4'h3 : _GEN_26431; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26433 = 10'h2b8 == _T_375[9:0] ? 4'h6 : _GEN_26432; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26434 = 10'h2b9 == _T_375[9:0] ? 4'h9 : _GEN_26433; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26435 = 10'h2ba == _T_375[9:0] ? 4'h3 : _GEN_26434; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26436 = 10'h2bb == _T_375[9:0] ? 4'h3 : _GEN_26435; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26437 = 10'h2bc == _T_375[9:0] ? 4'h3 : _GEN_26436; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26438 = 10'h2bd == _T_375[9:0] ? 4'h2 : _GEN_26437; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26439 = 10'h2be == _T_375[9:0] ? 4'h3 : _GEN_26438; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26440 = 10'h2bf == _T_375[9:0] ? 4'h3 : _GEN_26439; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26441 = 10'h2c0 == _T_375[9:0] ? 4'h5 : _GEN_26440; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26442 = 10'h2c1 == _T_375[9:0] ? 4'h5 : _GEN_26441; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26443 = 10'h2c2 == _T_375[9:0] ? 4'h5 : _GEN_26442; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26444 = 10'h2c3 == _T_375[9:0] ? 4'h5 : _GEN_26443; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26445 = 10'h2c4 == _T_375[9:0] ? 4'h5 : _GEN_26444; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26446 = 10'h2c5 == _T_375[9:0] ? 4'h5 : _GEN_26445; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26447 = 10'h2c6 == _T_375[9:0] ? 4'h6 : _GEN_26446; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26448 = 10'h2c7 == _T_375[9:0] ? 4'h7 : _GEN_26447; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26449 = 10'h2c8 == _T_375[9:0] ? 4'h5 : _GEN_26448; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26450 = 10'h2c9 == _T_375[9:0] ? 4'h2 : _GEN_26449; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26451 = 10'h2ca == _T_375[9:0] ? 4'h2 : _GEN_26450; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26452 = 10'h2cb == _T_375[9:0] ? 4'h3 : _GEN_26451; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26453 = 10'h2cc == _T_375[9:0] ? 4'h3 : _GEN_26452; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26454 = 10'h2cd == _T_375[9:0] ? 4'h2 : _GEN_26453; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26455 = 10'h2ce == _T_375[9:0] ? 4'h2 : _GEN_26454; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26456 = 10'h2cf == _T_375[9:0] ? 4'h2 : _GEN_26455; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26457 = 10'h2d0 == _T_375[9:0] ? 4'h2 : _GEN_26456; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26458 = 10'h2d1 == _T_375[9:0] ? 4'h2 : _GEN_26457; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26459 = 10'h2d2 == _T_375[9:0] ? 4'h7 : _GEN_26458; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26460 = 10'h2d3 == _T_375[9:0] ? 4'h7 : _GEN_26459; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26461 = 10'h2d4 == _T_375[9:0] ? 4'h8 : _GEN_26460; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26462 = 10'h2d5 == _T_375[9:0] ? 4'h8 : _GEN_26461; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26463 = 10'h2d6 == _T_375[9:0] ? 4'h8 : _GEN_26462; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26464 = 10'h2d7 == _T_375[9:0] ? 4'h8 : _GEN_26463; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26465 = 10'h2d8 == _T_375[9:0] ? 4'h7 : _GEN_26464; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26466 = 10'h2d9 == _T_375[9:0] ? 4'h6 : _GEN_26465; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26467 = 10'h2da == _T_375[9:0] ? 4'h4 : _GEN_26466; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26468 = 10'h2db == _T_375[9:0] ? 4'h2 : _GEN_26467; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26469 = 10'h2dc == _T_375[9:0] ? 4'h2 : _GEN_26468; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26470 = 10'h2dd == _T_375[9:0] ? 4'h3 : _GEN_26469; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26471 = 10'h2de == _T_375[9:0] ? 4'h3 : _GEN_26470; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26472 = 10'h2df == _T_375[9:0] ? 4'h3 : _GEN_26471; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26473 = 10'h2e0 == _T_375[9:0] ? 4'h3 : _GEN_26472; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26474 = 10'h2e1 == _T_375[9:0] ? 4'h3 : _GEN_26473; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26475 = 10'h2e2 == _T_375[9:0] ? 4'h3 : _GEN_26474; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26476 = 10'h2e3 == _T_375[9:0] ? 4'h2 : _GEN_26475; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26477 = 10'h2e4 == _T_375[9:0] ? 4'h3 : _GEN_26476; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26478 = 10'h2e5 == _T_375[9:0] ? 4'h2 : _GEN_26477; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26479 = 10'h2e6 == _T_375[9:0] ? 4'h5 : _GEN_26478; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26480 = 10'h2e7 == _T_375[9:0] ? 4'h5 : _GEN_26479; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26481 = 10'h2e8 == _T_375[9:0] ? 4'h5 : _GEN_26480; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26482 = 10'h2e9 == _T_375[9:0] ? 4'h5 : _GEN_26481; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26483 = 10'h2ea == _T_375[9:0] ? 4'h5 : _GEN_26482; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26484 = 10'h2eb == _T_375[9:0] ? 4'h5 : _GEN_26483; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26485 = 10'h2ec == _T_375[9:0] ? 4'h6 : _GEN_26484; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26486 = 10'h2ed == _T_375[9:0] ? 4'h7 : _GEN_26485; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26487 = 10'h2ee == _T_375[9:0] ? 4'h6 : _GEN_26486; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26488 = 10'h2ef == _T_375[9:0] ? 4'h2 : _GEN_26487; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26489 = 10'h2f0 == _T_375[9:0] ? 4'h2 : _GEN_26488; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26490 = 10'h2f1 == _T_375[9:0] ? 4'h2 : _GEN_26489; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26491 = 10'h2f2 == _T_375[9:0] ? 4'h2 : _GEN_26490; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26492 = 10'h2f3 == _T_375[9:0] ? 4'h2 : _GEN_26491; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26493 = 10'h2f4 == _T_375[9:0] ? 4'h2 : _GEN_26492; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26494 = 10'h2f5 == _T_375[9:0] ? 4'h2 : _GEN_26493; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26495 = 10'h2f6 == _T_375[9:0] ? 4'h2 : _GEN_26494; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26496 = 10'h2f7 == _T_375[9:0] ? 4'h2 : _GEN_26495; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26497 = 10'h2f8 == _T_375[9:0] ? 4'h7 : _GEN_26496; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26498 = 10'h2f9 == _T_375[9:0] ? 4'h7 : _GEN_26497; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26499 = 10'h2fa == _T_375[9:0] ? 4'h8 : _GEN_26498; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26500 = 10'h2fb == _T_375[9:0] ? 4'h8 : _GEN_26499; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26501 = 10'h2fc == _T_375[9:0] ? 4'h7 : _GEN_26500; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26502 = 10'h2fd == _T_375[9:0] ? 4'h7 : _GEN_26501; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26503 = 10'h2fe == _T_375[9:0] ? 4'h7 : _GEN_26502; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26504 = 10'h2ff == _T_375[9:0] ? 4'h7 : _GEN_26503; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26505 = 10'h300 == _T_375[9:0] ? 4'h8 : _GEN_26504; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26506 = 10'h301 == _T_375[9:0] ? 4'h7 : _GEN_26505; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26507 = 10'h302 == _T_375[9:0] ? 4'h3 : _GEN_26506; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26508 = 10'h303 == _T_375[9:0] ? 4'h3 : _GEN_26507; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26509 = 10'h304 == _T_375[9:0] ? 4'h2 : _GEN_26508; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26510 = 10'h305 == _T_375[9:0] ? 4'h2 : _GEN_26509; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26511 = 10'h306 == _T_375[9:0] ? 4'h2 : _GEN_26510; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26512 = 10'h307 == _T_375[9:0] ? 4'h2 : _GEN_26511; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26513 = 10'h308 == _T_375[9:0] ? 4'h2 : _GEN_26512; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26514 = 10'h309 == _T_375[9:0] ? 4'h2 : _GEN_26513; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26515 = 10'h30a == _T_375[9:0] ? 4'h2 : _GEN_26514; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26516 = 10'h30b == _T_375[9:0] ? 4'h3 : _GEN_26515; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26517 = 10'h30c == _T_375[9:0] ? 4'h4 : _GEN_26516; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26518 = 10'h30d == _T_375[9:0] ? 4'h5 : _GEN_26517; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26519 = 10'h30e == _T_375[9:0] ? 4'h5 : _GEN_26518; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26520 = 10'h30f == _T_375[9:0] ? 4'h5 : _GEN_26519; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26521 = 10'h310 == _T_375[9:0] ? 4'h5 : _GEN_26520; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26522 = 10'h311 == _T_375[9:0] ? 4'h5 : _GEN_26521; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26523 = 10'h312 == _T_375[9:0] ? 4'h6 : _GEN_26522; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26524 = 10'h313 == _T_375[9:0] ? 4'h7 : _GEN_26523; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26525 = 10'h314 == _T_375[9:0] ? 4'h7 : _GEN_26524; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26526 = 10'h315 == _T_375[9:0] ? 4'h3 : _GEN_26525; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26527 = 10'h316 == _T_375[9:0] ? 4'h2 : _GEN_26526; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26528 = 10'h317 == _T_375[9:0] ? 4'h2 : _GEN_26527; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26529 = 10'h318 == _T_375[9:0] ? 4'h2 : _GEN_26528; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26530 = 10'h319 == _T_375[9:0] ? 4'h2 : _GEN_26529; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26531 = 10'h31a == _T_375[9:0] ? 4'h2 : _GEN_26530; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26532 = 10'h31b == _T_375[9:0] ? 4'h2 : _GEN_26531; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26533 = 10'h31c == _T_375[9:0] ? 4'h2 : _GEN_26532; // @[Filter.scala 230:142]
  wire [3:0] _GEN_26534 = 10'h31d == _T_375[9:0] ? 4'h2 : _GEN_26533; // @[Filter.scala 230:142]
  wire [7:0] _T_389 = _GEN_26534 * 4'ha; // @[Filter.scala 230:142]
  wire [10:0] _GEN_39019 = {{3'd0}, _T_389}; // @[Filter.scala 230:109]
  wire [10:0] _T_391 = _T_384 + _GEN_39019; // @[Filter.scala 230:109]
  wire [10:0] _T_392 = _T_391 / 11'h64; // @[Filter.scala 230:150]
  wire  _T_394 = _T_365 >= 6'h20; // @[Filter.scala 233:31]
  wire  _T_398 = _T_372 >= 32'h12; // @[Filter.scala 233:63]
  wire  _T_399 = _T_394 | _T_398; // @[Filter.scala 233:58]
  wire [10:0] _GEN_27333 = io_SPI_distort ? _T_392 : {{7'd0}, _GEN_24938}; // @[Filter.scala 235:35]
  wire [10:0] _GEN_27334 = _T_399 ? 11'h0 : _GEN_27333; // @[Filter.scala 233:80]
  wire [10:0] _GEN_28133 = io_SPI_distort ? _T_392 : {{7'd0}, _GEN_25736}; // @[Filter.scala 235:35]
  wire [10:0] _GEN_28134 = _T_399 ? 11'h0 : _GEN_28133; // @[Filter.scala 233:80]
  wire [10:0] _GEN_28933 = io_SPI_distort ? _T_392 : {{7'd0}, _GEN_26534}; // @[Filter.scala 235:35]
  wire [10:0] _GEN_28934 = _T_399 ? 11'h0 : _GEN_28933; // @[Filter.scala 233:80]
  wire [31:0] _T_427 = pixelIndex + 32'h6; // @[Filter.scala 228:31]
  wire [31:0] _GEN_6 = _T_427 % 32'h20; // @[Filter.scala 228:38]
  wire [5:0] _T_428 = _GEN_6[5:0]; // @[Filter.scala 228:38]
  wire [5:0] _T_430 = _T_428 + _GEN_38951; // @[Filter.scala 228:53]
  wire [5:0] _T_432 = _T_430 - 6'h1; // @[Filter.scala 228:69]
  wire [31:0] _T_435 = _T_427 / 32'h20; // @[Filter.scala 229:38]
  wire [31:0] _T_437 = _T_435 + _GEN_38952; // @[Filter.scala 229:53]
  wire [31:0] _T_439 = _T_437 - 32'h1; // @[Filter.scala 229:69]
  wire [37:0] _T_440 = _T_439 * 32'h20; // @[Filter.scala 230:42]
  wire [37:0] _GEN_39025 = {{32'd0}, _T_432}; // @[Filter.scala 230:57]
  wire [37:0] _T_442 = _T_440 + _GEN_39025; // @[Filter.scala 230:57]
  wire [3:0] _GEN_28957 = 10'h16 == _T_442[9:0] ? 4'h9 : 4'ha; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28958 = 10'h17 == _T_442[9:0] ? 4'h3 : _GEN_28957; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28959 = 10'h18 == _T_442[9:0] ? 4'h6 : _GEN_28958; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28960 = 10'h19 == _T_442[9:0] ? 4'ha : _GEN_28959; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28961 = 10'h1a == _T_442[9:0] ? 4'ha : _GEN_28960; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28962 = 10'h1b == _T_442[9:0] ? 4'ha : _GEN_28961; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28963 = 10'h1c == _T_442[9:0] ? 4'ha : _GEN_28962; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28964 = 10'h1d == _T_442[9:0] ? 4'ha : _GEN_28963; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28965 = 10'h1e == _T_442[9:0] ? 4'ha : _GEN_28964; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28966 = 10'h1f == _T_442[9:0] ? 4'ha : _GEN_28965; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28967 = 10'h20 == _T_442[9:0] ? 4'ha : _GEN_28966; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28968 = 10'h21 == _T_442[9:0] ? 4'ha : _GEN_28967; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28969 = 10'h22 == _T_442[9:0] ? 4'ha : _GEN_28968; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28970 = 10'h23 == _T_442[9:0] ? 4'ha : _GEN_28969; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28971 = 10'h24 == _T_442[9:0] ? 4'ha : _GEN_28970; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28972 = 10'h25 == _T_442[9:0] ? 4'ha : _GEN_28971; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28973 = 10'h26 == _T_442[9:0] ? 4'ha : _GEN_28972; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28974 = 10'h27 == _T_442[9:0] ? 4'ha : _GEN_28973; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28975 = 10'h28 == _T_442[9:0] ? 4'ha : _GEN_28974; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28976 = 10'h29 == _T_442[9:0] ? 4'ha : _GEN_28975; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28977 = 10'h2a == _T_442[9:0] ? 4'ha : _GEN_28976; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28978 = 10'h2b == _T_442[9:0] ? 4'ha : _GEN_28977; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28979 = 10'h2c == _T_442[9:0] ? 4'ha : _GEN_28978; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28980 = 10'h2d == _T_442[9:0] ? 4'ha : _GEN_28979; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28981 = 10'h2e == _T_442[9:0] ? 4'ha : _GEN_28980; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28982 = 10'h2f == _T_442[9:0] ? 4'ha : _GEN_28981; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28983 = 10'h30 == _T_442[9:0] ? 4'ha : _GEN_28982; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28984 = 10'h31 == _T_442[9:0] ? 4'ha : _GEN_28983; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28985 = 10'h32 == _T_442[9:0] ? 4'ha : _GEN_28984; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28986 = 10'h33 == _T_442[9:0] ? 4'ha : _GEN_28985; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28987 = 10'h34 == _T_442[9:0] ? 4'ha : _GEN_28986; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28988 = 10'h35 == _T_442[9:0] ? 4'ha : _GEN_28987; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28989 = 10'h36 == _T_442[9:0] ? 4'ha : _GEN_28988; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28990 = 10'h37 == _T_442[9:0] ? 4'ha : _GEN_28989; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28991 = 10'h38 == _T_442[9:0] ? 4'ha : _GEN_28990; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28992 = 10'h39 == _T_442[9:0] ? 4'ha : _GEN_28991; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28993 = 10'h3a == _T_442[9:0] ? 4'ha : _GEN_28992; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28994 = 10'h3b == _T_442[9:0] ? 4'h9 : _GEN_28993; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28995 = 10'h3c == _T_442[9:0] ? 4'h4 : _GEN_28994; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28996 = 10'h3d == _T_442[9:0] ? 4'h3 : _GEN_28995; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28997 = 10'h3e == _T_442[9:0] ? 4'h4 : _GEN_28996; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28998 = 10'h3f == _T_442[9:0] ? 4'ha : _GEN_28997; // @[Filter.scala 230:62]
  wire [3:0] _GEN_28999 = 10'h40 == _T_442[9:0] ? 4'ha : _GEN_28998; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29000 = 10'h41 == _T_442[9:0] ? 4'ha : _GEN_28999; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29001 = 10'h42 == _T_442[9:0] ? 4'ha : _GEN_29000; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29002 = 10'h43 == _T_442[9:0] ? 4'ha : _GEN_29001; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29003 = 10'h44 == _T_442[9:0] ? 4'ha : _GEN_29002; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29004 = 10'h45 == _T_442[9:0] ? 4'ha : _GEN_29003; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29005 = 10'h46 == _T_442[9:0] ? 4'ha : _GEN_29004; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29006 = 10'h47 == _T_442[9:0] ? 4'ha : _GEN_29005; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29007 = 10'h48 == _T_442[9:0] ? 4'ha : _GEN_29006; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29008 = 10'h49 == _T_442[9:0] ? 4'ha : _GEN_29007; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29009 = 10'h4a == _T_442[9:0] ? 4'ha : _GEN_29008; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29010 = 10'h4b == _T_442[9:0] ? 4'ha : _GEN_29009; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29011 = 10'h4c == _T_442[9:0] ? 4'ha : _GEN_29010; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29012 = 10'h4d == _T_442[9:0] ? 4'ha : _GEN_29011; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29013 = 10'h4e == _T_442[9:0] ? 4'ha : _GEN_29012; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29014 = 10'h4f == _T_442[9:0] ? 4'ha : _GEN_29013; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29015 = 10'h50 == _T_442[9:0] ? 4'ha : _GEN_29014; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29016 = 10'h51 == _T_442[9:0] ? 4'ha : _GEN_29015; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29017 = 10'h52 == _T_442[9:0] ? 4'ha : _GEN_29016; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29018 = 10'h53 == _T_442[9:0] ? 4'ha : _GEN_29017; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29019 = 10'h54 == _T_442[9:0] ? 4'ha : _GEN_29018; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29020 = 10'h55 == _T_442[9:0] ? 4'ha : _GEN_29019; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29021 = 10'h56 == _T_442[9:0] ? 4'ha : _GEN_29020; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29022 = 10'h57 == _T_442[9:0] ? 4'ha : _GEN_29021; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29023 = 10'h58 == _T_442[9:0] ? 4'ha : _GEN_29022; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29024 = 10'h59 == _T_442[9:0] ? 4'ha : _GEN_29023; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29025 = 10'h5a == _T_442[9:0] ? 4'h7 : _GEN_29024; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29026 = 10'h5b == _T_442[9:0] ? 4'h7 : _GEN_29025; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29027 = 10'h5c == _T_442[9:0] ? 4'ha : _GEN_29026; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29028 = 10'h5d == _T_442[9:0] ? 4'ha : _GEN_29027; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29029 = 10'h5e == _T_442[9:0] ? 4'ha : _GEN_29028; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29030 = 10'h5f == _T_442[9:0] ? 4'ha : _GEN_29029; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29031 = 10'h60 == _T_442[9:0] ? 4'ha : _GEN_29030; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29032 = 10'h61 == _T_442[9:0] ? 4'h8 : _GEN_29031; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29033 = 10'h62 == _T_442[9:0] ? 4'h3 : _GEN_29032; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29034 = 10'h63 == _T_442[9:0] ? 4'h3 : _GEN_29033; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29035 = 10'h64 == _T_442[9:0] ? 4'h3 : _GEN_29034; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29036 = 10'h65 == _T_442[9:0] ? 4'h9 : _GEN_29035; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29037 = 10'h66 == _T_442[9:0] ? 4'ha : _GEN_29036; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29038 = 10'h67 == _T_442[9:0] ? 4'ha : _GEN_29037; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29039 = 10'h68 == _T_442[9:0] ? 4'ha : _GEN_29038; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29040 = 10'h69 == _T_442[9:0] ? 4'ha : _GEN_29039; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29041 = 10'h6a == _T_442[9:0] ? 4'ha : _GEN_29040; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29042 = 10'h6b == _T_442[9:0] ? 4'h8 : _GEN_29041; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29043 = 10'h6c == _T_442[9:0] ? 4'h5 : _GEN_29042; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29044 = 10'h6d == _T_442[9:0] ? 4'h8 : _GEN_29043; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29045 = 10'h6e == _T_442[9:0] ? 4'ha : _GEN_29044; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29046 = 10'h6f == _T_442[9:0] ? 4'ha : _GEN_29045; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29047 = 10'h70 == _T_442[9:0] ? 4'ha : _GEN_29046; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29048 = 10'h71 == _T_442[9:0] ? 4'ha : _GEN_29047; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29049 = 10'h72 == _T_442[9:0] ? 4'ha : _GEN_29048; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29050 = 10'h73 == _T_442[9:0] ? 4'ha : _GEN_29049; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29051 = 10'h74 == _T_442[9:0] ? 4'ha : _GEN_29050; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29052 = 10'h75 == _T_442[9:0] ? 4'ha : _GEN_29051; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29053 = 10'h76 == _T_442[9:0] ? 4'ha : _GEN_29052; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29054 = 10'h77 == _T_442[9:0] ? 4'ha : _GEN_29053; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29055 = 10'h78 == _T_442[9:0] ? 4'ha : _GEN_29054; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29056 = 10'h79 == _T_442[9:0] ? 4'ha : _GEN_29055; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29057 = 10'h7a == _T_442[9:0] ? 4'ha : _GEN_29056; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29058 = 10'h7b == _T_442[9:0] ? 4'ha : _GEN_29057; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29059 = 10'h7c == _T_442[9:0] ? 4'ha : _GEN_29058; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29060 = 10'h7d == _T_442[9:0] ? 4'ha : _GEN_29059; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29061 = 10'h7e == _T_442[9:0] ? 4'ha : _GEN_29060; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29062 = 10'h7f == _T_442[9:0] ? 4'ha : _GEN_29061; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29063 = 10'h80 == _T_442[9:0] ? 4'ha : _GEN_29062; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29064 = 10'h81 == _T_442[9:0] ? 4'h5 : _GEN_29063; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29065 = 10'h82 == _T_442[9:0] ? 4'h5 : _GEN_29064; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29066 = 10'h83 == _T_442[9:0] ? 4'h7 : _GEN_29065; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29067 = 10'h84 == _T_442[9:0] ? 4'ha : _GEN_29066; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29068 = 10'h85 == _T_442[9:0] ? 4'ha : _GEN_29067; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29069 = 10'h86 == _T_442[9:0] ? 4'ha : _GEN_29068; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29070 = 10'h87 == _T_442[9:0] ? 4'h5 : _GEN_29069; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29071 = 10'h88 == _T_442[9:0] ? 4'h3 : _GEN_29070; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29072 = 10'h89 == _T_442[9:0] ? 4'h3 : _GEN_29071; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29073 = 10'h8a == _T_442[9:0] ? 4'h4 : _GEN_29072; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29074 = 10'h8b == _T_442[9:0] ? 4'h9 : _GEN_29073; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29075 = 10'h8c == _T_442[9:0] ? 4'ha : _GEN_29074; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29076 = 10'h8d == _T_442[9:0] ? 4'ha : _GEN_29075; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29077 = 10'h8e == _T_442[9:0] ? 4'ha : _GEN_29076; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29078 = 10'h8f == _T_442[9:0] ? 4'h6 : _GEN_29077; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29079 = 10'h90 == _T_442[9:0] ? 4'h4 : _GEN_29078; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29080 = 10'h91 == _T_442[9:0] ? 4'h3 : _GEN_29079; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29081 = 10'h92 == _T_442[9:0] ? 4'h7 : _GEN_29080; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29082 = 10'h93 == _T_442[9:0] ? 4'ha : _GEN_29081; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29083 = 10'h94 == _T_442[9:0] ? 4'ha : _GEN_29082; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29084 = 10'h95 == _T_442[9:0] ? 4'ha : _GEN_29083; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29085 = 10'h96 == _T_442[9:0] ? 4'ha : _GEN_29084; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29086 = 10'h97 == _T_442[9:0] ? 4'ha : _GEN_29085; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29087 = 10'h98 == _T_442[9:0] ? 4'ha : _GEN_29086; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29088 = 10'h99 == _T_442[9:0] ? 4'ha : _GEN_29087; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29089 = 10'h9a == _T_442[9:0] ? 4'ha : _GEN_29088; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29090 = 10'h9b == _T_442[9:0] ? 4'ha : _GEN_29089; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29091 = 10'h9c == _T_442[9:0] ? 4'ha : _GEN_29090; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29092 = 10'h9d == _T_442[9:0] ? 4'ha : _GEN_29091; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29093 = 10'h9e == _T_442[9:0] ? 4'ha : _GEN_29092; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29094 = 10'h9f == _T_442[9:0] ? 4'ha : _GEN_29093; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29095 = 10'ha0 == _T_442[9:0] ? 4'ha : _GEN_29094; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29096 = 10'ha1 == _T_442[9:0] ? 4'ha : _GEN_29095; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29097 = 10'ha2 == _T_442[9:0] ? 4'ha : _GEN_29096; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29098 = 10'ha3 == _T_442[9:0] ? 4'ha : _GEN_29097; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29099 = 10'ha4 == _T_442[9:0] ? 4'ha : _GEN_29098; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29100 = 10'ha5 == _T_442[9:0] ? 4'ha : _GEN_29099; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29101 = 10'ha6 == _T_442[9:0] ? 4'ha : _GEN_29100; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29102 = 10'ha7 == _T_442[9:0] ? 4'h9 : _GEN_29101; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29103 = 10'ha8 == _T_442[9:0] ? 4'h4 : _GEN_29102; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29104 = 10'ha9 == _T_442[9:0] ? 4'h3 : _GEN_29103; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29105 = 10'haa == _T_442[9:0] ? 4'h4 : _GEN_29104; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29106 = 10'hab == _T_442[9:0] ? 4'h7 : _GEN_29105; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29107 = 10'hac == _T_442[9:0] ? 4'h8 : _GEN_29106; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29108 = 10'had == _T_442[9:0] ? 4'h3 : _GEN_29107; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29109 = 10'hae == _T_442[9:0] ? 4'h3 : _GEN_29108; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29110 = 10'haf == _T_442[9:0] ? 4'h3 : _GEN_29109; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29111 = 10'hb0 == _T_442[9:0] ? 4'h3 : _GEN_29110; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29112 = 10'hb1 == _T_442[9:0] ? 4'h7 : _GEN_29111; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29113 = 10'hb2 == _T_442[9:0] ? 4'h9 : _GEN_29112; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29114 = 10'hb3 == _T_442[9:0] ? 4'h6 : _GEN_29113; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29115 = 10'hb4 == _T_442[9:0] ? 4'h4 : _GEN_29114; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29116 = 10'hb5 == _T_442[9:0] ? 4'h3 : _GEN_29115; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29117 = 10'hb6 == _T_442[9:0] ? 4'h3 : _GEN_29116; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29118 = 10'hb7 == _T_442[9:0] ? 4'h6 : _GEN_29117; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29119 = 10'hb8 == _T_442[9:0] ? 4'ha : _GEN_29118; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29120 = 10'hb9 == _T_442[9:0] ? 4'ha : _GEN_29119; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29121 = 10'hba == _T_442[9:0] ? 4'ha : _GEN_29120; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29122 = 10'hbb == _T_442[9:0] ? 4'ha : _GEN_29121; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29123 = 10'hbc == _T_442[9:0] ? 4'ha : _GEN_29122; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29124 = 10'hbd == _T_442[9:0] ? 4'h9 : _GEN_29123; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29125 = 10'hbe == _T_442[9:0] ? 4'ha : _GEN_29124; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29126 = 10'hbf == _T_442[9:0] ? 4'ha : _GEN_29125; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29127 = 10'hc0 == _T_442[9:0] ? 4'ha : _GEN_29126; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29128 = 10'hc1 == _T_442[9:0] ? 4'ha : _GEN_29127; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29129 = 10'hc2 == _T_442[9:0] ? 4'ha : _GEN_29128; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29130 = 10'hc3 == _T_442[9:0] ? 4'ha : _GEN_29129; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29131 = 10'hc4 == _T_442[9:0] ? 4'ha : _GEN_29130; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29132 = 10'hc5 == _T_442[9:0] ? 4'ha : _GEN_29131; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29133 = 10'hc6 == _T_442[9:0] ? 4'ha : _GEN_29132; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29134 = 10'hc7 == _T_442[9:0] ? 4'h9 : _GEN_29133; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29135 = 10'hc8 == _T_442[9:0] ? 4'h8 : _GEN_29134; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29136 = 10'hc9 == _T_442[9:0] ? 4'h8 : _GEN_29135; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29137 = 10'hca == _T_442[9:0] ? 4'h9 : _GEN_29136; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29138 = 10'hcb == _T_442[9:0] ? 4'ha : _GEN_29137; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29139 = 10'hcc == _T_442[9:0] ? 4'ha : _GEN_29138; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29140 = 10'hcd == _T_442[9:0] ? 4'ha : _GEN_29139; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29141 = 10'hce == _T_442[9:0] ? 4'h8 : _GEN_29140; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29142 = 10'hcf == _T_442[9:0] ? 4'h3 : _GEN_29141; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29143 = 10'hd0 == _T_442[9:0] ? 4'h3 : _GEN_29142; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29144 = 10'hd1 == _T_442[9:0] ? 4'h3 : _GEN_29143; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29145 = 10'hd2 == _T_442[9:0] ? 4'h4 : _GEN_29144; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29146 = 10'hd3 == _T_442[9:0] ? 4'h3 : _GEN_29145; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29147 = 10'hd4 == _T_442[9:0] ? 4'h3 : _GEN_29146; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29148 = 10'hd5 == _T_442[9:0] ? 4'h3 : _GEN_29147; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29149 = 10'hd6 == _T_442[9:0] ? 4'h3 : _GEN_29148; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29150 = 10'hd7 == _T_442[9:0] ? 4'h5 : _GEN_29149; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29151 = 10'hd8 == _T_442[9:0] ? 4'h4 : _GEN_29150; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29152 = 10'hd9 == _T_442[9:0] ? 4'h3 : _GEN_29151; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29153 = 10'hda == _T_442[9:0] ? 4'h3 : _GEN_29152; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29154 = 10'hdb == _T_442[9:0] ? 4'h3 : _GEN_29153; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29155 = 10'hdc == _T_442[9:0] ? 4'h4 : _GEN_29154; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29156 = 10'hdd == _T_442[9:0] ? 4'ha : _GEN_29155; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29157 = 10'hde == _T_442[9:0] ? 4'ha : _GEN_29156; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29158 = 10'hdf == _T_442[9:0] ? 4'ha : _GEN_29157; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29159 = 10'he0 == _T_442[9:0] ? 4'ha : _GEN_29158; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29160 = 10'he1 == _T_442[9:0] ? 4'ha : _GEN_29159; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29161 = 10'he2 == _T_442[9:0] ? 4'ha : _GEN_29160; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29162 = 10'he3 == _T_442[9:0] ? 4'h5 : _GEN_29161; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29163 = 10'he4 == _T_442[9:0] ? 4'ha : _GEN_29162; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29164 = 10'he5 == _T_442[9:0] ? 4'ha : _GEN_29163; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29165 = 10'he6 == _T_442[9:0] ? 4'ha : _GEN_29164; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29166 = 10'he7 == _T_442[9:0] ? 4'ha : _GEN_29165; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29167 = 10'he8 == _T_442[9:0] ? 4'ha : _GEN_29166; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29168 = 10'he9 == _T_442[9:0] ? 4'ha : _GEN_29167; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29169 = 10'hea == _T_442[9:0] ? 4'ha : _GEN_29168; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29170 = 10'heb == _T_442[9:0] ? 4'h9 : _GEN_29169; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29171 = 10'hec == _T_442[9:0] ? 4'h7 : _GEN_29170; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29172 = 10'hed == _T_442[9:0] ? 4'h3 : _GEN_29171; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29173 = 10'hee == _T_442[9:0] ? 4'h3 : _GEN_29172; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29174 = 10'hef == _T_442[9:0] ? 4'h3 : _GEN_29173; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29175 = 10'hf0 == _T_442[9:0] ? 4'h4 : _GEN_29174; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29176 = 10'hf1 == _T_442[9:0] ? 4'h7 : _GEN_29175; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29177 = 10'hf2 == _T_442[9:0] ? 4'ha : _GEN_29176; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29178 = 10'hf3 == _T_442[9:0] ? 4'ha : _GEN_29177; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29179 = 10'hf4 == _T_442[9:0] ? 4'ha : _GEN_29178; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29180 = 10'hf5 == _T_442[9:0] ? 4'h7 : _GEN_29179; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29181 = 10'hf6 == _T_442[9:0] ? 4'h3 : _GEN_29180; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29182 = 10'hf7 == _T_442[9:0] ? 4'h3 : _GEN_29181; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29183 = 10'hf8 == _T_442[9:0] ? 4'h3 : _GEN_29182; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29184 = 10'hf9 == _T_442[9:0] ? 4'h3 : _GEN_29183; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29185 = 10'hfa == _T_442[9:0] ? 4'h3 : _GEN_29184; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29186 = 10'hfb == _T_442[9:0] ? 4'h3 : _GEN_29185; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29187 = 10'hfc == _T_442[9:0] ? 4'h3 : _GEN_29186; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29188 = 10'hfd == _T_442[9:0] ? 4'h3 : _GEN_29187; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29189 = 10'hfe == _T_442[9:0] ? 4'h3 : _GEN_29188; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29190 = 10'hff == _T_442[9:0] ? 4'h3 : _GEN_29189; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29191 = 10'h100 == _T_442[9:0] ? 4'h3 : _GEN_29190; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29192 = 10'h101 == _T_442[9:0] ? 4'h4 : _GEN_29191; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29193 = 10'h102 == _T_442[9:0] ? 4'h6 : _GEN_29192; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29194 = 10'h103 == _T_442[9:0] ? 4'ha : _GEN_29193; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29195 = 10'h104 == _T_442[9:0] ? 4'ha : _GEN_29194; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29196 = 10'h105 == _T_442[9:0] ? 4'h9 : _GEN_29195; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29197 = 10'h106 == _T_442[9:0] ? 4'h9 : _GEN_29196; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29198 = 10'h107 == _T_442[9:0] ? 4'h9 : _GEN_29197; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29199 = 10'h108 == _T_442[9:0] ? 4'h9 : _GEN_29198; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29200 = 10'h109 == _T_442[9:0] ? 4'h3 : _GEN_29199; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29201 = 10'h10a == _T_442[9:0] ? 4'ha : _GEN_29200; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29202 = 10'h10b == _T_442[9:0] ? 4'ha : _GEN_29201; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29203 = 10'h10c == _T_442[9:0] ? 4'ha : _GEN_29202; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29204 = 10'h10d == _T_442[9:0] ? 4'ha : _GEN_29203; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29205 = 10'h10e == _T_442[9:0] ? 4'ha : _GEN_29204; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29206 = 10'h10f == _T_442[9:0] ? 4'h9 : _GEN_29205; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29207 = 10'h110 == _T_442[9:0] ? 4'h9 : _GEN_29206; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29208 = 10'h111 == _T_442[9:0] ? 4'h4 : _GEN_29207; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29209 = 10'h112 == _T_442[9:0] ? 4'h8 : _GEN_29208; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29210 = 10'h113 == _T_442[9:0] ? 4'h3 : _GEN_29209; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29211 = 10'h114 == _T_442[9:0] ? 4'h3 : _GEN_29210; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29212 = 10'h115 == _T_442[9:0] ? 4'h4 : _GEN_29211; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29213 = 10'h116 == _T_442[9:0] ? 4'h4 : _GEN_29212; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29214 = 10'h117 == _T_442[9:0] ? 4'h3 : _GEN_29213; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29215 = 10'h118 == _T_442[9:0] ? 4'h8 : _GEN_29214; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29216 = 10'h119 == _T_442[9:0] ? 4'ha : _GEN_29215; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29217 = 10'h11a == _T_442[9:0] ? 4'ha : _GEN_29216; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29218 = 10'h11b == _T_442[9:0] ? 4'ha : _GEN_29217; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29219 = 10'h11c == _T_442[9:0] ? 4'h6 : _GEN_29218; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29220 = 10'h11d == _T_442[9:0] ? 4'h3 : _GEN_29219; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29221 = 10'h11e == _T_442[9:0] ? 4'h3 : _GEN_29220; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29222 = 10'h11f == _T_442[9:0] ? 4'h3 : _GEN_29221; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29223 = 10'h120 == _T_442[9:0] ? 4'h3 : _GEN_29222; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29224 = 10'h121 == _T_442[9:0] ? 4'h3 : _GEN_29223; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29225 = 10'h122 == _T_442[9:0] ? 4'h3 : _GEN_29224; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29226 = 10'h123 == _T_442[9:0] ? 4'h3 : _GEN_29225; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29227 = 10'h124 == _T_442[9:0] ? 4'h3 : _GEN_29226; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29228 = 10'h125 == _T_442[9:0] ? 4'h3 : _GEN_29227; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29229 = 10'h126 == _T_442[9:0] ? 4'h4 : _GEN_29228; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29230 = 10'h127 == _T_442[9:0] ? 4'h6 : _GEN_29229; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29231 = 10'h128 == _T_442[9:0] ? 4'h5 : _GEN_29230; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29232 = 10'h129 == _T_442[9:0] ? 4'h8 : _GEN_29231; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29233 = 10'h12a == _T_442[9:0] ? 4'h5 : _GEN_29232; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29234 = 10'h12b == _T_442[9:0] ? 4'h3 : _GEN_29233; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29235 = 10'h12c == _T_442[9:0] ? 4'h3 : _GEN_29234; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29236 = 10'h12d == _T_442[9:0] ? 4'h3 : _GEN_29235; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29237 = 10'h12e == _T_442[9:0] ? 4'h4 : _GEN_29236; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29238 = 10'h12f == _T_442[9:0] ? 4'h4 : _GEN_29237; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29239 = 10'h130 == _T_442[9:0] ? 4'ha : _GEN_29238; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29240 = 10'h131 == _T_442[9:0] ? 4'h9 : _GEN_29239; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29241 = 10'h132 == _T_442[9:0] ? 4'h9 : _GEN_29240; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29242 = 10'h133 == _T_442[9:0] ? 4'h8 : _GEN_29241; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29243 = 10'h134 == _T_442[9:0] ? 4'h9 : _GEN_29242; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29244 = 10'h135 == _T_442[9:0] ? 4'h8 : _GEN_29243; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29245 = 10'h136 == _T_442[9:0] ? 4'h7 : _GEN_29244; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29246 = 10'h137 == _T_442[9:0] ? 4'h6 : _GEN_29245; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29247 = 10'h138 == _T_442[9:0] ? 4'h8 : _GEN_29246; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29248 = 10'h139 == _T_442[9:0] ? 4'h3 : _GEN_29247; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29249 = 10'h13a == _T_442[9:0] ? 4'h3 : _GEN_29248; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29250 = 10'h13b == _T_442[9:0] ? 4'h4 : _GEN_29249; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29251 = 10'h13c == _T_442[9:0] ? 4'h4 : _GEN_29250; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29252 = 10'h13d == _T_442[9:0] ? 4'h3 : _GEN_29251; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29253 = 10'h13e == _T_442[9:0] ? 4'h5 : _GEN_29252; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29254 = 10'h13f == _T_442[9:0] ? 4'h9 : _GEN_29253; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29255 = 10'h140 == _T_442[9:0] ? 4'ha : _GEN_29254; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29256 = 10'h141 == _T_442[9:0] ? 4'ha : _GEN_29255; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29257 = 10'h142 == _T_442[9:0] ? 4'ha : _GEN_29256; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29258 = 10'h143 == _T_442[9:0] ? 4'h5 : _GEN_29257; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29259 = 10'h144 == _T_442[9:0] ? 4'h3 : _GEN_29258; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29260 = 10'h145 == _T_442[9:0] ? 4'h3 : _GEN_29259; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29261 = 10'h146 == _T_442[9:0] ? 4'h3 : _GEN_29260; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29262 = 10'h147 == _T_442[9:0] ? 4'h4 : _GEN_29261; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29263 = 10'h148 == _T_442[9:0] ? 4'h3 : _GEN_29262; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29264 = 10'h149 == _T_442[9:0] ? 4'h3 : _GEN_29263; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29265 = 10'h14a == _T_442[9:0] ? 4'h3 : _GEN_29264; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29266 = 10'h14b == _T_442[9:0] ? 4'h6 : _GEN_29265; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29267 = 10'h14c == _T_442[9:0] ? 4'h8 : _GEN_29266; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29268 = 10'h14d == _T_442[9:0] ? 4'h5 : _GEN_29267; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29269 = 10'h14e == _T_442[9:0] ? 4'h4 : _GEN_29268; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29270 = 10'h14f == _T_442[9:0] ? 4'h3 : _GEN_29269; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29271 = 10'h150 == _T_442[9:0] ? 4'h3 : _GEN_29270; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29272 = 10'h151 == _T_442[9:0] ? 4'h3 : _GEN_29271; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29273 = 10'h152 == _T_442[9:0] ? 4'h3 : _GEN_29272; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29274 = 10'h153 == _T_442[9:0] ? 4'h3 : _GEN_29273; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29275 = 10'h154 == _T_442[9:0] ? 4'h3 : _GEN_29274; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29276 = 10'h155 == _T_442[9:0] ? 4'h4 : _GEN_29275; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29277 = 10'h156 == _T_442[9:0] ? 4'h9 : _GEN_29276; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29278 = 10'h157 == _T_442[9:0] ? 4'h8 : _GEN_29277; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29279 = 10'h158 == _T_442[9:0] ? 4'h8 : _GEN_29278; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29280 = 10'h159 == _T_442[9:0] ? 4'h8 : _GEN_29279; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29281 = 10'h15a == _T_442[9:0] ? 4'h8 : _GEN_29280; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29282 = 10'h15b == _T_442[9:0] ? 4'h8 : _GEN_29281; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29283 = 10'h15c == _T_442[9:0] ? 4'h7 : _GEN_29282; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29284 = 10'h15d == _T_442[9:0] ? 4'h7 : _GEN_29283; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29285 = 10'h15e == _T_442[9:0] ? 4'h8 : _GEN_29284; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29286 = 10'h15f == _T_442[9:0] ? 4'h3 : _GEN_29285; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29287 = 10'h160 == _T_442[9:0] ? 4'h4 : _GEN_29286; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29288 = 10'h161 == _T_442[9:0] ? 4'h4 : _GEN_29287; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29289 = 10'h162 == _T_442[9:0] ? 4'h4 : _GEN_29288; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29290 = 10'h163 == _T_442[9:0] ? 4'h4 : _GEN_29289; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29291 = 10'h164 == _T_442[9:0] ? 4'h5 : _GEN_29290; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29292 = 10'h165 == _T_442[9:0] ? 4'ha : _GEN_29291; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29293 = 10'h166 == _T_442[9:0] ? 4'h9 : _GEN_29292; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29294 = 10'h167 == _T_442[9:0] ? 4'ha : _GEN_29293; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29295 = 10'h168 == _T_442[9:0] ? 4'ha : _GEN_29294; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29296 = 10'h169 == _T_442[9:0] ? 4'h6 : _GEN_29295; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29297 = 10'h16a == _T_442[9:0] ? 4'h3 : _GEN_29296; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29298 = 10'h16b == _T_442[9:0] ? 4'h3 : _GEN_29297; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29299 = 10'h16c == _T_442[9:0] ? 4'h3 : _GEN_29298; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29300 = 10'h16d == _T_442[9:0] ? 4'h4 : _GEN_29299; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29301 = 10'h16e == _T_442[9:0] ? 4'h3 : _GEN_29300; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29302 = 10'h16f == _T_442[9:0] ? 4'h3 : _GEN_29301; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29303 = 10'h170 == _T_442[9:0] ? 4'h3 : _GEN_29302; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29304 = 10'h171 == _T_442[9:0] ? 4'h7 : _GEN_29303; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29305 = 10'h172 == _T_442[9:0] ? 4'ha : _GEN_29304; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29306 = 10'h173 == _T_442[9:0] ? 4'h5 : _GEN_29305; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29307 = 10'h174 == _T_442[9:0] ? 4'h3 : _GEN_29306; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29308 = 10'h175 == _T_442[9:0] ? 4'h4 : _GEN_29307; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29309 = 10'h176 == _T_442[9:0] ? 4'h4 : _GEN_29308; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29310 = 10'h177 == _T_442[9:0] ? 4'h4 : _GEN_29309; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29311 = 10'h178 == _T_442[9:0] ? 4'h4 : _GEN_29310; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29312 = 10'h179 == _T_442[9:0] ? 4'h3 : _GEN_29311; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29313 = 10'h17a == _T_442[9:0] ? 4'h3 : _GEN_29312; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29314 = 10'h17b == _T_442[9:0] ? 4'h3 : _GEN_29313; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29315 = 10'h17c == _T_442[9:0] ? 4'h8 : _GEN_29314; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29316 = 10'h17d == _T_442[9:0] ? 4'h8 : _GEN_29315; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29317 = 10'h17e == _T_442[9:0] ? 4'h8 : _GEN_29316; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29318 = 10'h17f == _T_442[9:0] ? 4'h8 : _GEN_29317; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29319 = 10'h180 == _T_442[9:0] ? 4'h8 : _GEN_29318; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29320 = 10'h181 == _T_442[9:0] ? 4'h8 : _GEN_29319; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29321 = 10'h182 == _T_442[9:0] ? 4'h8 : _GEN_29320; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29322 = 10'h183 == _T_442[9:0] ? 4'h8 : _GEN_29321; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29323 = 10'h184 == _T_442[9:0] ? 4'h8 : _GEN_29322; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29324 = 10'h185 == _T_442[9:0] ? 4'h5 : _GEN_29323; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29325 = 10'h186 == _T_442[9:0] ? 4'h3 : _GEN_29324; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29326 = 10'h187 == _T_442[9:0] ? 4'h4 : _GEN_29325; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29327 = 10'h188 == _T_442[9:0] ? 4'h4 : _GEN_29326; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29328 = 10'h189 == _T_442[9:0] ? 4'h4 : _GEN_29327; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29329 = 10'h18a == _T_442[9:0] ? 4'h5 : _GEN_29328; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29330 = 10'h18b == _T_442[9:0] ? 4'ha : _GEN_29329; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29331 = 10'h18c == _T_442[9:0] ? 4'ha : _GEN_29330; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29332 = 10'h18d == _T_442[9:0] ? 4'h9 : _GEN_29331; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29333 = 10'h18e == _T_442[9:0] ? 4'ha : _GEN_29332; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29334 = 10'h18f == _T_442[9:0] ? 4'h4 : _GEN_29333; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29335 = 10'h190 == _T_442[9:0] ? 4'h3 : _GEN_29334; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29336 = 10'h191 == _T_442[9:0] ? 4'h3 : _GEN_29335; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29337 = 10'h192 == _T_442[9:0] ? 4'h5 : _GEN_29336; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29338 = 10'h193 == _T_442[9:0] ? 4'h6 : _GEN_29337; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29339 = 10'h194 == _T_442[9:0] ? 4'h5 : _GEN_29338; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29340 = 10'h195 == _T_442[9:0] ? 4'h3 : _GEN_29339; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29341 = 10'h196 == _T_442[9:0] ? 4'h3 : _GEN_29340; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29342 = 10'h197 == _T_442[9:0] ? 4'h5 : _GEN_29341; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29343 = 10'h198 == _T_442[9:0] ? 4'ha : _GEN_29342; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29344 = 10'h199 == _T_442[9:0] ? 4'h3 : _GEN_29343; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29345 = 10'h19a == _T_442[9:0] ? 4'h1 : _GEN_29344; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29346 = 10'h19b == _T_442[9:0] ? 4'h2 : _GEN_29345; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29347 = 10'h19c == _T_442[9:0] ? 4'h4 : _GEN_29346; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29348 = 10'h19d == _T_442[9:0] ? 4'h3 : _GEN_29347; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29349 = 10'h19e == _T_442[9:0] ? 4'h1 : _GEN_29348; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29350 = 10'h19f == _T_442[9:0] ? 4'h2 : _GEN_29349; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29351 = 10'h1a0 == _T_442[9:0] ? 4'h3 : _GEN_29350; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29352 = 10'h1a1 == _T_442[9:0] ? 4'h4 : _GEN_29351; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29353 = 10'h1a2 == _T_442[9:0] ? 4'h8 : _GEN_29352; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29354 = 10'h1a3 == _T_442[9:0] ? 4'h8 : _GEN_29353; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29355 = 10'h1a4 == _T_442[9:0] ? 4'h8 : _GEN_29354; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29356 = 10'h1a5 == _T_442[9:0] ? 4'h8 : _GEN_29355; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29357 = 10'h1a6 == _T_442[9:0] ? 4'h7 : _GEN_29356; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29358 = 10'h1a7 == _T_442[9:0] ? 4'h8 : _GEN_29357; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29359 = 10'h1a8 == _T_442[9:0] ? 4'h8 : _GEN_29358; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29360 = 10'h1a9 == _T_442[9:0] ? 4'h8 : _GEN_29359; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29361 = 10'h1aa == _T_442[9:0] ? 4'h7 : _GEN_29360; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29362 = 10'h1ab == _T_442[9:0] ? 4'h4 : _GEN_29361; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29363 = 10'h1ac == _T_442[9:0] ? 4'h4 : _GEN_29362; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29364 = 10'h1ad == _T_442[9:0] ? 4'h3 : _GEN_29363; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29365 = 10'h1ae == _T_442[9:0] ? 4'h3 : _GEN_29364; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29366 = 10'h1af == _T_442[9:0] ? 4'h4 : _GEN_29365; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29367 = 10'h1b0 == _T_442[9:0] ? 4'h6 : _GEN_29366; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29368 = 10'h1b1 == _T_442[9:0] ? 4'ha : _GEN_29367; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29369 = 10'h1b2 == _T_442[9:0] ? 4'ha : _GEN_29368; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29370 = 10'h1b3 == _T_442[9:0] ? 4'h9 : _GEN_29369; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29371 = 10'h1b4 == _T_442[9:0] ? 4'h9 : _GEN_29370; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29372 = 10'h1b5 == _T_442[9:0] ? 4'h3 : _GEN_29371; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29373 = 10'h1b6 == _T_442[9:0] ? 4'h3 : _GEN_29372; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29374 = 10'h1b7 == _T_442[9:0] ? 4'h4 : _GEN_29373; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29375 = 10'h1b8 == _T_442[9:0] ? 4'h5 : _GEN_29374; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29376 = 10'h1b9 == _T_442[9:0] ? 4'h6 : _GEN_29375; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29377 = 10'h1ba == _T_442[9:0] ? 4'h4 : _GEN_29376; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29378 = 10'h1bb == _T_442[9:0] ? 4'h3 : _GEN_29377; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29379 = 10'h1bc == _T_442[9:0] ? 4'h3 : _GEN_29378; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29380 = 10'h1bd == _T_442[9:0] ? 4'h4 : _GEN_29379; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29381 = 10'h1be == _T_442[9:0] ? 4'ha : _GEN_29380; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29382 = 10'h1bf == _T_442[9:0] ? 4'h4 : _GEN_29381; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29383 = 10'h1c0 == _T_442[9:0] ? 4'h5 : _GEN_29382; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29384 = 10'h1c1 == _T_442[9:0] ? 4'h5 : _GEN_29383; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29385 = 10'h1c2 == _T_442[9:0] ? 4'h4 : _GEN_29384; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29386 = 10'h1c3 == _T_442[9:0] ? 4'h5 : _GEN_29385; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29387 = 10'h1c4 == _T_442[9:0] ? 4'h4 : _GEN_29386; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29388 = 10'h1c5 == _T_442[9:0] ? 4'h3 : _GEN_29387; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29389 = 10'h1c6 == _T_442[9:0] ? 4'h4 : _GEN_29388; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29390 = 10'h1c7 == _T_442[9:0] ? 4'h3 : _GEN_29389; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29391 = 10'h1c8 == _T_442[9:0] ? 4'h8 : _GEN_29390; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29392 = 10'h1c9 == _T_442[9:0] ? 4'h8 : _GEN_29391; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29393 = 10'h1ca == _T_442[9:0] ? 4'h8 : _GEN_29392; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29394 = 10'h1cb == _T_442[9:0] ? 4'h8 : _GEN_29393; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29395 = 10'h1cc == _T_442[9:0] ? 4'h8 : _GEN_29394; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29396 = 10'h1cd == _T_442[9:0] ? 4'h8 : _GEN_29395; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29397 = 10'h1ce == _T_442[9:0] ? 4'h8 : _GEN_29396; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29398 = 10'h1cf == _T_442[9:0] ? 4'h8 : _GEN_29397; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29399 = 10'h1d0 == _T_442[9:0] ? 4'h5 : _GEN_29398; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29400 = 10'h1d1 == _T_442[9:0] ? 4'h4 : _GEN_29399; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29401 = 10'h1d2 == _T_442[9:0] ? 4'h6 : _GEN_29400; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29402 = 10'h1d3 == _T_442[9:0] ? 4'h6 : _GEN_29401; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29403 = 10'h1d4 == _T_442[9:0] ? 4'h6 : _GEN_29402; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29404 = 10'h1d5 == _T_442[9:0] ? 4'h5 : _GEN_29403; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29405 = 10'h1d6 == _T_442[9:0] ? 4'h8 : _GEN_29404; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29406 = 10'h1d7 == _T_442[9:0] ? 4'ha : _GEN_29405; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29407 = 10'h1d8 == _T_442[9:0] ? 4'ha : _GEN_29406; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29408 = 10'h1d9 == _T_442[9:0] ? 4'ha : _GEN_29407; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29409 = 10'h1da == _T_442[9:0] ? 4'h6 : _GEN_29408; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29410 = 10'h1db == _T_442[9:0] ? 4'h3 : _GEN_29409; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29411 = 10'h1dc == _T_442[9:0] ? 4'h5 : _GEN_29410; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29412 = 10'h1dd == _T_442[9:0] ? 4'h2 : _GEN_29411; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29413 = 10'h1de == _T_442[9:0] ? 4'h5 : _GEN_29412; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29414 = 10'h1df == _T_442[9:0] ? 4'h5 : _GEN_29413; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29415 = 10'h1e0 == _T_442[9:0] ? 4'h5 : _GEN_29414; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29416 = 10'h1e1 == _T_442[9:0] ? 4'h3 : _GEN_29415; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29417 = 10'h1e2 == _T_442[9:0] ? 4'h3 : _GEN_29416; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29418 = 10'h1e3 == _T_442[9:0] ? 4'h3 : _GEN_29417; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29419 = 10'h1e4 == _T_442[9:0] ? 4'h9 : _GEN_29418; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29420 = 10'h1e5 == _T_442[9:0] ? 4'h4 : _GEN_29419; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29421 = 10'h1e6 == _T_442[9:0] ? 4'h4 : _GEN_29420; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29422 = 10'h1e7 == _T_442[9:0] ? 4'h4 : _GEN_29421; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29423 = 10'h1e8 == _T_442[9:0] ? 4'h4 : _GEN_29422; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29424 = 10'h1e9 == _T_442[9:0] ? 4'h4 : _GEN_29423; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29425 = 10'h1ea == _T_442[9:0] ? 4'h4 : _GEN_29424; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29426 = 10'h1eb == _T_442[9:0] ? 4'h4 : _GEN_29425; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29427 = 10'h1ec == _T_442[9:0] ? 4'h4 : _GEN_29426; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29428 = 10'h1ed == _T_442[9:0] ? 4'h4 : _GEN_29427; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29429 = 10'h1ee == _T_442[9:0] ? 4'h8 : _GEN_29428; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29430 = 10'h1ef == _T_442[9:0] ? 4'h8 : _GEN_29429; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29431 = 10'h1f0 == _T_442[9:0] ? 4'h8 : _GEN_29430; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29432 = 10'h1f1 == _T_442[9:0] ? 4'h8 : _GEN_29431; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29433 = 10'h1f2 == _T_442[9:0] ? 4'h8 : _GEN_29432; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29434 = 10'h1f3 == _T_442[9:0] ? 4'h8 : _GEN_29433; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29435 = 10'h1f4 == _T_442[9:0] ? 4'h9 : _GEN_29434; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29436 = 10'h1f5 == _T_442[9:0] ? 4'h9 : _GEN_29435; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29437 = 10'h1f6 == _T_442[9:0] ? 4'ha : _GEN_29436; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29438 = 10'h1f7 == _T_442[9:0] ? 4'h5 : _GEN_29437; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29439 = 10'h1f8 == _T_442[9:0] ? 4'h5 : _GEN_29438; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29440 = 10'h1f9 == _T_442[9:0] ? 4'h7 : _GEN_29439; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29441 = 10'h1fa == _T_442[9:0] ? 4'h7 : _GEN_29440; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29442 = 10'h1fb == _T_442[9:0] ? 4'h5 : _GEN_29441; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29443 = 10'h1fc == _T_442[9:0] ? 4'ha : _GEN_29442; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29444 = 10'h1fd == _T_442[9:0] ? 4'hb : _GEN_29443; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29445 = 10'h1fe == _T_442[9:0] ? 4'hb : _GEN_29444; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29446 = 10'h1ff == _T_442[9:0] ? 4'ha : _GEN_29445; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29447 = 10'h200 == _T_442[9:0] ? 4'h4 : _GEN_29446; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29448 = 10'h201 == _T_442[9:0] ? 4'h3 : _GEN_29447; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29449 = 10'h202 == _T_442[9:0] ? 4'h2 : _GEN_29448; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29450 = 10'h203 == _T_442[9:0] ? 4'h2 : _GEN_29449; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29451 = 10'h204 == _T_442[9:0] ? 4'h2 : _GEN_29450; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29452 = 10'h205 == _T_442[9:0] ? 4'h2 : _GEN_29451; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29453 = 10'h206 == _T_442[9:0] ? 4'h2 : _GEN_29452; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29454 = 10'h207 == _T_442[9:0] ? 4'h2 : _GEN_29453; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29455 = 10'h208 == _T_442[9:0] ? 4'h3 : _GEN_29454; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29456 = 10'h209 == _T_442[9:0] ? 4'h3 : _GEN_29455; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29457 = 10'h20a == _T_442[9:0] ? 4'h8 : _GEN_29456; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29458 = 10'h20b == _T_442[9:0] ? 4'h4 : _GEN_29457; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29459 = 10'h20c == _T_442[9:0] ? 4'h4 : _GEN_29458; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29460 = 10'h20d == _T_442[9:0] ? 4'h4 : _GEN_29459; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29461 = 10'h20e == _T_442[9:0] ? 4'h4 : _GEN_29460; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29462 = 10'h20f == _T_442[9:0] ? 4'h4 : _GEN_29461; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29463 = 10'h210 == _T_442[9:0] ? 4'h4 : _GEN_29462; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29464 = 10'h211 == _T_442[9:0] ? 4'h4 : _GEN_29463; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29465 = 10'h212 == _T_442[9:0] ? 4'h4 : _GEN_29464; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29466 = 10'h213 == _T_442[9:0] ? 4'h6 : _GEN_29465; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29467 = 10'h214 == _T_442[9:0] ? 4'h7 : _GEN_29466; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29468 = 10'h215 == _T_442[9:0] ? 4'h8 : _GEN_29467; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29469 = 10'h216 == _T_442[9:0] ? 4'h8 : _GEN_29468; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29470 = 10'h217 == _T_442[9:0] ? 4'h8 : _GEN_29469; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29471 = 10'h218 == _T_442[9:0] ? 4'h8 : _GEN_29470; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29472 = 10'h219 == _T_442[9:0] ? 4'h8 : _GEN_29471; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29473 = 10'h21a == _T_442[9:0] ? 4'h8 : _GEN_29472; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29474 = 10'h21b == _T_442[9:0] ? 4'h8 : _GEN_29473; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29475 = 10'h21c == _T_442[9:0] ? 4'ha : _GEN_29474; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29476 = 10'h21d == _T_442[9:0] ? 4'h9 : _GEN_29475; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29477 = 10'h21e == _T_442[9:0] ? 4'h6 : _GEN_29476; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29478 = 10'h21f == _T_442[9:0] ? 4'h4 : _GEN_29477; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29479 = 10'h220 == _T_442[9:0] ? 4'h4 : _GEN_29478; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29480 = 10'h221 == _T_442[9:0] ? 4'h5 : _GEN_29479; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29481 = 10'h222 == _T_442[9:0] ? 4'ha : _GEN_29480; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29482 = 10'h223 == _T_442[9:0] ? 4'ha : _GEN_29481; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29483 = 10'h224 == _T_442[9:0] ? 4'ha : _GEN_29482; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29484 = 10'h225 == _T_442[9:0] ? 4'h8 : _GEN_29483; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29485 = 10'h226 == _T_442[9:0] ? 4'h4 : _GEN_29484; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29486 = 10'h227 == _T_442[9:0] ? 4'h2 : _GEN_29485; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29487 = 10'h228 == _T_442[9:0] ? 4'h2 : _GEN_29486; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29488 = 10'h229 == _T_442[9:0] ? 4'h2 : _GEN_29487; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29489 = 10'h22a == _T_442[9:0] ? 4'h2 : _GEN_29488; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29490 = 10'h22b == _T_442[9:0] ? 4'h2 : _GEN_29489; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29491 = 10'h22c == _T_442[9:0] ? 4'h2 : _GEN_29490; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29492 = 10'h22d == _T_442[9:0] ? 4'h2 : _GEN_29491; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29493 = 10'h22e == _T_442[9:0] ? 4'h2 : _GEN_29492; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29494 = 10'h22f == _T_442[9:0] ? 4'h3 : _GEN_29493; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29495 = 10'h230 == _T_442[9:0] ? 4'h3 : _GEN_29494; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29496 = 10'h231 == _T_442[9:0] ? 4'h3 : _GEN_29495; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29497 = 10'h232 == _T_442[9:0] ? 4'h4 : _GEN_29496; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29498 = 10'h233 == _T_442[9:0] ? 4'h6 : _GEN_29497; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29499 = 10'h234 == _T_442[9:0] ? 4'h6 : _GEN_29498; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29500 = 10'h235 == _T_442[9:0] ? 4'h4 : _GEN_29499; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29501 = 10'h236 == _T_442[9:0] ? 4'h4 : _GEN_29500; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29502 = 10'h237 == _T_442[9:0] ? 4'h4 : _GEN_29501; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29503 = 10'h238 == _T_442[9:0] ? 4'h4 : _GEN_29502; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29504 = 10'h239 == _T_442[9:0] ? 4'h3 : _GEN_29503; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29505 = 10'h23a == _T_442[9:0] ? 4'h7 : _GEN_29504; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29506 = 10'h23b == _T_442[9:0] ? 4'h7 : _GEN_29505; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29507 = 10'h23c == _T_442[9:0] ? 4'h7 : _GEN_29506; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29508 = 10'h23d == _T_442[9:0] ? 4'h7 : _GEN_29507; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29509 = 10'h23e == _T_442[9:0] ? 4'h7 : _GEN_29508; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29510 = 10'h23f == _T_442[9:0] ? 4'h7 : _GEN_29509; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29511 = 10'h240 == _T_442[9:0] ? 4'h7 : _GEN_29510; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29512 = 10'h241 == _T_442[9:0] ? 4'h8 : _GEN_29511; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29513 = 10'h242 == _T_442[9:0] ? 4'ha : _GEN_29512; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29514 = 10'h243 == _T_442[9:0] ? 4'ha : _GEN_29513; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29515 = 10'h244 == _T_442[9:0] ? 4'ha : _GEN_29514; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29516 = 10'h245 == _T_442[9:0] ? 4'h8 : _GEN_29515; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29517 = 10'h246 == _T_442[9:0] ? 4'h7 : _GEN_29516; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29518 = 10'h247 == _T_442[9:0] ? 4'h8 : _GEN_29517; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29519 = 10'h248 == _T_442[9:0] ? 4'ha : _GEN_29518; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29520 = 10'h249 == _T_442[9:0] ? 4'ha : _GEN_29519; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29521 = 10'h24a == _T_442[9:0] ? 4'ha : _GEN_29520; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29522 = 10'h24b == _T_442[9:0] ? 4'h4 : _GEN_29521; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29523 = 10'h24c == _T_442[9:0] ? 4'h4 : _GEN_29522; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29524 = 10'h24d == _T_442[9:0] ? 4'h2 : _GEN_29523; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29525 = 10'h24e == _T_442[9:0] ? 4'h2 : _GEN_29524; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29526 = 10'h24f == _T_442[9:0] ? 4'h2 : _GEN_29525; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29527 = 10'h250 == _T_442[9:0] ? 4'h2 : _GEN_29526; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29528 = 10'h251 == _T_442[9:0] ? 4'h2 : _GEN_29527; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29529 = 10'h252 == _T_442[9:0] ? 4'h2 : _GEN_29528; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29530 = 10'h253 == _T_442[9:0] ? 4'h2 : _GEN_29529; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29531 = 10'h254 == _T_442[9:0] ? 4'h2 : _GEN_29530; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29532 = 10'h255 == _T_442[9:0] ? 4'h3 : _GEN_29531; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29533 = 10'h256 == _T_442[9:0] ? 4'h4 : _GEN_29532; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29534 = 10'h257 == _T_442[9:0] ? 4'h3 : _GEN_29533; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29535 = 10'h258 == _T_442[9:0] ? 4'h4 : _GEN_29534; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29536 = 10'h259 == _T_442[9:0] ? 4'h4 : _GEN_29535; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29537 = 10'h25a == _T_442[9:0] ? 4'h4 : _GEN_29536; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29538 = 10'h25b == _T_442[9:0] ? 4'h3 : _GEN_29537; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29539 = 10'h25c == _T_442[9:0] ? 4'h4 : _GEN_29538; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29540 = 10'h25d == _T_442[9:0] ? 4'h4 : _GEN_29539; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29541 = 10'h25e == _T_442[9:0] ? 4'h3 : _GEN_29540; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29542 = 10'h25f == _T_442[9:0] ? 4'h3 : _GEN_29541; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29543 = 10'h260 == _T_442[9:0] ? 4'h8 : _GEN_29542; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29544 = 10'h261 == _T_442[9:0] ? 4'h7 : _GEN_29543; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29545 = 10'h262 == _T_442[9:0] ? 4'h6 : _GEN_29544; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29546 = 10'h263 == _T_442[9:0] ? 4'h5 : _GEN_29545; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29547 = 10'h264 == _T_442[9:0] ? 4'h6 : _GEN_29546; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29548 = 10'h265 == _T_442[9:0] ? 4'h5 : _GEN_29547; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29549 = 10'h266 == _T_442[9:0] ? 4'h5 : _GEN_29548; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29550 = 10'h267 == _T_442[9:0] ? 4'h7 : _GEN_29549; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29551 = 10'h268 == _T_442[9:0] ? 4'ha : _GEN_29550; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29552 = 10'h269 == _T_442[9:0] ? 4'ha : _GEN_29551; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29553 = 10'h26a == _T_442[9:0] ? 4'ha : _GEN_29552; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29554 = 10'h26b == _T_442[9:0] ? 4'ha : _GEN_29553; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29555 = 10'h26c == _T_442[9:0] ? 4'ha : _GEN_29554; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29556 = 10'h26d == _T_442[9:0] ? 4'ha : _GEN_29555; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29557 = 10'h26e == _T_442[9:0] ? 4'ha : _GEN_29556; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29558 = 10'h26f == _T_442[9:0] ? 4'ha : _GEN_29557; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29559 = 10'h270 == _T_442[9:0] ? 4'h5 : _GEN_29558; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29560 = 10'h271 == _T_442[9:0] ? 4'h4 : _GEN_29559; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29561 = 10'h272 == _T_442[9:0] ? 4'h3 : _GEN_29560; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29562 = 10'h273 == _T_442[9:0] ? 4'h2 : _GEN_29561; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29563 = 10'h274 == _T_442[9:0] ? 4'h2 : _GEN_29562; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29564 = 10'h275 == _T_442[9:0] ? 4'h2 : _GEN_29563; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29565 = 10'h276 == _T_442[9:0] ? 4'h2 : _GEN_29564; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29566 = 10'h277 == _T_442[9:0] ? 4'h2 : _GEN_29565; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29567 = 10'h278 == _T_442[9:0] ? 4'h2 : _GEN_29566; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29568 = 10'h279 == _T_442[9:0] ? 4'h2 : _GEN_29567; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29569 = 10'h27a == _T_442[9:0] ? 4'h2 : _GEN_29568; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29570 = 10'h27b == _T_442[9:0] ? 4'h4 : _GEN_29569; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29571 = 10'h27c == _T_442[9:0] ? 4'h3 : _GEN_29570; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29572 = 10'h27d == _T_442[9:0] ? 4'h4 : _GEN_29571; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29573 = 10'h27e == _T_442[9:0] ? 4'h5 : _GEN_29572; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29574 = 10'h27f == _T_442[9:0] ? 4'h4 : _GEN_29573; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29575 = 10'h280 == _T_442[9:0] ? 4'h4 : _GEN_29574; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29576 = 10'h281 == _T_442[9:0] ? 4'h4 : _GEN_29575; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29577 = 10'h282 == _T_442[9:0] ? 4'h4 : _GEN_29576; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29578 = 10'h283 == _T_442[9:0] ? 4'h3 : _GEN_29577; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29579 = 10'h284 == _T_442[9:0] ? 4'h3 : _GEN_29578; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29580 = 10'h285 == _T_442[9:0] ? 4'h3 : _GEN_29579; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29581 = 10'h286 == _T_442[9:0] ? 4'h8 : _GEN_29580; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29582 = 10'h287 == _T_442[9:0] ? 4'h6 : _GEN_29581; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29583 = 10'h288 == _T_442[9:0] ? 4'h6 : _GEN_29582; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29584 = 10'h289 == _T_442[9:0] ? 4'h6 : _GEN_29583; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29585 = 10'h28a == _T_442[9:0] ? 4'h7 : _GEN_29584; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29586 = 10'h28b == _T_442[9:0] ? 4'h7 : _GEN_29585; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29587 = 10'h28c == _T_442[9:0] ? 4'h6 : _GEN_29586; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29588 = 10'h28d == _T_442[9:0] ? 4'h6 : _GEN_29587; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29589 = 10'h28e == _T_442[9:0] ? 4'h4 : _GEN_29588; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29590 = 10'h28f == _T_442[9:0] ? 4'h7 : _GEN_29589; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29591 = 10'h290 == _T_442[9:0] ? 4'h9 : _GEN_29590; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29592 = 10'h291 == _T_442[9:0] ? 4'ha : _GEN_29591; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29593 = 10'h292 == _T_442[9:0] ? 4'ha : _GEN_29592; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29594 = 10'h293 == _T_442[9:0] ? 4'ha : _GEN_29593; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29595 = 10'h294 == _T_442[9:0] ? 4'h9 : _GEN_29594; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29596 = 10'h295 == _T_442[9:0] ? 4'h5 : _GEN_29595; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29597 = 10'h296 == _T_442[9:0] ? 4'h4 : _GEN_29596; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29598 = 10'h297 == _T_442[9:0] ? 4'h4 : _GEN_29597; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29599 = 10'h298 == _T_442[9:0] ? 4'h3 : _GEN_29598; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29600 = 10'h299 == _T_442[9:0] ? 4'h3 : _GEN_29599; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29601 = 10'h29a == _T_442[9:0] ? 4'h2 : _GEN_29600; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29602 = 10'h29b == _T_442[9:0] ? 4'h2 : _GEN_29601; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29603 = 10'h29c == _T_442[9:0] ? 4'h2 : _GEN_29602; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29604 = 10'h29d == _T_442[9:0] ? 4'h2 : _GEN_29603; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29605 = 10'h29e == _T_442[9:0] ? 4'h2 : _GEN_29604; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29606 = 10'h29f == _T_442[9:0] ? 4'h2 : _GEN_29605; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29607 = 10'h2a0 == _T_442[9:0] ? 4'h2 : _GEN_29606; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29608 = 10'h2a1 == _T_442[9:0] ? 4'h4 : _GEN_29607; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29609 = 10'h2a2 == _T_442[9:0] ? 4'h3 : _GEN_29608; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29610 = 10'h2a3 == _T_442[9:0] ? 4'h4 : _GEN_29609; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29611 = 10'h2a4 == _T_442[9:0] ? 4'h5 : _GEN_29610; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29612 = 10'h2a5 == _T_442[9:0] ? 4'h4 : _GEN_29611; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29613 = 10'h2a6 == _T_442[9:0] ? 4'h4 : _GEN_29612; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29614 = 10'h2a7 == _T_442[9:0] ? 4'h4 : _GEN_29613; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29615 = 10'h2a8 == _T_442[9:0] ? 4'h3 : _GEN_29614; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29616 = 10'h2a9 == _T_442[9:0] ? 4'h3 : _GEN_29615; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29617 = 10'h2aa == _T_442[9:0] ? 4'h3 : _GEN_29616; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29618 = 10'h2ab == _T_442[9:0] ? 4'h3 : _GEN_29617; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29619 = 10'h2ac == _T_442[9:0] ? 4'h8 : _GEN_29618; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29620 = 10'h2ad == _T_442[9:0] ? 4'h7 : _GEN_29619; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29621 = 10'h2ae == _T_442[9:0] ? 4'h5 : _GEN_29620; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29622 = 10'h2af == _T_442[9:0] ? 4'h6 : _GEN_29621; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29623 = 10'h2b0 == _T_442[9:0] ? 4'h7 : _GEN_29622; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29624 = 10'h2b1 == _T_442[9:0] ? 4'h6 : _GEN_29623; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29625 = 10'h2b2 == _T_442[9:0] ? 4'h6 : _GEN_29624; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29626 = 10'h2b3 == _T_442[9:0] ? 4'h6 : _GEN_29625; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29627 = 10'h2b4 == _T_442[9:0] ? 4'h3 : _GEN_29626; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29628 = 10'h2b5 == _T_442[9:0] ? 4'h3 : _GEN_29627; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29629 = 10'h2b6 == _T_442[9:0] ? 4'h3 : _GEN_29628; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29630 = 10'h2b7 == _T_442[9:0] ? 4'h4 : _GEN_29629; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29631 = 10'h2b8 == _T_442[9:0] ? 4'h6 : _GEN_29630; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29632 = 10'h2b9 == _T_442[9:0] ? 4'h9 : _GEN_29631; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29633 = 10'h2ba == _T_442[9:0] ? 4'h4 : _GEN_29632; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29634 = 10'h2bb == _T_442[9:0] ? 4'h3 : _GEN_29633; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29635 = 10'h2bc == _T_442[9:0] ? 4'h4 : _GEN_29634; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29636 = 10'h2bd == _T_442[9:0] ? 4'h3 : _GEN_29635; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29637 = 10'h2be == _T_442[9:0] ? 4'h3 : _GEN_29636; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29638 = 10'h2bf == _T_442[9:0] ? 4'h3 : _GEN_29637; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29639 = 10'h2c0 == _T_442[9:0] ? 4'h2 : _GEN_29638; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29640 = 10'h2c1 == _T_442[9:0] ? 4'h2 : _GEN_29639; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29641 = 10'h2c2 == _T_442[9:0] ? 4'h2 : _GEN_29640; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29642 = 10'h2c3 == _T_442[9:0] ? 4'h2 : _GEN_29641; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29643 = 10'h2c4 == _T_442[9:0] ? 4'h2 : _GEN_29642; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29644 = 10'h2c5 == _T_442[9:0] ? 4'h2 : _GEN_29643; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29645 = 10'h2c6 == _T_442[9:0] ? 4'h2 : _GEN_29644; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29646 = 10'h2c7 == _T_442[9:0] ? 4'h4 : _GEN_29645; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29647 = 10'h2c8 == _T_442[9:0] ? 4'h3 : _GEN_29646; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29648 = 10'h2c9 == _T_442[9:0] ? 4'h4 : _GEN_29647; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29649 = 10'h2ca == _T_442[9:0] ? 4'h5 : _GEN_29648; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29650 = 10'h2cb == _T_442[9:0] ? 4'h3 : _GEN_29649; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29651 = 10'h2cc == _T_442[9:0] ? 4'h3 : _GEN_29650; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29652 = 10'h2cd == _T_442[9:0] ? 4'h3 : _GEN_29651; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29653 = 10'h2ce == _T_442[9:0] ? 4'h3 : _GEN_29652; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29654 = 10'h2cf == _T_442[9:0] ? 4'h3 : _GEN_29653; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29655 = 10'h2d0 == _T_442[9:0] ? 4'h3 : _GEN_29654; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29656 = 10'h2d1 == _T_442[9:0] ? 4'h3 : _GEN_29655; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29657 = 10'h2d2 == _T_442[9:0] ? 4'h8 : _GEN_29656; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29658 = 10'h2d3 == _T_442[9:0] ? 4'h6 : _GEN_29657; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29659 = 10'h2d4 == _T_442[9:0] ? 4'h6 : _GEN_29658; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29660 = 10'h2d5 == _T_442[9:0] ? 4'h7 : _GEN_29659; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29661 = 10'h2d6 == _T_442[9:0] ? 4'h7 : _GEN_29660; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29662 = 10'h2d7 == _T_442[9:0] ? 4'h7 : _GEN_29661; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29663 = 10'h2d8 == _T_442[9:0] ? 4'h6 : _GEN_29662; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29664 = 10'h2d9 == _T_442[9:0] ? 4'h7 : _GEN_29663; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29665 = 10'h2da == _T_442[9:0] ? 4'h5 : _GEN_29664; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29666 = 10'h2db == _T_442[9:0] ? 4'h3 : _GEN_29665; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29667 = 10'h2dc == _T_442[9:0] ? 4'h3 : _GEN_29666; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29668 = 10'h2dd == _T_442[9:0] ? 4'h3 : _GEN_29667; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29669 = 10'h2de == _T_442[9:0] ? 4'h3 : _GEN_29668; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29670 = 10'h2df == _T_442[9:0] ? 4'h4 : _GEN_29669; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29671 = 10'h2e0 == _T_442[9:0] ? 4'h3 : _GEN_29670; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29672 = 10'h2e1 == _T_442[9:0] ? 4'h3 : _GEN_29671; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29673 = 10'h2e2 == _T_442[9:0] ? 4'h3 : _GEN_29672; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29674 = 10'h2e3 == _T_442[9:0] ? 4'h3 : _GEN_29673; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29675 = 10'h2e4 == _T_442[9:0] ? 4'h3 : _GEN_29674; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29676 = 10'h2e5 == _T_442[9:0] ? 4'h3 : _GEN_29675; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29677 = 10'h2e6 == _T_442[9:0] ? 4'h2 : _GEN_29676; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29678 = 10'h2e7 == _T_442[9:0] ? 4'h2 : _GEN_29677; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29679 = 10'h2e8 == _T_442[9:0] ? 4'h2 : _GEN_29678; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29680 = 10'h2e9 == _T_442[9:0] ? 4'h2 : _GEN_29679; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29681 = 10'h2ea == _T_442[9:0] ? 4'h2 : _GEN_29680; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29682 = 10'h2eb == _T_442[9:0] ? 4'h2 : _GEN_29681; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29683 = 10'h2ec == _T_442[9:0] ? 4'h3 : _GEN_29682; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29684 = 10'h2ed == _T_442[9:0] ? 4'h4 : _GEN_29683; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29685 = 10'h2ee == _T_442[9:0] ? 4'h3 : _GEN_29684; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29686 = 10'h2ef == _T_442[9:0] ? 4'h3 : _GEN_29685; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29687 = 10'h2f0 == _T_442[9:0] ? 4'h6 : _GEN_29686; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29688 = 10'h2f1 == _T_442[9:0] ? 4'h3 : _GEN_29687; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29689 = 10'h2f2 == _T_442[9:0] ? 4'h3 : _GEN_29688; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29690 = 10'h2f3 == _T_442[9:0] ? 4'h3 : _GEN_29689; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29691 = 10'h2f4 == _T_442[9:0] ? 4'h3 : _GEN_29690; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29692 = 10'h2f5 == _T_442[9:0] ? 4'h3 : _GEN_29691; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29693 = 10'h2f6 == _T_442[9:0] ? 4'h3 : _GEN_29692; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29694 = 10'h2f7 == _T_442[9:0] ? 4'h3 : _GEN_29693; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29695 = 10'h2f8 == _T_442[9:0] ? 4'h8 : _GEN_29694; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29696 = 10'h2f9 == _T_442[9:0] ? 4'h6 : _GEN_29695; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29697 = 10'h2fa == _T_442[9:0] ? 4'h7 : _GEN_29696; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29698 = 10'h2fb == _T_442[9:0] ? 4'h7 : _GEN_29697; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29699 = 10'h2fc == _T_442[9:0] ? 4'h6 : _GEN_29698; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29700 = 10'h2fd == _T_442[9:0] ? 4'h6 : _GEN_29699; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29701 = 10'h2fe == _T_442[9:0] ? 4'h6 : _GEN_29700; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29702 = 10'h2ff == _T_442[9:0] ? 4'h8 : _GEN_29701; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29703 = 10'h300 == _T_442[9:0] ? 4'h9 : _GEN_29702; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29704 = 10'h301 == _T_442[9:0] ? 4'h7 : _GEN_29703; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29705 = 10'h302 == _T_442[9:0] ? 4'h4 : _GEN_29704; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29706 = 10'h303 == _T_442[9:0] ? 4'h4 : _GEN_29705; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29707 = 10'h304 == _T_442[9:0] ? 4'h3 : _GEN_29706; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29708 = 10'h305 == _T_442[9:0] ? 4'h3 : _GEN_29707; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29709 = 10'h306 == _T_442[9:0] ? 4'h3 : _GEN_29708; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29710 = 10'h307 == _T_442[9:0] ? 4'h3 : _GEN_29709; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29711 = 10'h308 == _T_442[9:0] ? 4'h3 : _GEN_29710; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29712 = 10'h309 == _T_442[9:0] ? 4'h3 : _GEN_29711; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29713 = 10'h30a == _T_442[9:0] ? 4'h3 : _GEN_29712; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29714 = 10'h30b == _T_442[9:0] ? 4'h3 : _GEN_29713; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29715 = 10'h30c == _T_442[9:0] ? 4'h2 : _GEN_29714; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29716 = 10'h30d == _T_442[9:0] ? 4'h2 : _GEN_29715; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29717 = 10'h30e == _T_442[9:0] ? 4'h2 : _GEN_29716; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29718 = 10'h30f == _T_442[9:0] ? 4'h2 : _GEN_29717; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29719 = 10'h310 == _T_442[9:0] ? 4'h2 : _GEN_29718; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29720 = 10'h311 == _T_442[9:0] ? 4'h2 : _GEN_29719; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29721 = 10'h312 == _T_442[9:0] ? 4'h3 : _GEN_29720; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29722 = 10'h313 == _T_442[9:0] ? 4'h4 : _GEN_29721; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29723 = 10'h314 == _T_442[9:0] ? 4'h3 : _GEN_29722; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29724 = 10'h315 == _T_442[9:0] ? 4'h3 : _GEN_29723; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29725 = 10'h316 == _T_442[9:0] ? 4'h5 : _GEN_29724; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29726 = 10'h317 == _T_442[9:0] ? 4'h5 : _GEN_29725; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29727 = 10'h318 == _T_442[9:0] ? 4'h3 : _GEN_29726; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29728 = 10'h319 == _T_442[9:0] ? 4'h3 : _GEN_29727; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29729 = 10'h31a == _T_442[9:0] ? 4'h3 : _GEN_29728; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29730 = 10'h31b == _T_442[9:0] ? 4'h3 : _GEN_29729; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29731 = 10'h31c == _T_442[9:0] ? 4'h3 : _GEN_29730; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29732 = 10'h31d == _T_442[9:0] ? 4'h3 : _GEN_29731; // @[Filter.scala 230:62]
  wire [4:0] _GEN_39026 = {{1'd0}, _GEN_29732}; // @[Filter.scala 230:62]
  wire [8:0] _T_444 = _GEN_39026 * 5'h14; // @[Filter.scala 230:62]
  wire [3:0] _GEN_29756 = 10'h17 == _T_442[9:0] ? 4'hb : 4'he; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29757 = 10'h18 == _T_442[9:0] ? 4'hc : _GEN_29756; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29758 = 10'h19 == _T_442[9:0] ? 4'he : _GEN_29757; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29759 = 10'h1a == _T_442[9:0] ? 4'he : _GEN_29758; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29760 = 10'h1b == _T_442[9:0] ? 4'he : _GEN_29759; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29761 = 10'h1c == _T_442[9:0] ? 4'he : _GEN_29760; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29762 = 10'h1d == _T_442[9:0] ? 4'he : _GEN_29761; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29763 = 10'h1e == _T_442[9:0] ? 4'he : _GEN_29762; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29764 = 10'h1f == _T_442[9:0] ? 4'he : _GEN_29763; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29765 = 10'h20 == _T_442[9:0] ? 4'he : _GEN_29764; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29766 = 10'h21 == _T_442[9:0] ? 4'he : _GEN_29765; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29767 = 10'h22 == _T_442[9:0] ? 4'he : _GEN_29766; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29768 = 10'h23 == _T_442[9:0] ? 4'he : _GEN_29767; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29769 = 10'h24 == _T_442[9:0] ? 4'he : _GEN_29768; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29770 = 10'h25 == _T_442[9:0] ? 4'he : _GEN_29769; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29771 = 10'h26 == _T_442[9:0] ? 4'he : _GEN_29770; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29772 = 10'h27 == _T_442[9:0] ? 4'he : _GEN_29771; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29773 = 10'h28 == _T_442[9:0] ? 4'he : _GEN_29772; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29774 = 10'h29 == _T_442[9:0] ? 4'he : _GEN_29773; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29775 = 10'h2a == _T_442[9:0] ? 4'he : _GEN_29774; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29776 = 10'h2b == _T_442[9:0] ? 4'he : _GEN_29775; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29777 = 10'h2c == _T_442[9:0] ? 4'he : _GEN_29776; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29778 = 10'h2d == _T_442[9:0] ? 4'he : _GEN_29777; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29779 = 10'h2e == _T_442[9:0] ? 4'he : _GEN_29778; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29780 = 10'h2f == _T_442[9:0] ? 4'he : _GEN_29779; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29781 = 10'h30 == _T_442[9:0] ? 4'he : _GEN_29780; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29782 = 10'h31 == _T_442[9:0] ? 4'he : _GEN_29781; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29783 = 10'h32 == _T_442[9:0] ? 4'he : _GEN_29782; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29784 = 10'h33 == _T_442[9:0] ? 4'he : _GEN_29783; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29785 = 10'h34 == _T_442[9:0] ? 4'he : _GEN_29784; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29786 = 10'h35 == _T_442[9:0] ? 4'he : _GEN_29785; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29787 = 10'h36 == _T_442[9:0] ? 4'he : _GEN_29786; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29788 = 10'h37 == _T_442[9:0] ? 4'he : _GEN_29787; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29789 = 10'h38 == _T_442[9:0] ? 4'he : _GEN_29788; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29790 = 10'h39 == _T_442[9:0] ? 4'he : _GEN_29789; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29791 = 10'h3a == _T_442[9:0] ? 4'he : _GEN_29790; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29792 = 10'h3b == _T_442[9:0] ? 4'he : _GEN_29791; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29793 = 10'h3c == _T_442[9:0] ? 4'ha : _GEN_29792; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29794 = 10'h3d == _T_442[9:0] ? 4'hc : _GEN_29793; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29795 = 10'h3e == _T_442[9:0] ? 4'hb : _GEN_29794; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29796 = 10'h3f == _T_442[9:0] ? 4'he : _GEN_29795; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29797 = 10'h40 == _T_442[9:0] ? 4'he : _GEN_29796; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29798 = 10'h41 == _T_442[9:0] ? 4'he : _GEN_29797; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29799 = 10'h42 == _T_442[9:0] ? 4'he : _GEN_29798; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29800 = 10'h43 == _T_442[9:0] ? 4'he : _GEN_29799; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29801 = 10'h44 == _T_442[9:0] ? 4'he : _GEN_29800; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29802 = 10'h45 == _T_442[9:0] ? 4'he : _GEN_29801; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29803 = 10'h46 == _T_442[9:0] ? 4'he : _GEN_29802; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29804 = 10'h47 == _T_442[9:0] ? 4'he : _GEN_29803; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29805 = 10'h48 == _T_442[9:0] ? 4'he : _GEN_29804; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29806 = 10'h49 == _T_442[9:0] ? 4'he : _GEN_29805; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29807 = 10'h4a == _T_442[9:0] ? 4'he : _GEN_29806; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29808 = 10'h4b == _T_442[9:0] ? 4'he : _GEN_29807; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29809 = 10'h4c == _T_442[9:0] ? 4'he : _GEN_29808; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29810 = 10'h4d == _T_442[9:0] ? 4'he : _GEN_29809; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29811 = 10'h4e == _T_442[9:0] ? 4'he : _GEN_29810; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29812 = 10'h4f == _T_442[9:0] ? 4'he : _GEN_29811; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29813 = 10'h50 == _T_442[9:0] ? 4'he : _GEN_29812; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29814 = 10'h51 == _T_442[9:0] ? 4'he : _GEN_29813; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29815 = 10'h52 == _T_442[9:0] ? 4'he : _GEN_29814; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29816 = 10'h53 == _T_442[9:0] ? 4'he : _GEN_29815; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29817 = 10'h54 == _T_442[9:0] ? 4'he : _GEN_29816; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29818 = 10'h55 == _T_442[9:0] ? 4'he : _GEN_29817; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29819 = 10'h56 == _T_442[9:0] ? 4'he : _GEN_29818; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29820 = 10'h57 == _T_442[9:0] ? 4'he : _GEN_29819; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29821 = 10'h58 == _T_442[9:0] ? 4'he : _GEN_29820; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29822 = 10'h59 == _T_442[9:0] ? 4'he : _GEN_29821; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29823 = 10'h5a == _T_442[9:0] ? 4'hc : _GEN_29822; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29824 = 10'h5b == _T_442[9:0] ? 4'hd : _GEN_29823; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29825 = 10'h5c == _T_442[9:0] ? 4'he : _GEN_29824; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29826 = 10'h5d == _T_442[9:0] ? 4'he : _GEN_29825; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29827 = 10'h5e == _T_442[9:0] ? 4'he : _GEN_29826; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29828 = 10'h5f == _T_442[9:0] ? 4'he : _GEN_29827; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29829 = 10'h60 == _T_442[9:0] ? 4'he : _GEN_29828; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29830 = 10'h61 == _T_442[9:0] ? 4'hd : _GEN_29829; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29831 = 10'h62 == _T_442[9:0] ? 4'hb : _GEN_29830; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29832 = 10'h63 == _T_442[9:0] ? 4'hc : _GEN_29831; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29833 = 10'h64 == _T_442[9:0] ? 4'ha : _GEN_29832; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29834 = 10'h65 == _T_442[9:0] ? 4'hd : _GEN_29833; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29835 = 10'h66 == _T_442[9:0] ? 4'he : _GEN_29834; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29836 = 10'h67 == _T_442[9:0] ? 4'he : _GEN_29835; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29837 = 10'h68 == _T_442[9:0] ? 4'he : _GEN_29836; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29838 = 10'h69 == _T_442[9:0] ? 4'he : _GEN_29837; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29839 = 10'h6a == _T_442[9:0] ? 4'he : _GEN_29838; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29840 = 10'h6b == _T_442[9:0] ? 4'hd : _GEN_29839; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29841 = 10'h6c == _T_442[9:0] ? 4'hc : _GEN_29840; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29842 = 10'h6d == _T_442[9:0] ? 4'hc : _GEN_29841; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29843 = 10'h6e == _T_442[9:0] ? 4'he : _GEN_29842; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29844 = 10'h6f == _T_442[9:0] ? 4'he : _GEN_29843; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29845 = 10'h70 == _T_442[9:0] ? 4'he : _GEN_29844; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29846 = 10'h71 == _T_442[9:0] ? 4'he : _GEN_29845; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29847 = 10'h72 == _T_442[9:0] ? 4'he : _GEN_29846; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29848 = 10'h73 == _T_442[9:0] ? 4'he : _GEN_29847; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29849 = 10'h74 == _T_442[9:0] ? 4'he : _GEN_29848; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29850 = 10'h75 == _T_442[9:0] ? 4'he : _GEN_29849; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29851 = 10'h76 == _T_442[9:0] ? 4'he : _GEN_29850; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29852 = 10'h77 == _T_442[9:0] ? 4'he : _GEN_29851; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29853 = 10'h78 == _T_442[9:0] ? 4'he : _GEN_29852; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29854 = 10'h79 == _T_442[9:0] ? 4'he : _GEN_29853; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29855 = 10'h7a == _T_442[9:0] ? 4'he : _GEN_29854; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29856 = 10'h7b == _T_442[9:0] ? 4'he : _GEN_29855; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29857 = 10'h7c == _T_442[9:0] ? 4'he : _GEN_29856; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29858 = 10'h7d == _T_442[9:0] ? 4'he : _GEN_29857; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29859 = 10'h7e == _T_442[9:0] ? 4'he : _GEN_29858; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29860 = 10'h7f == _T_442[9:0] ? 4'he : _GEN_29859; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29861 = 10'h80 == _T_442[9:0] ? 4'he : _GEN_29860; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29862 = 10'h81 == _T_442[9:0] ? 4'hb : _GEN_29861; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29863 = 10'h82 == _T_442[9:0] ? 4'hc : _GEN_29862; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29864 = 10'h83 == _T_442[9:0] ? 4'hc : _GEN_29863; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29865 = 10'h84 == _T_442[9:0] ? 4'he : _GEN_29864; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29866 = 10'h85 == _T_442[9:0] ? 4'he : _GEN_29865; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29867 = 10'h86 == _T_442[9:0] ? 4'he : _GEN_29866; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29868 = 10'h87 == _T_442[9:0] ? 4'ha : _GEN_29867; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29869 = 10'h88 == _T_442[9:0] ? 4'hd : _GEN_29868; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29870 = 10'h89 == _T_442[9:0] ? 4'hd : _GEN_29869; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29871 = 10'h8a == _T_442[9:0] ? 4'hc : _GEN_29870; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29872 = 10'h8b == _T_442[9:0] ? 4'he : _GEN_29871; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29873 = 10'h8c == _T_442[9:0] ? 4'he : _GEN_29872; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29874 = 10'h8d == _T_442[9:0] ? 4'he : _GEN_29873; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29875 = 10'h8e == _T_442[9:0] ? 4'he : _GEN_29874; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29876 = 10'h8f == _T_442[9:0] ? 4'hb : _GEN_29875; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29877 = 10'h90 == _T_442[9:0] ? 4'hc : _GEN_29876; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29878 = 10'h91 == _T_442[9:0] ? 4'hc : _GEN_29877; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29879 = 10'h92 == _T_442[9:0] ? 4'hd : _GEN_29878; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29880 = 10'h93 == _T_442[9:0] ? 4'he : _GEN_29879; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29881 = 10'h94 == _T_442[9:0] ? 4'he : _GEN_29880; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29882 = 10'h95 == _T_442[9:0] ? 4'he : _GEN_29881; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29883 = 10'h96 == _T_442[9:0] ? 4'he : _GEN_29882; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29884 = 10'h97 == _T_442[9:0] ? 4'he : _GEN_29883; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29885 = 10'h98 == _T_442[9:0] ? 4'he : _GEN_29884; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29886 = 10'h99 == _T_442[9:0] ? 4'he : _GEN_29885; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29887 = 10'h9a == _T_442[9:0] ? 4'he : _GEN_29886; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29888 = 10'h9b == _T_442[9:0] ? 4'he : _GEN_29887; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29889 = 10'h9c == _T_442[9:0] ? 4'he : _GEN_29888; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29890 = 10'h9d == _T_442[9:0] ? 4'he : _GEN_29889; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29891 = 10'h9e == _T_442[9:0] ? 4'he : _GEN_29890; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29892 = 10'h9f == _T_442[9:0] ? 4'he : _GEN_29891; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29893 = 10'ha0 == _T_442[9:0] ? 4'he : _GEN_29892; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29894 = 10'ha1 == _T_442[9:0] ? 4'he : _GEN_29893; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29895 = 10'ha2 == _T_442[9:0] ? 4'he : _GEN_29894; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29896 = 10'ha3 == _T_442[9:0] ? 4'he : _GEN_29895; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29897 = 10'ha4 == _T_442[9:0] ? 4'he : _GEN_29896; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29898 = 10'ha5 == _T_442[9:0] ? 4'he : _GEN_29897; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29899 = 10'ha6 == _T_442[9:0] ? 4'he : _GEN_29898; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29900 = 10'ha7 == _T_442[9:0] ? 4'he : _GEN_29899; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29901 = 10'ha8 == _T_442[9:0] ? 4'hb : _GEN_29900; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29902 = 10'ha9 == _T_442[9:0] ? 4'hc : _GEN_29901; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29903 = 10'haa == _T_442[9:0] ? 4'hb : _GEN_29902; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29904 = 10'hab == _T_442[9:0] ? 4'hc : _GEN_29903; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29905 = 10'hac == _T_442[9:0] ? 4'hd : _GEN_29904; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29906 = 10'had == _T_442[9:0] ? 4'ha : _GEN_29905; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29907 = 10'hae == _T_442[9:0] ? 4'hd : _GEN_29906; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29908 = 10'haf == _T_442[9:0] ? 4'hd : _GEN_29907; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29909 = 10'hb0 == _T_442[9:0] ? 4'hb : _GEN_29908; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29910 = 10'hb1 == _T_442[9:0] ? 4'hc : _GEN_29909; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29911 = 10'hb2 == _T_442[9:0] ? 4'he : _GEN_29910; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29912 = 10'hb3 == _T_442[9:0] ? 4'hb : _GEN_29911; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29913 = 10'hb4 == _T_442[9:0] ? 4'hc : _GEN_29912; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29914 = 10'hb5 == _T_442[9:0] ? 4'hd : _GEN_29913; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29915 = 10'hb6 == _T_442[9:0] ? 4'hd : _GEN_29914; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29916 = 10'hb7 == _T_442[9:0] ? 4'hc : _GEN_29915; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29917 = 10'hb8 == _T_442[9:0] ? 4'he : _GEN_29916; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29918 = 10'hb9 == _T_442[9:0] ? 4'he : _GEN_29917; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29919 = 10'hba == _T_442[9:0] ? 4'he : _GEN_29918; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29920 = 10'hbb == _T_442[9:0] ? 4'he : _GEN_29919; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29921 = 10'hbc == _T_442[9:0] ? 4'he : _GEN_29920; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29922 = 10'hbd == _T_442[9:0] ? 4'he : _GEN_29921; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29923 = 10'hbe == _T_442[9:0] ? 4'he : _GEN_29922; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29924 = 10'hbf == _T_442[9:0] ? 4'he : _GEN_29923; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29925 = 10'hc0 == _T_442[9:0] ? 4'he : _GEN_29924; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29926 = 10'hc1 == _T_442[9:0] ? 4'he : _GEN_29925; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29927 = 10'hc2 == _T_442[9:0] ? 4'he : _GEN_29926; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29928 = 10'hc3 == _T_442[9:0] ? 4'he : _GEN_29927; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29929 = 10'hc4 == _T_442[9:0] ? 4'he : _GEN_29928; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29930 = 10'hc5 == _T_442[9:0] ? 4'he : _GEN_29929; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29931 = 10'hc6 == _T_442[9:0] ? 4'he : _GEN_29930; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29932 = 10'hc7 == _T_442[9:0] ? 4'hd : _GEN_29931; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29933 = 10'hc8 == _T_442[9:0] ? 4'hb : _GEN_29932; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29934 = 10'hc9 == _T_442[9:0] ? 4'hc : _GEN_29933; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29935 = 10'hca == _T_442[9:0] ? 4'he : _GEN_29934; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29936 = 10'hcb == _T_442[9:0] ? 4'he : _GEN_29935; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29937 = 10'hcc == _T_442[9:0] ? 4'he : _GEN_29936; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29938 = 10'hcd == _T_442[9:0] ? 4'he : _GEN_29937; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29939 = 10'hce == _T_442[9:0] ? 4'hd : _GEN_29938; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29940 = 10'hcf == _T_442[9:0] ? 4'hb : _GEN_29939; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29941 = 10'hd0 == _T_442[9:0] ? 4'hc : _GEN_29940; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29942 = 10'hd1 == _T_442[9:0] ? 4'hc : _GEN_29941; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29943 = 10'hd2 == _T_442[9:0] ? 4'hb : _GEN_29942; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29944 = 10'hd3 == _T_442[9:0] ? 4'hd : _GEN_29943; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29945 = 10'hd4 == _T_442[9:0] ? 4'hd : _GEN_29944; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29946 = 10'hd5 == _T_442[9:0] ? 4'hd : _GEN_29945; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29947 = 10'hd6 == _T_442[9:0] ? 4'hd : _GEN_29946; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29948 = 10'hd7 == _T_442[9:0] ? 4'hc : _GEN_29947; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29949 = 10'hd8 == _T_442[9:0] ? 4'hc : _GEN_29948; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29950 = 10'hd9 == _T_442[9:0] ? 4'hc : _GEN_29949; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29951 = 10'hda == _T_442[9:0] ? 4'hd : _GEN_29950; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29952 = 10'hdb == _T_442[9:0] ? 4'hc : _GEN_29951; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29953 = 10'hdc == _T_442[9:0] ? 4'h9 : _GEN_29952; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29954 = 10'hdd == _T_442[9:0] ? 4'he : _GEN_29953; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29955 = 10'hde == _T_442[9:0] ? 4'he : _GEN_29954; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29956 = 10'hdf == _T_442[9:0] ? 4'he : _GEN_29955; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29957 = 10'he0 == _T_442[9:0] ? 4'he : _GEN_29956; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29958 = 10'he1 == _T_442[9:0] ? 4'he : _GEN_29957; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29959 = 10'he2 == _T_442[9:0] ? 4'he : _GEN_29958; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29960 = 10'he3 == _T_442[9:0] ? 4'h9 : _GEN_29959; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29961 = 10'he4 == _T_442[9:0] ? 4'he : _GEN_29960; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29962 = 10'he5 == _T_442[9:0] ? 4'he : _GEN_29961; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29963 = 10'he6 == _T_442[9:0] ? 4'he : _GEN_29962; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29964 = 10'he7 == _T_442[9:0] ? 4'he : _GEN_29963; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29965 = 10'he8 == _T_442[9:0] ? 4'he : _GEN_29964; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29966 = 10'he9 == _T_442[9:0] ? 4'he : _GEN_29965; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29967 = 10'hea == _T_442[9:0] ? 4'he : _GEN_29966; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29968 = 10'heb == _T_442[9:0] ? 4'hc : _GEN_29967; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29969 = 10'hec == _T_442[9:0] ? 4'h7 : _GEN_29968; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29970 = 10'hed == _T_442[9:0] ? 4'h1 : _GEN_29969; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29971 = 10'hee == _T_442[9:0] ? 4'h0 : _GEN_29970; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29972 = 10'hef == _T_442[9:0] ? 4'h0 : _GEN_29971; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29973 = 10'hf0 == _T_442[9:0] ? 4'h2 : _GEN_29972; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29974 = 10'hf1 == _T_442[9:0] ? 4'h9 : _GEN_29973; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29975 = 10'hf2 == _T_442[9:0] ? 4'he : _GEN_29974; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29976 = 10'hf3 == _T_442[9:0] ? 4'he : _GEN_29975; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29977 = 10'hf4 == _T_442[9:0] ? 4'he : _GEN_29976; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29978 = 10'hf5 == _T_442[9:0] ? 4'hc : _GEN_29977; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29979 = 10'hf6 == _T_442[9:0] ? 4'hc : _GEN_29978; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29980 = 10'hf7 == _T_442[9:0] ? 4'hd : _GEN_29979; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29981 = 10'hf8 == _T_442[9:0] ? 4'hd : _GEN_29980; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29982 = 10'hf9 == _T_442[9:0] ? 4'hd : _GEN_29981; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29983 = 10'hfa == _T_442[9:0] ? 4'hd : _GEN_29982; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29984 = 10'hfb == _T_442[9:0] ? 4'hd : _GEN_29983; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29985 = 10'hfc == _T_442[9:0] ? 4'hd : _GEN_29984; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29986 = 10'hfd == _T_442[9:0] ? 4'hd : _GEN_29985; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29987 = 10'hfe == _T_442[9:0] ? 4'hd : _GEN_29986; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29988 = 10'hff == _T_442[9:0] ? 4'hd : _GEN_29987; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29989 = 10'h100 == _T_442[9:0] ? 4'hd : _GEN_29988; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29990 = 10'h101 == _T_442[9:0] ? 4'h9 : _GEN_29989; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29991 = 10'h102 == _T_442[9:0] ? 4'h9 : _GEN_29990; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29992 = 10'h103 == _T_442[9:0] ? 4'he : _GEN_29991; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29993 = 10'h104 == _T_442[9:0] ? 4'he : _GEN_29992; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29994 = 10'h105 == _T_442[9:0] ? 4'he : _GEN_29993; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29995 = 10'h106 == _T_442[9:0] ? 4'he : _GEN_29994; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29996 = 10'h107 == _T_442[9:0] ? 4'he : _GEN_29995; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29997 = 10'h108 == _T_442[9:0] ? 4'he : _GEN_29996; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29998 = 10'h109 == _T_442[9:0] ? 4'h6 : _GEN_29997; // @[Filter.scala 230:102]
  wire [3:0] _GEN_29999 = 10'h10a == _T_442[9:0] ? 4'he : _GEN_29998; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30000 = 10'h10b == _T_442[9:0] ? 4'he : _GEN_29999; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30001 = 10'h10c == _T_442[9:0] ? 4'he : _GEN_30000; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30002 = 10'h10d == _T_442[9:0] ? 4'he : _GEN_30001; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30003 = 10'h10e == _T_442[9:0] ? 4'he : _GEN_30002; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30004 = 10'h10f == _T_442[9:0] ? 4'ha : _GEN_30003; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30005 = 10'h110 == _T_442[9:0] ? 4'hd : _GEN_30004; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30006 = 10'h111 == _T_442[9:0] ? 4'h4 : _GEN_30005; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30007 = 10'h112 == _T_442[9:0] ? 4'h7 : _GEN_30006; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30008 = 10'h113 == _T_442[9:0] ? 4'h0 : _GEN_30007; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30009 = 10'h114 == _T_442[9:0] ? 4'h0 : _GEN_30008; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30010 = 10'h115 == _T_442[9:0] ? 4'h0 : _GEN_30009; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30011 = 10'h116 == _T_442[9:0] ? 4'h0 : _GEN_30010; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30012 = 10'h117 == _T_442[9:0] ? 4'h0 : _GEN_30011; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30013 = 10'h118 == _T_442[9:0] ? 4'ha : _GEN_30012; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30014 = 10'h119 == _T_442[9:0] ? 4'he : _GEN_30013; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30015 = 10'h11a == _T_442[9:0] ? 4'he : _GEN_30014; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30016 = 10'h11b == _T_442[9:0] ? 4'he : _GEN_30015; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30017 = 10'h11c == _T_442[9:0] ? 4'hb : _GEN_30016; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30018 = 10'h11d == _T_442[9:0] ? 4'hc : _GEN_30017; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30019 = 10'h11e == _T_442[9:0] ? 4'hd : _GEN_30018; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30020 = 10'h11f == _T_442[9:0] ? 4'hb : _GEN_30019; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30021 = 10'h120 == _T_442[9:0] ? 4'ha : _GEN_30020; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30022 = 10'h121 == _T_442[9:0] ? 4'hc : _GEN_30021; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30023 = 10'h122 == _T_442[9:0] ? 4'ha : _GEN_30022; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30024 = 10'h123 == _T_442[9:0] ? 4'ha : _GEN_30023; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30025 = 10'h124 == _T_442[9:0] ? 4'hd : _GEN_30024; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30026 = 10'h125 == _T_442[9:0] ? 4'hd : _GEN_30025; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30027 = 10'h126 == _T_442[9:0] ? 4'hb : _GEN_30026; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30028 = 10'h127 == _T_442[9:0] ? 4'h9 : _GEN_30027; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30029 = 10'h128 == _T_442[9:0] ? 4'h7 : _GEN_30028; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30030 = 10'h129 == _T_442[9:0] ? 4'hd : _GEN_30029; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30031 = 10'h12a == _T_442[9:0] ? 4'hc : _GEN_30030; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30032 = 10'h12b == _T_442[9:0] ? 4'hb : _GEN_30031; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30033 = 10'h12c == _T_442[9:0] ? 4'hc : _GEN_30032; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30034 = 10'h12d == _T_442[9:0] ? 4'hb : _GEN_30033; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30035 = 10'h12e == _T_442[9:0] ? 4'ha : _GEN_30034; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30036 = 10'h12f == _T_442[9:0] ? 4'h6 : _GEN_30035; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30037 = 10'h130 == _T_442[9:0] ? 4'he : _GEN_30036; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30038 = 10'h131 == _T_442[9:0] ? 4'hc : _GEN_30037; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30039 = 10'h132 == _T_442[9:0] ? 4'ha : _GEN_30038; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30040 = 10'h133 == _T_442[9:0] ? 4'h9 : _GEN_30039; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30041 = 10'h134 == _T_442[9:0] ? 4'hb : _GEN_30040; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30042 = 10'h135 == _T_442[9:0] ? 4'h8 : _GEN_30041; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30043 = 10'h136 == _T_442[9:0] ? 4'h8 : _GEN_30042; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30044 = 10'h137 == _T_442[9:0] ? 4'h4 : _GEN_30043; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30045 = 10'h138 == _T_442[9:0] ? 4'h7 : _GEN_30044; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30046 = 10'h139 == _T_442[9:0] ? 4'h0 : _GEN_30045; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30047 = 10'h13a == _T_442[9:0] ? 4'h0 : _GEN_30046; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30048 = 10'h13b == _T_442[9:0] ? 4'h0 : _GEN_30047; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30049 = 10'h13c == _T_442[9:0] ? 4'h0 : _GEN_30048; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30050 = 10'h13d == _T_442[9:0] ? 4'h0 : _GEN_30049; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30051 = 10'h13e == _T_442[9:0] ? 4'h4 : _GEN_30050; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30052 = 10'h13f == _T_442[9:0] ? 4'hc : _GEN_30051; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30053 = 10'h140 == _T_442[9:0] ? 4'he : _GEN_30052; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30054 = 10'h141 == _T_442[9:0] ? 4'he : _GEN_30053; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30055 = 10'h142 == _T_442[9:0] ? 4'he : _GEN_30054; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30056 = 10'h143 == _T_442[9:0] ? 4'hc : _GEN_30055; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30057 = 10'h144 == _T_442[9:0] ? 4'hd : _GEN_30056; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30058 = 10'h145 == _T_442[9:0] ? 4'hb : _GEN_30057; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30059 = 10'h146 == _T_442[9:0] ? 4'hb : _GEN_30058; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30060 = 10'h147 == _T_442[9:0] ? 4'ha : _GEN_30059; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30061 = 10'h148 == _T_442[9:0] ? 4'ha : _GEN_30060; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30062 = 10'h149 == _T_442[9:0] ? 4'hc : _GEN_30061; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30063 = 10'h14a == _T_442[9:0] ? 4'hd : _GEN_30062; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30064 = 10'h14b == _T_442[9:0] ? 4'hc : _GEN_30063; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30065 = 10'h14c == _T_442[9:0] ? 4'hd : _GEN_30064; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30066 = 10'h14d == _T_442[9:0] ? 4'h9 : _GEN_30065; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30067 = 10'h14e == _T_442[9:0] ? 4'h7 : _GEN_30066; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30068 = 10'h14f == _T_442[9:0] ? 4'ha : _GEN_30067; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30069 = 10'h150 == _T_442[9:0] ? 4'ha : _GEN_30068; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30070 = 10'h151 == _T_442[9:0] ? 4'hb : _GEN_30069; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30071 = 10'h152 == _T_442[9:0] ? 4'hb : _GEN_30070; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30072 = 10'h153 == _T_442[9:0] ? 4'hc : _GEN_30071; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30073 = 10'h154 == _T_442[9:0] ? 4'hb : _GEN_30072; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30074 = 10'h155 == _T_442[9:0] ? 4'h6 : _GEN_30073; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30075 = 10'h156 == _T_442[9:0] ? 4'hb : _GEN_30074; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30076 = 10'h157 == _T_442[9:0] ? 4'h7 : _GEN_30075; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30077 = 10'h158 == _T_442[9:0] ? 4'h7 : _GEN_30076; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30078 = 10'h159 == _T_442[9:0] ? 4'h7 : _GEN_30077; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30079 = 10'h15a == _T_442[9:0] ? 4'h7 : _GEN_30078; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30080 = 10'h15b == _T_442[9:0] ? 4'h7 : _GEN_30079; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30081 = 10'h15c == _T_442[9:0] ? 4'h7 : _GEN_30080; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30082 = 10'h15d == _T_442[9:0] ? 4'h6 : _GEN_30081; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30083 = 10'h15e == _T_442[9:0] ? 4'h7 : _GEN_30082; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30084 = 10'h15f == _T_442[9:0] ? 4'h0 : _GEN_30083; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30085 = 10'h160 == _T_442[9:0] ? 4'h0 : _GEN_30084; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30086 = 10'h161 == _T_442[9:0] ? 4'h0 : _GEN_30085; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30087 = 10'h162 == _T_442[9:0] ? 4'h0 : _GEN_30086; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30088 = 10'h163 == _T_442[9:0] ? 4'h2 : _GEN_30087; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30089 = 10'h164 == _T_442[9:0] ? 4'h4 : _GEN_30088; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30090 = 10'h165 == _T_442[9:0] ? 4'hb : _GEN_30089; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30091 = 10'h166 == _T_442[9:0] ? 4'hb : _GEN_30090; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30092 = 10'h167 == _T_442[9:0] ? 4'he : _GEN_30091; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30093 = 10'h168 == _T_442[9:0] ? 4'he : _GEN_30092; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30094 = 10'h169 == _T_442[9:0] ? 4'hc : _GEN_30093; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30095 = 10'h16a == _T_442[9:0] ? 4'hd : _GEN_30094; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30096 = 10'h16b == _T_442[9:0] ? 4'hd : _GEN_30095; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30097 = 10'h16c == _T_442[9:0] ? 4'ha : _GEN_30096; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30098 = 10'h16d == _T_442[9:0] ? 4'ha : _GEN_30097; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30099 = 10'h16e == _T_442[9:0] ? 4'ha : _GEN_30098; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30100 = 10'h16f == _T_442[9:0] ? 4'hd : _GEN_30099; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30101 = 10'h170 == _T_442[9:0] ? 4'hd : _GEN_30100; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30102 = 10'h171 == _T_442[9:0] ? 4'hd : _GEN_30101; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30103 = 10'h172 == _T_442[9:0] ? 4'he : _GEN_30102; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30104 = 10'h173 == _T_442[9:0] ? 4'h8 : _GEN_30103; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30105 = 10'h174 == _T_442[9:0] ? 4'h5 : _GEN_30104; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30106 = 10'h175 == _T_442[9:0] ? 4'h6 : _GEN_30105; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30107 = 10'h176 == _T_442[9:0] ? 4'h6 : _GEN_30106; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30108 = 10'h177 == _T_442[9:0] ? 4'h6 : _GEN_30107; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30109 = 10'h178 == _T_442[9:0] ? 4'h7 : _GEN_30108; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30110 = 10'h179 == _T_442[9:0] ? 4'h9 : _GEN_30109; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30111 = 10'h17a == _T_442[9:0] ? 4'h9 : _GEN_30110; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30112 = 10'h17b == _T_442[9:0] ? 4'h6 : _GEN_30111; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30113 = 10'h17c == _T_442[9:0] ? 4'h7 : _GEN_30112; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30114 = 10'h17d == _T_442[9:0] ? 4'h7 : _GEN_30113; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30115 = 10'h17e == _T_442[9:0] ? 4'h7 : _GEN_30114; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30116 = 10'h17f == _T_442[9:0] ? 4'h7 : _GEN_30115; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30117 = 10'h180 == _T_442[9:0] ? 4'h7 : _GEN_30116; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30118 = 10'h181 == _T_442[9:0] ? 4'h7 : _GEN_30117; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30119 = 10'h182 == _T_442[9:0] ? 4'h8 : _GEN_30118; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30120 = 10'h183 == _T_442[9:0] ? 4'h8 : _GEN_30119; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30121 = 10'h184 == _T_442[9:0] ? 4'h8 : _GEN_30120; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30122 = 10'h185 == _T_442[9:0] ? 4'h7 : _GEN_30121; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30123 = 10'h186 == _T_442[9:0] ? 4'h1 : _GEN_30122; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30124 = 10'h187 == _T_442[9:0] ? 4'h0 : _GEN_30123; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30125 = 10'h188 == _T_442[9:0] ? 4'h0 : _GEN_30124; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30126 = 10'h189 == _T_442[9:0] ? 4'h4 : _GEN_30125; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30127 = 10'h18a == _T_442[9:0] ? 4'h4 : _GEN_30126; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30128 = 10'h18b == _T_442[9:0] ? 4'hb : _GEN_30127; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30129 = 10'h18c == _T_442[9:0] ? 4'hb : _GEN_30128; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30130 = 10'h18d == _T_442[9:0] ? 4'hc : _GEN_30129; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30131 = 10'h18e == _T_442[9:0] ? 4'he : _GEN_30130; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30132 = 10'h18f == _T_442[9:0] ? 4'hb : _GEN_30131; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30133 = 10'h190 == _T_442[9:0] ? 4'hd : _GEN_30132; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30134 = 10'h191 == _T_442[9:0] ? 4'hc : _GEN_30133; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30135 = 10'h192 == _T_442[9:0] ? 4'h9 : _GEN_30134; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30136 = 10'h193 == _T_442[9:0] ? 4'ha : _GEN_30135; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30137 = 10'h194 == _T_442[9:0] ? 4'h9 : _GEN_30136; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30138 = 10'h195 == _T_442[9:0] ? 4'hd : _GEN_30137; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30139 = 10'h196 == _T_442[9:0] ? 4'hd : _GEN_30138; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30140 = 10'h197 == _T_442[9:0] ? 4'hb : _GEN_30139; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30141 = 10'h198 == _T_442[9:0] ? 4'he : _GEN_30140; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30142 = 10'h199 == _T_442[9:0] ? 4'h5 : _GEN_30141; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30143 = 10'h19a == _T_442[9:0] ? 4'h1 : _GEN_30142; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30144 = 10'h19b == _T_442[9:0] ? 4'h3 : _GEN_30143; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30145 = 10'h19c == _T_442[9:0] ? 4'h6 : _GEN_30144; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30146 = 10'h19d == _T_442[9:0] ? 4'h4 : _GEN_30145; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30147 = 10'h19e == _T_442[9:0] ? 4'h1 : _GEN_30146; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30148 = 10'h19f == _T_442[9:0] ? 4'h3 : _GEN_30147; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30149 = 10'h1a0 == _T_442[9:0] ? 4'h6 : _GEN_30148; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30150 = 10'h1a1 == _T_442[9:0] ? 4'h6 : _GEN_30149; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30151 = 10'h1a2 == _T_442[9:0] ? 4'h7 : _GEN_30150; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30152 = 10'h1a3 == _T_442[9:0] ? 4'h7 : _GEN_30151; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30153 = 10'h1a4 == _T_442[9:0] ? 4'h7 : _GEN_30152; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30154 = 10'h1a5 == _T_442[9:0] ? 4'h7 : _GEN_30153; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30155 = 10'h1a6 == _T_442[9:0] ? 4'h7 : _GEN_30154; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30156 = 10'h1a7 == _T_442[9:0] ? 4'h7 : _GEN_30155; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30157 = 10'h1a8 == _T_442[9:0] ? 4'h8 : _GEN_30156; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30158 = 10'h1a9 == _T_442[9:0] ? 4'h8 : _GEN_30157; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30159 = 10'h1aa == _T_442[9:0] ? 4'h7 : _GEN_30158; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30160 = 10'h1ab == _T_442[9:0] ? 4'h8 : _GEN_30159; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30161 = 10'h1ac == _T_442[9:0] ? 4'h8 : _GEN_30160; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30162 = 10'h1ad == _T_442[9:0] ? 4'h3 : _GEN_30161; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30163 = 10'h1ae == _T_442[9:0] ? 4'h2 : _GEN_30162; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30164 = 10'h1af == _T_442[9:0] ? 4'h8 : _GEN_30163; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30165 = 10'h1b0 == _T_442[9:0] ? 4'h6 : _GEN_30164; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30166 = 10'h1b1 == _T_442[9:0] ? 4'hb : _GEN_30165; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30167 = 10'h1b2 == _T_442[9:0] ? 4'hb : _GEN_30166; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30168 = 10'h1b3 == _T_442[9:0] ? 4'ha : _GEN_30167; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30169 = 10'h1b4 == _T_442[9:0] ? 4'he : _GEN_30168; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30170 = 10'h1b5 == _T_442[9:0] ? 4'hb : _GEN_30169; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30171 = 10'h1b6 == _T_442[9:0] ? 4'hc : _GEN_30170; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30172 = 10'h1b7 == _T_442[9:0] ? 4'ha : _GEN_30171; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30173 = 10'h1b8 == _T_442[9:0] ? 4'h9 : _GEN_30172; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30174 = 10'h1b9 == _T_442[9:0] ? 4'h9 : _GEN_30173; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30175 = 10'h1ba == _T_442[9:0] ? 4'h9 : _GEN_30174; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30176 = 10'h1bb == _T_442[9:0] ? 4'hb : _GEN_30175; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30177 = 10'h1bc == _T_442[9:0] ? 4'hd : _GEN_30176; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30178 = 10'h1bd == _T_442[9:0] ? 4'hd : _GEN_30177; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30179 = 10'h1be == _T_442[9:0] ? 4'he : _GEN_30178; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30180 = 10'h1bf == _T_442[9:0] ? 4'h7 : _GEN_30179; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30181 = 10'h1c0 == _T_442[9:0] ? 4'h6 : _GEN_30180; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30182 = 10'h1c1 == _T_442[9:0] ? 4'h6 : _GEN_30181; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30183 = 10'h1c2 == _T_442[9:0] ? 4'h5 : _GEN_30182; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30184 = 10'h1c3 == _T_442[9:0] ? 4'h5 : _GEN_30183; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30185 = 10'h1c4 == _T_442[9:0] ? 4'h4 : _GEN_30184; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30186 = 10'h1c5 == _T_442[9:0] ? 4'h5 : _GEN_30185; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30187 = 10'h1c6 == _T_442[9:0] ? 4'h6 : _GEN_30186; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30188 = 10'h1c7 == _T_442[9:0] ? 4'h6 : _GEN_30187; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30189 = 10'h1c8 == _T_442[9:0] ? 4'h7 : _GEN_30188; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30190 = 10'h1c9 == _T_442[9:0] ? 4'h7 : _GEN_30189; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30191 = 10'h1ca == _T_442[9:0] ? 4'h7 : _GEN_30190; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30192 = 10'h1cb == _T_442[9:0] ? 4'h7 : _GEN_30191; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30193 = 10'h1cc == _T_442[9:0] ? 4'h7 : _GEN_30192; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30194 = 10'h1cd == _T_442[9:0] ? 4'h8 : _GEN_30193; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30195 = 10'h1ce == _T_442[9:0] ? 4'h8 : _GEN_30194; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30196 = 10'h1cf == _T_442[9:0] ? 4'h8 : _GEN_30195; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30197 = 10'h1d0 == _T_442[9:0] ? 4'h5 : _GEN_30196; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30198 = 10'h1d1 == _T_442[9:0] ? 4'h8 : _GEN_30197; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30199 = 10'h1d2 == _T_442[9:0] ? 4'h8 : _GEN_30198; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30200 = 10'h1d3 == _T_442[9:0] ? 4'h8 : _GEN_30199; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30201 = 10'h1d4 == _T_442[9:0] ? 4'h8 : _GEN_30200; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30202 = 10'h1d5 == _T_442[9:0] ? 4'h7 : _GEN_30201; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30203 = 10'h1d6 == _T_442[9:0] ? 4'h9 : _GEN_30202; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30204 = 10'h1d7 == _T_442[9:0] ? 4'hb : _GEN_30203; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30205 = 10'h1d8 == _T_442[9:0] ? 4'hb : _GEN_30204; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30206 = 10'h1d9 == _T_442[9:0] ? 4'hb : _GEN_30205; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30207 = 10'h1da == _T_442[9:0] ? 4'ha : _GEN_30206; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30208 = 10'h1db == _T_442[9:0] ? 4'hc : _GEN_30207; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30209 = 10'h1dc == _T_442[9:0] ? 4'hb : _GEN_30208; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30210 = 10'h1dd == _T_442[9:0] ? 4'h5 : _GEN_30209; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30211 = 10'h1de == _T_442[9:0] ? 4'h9 : _GEN_30210; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30212 = 10'h1df == _T_442[9:0] ? 4'h9 : _GEN_30211; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30213 = 10'h1e0 == _T_442[9:0] ? 4'h9 : _GEN_30212; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30214 = 10'h1e1 == _T_442[9:0] ? 4'h7 : _GEN_30213; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30215 = 10'h1e2 == _T_442[9:0] ? 4'hc : _GEN_30214; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30216 = 10'h1e3 == _T_442[9:0] ? 4'hc : _GEN_30215; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30217 = 10'h1e4 == _T_442[9:0] ? 4'hd : _GEN_30216; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30218 = 10'h1e5 == _T_442[9:0] ? 4'h7 : _GEN_30217; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30219 = 10'h1e6 == _T_442[9:0] ? 4'h6 : _GEN_30218; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30220 = 10'h1e7 == _T_442[9:0] ? 4'h6 : _GEN_30219; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30221 = 10'h1e8 == _T_442[9:0] ? 4'h6 : _GEN_30220; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30222 = 10'h1e9 == _T_442[9:0] ? 4'h6 : _GEN_30221; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30223 = 10'h1ea == _T_442[9:0] ? 4'h6 : _GEN_30222; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30224 = 10'h1eb == _T_442[9:0] ? 4'h6 : _GEN_30223; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30225 = 10'h1ec == _T_442[9:0] ? 4'h6 : _GEN_30224; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30226 = 10'h1ed == _T_442[9:0] ? 4'h8 : _GEN_30225; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30227 = 10'h1ee == _T_442[9:0] ? 4'h7 : _GEN_30226; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30228 = 10'h1ef == _T_442[9:0] ? 4'h7 : _GEN_30227; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30229 = 10'h1f0 == _T_442[9:0] ? 4'h7 : _GEN_30228; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30230 = 10'h1f1 == _T_442[9:0] ? 4'h7 : _GEN_30229; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30231 = 10'h1f2 == _T_442[9:0] ? 4'h7 : _GEN_30230; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30232 = 10'h1f3 == _T_442[9:0] ? 4'h8 : _GEN_30231; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30233 = 10'h1f4 == _T_442[9:0] ? 4'h8 : _GEN_30232; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30234 = 10'h1f5 == _T_442[9:0] ? 4'h8 : _GEN_30233; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30235 = 10'h1f6 == _T_442[9:0] ? 4'ha : _GEN_30234; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30236 = 10'h1f7 == _T_442[9:0] ? 4'h8 : _GEN_30235; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30237 = 10'h1f8 == _T_442[9:0] ? 4'h8 : _GEN_30236; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30238 = 10'h1f9 == _T_442[9:0] ? 4'h9 : _GEN_30237; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30239 = 10'h1fa == _T_442[9:0] ? 4'h9 : _GEN_30238; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30240 = 10'h1fb == _T_442[9:0] ? 4'h8 : _GEN_30239; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30241 = 10'h1fc == _T_442[9:0] ? 4'hb : _GEN_30240; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30242 = 10'h1fd == _T_442[9:0] ? 4'hb : _GEN_30241; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30243 = 10'h1fe == _T_442[9:0] ? 4'hb : _GEN_30242; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30244 = 10'h1ff == _T_442[9:0] ? 4'ha : _GEN_30243; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30245 = 10'h200 == _T_442[9:0] ? 4'h3 : _GEN_30244; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30246 = 10'h201 == _T_442[9:0] ? 4'h9 : _GEN_30245; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30247 = 10'h202 == _T_442[9:0] ? 4'h5 : _GEN_30246; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30248 = 10'h203 == _T_442[9:0] ? 4'h3 : _GEN_30247; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30249 = 10'h204 == _T_442[9:0] ? 4'h4 : _GEN_30248; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30250 = 10'h205 == _T_442[9:0] ? 4'h4 : _GEN_30249; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30251 = 10'h206 == _T_442[9:0] ? 4'h4 : _GEN_30250; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30252 = 10'h207 == _T_442[9:0] ? 4'h4 : _GEN_30251; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30253 = 10'h208 == _T_442[9:0] ? 4'h8 : _GEN_30252; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30254 = 10'h209 == _T_442[9:0] ? 4'hc : _GEN_30253; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30255 = 10'h20a == _T_442[9:0] ? 4'hd : _GEN_30254; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30256 = 10'h20b == _T_442[9:0] ? 4'h7 : _GEN_30255; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30257 = 10'h20c == _T_442[9:0] ? 4'h6 : _GEN_30256; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30258 = 10'h20d == _T_442[9:0] ? 4'h6 : _GEN_30257; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30259 = 10'h20e == _T_442[9:0] ? 4'h6 : _GEN_30258; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30260 = 10'h20f == _T_442[9:0] ? 4'h5 : _GEN_30259; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30261 = 10'h210 == _T_442[9:0] ? 4'h6 : _GEN_30260; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30262 = 10'h211 == _T_442[9:0] ? 4'h6 : _GEN_30261; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30263 = 10'h212 == _T_442[9:0] ? 4'h7 : _GEN_30262; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30264 = 10'h213 == _T_442[9:0] ? 4'ha : _GEN_30263; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30265 = 10'h214 == _T_442[9:0] ? 4'h6 : _GEN_30264; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30266 = 10'h215 == _T_442[9:0] ? 4'h7 : _GEN_30265; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30267 = 10'h216 == _T_442[9:0] ? 4'h7 : _GEN_30266; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30268 = 10'h217 == _T_442[9:0] ? 4'h7 : _GEN_30267; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30269 = 10'h218 == _T_442[9:0] ? 4'h7 : _GEN_30268; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30270 = 10'h219 == _T_442[9:0] ? 4'h8 : _GEN_30269; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30271 = 10'h21a == _T_442[9:0] ? 4'h7 : _GEN_30270; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30272 = 10'h21b == _T_442[9:0] ? 4'h8 : _GEN_30271; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30273 = 10'h21c == _T_442[9:0] ? 4'hb : _GEN_30272; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30274 = 10'h21d == _T_442[9:0] ? 4'ha : _GEN_30273; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30275 = 10'h21e == _T_442[9:0] ? 4'h9 : _GEN_30274; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30276 = 10'h21f == _T_442[9:0] ? 4'h9 : _GEN_30275; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30277 = 10'h220 == _T_442[9:0] ? 4'h8 : _GEN_30276; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30278 = 10'h221 == _T_442[9:0] ? 4'h9 : _GEN_30277; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30279 = 10'h222 == _T_442[9:0] ? 4'hb : _GEN_30278; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30280 = 10'h223 == _T_442[9:0] ? 4'hb : _GEN_30279; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30281 = 10'h224 == _T_442[9:0] ? 4'hb : _GEN_30280; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30282 = 10'h225 == _T_442[9:0] ? 4'h8 : _GEN_30281; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30283 = 10'h226 == _T_442[9:0] ? 4'h1 : _GEN_30282; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30284 = 10'h227 == _T_442[9:0] ? 4'h3 : _GEN_30283; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30285 = 10'h228 == _T_442[9:0] ? 4'h3 : _GEN_30284; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30286 = 10'h229 == _T_442[9:0] ? 4'h3 : _GEN_30285; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30287 = 10'h22a == _T_442[9:0] ? 4'h3 : _GEN_30286; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30288 = 10'h22b == _T_442[9:0] ? 4'h3 : _GEN_30287; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30289 = 10'h22c == _T_442[9:0] ? 4'h3 : _GEN_30288; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30290 = 10'h22d == _T_442[9:0] ? 4'h3 : _GEN_30289; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30291 = 10'h22e == _T_442[9:0] ? 4'h3 : _GEN_30290; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30292 = 10'h22f == _T_442[9:0] ? 4'h9 : _GEN_30291; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30293 = 10'h230 == _T_442[9:0] ? 4'h6 : _GEN_30292; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30294 = 10'h231 == _T_442[9:0] ? 4'h7 : _GEN_30293; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30295 = 10'h232 == _T_442[9:0] ? 4'h6 : _GEN_30294; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30296 = 10'h233 == _T_442[9:0] ? 4'h7 : _GEN_30295; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30297 = 10'h234 == _T_442[9:0] ? 4'h7 : _GEN_30296; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30298 = 10'h235 == _T_442[9:0] ? 4'h6 : _GEN_30297; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30299 = 10'h236 == _T_442[9:0] ? 4'h6 : _GEN_30298; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30300 = 10'h237 == _T_442[9:0] ? 4'h6 : _GEN_30299; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30301 = 10'h238 == _T_442[9:0] ? 4'h6 : _GEN_30300; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30302 = 10'h239 == _T_442[9:0] ? 4'h8 : _GEN_30301; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30303 = 10'h23a == _T_442[9:0] ? 4'h6 : _GEN_30302; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30304 = 10'h23b == _T_442[9:0] ? 4'h7 : _GEN_30303; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30305 = 10'h23c == _T_442[9:0] ? 4'h7 : _GEN_30304; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30306 = 10'h23d == _T_442[9:0] ? 4'h7 : _GEN_30305; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30307 = 10'h23e == _T_442[9:0] ? 4'h7 : _GEN_30306; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30308 = 10'h23f == _T_442[9:0] ? 4'h7 : _GEN_30307; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30309 = 10'h240 == _T_442[9:0] ? 4'h7 : _GEN_30308; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30310 = 10'h241 == _T_442[9:0] ? 4'h8 : _GEN_30309; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30311 = 10'h242 == _T_442[9:0] ? 4'hb : _GEN_30310; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30312 = 10'h243 == _T_442[9:0] ? 4'hb : _GEN_30311; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30313 = 10'h244 == _T_442[9:0] ? 4'hb : _GEN_30312; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30314 = 10'h245 == _T_442[9:0] ? 4'ha : _GEN_30313; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30315 = 10'h246 == _T_442[9:0] ? 4'h9 : _GEN_30314; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30316 = 10'h247 == _T_442[9:0] ? 4'ha : _GEN_30315; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30317 = 10'h248 == _T_442[9:0] ? 4'hb : _GEN_30316; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30318 = 10'h249 == _T_442[9:0] ? 4'hb : _GEN_30317; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30319 = 10'h24a == _T_442[9:0] ? 4'ha : _GEN_30318; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30320 = 10'h24b == _T_442[9:0] ? 4'h2 : _GEN_30319; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30321 = 10'h24c == _T_442[9:0] ? 4'h0 : _GEN_30320; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30322 = 10'h24d == _T_442[9:0] ? 4'h2 : _GEN_30321; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30323 = 10'h24e == _T_442[9:0] ? 4'h3 : _GEN_30322; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30324 = 10'h24f == _T_442[9:0] ? 4'h3 : _GEN_30323; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30325 = 10'h250 == _T_442[9:0] ? 4'h3 : _GEN_30324; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30326 = 10'h251 == _T_442[9:0] ? 4'h3 : _GEN_30325; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30327 = 10'h252 == _T_442[9:0] ? 4'h3 : _GEN_30326; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30328 = 10'h253 == _T_442[9:0] ? 4'h3 : _GEN_30327; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30329 = 10'h254 == _T_442[9:0] ? 4'h3 : _GEN_30328; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30330 = 10'h255 == _T_442[9:0] ? 4'h5 : _GEN_30329; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30331 = 10'h256 == _T_442[9:0] ? 4'h6 : _GEN_30330; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30332 = 10'h257 == _T_442[9:0] ? 4'h8 : _GEN_30331; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30333 = 10'h258 == _T_442[9:0] ? 4'h5 : _GEN_30332; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30334 = 10'h259 == _T_442[9:0] ? 4'h6 : _GEN_30333; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30335 = 10'h25a == _T_442[9:0] ? 4'h6 : _GEN_30334; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30336 = 10'h25b == _T_442[9:0] ? 4'h5 : _GEN_30335; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30337 = 10'h25c == _T_442[9:0] ? 4'h6 : _GEN_30336; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30338 = 10'h25d == _T_442[9:0] ? 4'h6 : _GEN_30337; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30339 = 10'h25e == _T_442[9:0] ? 4'h9 : _GEN_30338; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30340 = 10'h25f == _T_442[9:0] ? 4'hc : _GEN_30339; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30341 = 10'h260 == _T_442[9:0] ? 4'h7 : _GEN_30340; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30342 = 10'h261 == _T_442[9:0] ? 4'h9 : _GEN_30341; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30343 = 10'h262 == _T_442[9:0] ? 4'ha : _GEN_30342; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30344 = 10'h263 == _T_442[9:0] ? 4'h8 : _GEN_30343; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30345 = 10'h264 == _T_442[9:0] ? 4'ha : _GEN_30344; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30346 = 10'h265 == _T_442[9:0] ? 4'h9 : _GEN_30345; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30347 = 10'h266 == _T_442[9:0] ? 4'h8 : _GEN_30346; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30348 = 10'h267 == _T_442[9:0] ? 4'h8 : _GEN_30347; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30349 = 10'h268 == _T_442[9:0] ? 4'ha : _GEN_30348; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30350 = 10'h269 == _T_442[9:0] ? 4'ha : _GEN_30349; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30351 = 10'h26a == _T_442[9:0] ? 4'hb : _GEN_30350; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30352 = 10'h26b == _T_442[9:0] ? 4'hb : _GEN_30351; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30353 = 10'h26c == _T_442[9:0] ? 4'hb : _GEN_30352; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30354 = 10'h26d == _T_442[9:0] ? 4'hb : _GEN_30353; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30355 = 10'h26e == _T_442[9:0] ? 4'hb : _GEN_30354; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30356 = 10'h26f == _T_442[9:0] ? 4'ha : _GEN_30355; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30357 = 10'h270 == _T_442[9:0] ? 4'h3 : _GEN_30356; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30358 = 10'h271 == _T_442[9:0] ? 4'h0 : _GEN_30357; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30359 = 10'h272 == _T_442[9:0] ? 4'h0 : _GEN_30358; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30360 = 10'h273 == _T_442[9:0] ? 4'h2 : _GEN_30359; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30361 = 10'h274 == _T_442[9:0] ? 4'h3 : _GEN_30360; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30362 = 10'h275 == _T_442[9:0] ? 4'h3 : _GEN_30361; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30363 = 10'h276 == _T_442[9:0] ? 4'h3 : _GEN_30362; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30364 = 10'h277 == _T_442[9:0] ? 4'h3 : _GEN_30363; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30365 = 10'h278 == _T_442[9:0] ? 4'h3 : _GEN_30364; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30366 = 10'h279 == _T_442[9:0] ? 4'h3 : _GEN_30365; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30367 = 10'h27a == _T_442[9:0] ? 4'h3 : _GEN_30366; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30368 = 10'h27b == _T_442[9:0] ? 4'h6 : _GEN_30367; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30369 = 10'h27c == _T_442[9:0] ? 4'h7 : _GEN_30368; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30370 = 10'h27d == _T_442[9:0] ? 4'h7 : _GEN_30369; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30371 = 10'h27e == _T_442[9:0] ? 4'h4 : _GEN_30370; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30372 = 10'h27f == _T_442[9:0] ? 4'h6 : _GEN_30371; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30373 = 10'h280 == _T_442[9:0] ? 4'h6 : _GEN_30372; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30374 = 10'h281 == _T_442[9:0] ? 4'h6 : _GEN_30373; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30375 = 10'h282 == _T_442[9:0] ? 4'h6 : _GEN_30374; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30376 = 10'h283 == _T_442[9:0] ? 4'ha : _GEN_30375; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30377 = 10'h284 == _T_442[9:0] ? 4'hc : _GEN_30376; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30378 = 10'h285 == _T_442[9:0] ? 4'hc : _GEN_30377; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30379 = 10'h286 == _T_442[9:0] ? 4'h8 : _GEN_30378; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30380 = 10'h287 == _T_442[9:0] ? 4'ha : _GEN_30379; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30381 = 10'h288 == _T_442[9:0] ? 4'ha : _GEN_30380; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30382 = 10'h289 == _T_442[9:0] ? 4'ha : _GEN_30381; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30383 = 10'h28a == _T_442[9:0] ? 4'hc : _GEN_30382; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30384 = 10'h28b == _T_442[9:0] ? 4'hb : _GEN_30383; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30385 = 10'h28c == _T_442[9:0] ? 4'ha : _GEN_30384; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30386 = 10'h28d == _T_442[9:0] ? 4'h7 : _GEN_30385; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30387 = 10'h28e == _T_442[9:0] ? 4'h2 : _GEN_30386; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30388 = 10'h28f == _T_442[9:0] ? 4'h5 : _GEN_30387; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30389 = 10'h290 == _T_442[9:0] ? 4'h8 : _GEN_30388; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30390 = 10'h291 == _T_442[9:0] ? 4'ha : _GEN_30389; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30391 = 10'h292 == _T_442[9:0] ? 4'ha : _GEN_30390; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30392 = 10'h293 == _T_442[9:0] ? 4'ha : _GEN_30391; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30393 = 10'h294 == _T_442[9:0] ? 4'h9 : _GEN_30392; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30394 = 10'h295 == _T_442[9:0] ? 4'h3 : _GEN_30393; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30395 = 10'h296 == _T_442[9:0] ? 4'h0 : _GEN_30394; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30396 = 10'h297 == _T_442[9:0] ? 4'h0 : _GEN_30395; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30397 = 10'h298 == _T_442[9:0] ? 4'h0 : _GEN_30396; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30398 = 10'h299 == _T_442[9:0] ? 4'h1 : _GEN_30397; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30399 = 10'h29a == _T_442[9:0] ? 4'h3 : _GEN_30398; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30400 = 10'h29b == _T_442[9:0] ? 4'h3 : _GEN_30399; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30401 = 10'h29c == _T_442[9:0] ? 4'h3 : _GEN_30400; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30402 = 10'h29d == _T_442[9:0] ? 4'h3 : _GEN_30401; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30403 = 10'h29e == _T_442[9:0] ? 4'h3 : _GEN_30402; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30404 = 10'h29f == _T_442[9:0] ? 4'h3 : _GEN_30403; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30405 = 10'h2a0 == _T_442[9:0] ? 4'h4 : _GEN_30404; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30406 = 10'h2a1 == _T_442[9:0] ? 4'h6 : _GEN_30405; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30407 = 10'h2a2 == _T_442[9:0] ? 4'h7 : _GEN_30406; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30408 = 10'h2a3 == _T_442[9:0] ? 4'h6 : _GEN_30407; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30409 = 10'h2a4 == _T_442[9:0] ? 4'h4 : _GEN_30408; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30410 = 10'h2a5 == _T_442[9:0] ? 4'h6 : _GEN_30409; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30411 = 10'h2a6 == _T_442[9:0] ? 4'h6 : _GEN_30410; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30412 = 10'h2a7 == _T_442[9:0] ? 4'h7 : _GEN_30411; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30413 = 10'h2a8 == _T_442[9:0] ? 4'ha : _GEN_30412; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30414 = 10'h2a9 == _T_442[9:0] ? 4'hb : _GEN_30413; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30415 = 10'h2aa == _T_442[9:0] ? 4'hb : _GEN_30414; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30416 = 10'h2ab == _T_442[9:0] ? 4'hb : _GEN_30415; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30417 = 10'h2ac == _T_442[9:0] ? 4'h8 : _GEN_30416; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30418 = 10'h2ad == _T_442[9:0] ? 4'hb : _GEN_30417; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30419 = 10'h2ae == _T_442[9:0] ? 4'ha : _GEN_30418; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30420 = 10'h2af == _T_442[9:0] ? 4'hb : _GEN_30419; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30421 = 10'h2b0 == _T_442[9:0] ? 4'hc : _GEN_30420; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30422 = 10'h2b1 == _T_442[9:0] ? 4'hb : _GEN_30421; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30423 = 10'h2b2 == _T_442[9:0] ? 4'ha : _GEN_30422; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30424 = 10'h2b3 == _T_442[9:0] ? 4'h6 : _GEN_30423; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30425 = 10'h2b4 == _T_442[9:0] ? 4'h0 : _GEN_30424; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30426 = 10'h2b5 == _T_442[9:0] ? 4'h0 : _GEN_30425; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30427 = 10'h2b6 == _T_442[9:0] ? 4'h0 : _GEN_30426; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30428 = 10'h2b7 == _T_442[9:0] ? 4'h1 : _GEN_30427; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30429 = 10'h2b8 == _T_442[9:0] ? 4'h5 : _GEN_30428; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30430 = 10'h2b9 == _T_442[9:0] ? 4'h9 : _GEN_30429; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30431 = 10'h2ba == _T_442[9:0] ? 4'h1 : _GEN_30430; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30432 = 10'h2bb == _T_442[9:0] ? 4'h0 : _GEN_30431; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30433 = 10'h2bc == _T_442[9:0] ? 4'h0 : _GEN_30432; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30434 = 10'h2bd == _T_442[9:0] ? 4'h0 : _GEN_30433; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30435 = 10'h2be == _T_442[9:0] ? 4'h0 : _GEN_30434; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30436 = 10'h2bf == _T_442[9:0] ? 4'h0 : _GEN_30435; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30437 = 10'h2c0 == _T_442[9:0] ? 4'h3 : _GEN_30436; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30438 = 10'h2c1 == _T_442[9:0] ? 4'h3 : _GEN_30437; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30439 = 10'h2c2 == _T_442[9:0] ? 4'h3 : _GEN_30438; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30440 = 10'h2c3 == _T_442[9:0] ? 4'h3 : _GEN_30439; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30441 = 10'h2c4 == _T_442[9:0] ? 4'h3 : _GEN_30440; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30442 = 10'h2c5 == _T_442[9:0] ? 4'h3 : _GEN_30441; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30443 = 10'h2c6 == _T_442[9:0] ? 4'h4 : _GEN_30442; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30444 = 10'h2c7 == _T_442[9:0] ? 4'h5 : _GEN_30443; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30445 = 10'h2c8 == _T_442[9:0] ? 4'h7 : _GEN_30444; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30446 = 10'h2c9 == _T_442[9:0] ? 4'h7 : _GEN_30445; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30447 = 10'h2ca == _T_442[9:0] ? 4'h4 : _GEN_30446; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30448 = 10'h2cb == _T_442[9:0] ? 4'h9 : _GEN_30447; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30449 = 10'h2cc == _T_442[9:0] ? 4'h9 : _GEN_30448; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30450 = 10'h2cd == _T_442[9:0] ? 4'hb : _GEN_30449; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30451 = 10'h2ce == _T_442[9:0] ? 4'hb : _GEN_30450; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30452 = 10'h2cf == _T_442[9:0] ? 4'hb : _GEN_30451; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30453 = 10'h2d0 == _T_442[9:0] ? 4'hb : _GEN_30452; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30454 = 10'h2d1 == _T_442[9:0] ? 4'hb : _GEN_30453; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30455 = 10'h2d2 == _T_442[9:0] ? 4'h8 : _GEN_30454; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30456 = 10'h2d3 == _T_442[9:0] ? 4'ha : _GEN_30455; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30457 = 10'h2d4 == _T_442[9:0] ? 4'hb : _GEN_30456; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30458 = 10'h2d5 == _T_442[9:0] ? 4'ha : _GEN_30457; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30459 = 10'h2d6 == _T_442[9:0] ? 4'ha : _GEN_30458; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30460 = 10'h2d7 == _T_442[9:0] ? 4'ha : _GEN_30459; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30461 = 10'h2d8 == _T_442[9:0] ? 4'ha : _GEN_30460; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30462 = 10'h2d9 == _T_442[9:0] ? 4'h7 : _GEN_30461; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30463 = 10'h2da == _T_442[9:0] ? 4'h2 : _GEN_30462; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30464 = 10'h2db == _T_442[9:0] ? 4'h0 : _GEN_30463; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30465 = 10'h2dc == _T_442[9:0] ? 4'h0 : _GEN_30464; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30466 = 10'h2dd == _T_442[9:0] ? 4'h0 : _GEN_30465; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30467 = 10'h2de == _T_442[9:0] ? 4'h0 : _GEN_30466; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30468 = 10'h2df == _T_442[9:0] ? 4'h2 : _GEN_30467; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30469 = 10'h2e0 == _T_442[9:0] ? 4'h0 : _GEN_30468; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30470 = 10'h2e1 == _T_442[9:0] ? 4'h0 : _GEN_30469; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30471 = 10'h2e2 == _T_442[9:0] ? 4'h0 : _GEN_30470; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30472 = 10'h2e3 == _T_442[9:0] ? 4'h0 : _GEN_30471; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30473 = 10'h2e4 == _T_442[9:0] ? 4'h0 : _GEN_30472; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30474 = 10'h2e5 == _T_442[9:0] ? 4'h0 : _GEN_30473; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30475 = 10'h2e6 == _T_442[9:0] ? 4'h2 : _GEN_30474; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30476 = 10'h2e7 == _T_442[9:0] ? 4'h3 : _GEN_30475; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30477 = 10'h2e8 == _T_442[9:0] ? 4'h3 : _GEN_30476; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30478 = 10'h2e9 == _T_442[9:0] ? 4'h3 : _GEN_30477; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30479 = 10'h2ea == _T_442[9:0] ? 4'h3 : _GEN_30478; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30480 = 10'h2eb == _T_442[9:0] ? 4'h3 : _GEN_30479; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30481 = 10'h2ec == _T_442[9:0] ? 4'h4 : _GEN_30480; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30482 = 10'h2ed == _T_442[9:0] ? 4'h5 : _GEN_30481; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30483 = 10'h2ee == _T_442[9:0] ? 4'h6 : _GEN_30482; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30484 = 10'h2ef == _T_442[9:0] ? 4'h8 : _GEN_30483; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30485 = 10'h2f0 == _T_442[9:0] ? 4'h4 : _GEN_30484; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30486 = 10'h2f1 == _T_442[9:0] ? 4'h9 : _GEN_30485; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30487 = 10'h2f2 == _T_442[9:0] ? 4'hb : _GEN_30486; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30488 = 10'h2f3 == _T_442[9:0] ? 4'hb : _GEN_30487; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30489 = 10'h2f4 == _T_442[9:0] ? 4'hb : _GEN_30488; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30490 = 10'h2f5 == _T_442[9:0] ? 4'hb : _GEN_30489; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30491 = 10'h2f6 == _T_442[9:0] ? 4'hb : _GEN_30490; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30492 = 10'h2f7 == _T_442[9:0] ? 4'hb : _GEN_30491; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30493 = 10'h2f8 == _T_442[9:0] ? 4'h8 : _GEN_30492; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30494 = 10'h2f9 == _T_442[9:0] ? 4'h9 : _GEN_30493; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30495 = 10'h2fa == _T_442[9:0] ? 4'hb : _GEN_30494; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30496 = 10'h2fb == _T_442[9:0] ? 4'hb : _GEN_30495; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30497 = 10'h2fc == _T_442[9:0] ? 4'ha : _GEN_30496; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30498 = 10'h2fd == _T_442[9:0] ? 4'ha : _GEN_30497; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30499 = 10'h2fe == _T_442[9:0] ? 4'h9 : _GEN_30498; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30500 = 10'h2ff == _T_442[9:0] ? 4'h8 : _GEN_30499; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30501 = 10'h300 == _T_442[9:0] ? 4'h8 : _GEN_30500; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30502 = 10'h301 == _T_442[9:0] ? 4'h6 : _GEN_30501; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30503 = 10'h302 == _T_442[9:0] ? 4'h1 : _GEN_30502; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30504 = 10'h303 == _T_442[9:0] ? 4'h0 : _GEN_30503; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30505 = 10'h304 == _T_442[9:0] ? 4'h0 : _GEN_30504; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30506 = 10'h305 == _T_442[9:0] ? 4'h0 : _GEN_30505; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30507 = 10'h306 == _T_442[9:0] ? 4'h0 : _GEN_30506; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30508 = 10'h307 == _T_442[9:0] ? 4'h0 : _GEN_30507; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30509 = 10'h308 == _T_442[9:0] ? 4'h0 : _GEN_30508; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30510 = 10'h309 == _T_442[9:0] ? 4'h0 : _GEN_30509; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30511 = 10'h30a == _T_442[9:0] ? 4'h0 : _GEN_30510; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30512 = 10'h30b == _T_442[9:0] ? 4'h0 : _GEN_30511; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30513 = 10'h30c == _T_442[9:0] ? 4'h2 : _GEN_30512; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30514 = 10'h30d == _T_442[9:0] ? 4'h3 : _GEN_30513; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30515 = 10'h30e == _T_442[9:0] ? 4'h3 : _GEN_30514; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30516 = 10'h30f == _T_442[9:0] ? 4'h3 : _GEN_30515; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30517 = 10'h310 == _T_442[9:0] ? 4'h3 : _GEN_30516; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30518 = 10'h311 == _T_442[9:0] ? 4'h3 : _GEN_30517; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30519 = 10'h312 == _T_442[9:0] ? 4'h4 : _GEN_30518; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30520 = 10'h313 == _T_442[9:0] ? 4'h5 : _GEN_30519; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30521 = 10'h314 == _T_442[9:0] ? 4'h5 : _GEN_30520; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30522 = 10'h315 == _T_442[9:0] ? 4'h8 : _GEN_30521; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30523 = 10'h316 == _T_442[9:0] ? 4'h4 : _GEN_30522; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30524 = 10'h317 == _T_442[9:0] ? 4'h6 : _GEN_30523; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30525 = 10'h318 == _T_442[9:0] ? 4'hb : _GEN_30524; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30526 = 10'h319 == _T_442[9:0] ? 4'hb : _GEN_30525; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30527 = 10'h31a == _T_442[9:0] ? 4'hb : _GEN_30526; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30528 = 10'h31b == _T_442[9:0] ? 4'hb : _GEN_30527; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30529 = 10'h31c == _T_442[9:0] ? 4'hb : _GEN_30528; // @[Filter.scala 230:102]
  wire [3:0] _GEN_30530 = 10'h31d == _T_442[9:0] ? 4'hb : _GEN_30529; // @[Filter.scala 230:102]
  wire [6:0] _GEN_39028 = {{3'd0}, _GEN_30530}; // @[Filter.scala 230:102]
  wire [10:0] _T_449 = _GEN_39028 * 7'h46; // @[Filter.scala 230:102]
  wire [10:0] _GEN_39029 = {{2'd0}, _T_444}; // @[Filter.scala 230:69]
  wire [10:0] _T_451 = _GEN_39029 + _T_449; // @[Filter.scala 230:69]
  wire [3:0] _GEN_30553 = 10'h16 == _T_442[9:0] ? 4'hb : 4'hc; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30554 = 10'h17 == _T_442[9:0] ? 4'h8 : _GEN_30553; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30555 = 10'h18 == _T_442[9:0] ? 4'ha : _GEN_30554; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30556 = 10'h19 == _T_442[9:0] ? 4'hc : _GEN_30555; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30557 = 10'h1a == _T_442[9:0] ? 4'hc : _GEN_30556; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30558 = 10'h1b == _T_442[9:0] ? 4'hc : _GEN_30557; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30559 = 10'h1c == _T_442[9:0] ? 4'hc : _GEN_30558; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30560 = 10'h1d == _T_442[9:0] ? 4'hc : _GEN_30559; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30561 = 10'h1e == _T_442[9:0] ? 4'hc : _GEN_30560; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30562 = 10'h1f == _T_442[9:0] ? 4'hc : _GEN_30561; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30563 = 10'h20 == _T_442[9:0] ? 4'hc : _GEN_30562; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30564 = 10'h21 == _T_442[9:0] ? 4'hc : _GEN_30563; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30565 = 10'h22 == _T_442[9:0] ? 4'hc : _GEN_30564; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30566 = 10'h23 == _T_442[9:0] ? 4'hc : _GEN_30565; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30567 = 10'h24 == _T_442[9:0] ? 4'hc : _GEN_30566; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30568 = 10'h25 == _T_442[9:0] ? 4'hc : _GEN_30567; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30569 = 10'h26 == _T_442[9:0] ? 4'hc : _GEN_30568; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30570 = 10'h27 == _T_442[9:0] ? 4'hc : _GEN_30569; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30571 = 10'h28 == _T_442[9:0] ? 4'hc : _GEN_30570; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30572 = 10'h29 == _T_442[9:0] ? 4'hc : _GEN_30571; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30573 = 10'h2a == _T_442[9:0] ? 4'hc : _GEN_30572; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30574 = 10'h2b == _T_442[9:0] ? 4'hc : _GEN_30573; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30575 = 10'h2c == _T_442[9:0] ? 4'hc : _GEN_30574; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30576 = 10'h2d == _T_442[9:0] ? 4'hc : _GEN_30575; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30577 = 10'h2e == _T_442[9:0] ? 4'hc : _GEN_30576; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30578 = 10'h2f == _T_442[9:0] ? 4'hc : _GEN_30577; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30579 = 10'h30 == _T_442[9:0] ? 4'hc : _GEN_30578; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30580 = 10'h31 == _T_442[9:0] ? 4'hc : _GEN_30579; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30581 = 10'h32 == _T_442[9:0] ? 4'hc : _GEN_30580; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30582 = 10'h33 == _T_442[9:0] ? 4'hc : _GEN_30581; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30583 = 10'h34 == _T_442[9:0] ? 4'hc : _GEN_30582; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30584 = 10'h35 == _T_442[9:0] ? 4'hc : _GEN_30583; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30585 = 10'h36 == _T_442[9:0] ? 4'hc : _GEN_30584; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30586 = 10'h37 == _T_442[9:0] ? 4'hc : _GEN_30585; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30587 = 10'h38 == _T_442[9:0] ? 4'hc : _GEN_30586; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30588 = 10'h39 == _T_442[9:0] ? 4'hc : _GEN_30587; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30589 = 10'h3a == _T_442[9:0] ? 4'hc : _GEN_30588; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30590 = 10'h3b == _T_442[9:0] ? 4'hc : _GEN_30589; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30591 = 10'h3c == _T_442[9:0] ? 4'h7 : _GEN_30590; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30592 = 10'h3d == _T_442[9:0] ? 4'h9 : _GEN_30591; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30593 = 10'h3e == _T_442[9:0] ? 4'h8 : _GEN_30592; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30594 = 10'h3f == _T_442[9:0] ? 4'hc : _GEN_30593; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30595 = 10'h40 == _T_442[9:0] ? 4'hc : _GEN_30594; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30596 = 10'h41 == _T_442[9:0] ? 4'hc : _GEN_30595; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30597 = 10'h42 == _T_442[9:0] ? 4'hc : _GEN_30596; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30598 = 10'h43 == _T_442[9:0] ? 4'hc : _GEN_30597; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30599 = 10'h44 == _T_442[9:0] ? 4'hc : _GEN_30598; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30600 = 10'h45 == _T_442[9:0] ? 4'hc : _GEN_30599; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30601 = 10'h46 == _T_442[9:0] ? 4'hc : _GEN_30600; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30602 = 10'h47 == _T_442[9:0] ? 4'hc : _GEN_30601; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30603 = 10'h48 == _T_442[9:0] ? 4'hc : _GEN_30602; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30604 = 10'h49 == _T_442[9:0] ? 4'hc : _GEN_30603; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30605 = 10'h4a == _T_442[9:0] ? 4'hc : _GEN_30604; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30606 = 10'h4b == _T_442[9:0] ? 4'hc : _GEN_30605; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30607 = 10'h4c == _T_442[9:0] ? 4'hc : _GEN_30606; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30608 = 10'h4d == _T_442[9:0] ? 4'hc : _GEN_30607; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30609 = 10'h4e == _T_442[9:0] ? 4'hc : _GEN_30608; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30610 = 10'h4f == _T_442[9:0] ? 4'hc : _GEN_30609; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30611 = 10'h50 == _T_442[9:0] ? 4'hc : _GEN_30610; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30612 = 10'h51 == _T_442[9:0] ? 4'hc : _GEN_30611; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30613 = 10'h52 == _T_442[9:0] ? 4'hc : _GEN_30612; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30614 = 10'h53 == _T_442[9:0] ? 4'hc : _GEN_30613; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30615 = 10'h54 == _T_442[9:0] ? 4'hc : _GEN_30614; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30616 = 10'h55 == _T_442[9:0] ? 4'hc : _GEN_30615; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30617 = 10'h56 == _T_442[9:0] ? 4'hc : _GEN_30616; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30618 = 10'h57 == _T_442[9:0] ? 4'hc : _GEN_30617; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30619 = 10'h58 == _T_442[9:0] ? 4'hc : _GEN_30618; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30620 = 10'h59 == _T_442[9:0] ? 4'hc : _GEN_30619; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30621 = 10'h5a == _T_442[9:0] ? 4'h9 : _GEN_30620; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30622 = 10'h5b == _T_442[9:0] ? 4'ha : _GEN_30621; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30623 = 10'h5c == _T_442[9:0] ? 4'hc : _GEN_30622; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30624 = 10'h5d == _T_442[9:0] ? 4'hc : _GEN_30623; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30625 = 10'h5e == _T_442[9:0] ? 4'hc : _GEN_30624; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30626 = 10'h5f == _T_442[9:0] ? 4'hc : _GEN_30625; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30627 = 10'h60 == _T_442[9:0] ? 4'hc : _GEN_30626; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30628 = 10'h61 == _T_442[9:0] ? 4'hb : _GEN_30627; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30629 = 10'h62 == _T_442[9:0] ? 4'h8 : _GEN_30628; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30630 = 10'h63 == _T_442[9:0] ? 4'h9 : _GEN_30629; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30631 = 10'h64 == _T_442[9:0] ? 4'h7 : _GEN_30630; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30632 = 10'h65 == _T_442[9:0] ? 4'hb : _GEN_30631; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30633 = 10'h66 == _T_442[9:0] ? 4'hc : _GEN_30632; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30634 = 10'h67 == _T_442[9:0] ? 4'hc : _GEN_30633; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30635 = 10'h68 == _T_442[9:0] ? 4'hc : _GEN_30634; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30636 = 10'h69 == _T_442[9:0] ? 4'hc : _GEN_30635; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30637 = 10'h6a == _T_442[9:0] ? 4'hc : _GEN_30636; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30638 = 10'h6b == _T_442[9:0] ? 4'hb : _GEN_30637; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30639 = 10'h6c == _T_442[9:0] ? 4'h9 : _GEN_30638; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30640 = 10'h6d == _T_442[9:0] ? 4'ha : _GEN_30639; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30641 = 10'h6e == _T_442[9:0] ? 4'hc : _GEN_30640; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30642 = 10'h6f == _T_442[9:0] ? 4'hc : _GEN_30641; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30643 = 10'h70 == _T_442[9:0] ? 4'hc : _GEN_30642; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30644 = 10'h71 == _T_442[9:0] ? 4'hc : _GEN_30643; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30645 = 10'h72 == _T_442[9:0] ? 4'hc : _GEN_30644; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30646 = 10'h73 == _T_442[9:0] ? 4'hc : _GEN_30645; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30647 = 10'h74 == _T_442[9:0] ? 4'hc : _GEN_30646; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30648 = 10'h75 == _T_442[9:0] ? 4'hc : _GEN_30647; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30649 = 10'h76 == _T_442[9:0] ? 4'hc : _GEN_30648; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30650 = 10'h77 == _T_442[9:0] ? 4'hc : _GEN_30649; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30651 = 10'h78 == _T_442[9:0] ? 4'hc : _GEN_30650; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30652 = 10'h79 == _T_442[9:0] ? 4'hc : _GEN_30651; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30653 = 10'h7a == _T_442[9:0] ? 4'hc : _GEN_30652; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30654 = 10'h7b == _T_442[9:0] ? 4'hc : _GEN_30653; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30655 = 10'h7c == _T_442[9:0] ? 4'hc : _GEN_30654; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30656 = 10'h7d == _T_442[9:0] ? 4'hc : _GEN_30655; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30657 = 10'h7e == _T_442[9:0] ? 4'hc : _GEN_30656; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30658 = 10'h7f == _T_442[9:0] ? 4'hc : _GEN_30657; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30659 = 10'h80 == _T_442[9:0] ? 4'hc : _GEN_30658; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30660 = 10'h81 == _T_442[9:0] ? 4'h9 : _GEN_30659; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30661 = 10'h82 == _T_442[9:0] ? 4'h9 : _GEN_30660; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30662 = 10'h83 == _T_442[9:0] ? 4'h9 : _GEN_30661; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30663 = 10'h84 == _T_442[9:0] ? 4'hc : _GEN_30662; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30664 = 10'h85 == _T_442[9:0] ? 4'hc : _GEN_30663; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30665 = 10'h86 == _T_442[9:0] ? 4'hc : _GEN_30664; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30666 = 10'h87 == _T_442[9:0] ? 4'h8 : _GEN_30665; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30667 = 10'h88 == _T_442[9:0] ? 4'h9 : _GEN_30666; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30668 = 10'h89 == _T_442[9:0] ? 4'h9 : _GEN_30667; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30669 = 10'h8a == _T_442[9:0] ? 4'h9 : _GEN_30668; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30670 = 10'h8b == _T_442[9:0] ? 4'hc : _GEN_30669; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30671 = 10'h8c == _T_442[9:0] ? 4'hc : _GEN_30670; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30672 = 10'h8d == _T_442[9:0] ? 4'hc : _GEN_30671; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30673 = 10'h8e == _T_442[9:0] ? 4'hc : _GEN_30672; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30674 = 10'h8f == _T_442[9:0] ? 4'h9 : _GEN_30673; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30675 = 10'h90 == _T_442[9:0] ? 4'h9 : _GEN_30674; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30676 = 10'h91 == _T_442[9:0] ? 4'h9 : _GEN_30675; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30677 = 10'h92 == _T_442[9:0] ? 4'ha : _GEN_30676; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30678 = 10'h93 == _T_442[9:0] ? 4'hc : _GEN_30677; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30679 = 10'h94 == _T_442[9:0] ? 4'hc : _GEN_30678; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30680 = 10'h95 == _T_442[9:0] ? 4'hc : _GEN_30679; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30681 = 10'h96 == _T_442[9:0] ? 4'hc : _GEN_30680; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30682 = 10'h97 == _T_442[9:0] ? 4'hc : _GEN_30681; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30683 = 10'h98 == _T_442[9:0] ? 4'hc : _GEN_30682; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30684 = 10'h99 == _T_442[9:0] ? 4'hc : _GEN_30683; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30685 = 10'h9a == _T_442[9:0] ? 4'hc : _GEN_30684; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30686 = 10'h9b == _T_442[9:0] ? 4'hc : _GEN_30685; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30687 = 10'h9c == _T_442[9:0] ? 4'hc : _GEN_30686; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30688 = 10'h9d == _T_442[9:0] ? 4'hc : _GEN_30687; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30689 = 10'h9e == _T_442[9:0] ? 4'hc : _GEN_30688; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30690 = 10'h9f == _T_442[9:0] ? 4'hc : _GEN_30689; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30691 = 10'ha0 == _T_442[9:0] ? 4'hc : _GEN_30690; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30692 = 10'ha1 == _T_442[9:0] ? 4'hc : _GEN_30691; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30693 = 10'ha2 == _T_442[9:0] ? 4'hc : _GEN_30692; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30694 = 10'ha3 == _T_442[9:0] ? 4'hc : _GEN_30693; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30695 = 10'ha4 == _T_442[9:0] ? 4'hc : _GEN_30694; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30696 = 10'ha5 == _T_442[9:0] ? 4'hc : _GEN_30695; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30697 = 10'ha6 == _T_442[9:0] ? 4'hc : _GEN_30696; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30698 = 10'ha7 == _T_442[9:0] ? 4'hc : _GEN_30697; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30699 = 10'ha8 == _T_442[9:0] ? 4'h9 : _GEN_30698; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30700 = 10'ha9 == _T_442[9:0] ? 4'h8 : _GEN_30699; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30701 = 10'haa == _T_442[9:0] ? 4'h8 : _GEN_30700; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30702 = 10'hab == _T_442[9:0] ? 4'ha : _GEN_30701; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30703 = 10'hac == _T_442[9:0] ? 4'hb : _GEN_30702; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30704 = 10'had == _T_442[9:0] ? 4'h7 : _GEN_30703; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30705 = 10'hae == _T_442[9:0] ? 4'h9 : _GEN_30704; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30706 = 10'haf == _T_442[9:0] ? 4'h9 : _GEN_30705; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30707 = 10'hb0 == _T_442[9:0] ? 4'h8 : _GEN_30706; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30708 = 10'hb1 == _T_442[9:0] ? 4'h9 : _GEN_30707; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30709 = 10'hb2 == _T_442[9:0] ? 4'hc : _GEN_30708; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30710 = 10'hb3 == _T_442[9:0] ? 4'h9 : _GEN_30709; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30711 = 10'hb4 == _T_442[9:0] ? 4'h9 : _GEN_30710; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30712 = 10'hb5 == _T_442[9:0] ? 4'h9 : _GEN_30711; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30713 = 10'hb6 == _T_442[9:0] ? 4'h9 : _GEN_30712; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30714 = 10'hb7 == _T_442[9:0] ? 4'ha : _GEN_30713; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30715 = 10'hb8 == _T_442[9:0] ? 4'hc : _GEN_30714; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30716 = 10'hb9 == _T_442[9:0] ? 4'hc : _GEN_30715; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30717 = 10'hba == _T_442[9:0] ? 4'hc : _GEN_30716; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30718 = 10'hbb == _T_442[9:0] ? 4'hc : _GEN_30717; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30719 = 10'hbc == _T_442[9:0] ? 4'hc : _GEN_30718; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30720 = 10'hbd == _T_442[9:0] ? 4'hb : _GEN_30719; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30721 = 10'hbe == _T_442[9:0] ? 4'hc : _GEN_30720; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30722 = 10'hbf == _T_442[9:0] ? 4'hc : _GEN_30721; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30723 = 10'hc0 == _T_442[9:0] ? 4'hc : _GEN_30722; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30724 = 10'hc1 == _T_442[9:0] ? 4'hc : _GEN_30723; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30725 = 10'hc2 == _T_442[9:0] ? 4'hc : _GEN_30724; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30726 = 10'hc3 == _T_442[9:0] ? 4'hc : _GEN_30725; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30727 = 10'hc4 == _T_442[9:0] ? 4'hc : _GEN_30726; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30728 = 10'hc5 == _T_442[9:0] ? 4'hc : _GEN_30727; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30729 = 10'hc6 == _T_442[9:0] ? 4'hb : _GEN_30728; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30730 = 10'hc7 == _T_442[9:0] ? 4'hb : _GEN_30729; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30731 = 10'hc8 == _T_442[9:0] ? 4'ha : _GEN_30730; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30732 = 10'hc9 == _T_442[9:0] ? 4'ha : _GEN_30731; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30733 = 10'hca == _T_442[9:0] ? 4'hb : _GEN_30732; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30734 = 10'hcb == _T_442[9:0] ? 4'hc : _GEN_30733; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30735 = 10'hcc == _T_442[9:0] ? 4'hc : _GEN_30734; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30736 = 10'hcd == _T_442[9:0] ? 4'hc : _GEN_30735; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30737 = 10'hce == _T_442[9:0] ? 4'ha : _GEN_30736; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30738 = 10'hcf == _T_442[9:0] ? 4'h8 : _GEN_30737; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30739 = 10'hd0 == _T_442[9:0] ? 4'h9 : _GEN_30738; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30740 = 10'hd1 == _T_442[9:0] ? 4'h8 : _GEN_30739; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30741 = 10'hd2 == _T_442[9:0] ? 4'h9 : _GEN_30740; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30742 = 10'hd3 == _T_442[9:0] ? 4'h9 : _GEN_30741; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30743 = 10'hd4 == _T_442[9:0] ? 4'h9 : _GEN_30742; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30744 = 10'hd5 == _T_442[9:0] ? 4'h9 : _GEN_30743; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30745 = 10'hd6 == _T_442[9:0] ? 4'ha : _GEN_30744; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30746 = 10'hd7 == _T_442[9:0] ? 4'h9 : _GEN_30745; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30747 = 10'hd8 == _T_442[9:0] ? 4'h9 : _GEN_30746; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30748 = 10'hd9 == _T_442[9:0] ? 4'h9 : _GEN_30747; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30749 = 10'hda == _T_442[9:0] ? 4'ha : _GEN_30748; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30750 = 10'hdb == _T_442[9:0] ? 4'h9 : _GEN_30749; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30751 = 10'hdc == _T_442[9:0] ? 4'h7 : _GEN_30750; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30752 = 10'hdd == _T_442[9:0] ? 4'hc : _GEN_30751; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30753 = 10'hde == _T_442[9:0] ? 4'hc : _GEN_30752; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30754 = 10'hdf == _T_442[9:0] ? 4'hc : _GEN_30753; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30755 = 10'he0 == _T_442[9:0] ? 4'hc : _GEN_30754; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30756 = 10'he1 == _T_442[9:0] ? 4'hc : _GEN_30755; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30757 = 10'he2 == _T_442[9:0] ? 4'hc : _GEN_30756; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30758 = 10'he3 == _T_442[9:0] ? 4'h8 : _GEN_30757; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30759 = 10'he4 == _T_442[9:0] ? 4'hc : _GEN_30758; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30760 = 10'he5 == _T_442[9:0] ? 4'hc : _GEN_30759; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30761 = 10'he6 == _T_442[9:0] ? 4'hc : _GEN_30760; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30762 = 10'he7 == _T_442[9:0] ? 4'hc : _GEN_30761; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30763 = 10'he8 == _T_442[9:0] ? 4'hc : _GEN_30762; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30764 = 10'he9 == _T_442[9:0] ? 4'hc : _GEN_30763; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30765 = 10'hea == _T_442[9:0] ? 4'hc : _GEN_30764; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30766 = 10'heb == _T_442[9:0] ? 4'ha : _GEN_30765; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30767 = 10'hec == _T_442[9:0] ? 4'h7 : _GEN_30766; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30768 = 10'hed == _T_442[9:0] ? 4'h3 : _GEN_30767; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30769 = 10'hee == _T_442[9:0] ? 4'h3 : _GEN_30768; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30770 = 10'hef == _T_442[9:0] ? 4'h3 : _GEN_30769; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30771 = 10'hf0 == _T_442[9:0] ? 4'h3 : _GEN_30770; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30772 = 10'hf1 == _T_442[9:0] ? 4'h8 : _GEN_30771; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30773 = 10'hf2 == _T_442[9:0] ? 4'hc : _GEN_30772; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30774 = 10'hf3 == _T_442[9:0] ? 4'hc : _GEN_30773; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30775 = 10'hf4 == _T_442[9:0] ? 4'hc : _GEN_30774; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30776 = 10'hf5 == _T_442[9:0] ? 4'h9 : _GEN_30775; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30777 = 10'hf6 == _T_442[9:0] ? 4'h9 : _GEN_30776; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30778 = 10'hf7 == _T_442[9:0] ? 4'h9 : _GEN_30777; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30779 = 10'hf8 == _T_442[9:0] ? 4'h9 : _GEN_30778; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30780 = 10'hf9 == _T_442[9:0] ? 4'ha : _GEN_30779; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30781 = 10'hfa == _T_442[9:0] ? 4'h9 : _GEN_30780; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30782 = 10'hfb == _T_442[9:0] ? 4'h9 : _GEN_30781; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30783 = 10'hfc == _T_442[9:0] ? 4'h9 : _GEN_30782; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30784 = 10'hfd == _T_442[9:0] ? 4'h9 : _GEN_30783; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30785 = 10'hfe == _T_442[9:0] ? 4'h9 : _GEN_30784; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30786 = 10'hff == _T_442[9:0] ? 4'ha : _GEN_30785; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30787 = 10'h100 == _T_442[9:0] ? 4'ha : _GEN_30786; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30788 = 10'h101 == _T_442[9:0] ? 4'h7 : _GEN_30787; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30789 = 10'h102 == _T_442[9:0] ? 4'h9 : _GEN_30788; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30790 = 10'h103 == _T_442[9:0] ? 4'hc : _GEN_30789; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30791 = 10'h104 == _T_442[9:0] ? 4'hc : _GEN_30790; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30792 = 10'h105 == _T_442[9:0] ? 4'hb : _GEN_30791; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30793 = 10'h106 == _T_442[9:0] ? 4'hb : _GEN_30792; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30794 = 10'h107 == _T_442[9:0] ? 4'hb : _GEN_30793; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30795 = 10'h108 == _T_442[9:0] ? 4'hb : _GEN_30794; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30796 = 10'h109 == _T_442[9:0] ? 4'h7 : _GEN_30795; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30797 = 10'h10a == _T_442[9:0] ? 4'hc : _GEN_30796; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30798 = 10'h10b == _T_442[9:0] ? 4'hc : _GEN_30797; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30799 = 10'h10c == _T_442[9:0] ? 4'hc : _GEN_30798; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30800 = 10'h10d == _T_442[9:0] ? 4'hc : _GEN_30799; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30801 = 10'h10e == _T_442[9:0] ? 4'hc : _GEN_30800; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30802 = 10'h10f == _T_442[9:0] ? 4'h9 : _GEN_30801; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30803 = 10'h110 == _T_442[9:0] ? 4'hb : _GEN_30802; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30804 = 10'h111 == _T_442[9:0] ? 4'h4 : _GEN_30803; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30805 = 10'h112 == _T_442[9:0] ? 4'h7 : _GEN_30804; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30806 = 10'h113 == _T_442[9:0] ? 4'h3 : _GEN_30805; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30807 = 10'h114 == _T_442[9:0] ? 4'h3 : _GEN_30806; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30808 = 10'h115 == _T_442[9:0] ? 4'h3 : _GEN_30807; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30809 = 10'h116 == _T_442[9:0] ? 4'h3 : _GEN_30808; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30810 = 10'h117 == _T_442[9:0] ? 4'h2 : _GEN_30809; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30811 = 10'h118 == _T_442[9:0] ? 4'h9 : _GEN_30810; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30812 = 10'h119 == _T_442[9:0] ? 4'hc : _GEN_30811; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30813 = 10'h11a == _T_442[9:0] ? 4'hc : _GEN_30812; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30814 = 10'h11b == _T_442[9:0] ? 4'hc : _GEN_30813; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30815 = 10'h11c == _T_442[9:0] ? 4'h9 : _GEN_30814; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30816 = 10'h11d == _T_442[9:0] ? 4'h9 : _GEN_30815; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30817 = 10'h11e == _T_442[9:0] ? 4'h9 : _GEN_30816; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30818 = 10'h11f == _T_442[9:0] ? 4'h8 : _GEN_30817; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30819 = 10'h120 == _T_442[9:0] ? 4'h7 : _GEN_30818; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30820 = 10'h121 == _T_442[9:0] ? 4'h9 : _GEN_30819; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30821 = 10'h122 == _T_442[9:0] ? 4'h7 : _GEN_30820; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30822 = 10'h123 == _T_442[9:0] ? 4'h7 : _GEN_30821; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30823 = 10'h124 == _T_442[9:0] ? 4'h9 : _GEN_30822; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30824 = 10'h125 == _T_442[9:0] ? 4'h9 : _GEN_30823; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30825 = 10'h126 == _T_442[9:0] ? 4'h8 : _GEN_30824; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30826 = 10'h127 == _T_442[9:0] ? 4'h9 : _GEN_30825; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30827 = 10'h128 == _T_442[9:0] ? 4'h8 : _GEN_30826; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30828 = 10'h129 == _T_442[9:0] ? 4'ha : _GEN_30827; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30829 = 10'h12a == _T_442[9:0] ? 4'h5 : _GEN_30828; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30830 = 10'h12b == _T_442[9:0] ? 4'h3 : _GEN_30829; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30831 = 10'h12c == _T_442[9:0] ? 4'h3 : _GEN_30830; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30832 = 10'h12d == _T_442[9:0] ? 4'h3 : _GEN_30831; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30833 = 10'h12e == _T_442[9:0] ? 4'h5 : _GEN_30832; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30834 = 10'h12f == _T_442[9:0] ? 4'h8 : _GEN_30833; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30835 = 10'h130 == _T_442[9:0] ? 4'hc : _GEN_30834; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30836 = 10'h131 == _T_442[9:0] ? 4'hb : _GEN_30835; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30837 = 10'h132 == _T_442[9:0] ? 4'h9 : _GEN_30836; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30838 = 10'h133 == _T_442[9:0] ? 4'h8 : _GEN_30837; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30839 = 10'h134 == _T_442[9:0] ? 4'h9 : _GEN_30838; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30840 = 10'h135 == _T_442[9:0] ? 4'h7 : _GEN_30839; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30841 = 10'h136 == _T_442[9:0] ? 4'h7 : _GEN_30840; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30842 = 10'h137 == _T_442[9:0] ? 4'h5 : _GEN_30841; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30843 = 10'h138 == _T_442[9:0] ? 4'h7 : _GEN_30842; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30844 = 10'h139 == _T_442[9:0] ? 4'h3 : _GEN_30843; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30845 = 10'h13a == _T_442[9:0] ? 4'h3 : _GEN_30844; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30846 = 10'h13b == _T_442[9:0] ? 4'h3 : _GEN_30845; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30847 = 10'h13c == _T_442[9:0] ? 4'h3 : _GEN_30846; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30848 = 10'h13d == _T_442[9:0] ? 4'h3 : _GEN_30847; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30849 = 10'h13e == _T_442[9:0] ? 4'h5 : _GEN_30848; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30850 = 10'h13f == _T_442[9:0] ? 4'ha : _GEN_30849; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30851 = 10'h140 == _T_442[9:0] ? 4'hc : _GEN_30850; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30852 = 10'h141 == _T_442[9:0] ? 4'hc : _GEN_30851; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30853 = 10'h142 == _T_442[9:0] ? 4'hc : _GEN_30852; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30854 = 10'h143 == _T_442[9:0] ? 4'h9 : _GEN_30853; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30855 = 10'h144 == _T_442[9:0] ? 4'h9 : _GEN_30854; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30856 = 10'h145 == _T_442[9:0] ? 4'h8 : _GEN_30855; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30857 = 10'h146 == _T_442[9:0] ? 4'h8 : _GEN_30856; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30858 = 10'h147 == _T_442[9:0] ? 4'h7 : _GEN_30857; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30859 = 10'h148 == _T_442[9:0] ? 4'h8 : _GEN_30858; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30860 = 10'h149 == _T_442[9:0] ? 4'h9 : _GEN_30859; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30861 = 10'h14a == _T_442[9:0] ? 4'ha : _GEN_30860; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30862 = 10'h14b == _T_442[9:0] ? 4'h9 : _GEN_30861; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30863 = 10'h14c == _T_442[9:0] ? 4'ha : _GEN_30862; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30864 = 10'h14d == _T_442[9:0] ? 4'h9 : _GEN_30863; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30865 = 10'h14e == _T_442[9:0] ? 4'h7 : _GEN_30864; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30866 = 10'h14f == _T_442[9:0] ? 4'h3 : _GEN_30865; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30867 = 10'h150 == _T_442[9:0] ? 4'h3 : _GEN_30866; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30868 = 10'h151 == _T_442[9:0] ? 4'h3 : _GEN_30867; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30869 = 10'h152 == _T_442[9:0] ? 4'h3 : _GEN_30868; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30870 = 10'h153 == _T_442[9:0] ? 4'h3 : _GEN_30869; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30871 = 10'h154 == _T_442[9:0] ? 4'h3 : _GEN_30870; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30872 = 10'h155 == _T_442[9:0] ? 4'h8 : _GEN_30871; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30873 = 10'h156 == _T_442[9:0] ? 4'ha : _GEN_30872; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30874 = 10'h157 == _T_442[9:0] ? 4'h7 : _GEN_30873; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30875 = 10'h158 == _T_442[9:0] ? 4'h7 : _GEN_30874; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30876 = 10'h159 == _T_442[9:0] ? 4'h7 : _GEN_30875; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30877 = 10'h15a == _T_442[9:0] ? 4'h7 : _GEN_30876; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30878 = 10'h15b == _T_442[9:0] ? 4'h7 : _GEN_30877; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30879 = 10'h15c == _T_442[9:0] ? 4'h7 : _GEN_30878; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30880 = 10'h15d == _T_442[9:0] ? 4'h7 : _GEN_30879; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30881 = 10'h15e == _T_442[9:0] ? 4'h7 : _GEN_30880; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30882 = 10'h15f == _T_442[9:0] ? 4'h3 : _GEN_30881; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30883 = 10'h160 == _T_442[9:0] ? 4'h3 : _GEN_30882; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30884 = 10'h161 == _T_442[9:0] ? 4'h3 : _GEN_30883; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30885 = 10'h162 == _T_442[9:0] ? 4'h3 : _GEN_30884; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30886 = 10'h163 == _T_442[9:0] ? 4'h3 : _GEN_30885; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30887 = 10'h164 == _T_442[9:0] ? 4'h4 : _GEN_30886; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30888 = 10'h165 == _T_442[9:0] ? 4'ha : _GEN_30887; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30889 = 10'h166 == _T_442[9:0] ? 4'ha : _GEN_30888; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30890 = 10'h167 == _T_442[9:0] ? 4'hc : _GEN_30889; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30891 = 10'h168 == _T_442[9:0] ? 4'hc : _GEN_30890; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30892 = 10'h169 == _T_442[9:0] ? 4'h9 : _GEN_30891; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30893 = 10'h16a == _T_442[9:0] ? 4'h9 : _GEN_30892; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30894 = 10'h16b == _T_442[9:0] ? 4'ha : _GEN_30893; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30895 = 10'h16c == _T_442[9:0] ? 4'h7 : _GEN_30894; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30896 = 10'h16d == _T_442[9:0] ? 4'h7 : _GEN_30895; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30897 = 10'h16e == _T_442[9:0] ? 4'h7 : _GEN_30896; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30898 = 10'h16f == _T_442[9:0] ? 4'ha : _GEN_30897; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30899 = 10'h170 == _T_442[9:0] ? 4'ha : _GEN_30898; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30900 = 10'h171 == _T_442[9:0] ? 4'ha : _GEN_30899; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30901 = 10'h172 == _T_442[9:0] ? 4'hc : _GEN_30900; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30902 = 10'h173 == _T_442[9:0] ? 4'h8 : _GEN_30901; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30903 = 10'h174 == _T_442[9:0] ? 4'h5 : _GEN_30902; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30904 = 10'h175 == _T_442[9:0] ? 4'h8 : _GEN_30903; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30905 = 10'h176 == _T_442[9:0] ? 4'h7 : _GEN_30904; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30906 = 10'h177 == _T_442[9:0] ? 4'h8 : _GEN_30905; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30907 = 10'h178 == _T_442[9:0] ? 4'h7 : _GEN_30906; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30908 = 10'h179 == _T_442[9:0] ? 4'h5 : _GEN_30907; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30909 = 10'h17a == _T_442[9:0] ? 4'h5 : _GEN_30908; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30910 = 10'h17b == _T_442[9:0] ? 4'h7 : _GEN_30909; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30911 = 10'h17c == _T_442[9:0] ? 4'h7 : _GEN_30910; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30912 = 10'h17d == _T_442[9:0] ? 4'h7 : _GEN_30911; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30913 = 10'h17e == _T_442[9:0] ? 4'h7 : _GEN_30912; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30914 = 10'h17f == _T_442[9:0] ? 4'h7 : _GEN_30913; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30915 = 10'h180 == _T_442[9:0] ? 4'h7 : _GEN_30914; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30916 = 10'h181 == _T_442[9:0] ? 4'h7 : _GEN_30915; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30917 = 10'h182 == _T_442[9:0] ? 4'h7 : _GEN_30916; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30918 = 10'h183 == _T_442[9:0] ? 4'h7 : _GEN_30917; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30919 = 10'h184 == _T_442[9:0] ? 4'h7 : _GEN_30918; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30920 = 10'h185 == _T_442[9:0] ? 4'h5 : _GEN_30919; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30921 = 10'h186 == _T_442[9:0] ? 4'h3 : _GEN_30920; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30922 = 10'h187 == _T_442[9:0] ? 4'h3 : _GEN_30921; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30923 = 10'h188 == _T_442[9:0] ? 4'h3 : _GEN_30922; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30924 = 10'h189 == _T_442[9:0] ? 4'h4 : _GEN_30923; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30925 = 10'h18a == _T_442[9:0] ? 4'h5 : _GEN_30924; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30926 = 10'h18b == _T_442[9:0] ? 4'ha : _GEN_30925; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30927 = 10'h18c == _T_442[9:0] ? 4'ha : _GEN_30926; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30928 = 10'h18d == _T_442[9:0] ? 4'ha : _GEN_30927; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30929 = 10'h18e == _T_442[9:0] ? 4'hc : _GEN_30928; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30930 = 10'h18f == _T_442[9:0] ? 4'h8 : _GEN_30929; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30931 = 10'h190 == _T_442[9:0] ? 4'h9 : _GEN_30930; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30932 = 10'h191 == _T_442[9:0] ? 4'h8 : _GEN_30931; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30933 = 10'h192 == _T_442[9:0] ? 4'h7 : _GEN_30932; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30934 = 10'h193 == _T_442[9:0] ? 4'h7 : _GEN_30933; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30935 = 10'h194 == _T_442[9:0] ? 4'h7 : _GEN_30934; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30936 = 10'h195 == _T_442[9:0] ? 4'h9 : _GEN_30935; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30937 = 10'h196 == _T_442[9:0] ? 4'ha : _GEN_30936; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30938 = 10'h197 == _T_442[9:0] ? 4'h8 : _GEN_30937; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30939 = 10'h198 == _T_442[9:0] ? 4'hc : _GEN_30938; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30940 = 10'h199 == _T_442[9:0] ? 4'h5 : _GEN_30939; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30941 = 10'h19a == _T_442[9:0] ? 4'h1 : _GEN_30940; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30942 = 10'h19b == _T_442[9:0] ? 4'h4 : _GEN_30941; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30943 = 10'h19c == _T_442[9:0] ? 4'h7 : _GEN_30942; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30944 = 10'h19d == _T_442[9:0] ? 4'h5 : _GEN_30943; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30945 = 10'h19e == _T_442[9:0] ? 4'h2 : _GEN_30944; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30946 = 10'h19f == _T_442[9:0] ? 4'h3 : _GEN_30945; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30947 = 10'h1a0 == _T_442[9:0] ? 4'h7 : _GEN_30946; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30948 = 10'h1a1 == _T_442[9:0] ? 4'h7 : _GEN_30947; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30949 = 10'h1a2 == _T_442[9:0] ? 4'h7 : _GEN_30948; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30950 = 10'h1a3 == _T_442[9:0] ? 4'h7 : _GEN_30949; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30951 = 10'h1a4 == _T_442[9:0] ? 4'h7 : _GEN_30950; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30952 = 10'h1a5 == _T_442[9:0] ? 4'h7 : _GEN_30951; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30953 = 10'h1a6 == _T_442[9:0] ? 4'h7 : _GEN_30952; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30954 = 10'h1a7 == _T_442[9:0] ? 4'h7 : _GEN_30953; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30955 = 10'h1a8 == _T_442[9:0] ? 4'h8 : _GEN_30954; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30956 = 10'h1a9 == _T_442[9:0] ? 4'h8 : _GEN_30955; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30957 = 10'h1aa == _T_442[9:0] ? 4'h6 : _GEN_30956; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30958 = 10'h1ab == _T_442[9:0] ? 4'h6 : _GEN_30957; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30959 = 10'h1ac == _T_442[9:0] ? 4'h5 : _GEN_30958; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30960 = 10'h1ad == _T_442[9:0] ? 4'h4 : _GEN_30959; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30961 = 10'h1ae == _T_442[9:0] ? 4'h3 : _GEN_30960; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30962 = 10'h1af == _T_442[9:0] ? 4'h6 : _GEN_30961; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30963 = 10'h1b0 == _T_442[9:0] ? 4'h6 : _GEN_30962; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30964 = 10'h1b1 == _T_442[9:0] ? 4'ha : _GEN_30963; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30965 = 10'h1b2 == _T_442[9:0] ? 4'ha : _GEN_30964; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30966 = 10'h1b3 == _T_442[9:0] ? 4'h9 : _GEN_30965; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30967 = 10'h1b4 == _T_442[9:0] ? 4'hb : _GEN_30966; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30968 = 10'h1b5 == _T_442[9:0] ? 4'h8 : _GEN_30967; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30969 = 10'h1b6 == _T_442[9:0] ? 4'h8 : _GEN_30968; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30970 = 10'h1b7 == _T_442[9:0] ? 4'h7 : _GEN_30969; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30971 = 10'h1b8 == _T_442[9:0] ? 4'h6 : _GEN_30970; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30972 = 10'h1b9 == _T_442[9:0] ? 4'h7 : _GEN_30971; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30973 = 10'h1ba == _T_442[9:0] ? 4'h6 : _GEN_30972; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30974 = 10'h1bb == _T_442[9:0] ? 4'h8 : _GEN_30973; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30975 = 10'h1bc == _T_442[9:0] ? 4'ha : _GEN_30974; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30976 = 10'h1bd == _T_442[9:0] ? 4'h9 : _GEN_30975; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30977 = 10'h1be == _T_442[9:0] ? 4'hc : _GEN_30976; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30978 = 10'h1bf == _T_442[9:0] ? 4'h7 : _GEN_30977; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30979 = 10'h1c0 == _T_442[9:0] ? 4'h6 : _GEN_30978; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30980 = 10'h1c1 == _T_442[9:0] ? 4'h7 : _GEN_30979; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30981 = 10'h1c2 == _T_442[9:0] ? 4'h7 : _GEN_30980; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30982 = 10'h1c3 == _T_442[9:0] ? 4'h6 : _GEN_30981; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30983 = 10'h1c4 == _T_442[9:0] ? 4'h5 : _GEN_30982; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30984 = 10'h1c5 == _T_442[9:0] ? 4'h6 : _GEN_30983; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30985 = 10'h1c6 == _T_442[9:0] ? 4'h8 : _GEN_30984; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30986 = 10'h1c7 == _T_442[9:0] ? 4'h7 : _GEN_30985; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30987 = 10'h1c8 == _T_442[9:0] ? 4'h7 : _GEN_30986; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30988 = 10'h1c9 == _T_442[9:0] ? 4'h7 : _GEN_30987; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30989 = 10'h1ca == _T_442[9:0] ? 4'h7 : _GEN_30988; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30990 = 10'h1cb == _T_442[9:0] ? 4'h7 : _GEN_30989; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30991 = 10'h1cc == _T_442[9:0] ? 4'h7 : _GEN_30990; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30992 = 10'h1cd == _T_442[9:0] ? 4'h8 : _GEN_30991; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30993 = 10'h1ce == _T_442[9:0] ? 4'h8 : _GEN_30992; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30994 = 10'h1cf == _T_442[9:0] ? 4'h8 : _GEN_30993; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30995 = 10'h1d0 == _T_442[9:0] ? 4'h5 : _GEN_30994; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30996 = 10'h1d1 == _T_442[9:0] ? 4'h6 : _GEN_30995; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30997 = 10'h1d2 == _T_442[9:0] ? 4'h7 : _GEN_30996; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30998 = 10'h1d3 == _T_442[9:0] ? 4'h7 : _GEN_30997; // @[Filter.scala 230:142]
  wire [3:0] _GEN_30999 = 10'h1d4 == _T_442[9:0] ? 4'h7 : _GEN_30998; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31000 = 10'h1d5 == _T_442[9:0] ? 4'h6 : _GEN_30999; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31001 = 10'h1d6 == _T_442[9:0] ? 4'h8 : _GEN_31000; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31002 = 10'h1d7 == _T_442[9:0] ? 4'ha : _GEN_31001; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31003 = 10'h1d8 == _T_442[9:0] ? 4'ha : _GEN_31002; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31004 = 10'h1d9 == _T_442[9:0] ? 4'ha : _GEN_31003; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31005 = 10'h1da == _T_442[9:0] ? 4'h8 : _GEN_31004; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31006 = 10'h1db == _T_442[9:0] ? 4'h9 : _GEN_31005; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31007 = 10'h1dc == _T_442[9:0] ? 4'h9 : _GEN_31006; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31008 = 10'h1dd == _T_442[9:0] ? 4'h5 : _GEN_31007; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31009 = 10'h1de == _T_442[9:0] ? 4'h7 : _GEN_31008; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31010 = 10'h1df == _T_442[9:0] ? 4'h7 : _GEN_31009; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31011 = 10'h1e0 == _T_442[9:0] ? 4'h7 : _GEN_31010; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31012 = 10'h1e1 == _T_442[9:0] ? 4'h6 : _GEN_31011; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31013 = 10'h1e2 == _T_442[9:0] ? 4'h9 : _GEN_31012; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31014 = 10'h1e3 == _T_442[9:0] ? 4'h9 : _GEN_31013; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31015 = 10'h1e4 == _T_442[9:0] ? 4'hb : _GEN_31014; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31016 = 10'h1e5 == _T_442[9:0] ? 4'h8 : _GEN_31015; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31017 = 10'h1e6 == _T_442[9:0] ? 4'h7 : _GEN_31016; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31018 = 10'h1e7 == _T_442[9:0] ? 4'h8 : _GEN_31017; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31019 = 10'h1e8 == _T_442[9:0] ? 4'h8 : _GEN_31018; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31020 = 10'h1e9 == _T_442[9:0] ? 4'h8 : _GEN_31019; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31021 = 10'h1ea == _T_442[9:0] ? 4'h8 : _GEN_31020; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31022 = 10'h1eb == _T_442[9:0] ? 4'h8 : _GEN_31021; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31023 = 10'h1ec == _T_442[9:0] ? 4'h8 : _GEN_31022; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31024 = 10'h1ed == _T_442[9:0] ? 4'h6 : _GEN_31023; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31025 = 10'h1ee == _T_442[9:0] ? 4'h7 : _GEN_31024; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31026 = 10'h1ef == _T_442[9:0] ? 4'h7 : _GEN_31025; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31027 = 10'h1f0 == _T_442[9:0] ? 4'h7 : _GEN_31026; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31028 = 10'h1f1 == _T_442[9:0] ? 4'h7 : _GEN_31027; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31029 = 10'h1f2 == _T_442[9:0] ? 4'h7 : _GEN_31028; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31030 = 10'h1f3 == _T_442[9:0] ? 4'h8 : _GEN_31029; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31031 = 10'h1f4 == _T_442[9:0] ? 4'h8 : _GEN_31030; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31032 = 10'h1f5 == _T_442[9:0] ? 4'h8 : _GEN_31031; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31033 = 10'h1f6 == _T_442[9:0] ? 4'ha : _GEN_31032; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31034 = 10'h1f7 == _T_442[9:0] ? 4'h6 : _GEN_31033; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31035 = 10'h1f8 == _T_442[9:0] ? 4'h6 : _GEN_31034; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31036 = 10'h1f9 == _T_442[9:0] ? 4'h8 : _GEN_31035; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31037 = 10'h1fa == _T_442[9:0] ? 4'h8 : _GEN_31036; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31038 = 10'h1fb == _T_442[9:0] ? 4'h6 : _GEN_31037; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31039 = 10'h1fc == _T_442[9:0] ? 4'ha : _GEN_31038; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31040 = 10'h1fd == _T_442[9:0] ? 4'hb : _GEN_31039; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31041 = 10'h1fe == _T_442[9:0] ? 4'ha : _GEN_31040; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31042 = 10'h1ff == _T_442[9:0] ? 4'ha : _GEN_31041; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31043 = 10'h200 == _T_442[9:0] ? 4'h4 : _GEN_31042; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31044 = 10'h201 == _T_442[9:0] ? 4'h7 : _GEN_31043; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31045 = 10'h202 == _T_442[9:0] ? 4'h6 : _GEN_31044; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31046 = 10'h203 == _T_442[9:0] ? 4'h6 : _GEN_31045; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31047 = 10'h204 == _T_442[9:0] ? 4'h5 : _GEN_31046; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31048 = 10'h205 == _T_442[9:0] ? 4'h6 : _GEN_31047; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31049 = 10'h206 == _T_442[9:0] ? 4'h6 : _GEN_31048; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31050 = 10'h207 == _T_442[9:0] ? 4'h5 : _GEN_31049; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31051 = 10'h208 == _T_442[9:0] ? 4'h7 : _GEN_31050; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31052 = 10'h209 == _T_442[9:0] ? 4'h9 : _GEN_31051; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31053 = 10'h20a == _T_442[9:0] ? 4'hb : _GEN_31052; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31054 = 10'h20b == _T_442[9:0] ? 4'h7 : _GEN_31053; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31055 = 10'h20c == _T_442[9:0] ? 4'h7 : _GEN_31054; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31056 = 10'h20d == _T_442[9:0] ? 4'h7 : _GEN_31055; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31057 = 10'h20e == _T_442[9:0] ? 4'h7 : _GEN_31056; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31058 = 10'h20f == _T_442[9:0] ? 4'h7 : _GEN_31057; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31059 = 10'h210 == _T_442[9:0] ? 4'h7 : _GEN_31058; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31060 = 10'h211 == _T_442[9:0] ? 4'h8 : _GEN_31059; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31061 = 10'h212 == _T_442[9:0] ? 4'h8 : _GEN_31060; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31062 = 10'h213 == _T_442[9:0] ? 4'h9 : _GEN_31061; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31063 = 10'h214 == _T_442[9:0] ? 4'h6 : _GEN_31062; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31064 = 10'h215 == _T_442[9:0] ? 4'h7 : _GEN_31063; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31065 = 10'h216 == _T_442[9:0] ? 4'h7 : _GEN_31064; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31066 = 10'h217 == _T_442[9:0] ? 4'h7 : _GEN_31065; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31067 = 10'h218 == _T_442[9:0] ? 4'h7 : _GEN_31066; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31068 = 10'h219 == _T_442[9:0] ? 4'h8 : _GEN_31067; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31069 = 10'h21a == _T_442[9:0] ? 4'h7 : _GEN_31068; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31070 = 10'h21b == _T_442[9:0] ? 4'h8 : _GEN_31069; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31071 = 10'h21c == _T_442[9:0] ? 4'ha : _GEN_31070; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31072 = 10'h21d == _T_442[9:0] ? 4'ha : _GEN_31071; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31073 = 10'h21e == _T_442[9:0] ? 4'h7 : _GEN_31072; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31074 = 10'h21f == _T_442[9:0] ? 4'h6 : _GEN_31073; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31075 = 10'h220 == _T_442[9:0] ? 4'h6 : _GEN_31074; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31076 = 10'h221 == _T_442[9:0] ? 4'h7 : _GEN_31075; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31077 = 10'h222 == _T_442[9:0] ? 4'ha : _GEN_31076; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31078 = 10'h223 == _T_442[9:0] ? 4'ha : _GEN_31077; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31079 = 10'h224 == _T_442[9:0] ? 4'ha : _GEN_31078; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31080 = 10'h225 == _T_442[9:0] ? 4'h8 : _GEN_31079; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31081 = 10'h226 == _T_442[9:0] ? 4'h3 : _GEN_31080; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31082 = 10'h227 == _T_442[9:0] ? 4'h4 : _GEN_31081; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31083 = 10'h228 == _T_442[9:0] ? 4'h6 : _GEN_31082; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31084 = 10'h229 == _T_442[9:0] ? 4'h6 : _GEN_31083; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31085 = 10'h22a == _T_442[9:0] ? 4'h6 : _GEN_31084; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31086 = 10'h22b == _T_442[9:0] ? 4'h6 : _GEN_31085; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31087 = 10'h22c == _T_442[9:0] ? 4'h5 : _GEN_31086; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31088 = 10'h22d == _T_442[9:0] ? 4'h6 : _GEN_31087; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31089 = 10'h22e == _T_442[9:0] ? 4'h6 : _GEN_31088; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31090 = 10'h22f == _T_442[9:0] ? 4'h8 : _GEN_31089; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31091 = 10'h230 == _T_442[9:0] ? 4'h7 : _GEN_31090; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31092 = 10'h231 == _T_442[9:0] ? 4'h5 : _GEN_31091; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31093 = 10'h232 == _T_442[9:0] ? 4'h6 : _GEN_31092; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31094 = 10'h233 == _T_442[9:0] ? 4'h8 : _GEN_31093; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31095 = 10'h234 == _T_442[9:0] ? 4'h8 : _GEN_31094; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31096 = 10'h235 == _T_442[9:0] ? 4'h8 : _GEN_31095; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31097 = 10'h236 == _T_442[9:0] ? 4'h8 : _GEN_31096; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31098 = 10'h237 == _T_442[9:0] ? 4'h8 : _GEN_31097; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31099 = 10'h238 == _T_442[9:0] ? 4'h8 : _GEN_31098; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31100 = 10'h239 == _T_442[9:0] ? 4'h6 : _GEN_31099; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31101 = 10'h23a == _T_442[9:0] ? 4'h6 : _GEN_31100; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31102 = 10'h23b == _T_442[9:0] ? 4'h7 : _GEN_31101; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31103 = 10'h23c == _T_442[9:0] ? 4'h6 : _GEN_31102; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31104 = 10'h23d == _T_442[9:0] ? 4'h7 : _GEN_31103; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31105 = 10'h23e == _T_442[9:0] ? 4'h7 : _GEN_31104; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31106 = 10'h23f == _T_442[9:0] ? 4'h6 : _GEN_31105; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31107 = 10'h240 == _T_442[9:0] ? 4'h6 : _GEN_31106; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31108 = 10'h241 == _T_442[9:0] ? 4'h8 : _GEN_31107; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31109 = 10'h242 == _T_442[9:0] ? 4'ha : _GEN_31108; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31110 = 10'h243 == _T_442[9:0] ? 4'ha : _GEN_31109; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31111 = 10'h244 == _T_442[9:0] ? 4'ha : _GEN_31110; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31112 = 10'h245 == _T_442[9:0] ? 4'h8 : _GEN_31111; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31113 = 10'h246 == _T_442[9:0] ? 4'h8 : _GEN_31112; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31114 = 10'h247 == _T_442[9:0] ? 4'h9 : _GEN_31113; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31115 = 10'h248 == _T_442[9:0] ? 4'ha : _GEN_31114; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31116 = 10'h249 == _T_442[9:0] ? 4'ha : _GEN_31115; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31117 = 10'h24a == _T_442[9:0] ? 4'ha : _GEN_31116; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31118 = 10'h24b == _T_442[9:0] ? 4'h4 : _GEN_31117; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31119 = 10'h24c == _T_442[9:0] ? 4'h3 : _GEN_31118; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31120 = 10'h24d == _T_442[9:0] ? 4'h4 : _GEN_31119; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31121 = 10'h24e == _T_442[9:0] ? 4'h5 : _GEN_31120; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31122 = 10'h24f == _T_442[9:0] ? 4'h5 : _GEN_31121; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31123 = 10'h250 == _T_442[9:0] ? 4'h5 : _GEN_31122; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31124 = 10'h251 == _T_442[9:0] ? 4'h5 : _GEN_31123; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31125 = 10'h252 == _T_442[9:0] ? 4'h5 : _GEN_31124; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31126 = 10'h253 == _T_442[9:0] ? 4'h5 : _GEN_31125; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31127 = 10'h254 == _T_442[9:0] ? 4'h5 : _GEN_31126; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31128 = 10'h255 == _T_442[9:0] ? 4'h6 : _GEN_31127; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31129 = 10'h256 == _T_442[9:0] ? 4'h7 : _GEN_31128; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31130 = 10'h257 == _T_442[9:0] ? 4'h3 : _GEN_31129; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31131 = 10'h258 == _T_442[9:0] ? 4'h6 : _GEN_31130; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31132 = 10'h259 == _T_442[9:0] ? 4'h7 : _GEN_31131; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31133 = 10'h25a == _T_442[9:0] ? 4'h7 : _GEN_31132; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31134 = 10'h25b == _T_442[9:0] ? 4'h7 : _GEN_31133; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31135 = 10'h25c == _T_442[9:0] ? 4'h8 : _GEN_31134; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31136 = 10'h25d == _T_442[9:0] ? 4'h8 : _GEN_31135; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31137 = 10'h25e == _T_442[9:0] ? 4'h4 : _GEN_31136; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31138 = 10'h25f == _T_442[9:0] ? 4'h3 : _GEN_31137; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31139 = 10'h260 == _T_442[9:0] ? 4'h7 : _GEN_31138; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31140 = 10'h261 == _T_442[9:0] ? 4'h7 : _GEN_31139; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31141 = 10'h262 == _T_442[9:0] ? 4'h7 : _GEN_31140; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31142 = 10'h263 == _T_442[9:0] ? 4'h6 : _GEN_31141; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31143 = 10'h264 == _T_442[9:0] ? 4'h7 : _GEN_31142; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31144 = 10'h265 == _T_442[9:0] ? 4'h6 : _GEN_31143; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31145 = 10'h266 == _T_442[9:0] ? 4'h5 : _GEN_31144; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31146 = 10'h267 == _T_442[9:0] ? 4'h7 : _GEN_31145; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31147 = 10'h268 == _T_442[9:0] ? 4'ha : _GEN_31146; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31148 = 10'h269 == _T_442[9:0] ? 4'ha : _GEN_31147; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31149 = 10'h26a == _T_442[9:0] ? 4'ha : _GEN_31148; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31150 = 10'h26b == _T_442[9:0] ? 4'ha : _GEN_31149; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31151 = 10'h26c == _T_442[9:0] ? 4'ha : _GEN_31150; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31152 = 10'h26d == _T_442[9:0] ? 4'ha : _GEN_31151; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31153 = 10'h26e == _T_442[9:0] ? 4'ha : _GEN_31152; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31154 = 10'h26f == _T_442[9:0] ? 4'ha : _GEN_31153; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31155 = 10'h270 == _T_442[9:0] ? 4'h5 : _GEN_31154; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31156 = 10'h271 == _T_442[9:0] ? 4'h3 : _GEN_31155; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31157 = 10'h272 == _T_442[9:0] ? 4'h3 : _GEN_31156; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31158 = 10'h273 == _T_442[9:0] ? 4'h4 : _GEN_31157; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31159 = 10'h274 == _T_442[9:0] ? 4'h6 : _GEN_31158; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31160 = 10'h275 == _T_442[9:0] ? 4'h5 : _GEN_31159; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31161 = 10'h276 == _T_442[9:0] ? 4'h6 : _GEN_31160; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31162 = 10'h277 == _T_442[9:0] ? 4'h5 : _GEN_31161; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31163 = 10'h278 == _T_442[9:0] ? 4'h6 : _GEN_31162; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31164 = 10'h279 == _T_442[9:0] ? 4'h6 : _GEN_31163; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31165 = 10'h27a == _T_442[9:0] ? 4'h6 : _GEN_31164; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31166 = 10'h27b == _T_442[9:0] ? 4'h8 : _GEN_31165; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31167 = 10'h27c == _T_442[9:0] ? 4'h6 : _GEN_31166; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31168 = 10'h27d == _T_442[9:0] ? 4'h2 : _GEN_31167; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31169 = 10'h27e == _T_442[9:0] ? 4'h5 : _GEN_31168; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31170 = 10'h27f == _T_442[9:0] ? 4'h7 : _GEN_31169; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31171 = 10'h280 == _T_442[9:0] ? 4'h7 : _GEN_31170; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31172 = 10'h281 == _T_442[9:0] ? 4'h8 : _GEN_31171; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31173 = 10'h282 == _T_442[9:0] ? 4'h7 : _GEN_31172; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31174 = 10'h283 == _T_442[9:0] ? 4'h3 : _GEN_31173; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31175 = 10'h284 == _T_442[9:0] ? 4'h3 : _GEN_31174; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31176 = 10'h285 == _T_442[9:0] ? 4'h3 : _GEN_31175; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31177 = 10'h286 == _T_442[9:0] ? 4'h7 : _GEN_31176; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31178 = 10'h287 == _T_442[9:0] ? 4'h7 : _GEN_31177; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31179 = 10'h288 == _T_442[9:0] ? 4'h7 : _GEN_31178; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31180 = 10'h289 == _T_442[9:0] ? 4'h7 : _GEN_31179; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31181 = 10'h28a == _T_442[9:0] ? 4'h8 : _GEN_31180; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31182 = 10'h28b == _T_442[9:0] ? 4'h8 : _GEN_31181; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31183 = 10'h28c == _T_442[9:0] ? 4'h7 : _GEN_31182; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31184 = 10'h28d == _T_442[9:0] ? 4'h6 : _GEN_31183; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31185 = 10'h28e == _T_442[9:0] ? 4'h3 : _GEN_31184; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31186 = 10'h28f == _T_442[9:0] ? 4'h6 : _GEN_31185; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31187 = 10'h290 == _T_442[9:0] ? 4'h8 : _GEN_31186; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31188 = 10'h291 == _T_442[9:0] ? 4'ha : _GEN_31187; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31189 = 10'h292 == _T_442[9:0] ? 4'ha : _GEN_31188; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31190 = 10'h293 == _T_442[9:0] ? 4'ha : _GEN_31189; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31191 = 10'h294 == _T_442[9:0] ? 4'h9 : _GEN_31190; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31192 = 10'h295 == _T_442[9:0] ? 4'h4 : _GEN_31191; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31193 = 10'h296 == _T_442[9:0] ? 4'h3 : _GEN_31192; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31194 = 10'h297 == _T_442[9:0] ? 4'h3 : _GEN_31193; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31195 = 10'h298 == _T_442[9:0] ? 4'h3 : _GEN_31194; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31196 = 10'h299 == _T_442[9:0] ? 4'h4 : _GEN_31195; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31197 = 10'h29a == _T_442[9:0] ? 4'h5 : _GEN_31196; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31198 = 10'h29b == _T_442[9:0] ? 4'h5 : _GEN_31197; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31199 = 10'h29c == _T_442[9:0] ? 4'h5 : _GEN_31198; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31200 = 10'h29d == _T_442[9:0] ? 4'h5 : _GEN_31199; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31201 = 10'h29e == _T_442[9:0] ? 4'h5 : _GEN_31200; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31202 = 10'h29f == _T_442[9:0] ? 4'h5 : _GEN_31201; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31203 = 10'h2a0 == _T_442[9:0] ? 4'h6 : _GEN_31202; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31204 = 10'h2a1 == _T_442[9:0] ? 4'h7 : _GEN_31203; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31205 = 10'h2a2 == _T_442[9:0] ? 4'h5 : _GEN_31204; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31206 = 10'h2a3 == _T_442[9:0] ? 4'h2 : _GEN_31205; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31207 = 10'h2a4 == _T_442[9:0] ? 4'h3 : _GEN_31206; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31208 = 10'h2a5 == _T_442[9:0] ? 4'h7 : _GEN_31207; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31209 = 10'h2a6 == _T_442[9:0] ? 4'h8 : _GEN_31208; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31210 = 10'h2a7 == _T_442[9:0] ? 4'h7 : _GEN_31209; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31211 = 10'h2a8 == _T_442[9:0] ? 4'h3 : _GEN_31210; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31212 = 10'h2a9 == _T_442[9:0] ? 4'h2 : _GEN_31211; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31213 = 10'h2aa == _T_442[9:0] ? 4'h3 : _GEN_31212; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31214 = 10'h2ab == _T_442[9:0] ? 4'h3 : _GEN_31213; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31215 = 10'h2ac == _T_442[9:0] ? 4'h7 : _GEN_31214; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31216 = 10'h2ad == _T_442[9:0] ? 4'h8 : _GEN_31215; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31217 = 10'h2ae == _T_442[9:0] ? 4'h7 : _GEN_31216; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31218 = 10'h2af == _T_442[9:0] ? 4'h8 : _GEN_31217; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31219 = 10'h2b0 == _T_442[9:0] ? 4'h8 : _GEN_31218; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31220 = 10'h2b1 == _T_442[9:0] ? 4'h8 : _GEN_31219; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31221 = 10'h2b2 == _T_442[9:0] ? 4'h7 : _GEN_31220; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31222 = 10'h2b3 == _T_442[9:0] ? 4'h6 : _GEN_31221; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31223 = 10'h2b4 == _T_442[9:0] ? 4'h2 : _GEN_31222; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31224 = 10'h2b5 == _T_442[9:0] ? 4'h2 : _GEN_31223; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31225 = 10'h2b6 == _T_442[9:0] ? 4'h3 : _GEN_31224; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31226 = 10'h2b7 == _T_442[9:0] ? 4'h3 : _GEN_31225; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31227 = 10'h2b8 == _T_442[9:0] ? 4'h6 : _GEN_31226; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31228 = 10'h2b9 == _T_442[9:0] ? 4'h9 : _GEN_31227; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31229 = 10'h2ba == _T_442[9:0] ? 4'h3 : _GEN_31228; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31230 = 10'h2bb == _T_442[9:0] ? 4'h3 : _GEN_31229; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31231 = 10'h2bc == _T_442[9:0] ? 4'h3 : _GEN_31230; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31232 = 10'h2bd == _T_442[9:0] ? 4'h2 : _GEN_31231; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31233 = 10'h2be == _T_442[9:0] ? 4'h3 : _GEN_31232; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31234 = 10'h2bf == _T_442[9:0] ? 4'h3 : _GEN_31233; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31235 = 10'h2c0 == _T_442[9:0] ? 4'h5 : _GEN_31234; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31236 = 10'h2c1 == _T_442[9:0] ? 4'h5 : _GEN_31235; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31237 = 10'h2c2 == _T_442[9:0] ? 4'h5 : _GEN_31236; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31238 = 10'h2c3 == _T_442[9:0] ? 4'h5 : _GEN_31237; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31239 = 10'h2c4 == _T_442[9:0] ? 4'h5 : _GEN_31238; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31240 = 10'h2c5 == _T_442[9:0] ? 4'h5 : _GEN_31239; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31241 = 10'h2c6 == _T_442[9:0] ? 4'h6 : _GEN_31240; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31242 = 10'h2c7 == _T_442[9:0] ? 4'h7 : _GEN_31241; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31243 = 10'h2c8 == _T_442[9:0] ? 4'h5 : _GEN_31242; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31244 = 10'h2c9 == _T_442[9:0] ? 4'h2 : _GEN_31243; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31245 = 10'h2ca == _T_442[9:0] ? 4'h2 : _GEN_31244; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31246 = 10'h2cb == _T_442[9:0] ? 4'h3 : _GEN_31245; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31247 = 10'h2cc == _T_442[9:0] ? 4'h3 : _GEN_31246; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31248 = 10'h2cd == _T_442[9:0] ? 4'h2 : _GEN_31247; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31249 = 10'h2ce == _T_442[9:0] ? 4'h2 : _GEN_31248; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31250 = 10'h2cf == _T_442[9:0] ? 4'h2 : _GEN_31249; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31251 = 10'h2d0 == _T_442[9:0] ? 4'h2 : _GEN_31250; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31252 = 10'h2d1 == _T_442[9:0] ? 4'h2 : _GEN_31251; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31253 = 10'h2d2 == _T_442[9:0] ? 4'h7 : _GEN_31252; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31254 = 10'h2d3 == _T_442[9:0] ? 4'h7 : _GEN_31253; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31255 = 10'h2d4 == _T_442[9:0] ? 4'h8 : _GEN_31254; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31256 = 10'h2d5 == _T_442[9:0] ? 4'h8 : _GEN_31255; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31257 = 10'h2d6 == _T_442[9:0] ? 4'h8 : _GEN_31256; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31258 = 10'h2d7 == _T_442[9:0] ? 4'h8 : _GEN_31257; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31259 = 10'h2d8 == _T_442[9:0] ? 4'h7 : _GEN_31258; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31260 = 10'h2d9 == _T_442[9:0] ? 4'h6 : _GEN_31259; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31261 = 10'h2da == _T_442[9:0] ? 4'h4 : _GEN_31260; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31262 = 10'h2db == _T_442[9:0] ? 4'h2 : _GEN_31261; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31263 = 10'h2dc == _T_442[9:0] ? 4'h2 : _GEN_31262; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31264 = 10'h2dd == _T_442[9:0] ? 4'h3 : _GEN_31263; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31265 = 10'h2de == _T_442[9:0] ? 4'h3 : _GEN_31264; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31266 = 10'h2df == _T_442[9:0] ? 4'h3 : _GEN_31265; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31267 = 10'h2e0 == _T_442[9:0] ? 4'h3 : _GEN_31266; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31268 = 10'h2e1 == _T_442[9:0] ? 4'h3 : _GEN_31267; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31269 = 10'h2e2 == _T_442[9:0] ? 4'h3 : _GEN_31268; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31270 = 10'h2e3 == _T_442[9:0] ? 4'h2 : _GEN_31269; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31271 = 10'h2e4 == _T_442[9:0] ? 4'h3 : _GEN_31270; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31272 = 10'h2e5 == _T_442[9:0] ? 4'h2 : _GEN_31271; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31273 = 10'h2e6 == _T_442[9:0] ? 4'h5 : _GEN_31272; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31274 = 10'h2e7 == _T_442[9:0] ? 4'h5 : _GEN_31273; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31275 = 10'h2e8 == _T_442[9:0] ? 4'h5 : _GEN_31274; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31276 = 10'h2e9 == _T_442[9:0] ? 4'h5 : _GEN_31275; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31277 = 10'h2ea == _T_442[9:0] ? 4'h5 : _GEN_31276; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31278 = 10'h2eb == _T_442[9:0] ? 4'h5 : _GEN_31277; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31279 = 10'h2ec == _T_442[9:0] ? 4'h6 : _GEN_31278; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31280 = 10'h2ed == _T_442[9:0] ? 4'h7 : _GEN_31279; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31281 = 10'h2ee == _T_442[9:0] ? 4'h6 : _GEN_31280; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31282 = 10'h2ef == _T_442[9:0] ? 4'h2 : _GEN_31281; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31283 = 10'h2f0 == _T_442[9:0] ? 4'h2 : _GEN_31282; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31284 = 10'h2f1 == _T_442[9:0] ? 4'h2 : _GEN_31283; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31285 = 10'h2f2 == _T_442[9:0] ? 4'h2 : _GEN_31284; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31286 = 10'h2f3 == _T_442[9:0] ? 4'h2 : _GEN_31285; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31287 = 10'h2f4 == _T_442[9:0] ? 4'h2 : _GEN_31286; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31288 = 10'h2f5 == _T_442[9:0] ? 4'h2 : _GEN_31287; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31289 = 10'h2f6 == _T_442[9:0] ? 4'h2 : _GEN_31288; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31290 = 10'h2f7 == _T_442[9:0] ? 4'h2 : _GEN_31289; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31291 = 10'h2f8 == _T_442[9:0] ? 4'h7 : _GEN_31290; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31292 = 10'h2f9 == _T_442[9:0] ? 4'h7 : _GEN_31291; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31293 = 10'h2fa == _T_442[9:0] ? 4'h8 : _GEN_31292; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31294 = 10'h2fb == _T_442[9:0] ? 4'h8 : _GEN_31293; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31295 = 10'h2fc == _T_442[9:0] ? 4'h7 : _GEN_31294; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31296 = 10'h2fd == _T_442[9:0] ? 4'h7 : _GEN_31295; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31297 = 10'h2fe == _T_442[9:0] ? 4'h7 : _GEN_31296; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31298 = 10'h2ff == _T_442[9:0] ? 4'h7 : _GEN_31297; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31299 = 10'h300 == _T_442[9:0] ? 4'h8 : _GEN_31298; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31300 = 10'h301 == _T_442[9:0] ? 4'h7 : _GEN_31299; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31301 = 10'h302 == _T_442[9:0] ? 4'h3 : _GEN_31300; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31302 = 10'h303 == _T_442[9:0] ? 4'h3 : _GEN_31301; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31303 = 10'h304 == _T_442[9:0] ? 4'h2 : _GEN_31302; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31304 = 10'h305 == _T_442[9:0] ? 4'h2 : _GEN_31303; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31305 = 10'h306 == _T_442[9:0] ? 4'h2 : _GEN_31304; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31306 = 10'h307 == _T_442[9:0] ? 4'h2 : _GEN_31305; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31307 = 10'h308 == _T_442[9:0] ? 4'h2 : _GEN_31306; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31308 = 10'h309 == _T_442[9:0] ? 4'h2 : _GEN_31307; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31309 = 10'h30a == _T_442[9:0] ? 4'h2 : _GEN_31308; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31310 = 10'h30b == _T_442[9:0] ? 4'h3 : _GEN_31309; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31311 = 10'h30c == _T_442[9:0] ? 4'h4 : _GEN_31310; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31312 = 10'h30d == _T_442[9:0] ? 4'h5 : _GEN_31311; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31313 = 10'h30e == _T_442[9:0] ? 4'h5 : _GEN_31312; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31314 = 10'h30f == _T_442[9:0] ? 4'h5 : _GEN_31313; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31315 = 10'h310 == _T_442[9:0] ? 4'h5 : _GEN_31314; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31316 = 10'h311 == _T_442[9:0] ? 4'h5 : _GEN_31315; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31317 = 10'h312 == _T_442[9:0] ? 4'h6 : _GEN_31316; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31318 = 10'h313 == _T_442[9:0] ? 4'h7 : _GEN_31317; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31319 = 10'h314 == _T_442[9:0] ? 4'h7 : _GEN_31318; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31320 = 10'h315 == _T_442[9:0] ? 4'h3 : _GEN_31319; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31321 = 10'h316 == _T_442[9:0] ? 4'h2 : _GEN_31320; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31322 = 10'h317 == _T_442[9:0] ? 4'h2 : _GEN_31321; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31323 = 10'h318 == _T_442[9:0] ? 4'h2 : _GEN_31322; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31324 = 10'h319 == _T_442[9:0] ? 4'h2 : _GEN_31323; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31325 = 10'h31a == _T_442[9:0] ? 4'h2 : _GEN_31324; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31326 = 10'h31b == _T_442[9:0] ? 4'h2 : _GEN_31325; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31327 = 10'h31c == _T_442[9:0] ? 4'h2 : _GEN_31326; // @[Filter.scala 230:142]
  wire [3:0] _GEN_31328 = 10'h31d == _T_442[9:0] ? 4'h2 : _GEN_31327; // @[Filter.scala 230:142]
  wire [7:0] _T_456 = _GEN_31328 * 4'ha; // @[Filter.scala 230:142]
  wire [10:0] _GEN_39031 = {{3'd0}, _T_456}; // @[Filter.scala 230:109]
  wire [10:0] _T_458 = _T_451 + _GEN_39031; // @[Filter.scala 230:109]
  wire [10:0] _T_459 = _T_458 / 11'h64; // @[Filter.scala 230:150]
  wire  _T_461 = _T_432 >= 6'h20; // @[Filter.scala 233:31]
  wire  _T_465 = _T_439 >= 32'h12; // @[Filter.scala 233:63]
  wire  _T_466 = _T_461 | _T_465; // @[Filter.scala 233:58]
  wire [10:0] _GEN_32127 = io_SPI_distort ? _T_459 : {{7'd0}, _GEN_29732}; // @[Filter.scala 235:35]
  wire [10:0] _GEN_32128 = _T_466 ? 11'h0 : _GEN_32127; // @[Filter.scala 233:80]
  wire [10:0] _GEN_32927 = io_SPI_distort ? _T_459 : {{7'd0}, _GEN_30530}; // @[Filter.scala 235:35]
  wire [10:0] _GEN_32928 = _T_466 ? 11'h0 : _GEN_32927; // @[Filter.scala 233:80]
  wire [10:0] _GEN_33727 = io_SPI_distort ? _T_459 : {{7'd0}, _GEN_31328}; // @[Filter.scala 235:35]
  wire [10:0] _GEN_33728 = _T_466 ? 11'h0 : _GEN_33727; // @[Filter.scala 233:80]
  wire [31:0] _T_494 = pixelIndex + 32'h7; // @[Filter.scala 228:31]
  wire [31:0] _GEN_56 = _T_494 % 32'h20; // @[Filter.scala 228:38]
  wire [5:0] _T_495 = _GEN_56[5:0]; // @[Filter.scala 228:38]
  wire [5:0] _T_497 = _T_495 + _GEN_38951; // @[Filter.scala 228:53]
  wire [5:0] _T_499 = _T_497 - 6'h1; // @[Filter.scala 228:69]
  wire [31:0] _T_502 = _T_494 / 32'h20; // @[Filter.scala 229:38]
  wire [31:0] _T_504 = _T_502 + _GEN_38952; // @[Filter.scala 229:53]
  wire [31:0] _T_506 = _T_504 - 32'h1; // @[Filter.scala 229:69]
  wire [37:0] _T_507 = _T_506 * 32'h20; // @[Filter.scala 230:42]
  wire [37:0] _GEN_39037 = {{32'd0}, _T_499}; // @[Filter.scala 230:57]
  wire [37:0] _T_509 = _T_507 + _GEN_39037; // @[Filter.scala 230:57]
  wire [3:0] _GEN_33751 = 10'h16 == _T_509[9:0] ? 4'h9 : 4'ha; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33752 = 10'h17 == _T_509[9:0] ? 4'h3 : _GEN_33751; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33753 = 10'h18 == _T_509[9:0] ? 4'h6 : _GEN_33752; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33754 = 10'h19 == _T_509[9:0] ? 4'ha : _GEN_33753; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33755 = 10'h1a == _T_509[9:0] ? 4'ha : _GEN_33754; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33756 = 10'h1b == _T_509[9:0] ? 4'ha : _GEN_33755; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33757 = 10'h1c == _T_509[9:0] ? 4'ha : _GEN_33756; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33758 = 10'h1d == _T_509[9:0] ? 4'ha : _GEN_33757; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33759 = 10'h1e == _T_509[9:0] ? 4'ha : _GEN_33758; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33760 = 10'h1f == _T_509[9:0] ? 4'ha : _GEN_33759; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33761 = 10'h20 == _T_509[9:0] ? 4'ha : _GEN_33760; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33762 = 10'h21 == _T_509[9:0] ? 4'ha : _GEN_33761; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33763 = 10'h22 == _T_509[9:0] ? 4'ha : _GEN_33762; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33764 = 10'h23 == _T_509[9:0] ? 4'ha : _GEN_33763; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33765 = 10'h24 == _T_509[9:0] ? 4'ha : _GEN_33764; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33766 = 10'h25 == _T_509[9:0] ? 4'ha : _GEN_33765; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33767 = 10'h26 == _T_509[9:0] ? 4'ha : _GEN_33766; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33768 = 10'h27 == _T_509[9:0] ? 4'ha : _GEN_33767; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33769 = 10'h28 == _T_509[9:0] ? 4'ha : _GEN_33768; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33770 = 10'h29 == _T_509[9:0] ? 4'ha : _GEN_33769; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33771 = 10'h2a == _T_509[9:0] ? 4'ha : _GEN_33770; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33772 = 10'h2b == _T_509[9:0] ? 4'ha : _GEN_33771; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33773 = 10'h2c == _T_509[9:0] ? 4'ha : _GEN_33772; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33774 = 10'h2d == _T_509[9:0] ? 4'ha : _GEN_33773; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33775 = 10'h2e == _T_509[9:0] ? 4'ha : _GEN_33774; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33776 = 10'h2f == _T_509[9:0] ? 4'ha : _GEN_33775; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33777 = 10'h30 == _T_509[9:0] ? 4'ha : _GEN_33776; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33778 = 10'h31 == _T_509[9:0] ? 4'ha : _GEN_33777; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33779 = 10'h32 == _T_509[9:0] ? 4'ha : _GEN_33778; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33780 = 10'h33 == _T_509[9:0] ? 4'ha : _GEN_33779; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33781 = 10'h34 == _T_509[9:0] ? 4'ha : _GEN_33780; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33782 = 10'h35 == _T_509[9:0] ? 4'ha : _GEN_33781; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33783 = 10'h36 == _T_509[9:0] ? 4'ha : _GEN_33782; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33784 = 10'h37 == _T_509[9:0] ? 4'ha : _GEN_33783; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33785 = 10'h38 == _T_509[9:0] ? 4'ha : _GEN_33784; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33786 = 10'h39 == _T_509[9:0] ? 4'ha : _GEN_33785; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33787 = 10'h3a == _T_509[9:0] ? 4'ha : _GEN_33786; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33788 = 10'h3b == _T_509[9:0] ? 4'h9 : _GEN_33787; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33789 = 10'h3c == _T_509[9:0] ? 4'h4 : _GEN_33788; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33790 = 10'h3d == _T_509[9:0] ? 4'h3 : _GEN_33789; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33791 = 10'h3e == _T_509[9:0] ? 4'h4 : _GEN_33790; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33792 = 10'h3f == _T_509[9:0] ? 4'ha : _GEN_33791; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33793 = 10'h40 == _T_509[9:0] ? 4'ha : _GEN_33792; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33794 = 10'h41 == _T_509[9:0] ? 4'ha : _GEN_33793; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33795 = 10'h42 == _T_509[9:0] ? 4'ha : _GEN_33794; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33796 = 10'h43 == _T_509[9:0] ? 4'ha : _GEN_33795; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33797 = 10'h44 == _T_509[9:0] ? 4'ha : _GEN_33796; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33798 = 10'h45 == _T_509[9:0] ? 4'ha : _GEN_33797; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33799 = 10'h46 == _T_509[9:0] ? 4'ha : _GEN_33798; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33800 = 10'h47 == _T_509[9:0] ? 4'ha : _GEN_33799; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33801 = 10'h48 == _T_509[9:0] ? 4'ha : _GEN_33800; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33802 = 10'h49 == _T_509[9:0] ? 4'ha : _GEN_33801; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33803 = 10'h4a == _T_509[9:0] ? 4'ha : _GEN_33802; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33804 = 10'h4b == _T_509[9:0] ? 4'ha : _GEN_33803; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33805 = 10'h4c == _T_509[9:0] ? 4'ha : _GEN_33804; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33806 = 10'h4d == _T_509[9:0] ? 4'ha : _GEN_33805; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33807 = 10'h4e == _T_509[9:0] ? 4'ha : _GEN_33806; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33808 = 10'h4f == _T_509[9:0] ? 4'ha : _GEN_33807; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33809 = 10'h50 == _T_509[9:0] ? 4'ha : _GEN_33808; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33810 = 10'h51 == _T_509[9:0] ? 4'ha : _GEN_33809; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33811 = 10'h52 == _T_509[9:0] ? 4'ha : _GEN_33810; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33812 = 10'h53 == _T_509[9:0] ? 4'ha : _GEN_33811; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33813 = 10'h54 == _T_509[9:0] ? 4'ha : _GEN_33812; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33814 = 10'h55 == _T_509[9:0] ? 4'ha : _GEN_33813; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33815 = 10'h56 == _T_509[9:0] ? 4'ha : _GEN_33814; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33816 = 10'h57 == _T_509[9:0] ? 4'ha : _GEN_33815; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33817 = 10'h58 == _T_509[9:0] ? 4'ha : _GEN_33816; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33818 = 10'h59 == _T_509[9:0] ? 4'ha : _GEN_33817; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33819 = 10'h5a == _T_509[9:0] ? 4'h7 : _GEN_33818; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33820 = 10'h5b == _T_509[9:0] ? 4'h7 : _GEN_33819; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33821 = 10'h5c == _T_509[9:0] ? 4'ha : _GEN_33820; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33822 = 10'h5d == _T_509[9:0] ? 4'ha : _GEN_33821; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33823 = 10'h5e == _T_509[9:0] ? 4'ha : _GEN_33822; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33824 = 10'h5f == _T_509[9:0] ? 4'ha : _GEN_33823; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33825 = 10'h60 == _T_509[9:0] ? 4'ha : _GEN_33824; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33826 = 10'h61 == _T_509[9:0] ? 4'h8 : _GEN_33825; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33827 = 10'h62 == _T_509[9:0] ? 4'h3 : _GEN_33826; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33828 = 10'h63 == _T_509[9:0] ? 4'h3 : _GEN_33827; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33829 = 10'h64 == _T_509[9:0] ? 4'h3 : _GEN_33828; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33830 = 10'h65 == _T_509[9:0] ? 4'h9 : _GEN_33829; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33831 = 10'h66 == _T_509[9:0] ? 4'ha : _GEN_33830; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33832 = 10'h67 == _T_509[9:0] ? 4'ha : _GEN_33831; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33833 = 10'h68 == _T_509[9:0] ? 4'ha : _GEN_33832; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33834 = 10'h69 == _T_509[9:0] ? 4'ha : _GEN_33833; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33835 = 10'h6a == _T_509[9:0] ? 4'ha : _GEN_33834; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33836 = 10'h6b == _T_509[9:0] ? 4'h8 : _GEN_33835; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33837 = 10'h6c == _T_509[9:0] ? 4'h5 : _GEN_33836; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33838 = 10'h6d == _T_509[9:0] ? 4'h8 : _GEN_33837; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33839 = 10'h6e == _T_509[9:0] ? 4'ha : _GEN_33838; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33840 = 10'h6f == _T_509[9:0] ? 4'ha : _GEN_33839; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33841 = 10'h70 == _T_509[9:0] ? 4'ha : _GEN_33840; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33842 = 10'h71 == _T_509[9:0] ? 4'ha : _GEN_33841; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33843 = 10'h72 == _T_509[9:0] ? 4'ha : _GEN_33842; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33844 = 10'h73 == _T_509[9:0] ? 4'ha : _GEN_33843; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33845 = 10'h74 == _T_509[9:0] ? 4'ha : _GEN_33844; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33846 = 10'h75 == _T_509[9:0] ? 4'ha : _GEN_33845; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33847 = 10'h76 == _T_509[9:0] ? 4'ha : _GEN_33846; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33848 = 10'h77 == _T_509[9:0] ? 4'ha : _GEN_33847; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33849 = 10'h78 == _T_509[9:0] ? 4'ha : _GEN_33848; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33850 = 10'h79 == _T_509[9:0] ? 4'ha : _GEN_33849; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33851 = 10'h7a == _T_509[9:0] ? 4'ha : _GEN_33850; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33852 = 10'h7b == _T_509[9:0] ? 4'ha : _GEN_33851; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33853 = 10'h7c == _T_509[9:0] ? 4'ha : _GEN_33852; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33854 = 10'h7d == _T_509[9:0] ? 4'ha : _GEN_33853; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33855 = 10'h7e == _T_509[9:0] ? 4'ha : _GEN_33854; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33856 = 10'h7f == _T_509[9:0] ? 4'ha : _GEN_33855; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33857 = 10'h80 == _T_509[9:0] ? 4'ha : _GEN_33856; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33858 = 10'h81 == _T_509[9:0] ? 4'h5 : _GEN_33857; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33859 = 10'h82 == _T_509[9:0] ? 4'h5 : _GEN_33858; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33860 = 10'h83 == _T_509[9:0] ? 4'h7 : _GEN_33859; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33861 = 10'h84 == _T_509[9:0] ? 4'ha : _GEN_33860; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33862 = 10'h85 == _T_509[9:0] ? 4'ha : _GEN_33861; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33863 = 10'h86 == _T_509[9:0] ? 4'ha : _GEN_33862; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33864 = 10'h87 == _T_509[9:0] ? 4'h5 : _GEN_33863; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33865 = 10'h88 == _T_509[9:0] ? 4'h3 : _GEN_33864; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33866 = 10'h89 == _T_509[9:0] ? 4'h3 : _GEN_33865; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33867 = 10'h8a == _T_509[9:0] ? 4'h4 : _GEN_33866; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33868 = 10'h8b == _T_509[9:0] ? 4'h9 : _GEN_33867; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33869 = 10'h8c == _T_509[9:0] ? 4'ha : _GEN_33868; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33870 = 10'h8d == _T_509[9:0] ? 4'ha : _GEN_33869; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33871 = 10'h8e == _T_509[9:0] ? 4'ha : _GEN_33870; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33872 = 10'h8f == _T_509[9:0] ? 4'h6 : _GEN_33871; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33873 = 10'h90 == _T_509[9:0] ? 4'h4 : _GEN_33872; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33874 = 10'h91 == _T_509[9:0] ? 4'h3 : _GEN_33873; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33875 = 10'h92 == _T_509[9:0] ? 4'h7 : _GEN_33874; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33876 = 10'h93 == _T_509[9:0] ? 4'ha : _GEN_33875; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33877 = 10'h94 == _T_509[9:0] ? 4'ha : _GEN_33876; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33878 = 10'h95 == _T_509[9:0] ? 4'ha : _GEN_33877; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33879 = 10'h96 == _T_509[9:0] ? 4'ha : _GEN_33878; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33880 = 10'h97 == _T_509[9:0] ? 4'ha : _GEN_33879; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33881 = 10'h98 == _T_509[9:0] ? 4'ha : _GEN_33880; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33882 = 10'h99 == _T_509[9:0] ? 4'ha : _GEN_33881; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33883 = 10'h9a == _T_509[9:0] ? 4'ha : _GEN_33882; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33884 = 10'h9b == _T_509[9:0] ? 4'ha : _GEN_33883; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33885 = 10'h9c == _T_509[9:0] ? 4'ha : _GEN_33884; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33886 = 10'h9d == _T_509[9:0] ? 4'ha : _GEN_33885; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33887 = 10'h9e == _T_509[9:0] ? 4'ha : _GEN_33886; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33888 = 10'h9f == _T_509[9:0] ? 4'ha : _GEN_33887; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33889 = 10'ha0 == _T_509[9:0] ? 4'ha : _GEN_33888; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33890 = 10'ha1 == _T_509[9:0] ? 4'ha : _GEN_33889; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33891 = 10'ha2 == _T_509[9:0] ? 4'ha : _GEN_33890; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33892 = 10'ha3 == _T_509[9:0] ? 4'ha : _GEN_33891; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33893 = 10'ha4 == _T_509[9:0] ? 4'ha : _GEN_33892; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33894 = 10'ha5 == _T_509[9:0] ? 4'ha : _GEN_33893; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33895 = 10'ha6 == _T_509[9:0] ? 4'ha : _GEN_33894; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33896 = 10'ha7 == _T_509[9:0] ? 4'h9 : _GEN_33895; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33897 = 10'ha8 == _T_509[9:0] ? 4'h4 : _GEN_33896; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33898 = 10'ha9 == _T_509[9:0] ? 4'h3 : _GEN_33897; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33899 = 10'haa == _T_509[9:0] ? 4'h4 : _GEN_33898; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33900 = 10'hab == _T_509[9:0] ? 4'h7 : _GEN_33899; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33901 = 10'hac == _T_509[9:0] ? 4'h8 : _GEN_33900; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33902 = 10'had == _T_509[9:0] ? 4'h3 : _GEN_33901; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33903 = 10'hae == _T_509[9:0] ? 4'h3 : _GEN_33902; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33904 = 10'haf == _T_509[9:0] ? 4'h3 : _GEN_33903; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33905 = 10'hb0 == _T_509[9:0] ? 4'h3 : _GEN_33904; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33906 = 10'hb1 == _T_509[9:0] ? 4'h7 : _GEN_33905; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33907 = 10'hb2 == _T_509[9:0] ? 4'h9 : _GEN_33906; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33908 = 10'hb3 == _T_509[9:0] ? 4'h6 : _GEN_33907; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33909 = 10'hb4 == _T_509[9:0] ? 4'h4 : _GEN_33908; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33910 = 10'hb5 == _T_509[9:0] ? 4'h3 : _GEN_33909; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33911 = 10'hb6 == _T_509[9:0] ? 4'h3 : _GEN_33910; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33912 = 10'hb7 == _T_509[9:0] ? 4'h6 : _GEN_33911; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33913 = 10'hb8 == _T_509[9:0] ? 4'ha : _GEN_33912; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33914 = 10'hb9 == _T_509[9:0] ? 4'ha : _GEN_33913; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33915 = 10'hba == _T_509[9:0] ? 4'ha : _GEN_33914; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33916 = 10'hbb == _T_509[9:0] ? 4'ha : _GEN_33915; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33917 = 10'hbc == _T_509[9:0] ? 4'ha : _GEN_33916; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33918 = 10'hbd == _T_509[9:0] ? 4'h9 : _GEN_33917; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33919 = 10'hbe == _T_509[9:0] ? 4'ha : _GEN_33918; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33920 = 10'hbf == _T_509[9:0] ? 4'ha : _GEN_33919; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33921 = 10'hc0 == _T_509[9:0] ? 4'ha : _GEN_33920; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33922 = 10'hc1 == _T_509[9:0] ? 4'ha : _GEN_33921; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33923 = 10'hc2 == _T_509[9:0] ? 4'ha : _GEN_33922; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33924 = 10'hc3 == _T_509[9:0] ? 4'ha : _GEN_33923; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33925 = 10'hc4 == _T_509[9:0] ? 4'ha : _GEN_33924; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33926 = 10'hc5 == _T_509[9:0] ? 4'ha : _GEN_33925; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33927 = 10'hc6 == _T_509[9:0] ? 4'ha : _GEN_33926; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33928 = 10'hc7 == _T_509[9:0] ? 4'h9 : _GEN_33927; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33929 = 10'hc8 == _T_509[9:0] ? 4'h8 : _GEN_33928; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33930 = 10'hc9 == _T_509[9:0] ? 4'h8 : _GEN_33929; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33931 = 10'hca == _T_509[9:0] ? 4'h9 : _GEN_33930; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33932 = 10'hcb == _T_509[9:0] ? 4'ha : _GEN_33931; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33933 = 10'hcc == _T_509[9:0] ? 4'ha : _GEN_33932; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33934 = 10'hcd == _T_509[9:0] ? 4'ha : _GEN_33933; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33935 = 10'hce == _T_509[9:0] ? 4'h8 : _GEN_33934; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33936 = 10'hcf == _T_509[9:0] ? 4'h3 : _GEN_33935; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33937 = 10'hd0 == _T_509[9:0] ? 4'h3 : _GEN_33936; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33938 = 10'hd1 == _T_509[9:0] ? 4'h3 : _GEN_33937; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33939 = 10'hd2 == _T_509[9:0] ? 4'h4 : _GEN_33938; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33940 = 10'hd3 == _T_509[9:0] ? 4'h3 : _GEN_33939; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33941 = 10'hd4 == _T_509[9:0] ? 4'h3 : _GEN_33940; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33942 = 10'hd5 == _T_509[9:0] ? 4'h3 : _GEN_33941; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33943 = 10'hd6 == _T_509[9:0] ? 4'h3 : _GEN_33942; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33944 = 10'hd7 == _T_509[9:0] ? 4'h5 : _GEN_33943; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33945 = 10'hd8 == _T_509[9:0] ? 4'h4 : _GEN_33944; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33946 = 10'hd9 == _T_509[9:0] ? 4'h3 : _GEN_33945; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33947 = 10'hda == _T_509[9:0] ? 4'h3 : _GEN_33946; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33948 = 10'hdb == _T_509[9:0] ? 4'h3 : _GEN_33947; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33949 = 10'hdc == _T_509[9:0] ? 4'h4 : _GEN_33948; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33950 = 10'hdd == _T_509[9:0] ? 4'ha : _GEN_33949; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33951 = 10'hde == _T_509[9:0] ? 4'ha : _GEN_33950; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33952 = 10'hdf == _T_509[9:0] ? 4'ha : _GEN_33951; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33953 = 10'he0 == _T_509[9:0] ? 4'ha : _GEN_33952; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33954 = 10'he1 == _T_509[9:0] ? 4'ha : _GEN_33953; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33955 = 10'he2 == _T_509[9:0] ? 4'ha : _GEN_33954; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33956 = 10'he3 == _T_509[9:0] ? 4'h5 : _GEN_33955; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33957 = 10'he4 == _T_509[9:0] ? 4'ha : _GEN_33956; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33958 = 10'he5 == _T_509[9:0] ? 4'ha : _GEN_33957; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33959 = 10'he6 == _T_509[9:0] ? 4'ha : _GEN_33958; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33960 = 10'he7 == _T_509[9:0] ? 4'ha : _GEN_33959; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33961 = 10'he8 == _T_509[9:0] ? 4'ha : _GEN_33960; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33962 = 10'he9 == _T_509[9:0] ? 4'ha : _GEN_33961; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33963 = 10'hea == _T_509[9:0] ? 4'ha : _GEN_33962; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33964 = 10'heb == _T_509[9:0] ? 4'h9 : _GEN_33963; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33965 = 10'hec == _T_509[9:0] ? 4'h7 : _GEN_33964; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33966 = 10'hed == _T_509[9:0] ? 4'h3 : _GEN_33965; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33967 = 10'hee == _T_509[9:0] ? 4'h3 : _GEN_33966; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33968 = 10'hef == _T_509[9:0] ? 4'h3 : _GEN_33967; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33969 = 10'hf0 == _T_509[9:0] ? 4'h4 : _GEN_33968; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33970 = 10'hf1 == _T_509[9:0] ? 4'h7 : _GEN_33969; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33971 = 10'hf2 == _T_509[9:0] ? 4'ha : _GEN_33970; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33972 = 10'hf3 == _T_509[9:0] ? 4'ha : _GEN_33971; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33973 = 10'hf4 == _T_509[9:0] ? 4'ha : _GEN_33972; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33974 = 10'hf5 == _T_509[9:0] ? 4'h7 : _GEN_33973; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33975 = 10'hf6 == _T_509[9:0] ? 4'h3 : _GEN_33974; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33976 = 10'hf7 == _T_509[9:0] ? 4'h3 : _GEN_33975; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33977 = 10'hf8 == _T_509[9:0] ? 4'h3 : _GEN_33976; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33978 = 10'hf9 == _T_509[9:0] ? 4'h3 : _GEN_33977; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33979 = 10'hfa == _T_509[9:0] ? 4'h3 : _GEN_33978; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33980 = 10'hfb == _T_509[9:0] ? 4'h3 : _GEN_33979; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33981 = 10'hfc == _T_509[9:0] ? 4'h3 : _GEN_33980; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33982 = 10'hfd == _T_509[9:0] ? 4'h3 : _GEN_33981; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33983 = 10'hfe == _T_509[9:0] ? 4'h3 : _GEN_33982; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33984 = 10'hff == _T_509[9:0] ? 4'h3 : _GEN_33983; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33985 = 10'h100 == _T_509[9:0] ? 4'h3 : _GEN_33984; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33986 = 10'h101 == _T_509[9:0] ? 4'h4 : _GEN_33985; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33987 = 10'h102 == _T_509[9:0] ? 4'h6 : _GEN_33986; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33988 = 10'h103 == _T_509[9:0] ? 4'ha : _GEN_33987; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33989 = 10'h104 == _T_509[9:0] ? 4'ha : _GEN_33988; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33990 = 10'h105 == _T_509[9:0] ? 4'h9 : _GEN_33989; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33991 = 10'h106 == _T_509[9:0] ? 4'h9 : _GEN_33990; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33992 = 10'h107 == _T_509[9:0] ? 4'h9 : _GEN_33991; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33993 = 10'h108 == _T_509[9:0] ? 4'h9 : _GEN_33992; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33994 = 10'h109 == _T_509[9:0] ? 4'h3 : _GEN_33993; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33995 = 10'h10a == _T_509[9:0] ? 4'ha : _GEN_33994; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33996 = 10'h10b == _T_509[9:0] ? 4'ha : _GEN_33995; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33997 = 10'h10c == _T_509[9:0] ? 4'ha : _GEN_33996; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33998 = 10'h10d == _T_509[9:0] ? 4'ha : _GEN_33997; // @[Filter.scala 230:62]
  wire [3:0] _GEN_33999 = 10'h10e == _T_509[9:0] ? 4'ha : _GEN_33998; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34000 = 10'h10f == _T_509[9:0] ? 4'h9 : _GEN_33999; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34001 = 10'h110 == _T_509[9:0] ? 4'h9 : _GEN_34000; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34002 = 10'h111 == _T_509[9:0] ? 4'h4 : _GEN_34001; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34003 = 10'h112 == _T_509[9:0] ? 4'h8 : _GEN_34002; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34004 = 10'h113 == _T_509[9:0] ? 4'h3 : _GEN_34003; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34005 = 10'h114 == _T_509[9:0] ? 4'h3 : _GEN_34004; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34006 = 10'h115 == _T_509[9:0] ? 4'h4 : _GEN_34005; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34007 = 10'h116 == _T_509[9:0] ? 4'h4 : _GEN_34006; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34008 = 10'h117 == _T_509[9:0] ? 4'h3 : _GEN_34007; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34009 = 10'h118 == _T_509[9:0] ? 4'h8 : _GEN_34008; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34010 = 10'h119 == _T_509[9:0] ? 4'ha : _GEN_34009; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34011 = 10'h11a == _T_509[9:0] ? 4'ha : _GEN_34010; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34012 = 10'h11b == _T_509[9:0] ? 4'ha : _GEN_34011; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34013 = 10'h11c == _T_509[9:0] ? 4'h6 : _GEN_34012; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34014 = 10'h11d == _T_509[9:0] ? 4'h3 : _GEN_34013; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34015 = 10'h11e == _T_509[9:0] ? 4'h3 : _GEN_34014; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34016 = 10'h11f == _T_509[9:0] ? 4'h3 : _GEN_34015; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34017 = 10'h120 == _T_509[9:0] ? 4'h3 : _GEN_34016; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34018 = 10'h121 == _T_509[9:0] ? 4'h3 : _GEN_34017; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34019 = 10'h122 == _T_509[9:0] ? 4'h3 : _GEN_34018; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34020 = 10'h123 == _T_509[9:0] ? 4'h3 : _GEN_34019; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34021 = 10'h124 == _T_509[9:0] ? 4'h3 : _GEN_34020; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34022 = 10'h125 == _T_509[9:0] ? 4'h3 : _GEN_34021; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34023 = 10'h126 == _T_509[9:0] ? 4'h4 : _GEN_34022; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34024 = 10'h127 == _T_509[9:0] ? 4'h6 : _GEN_34023; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34025 = 10'h128 == _T_509[9:0] ? 4'h5 : _GEN_34024; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34026 = 10'h129 == _T_509[9:0] ? 4'h8 : _GEN_34025; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34027 = 10'h12a == _T_509[9:0] ? 4'h5 : _GEN_34026; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34028 = 10'h12b == _T_509[9:0] ? 4'h3 : _GEN_34027; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34029 = 10'h12c == _T_509[9:0] ? 4'h3 : _GEN_34028; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34030 = 10'h12d == _T_509[9:0] ? 4'h3 : _GEN_34029; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34031 = 10'h12e == _T_509[9:0] ? 4'h4 : _GEN_34030; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34032 = 10'h12f == _T_509[9:0] ? 4'h4 : _GEN_34031; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34033 = 10'h130 == _T_509[9:0] ? 4'ha : _GEN_34032; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34034 = 10'h131 == _T_509[9:0] ? 4'h9 : _GEN_34033; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34035 = 10'h132 == _T_509[9:0] ? 4'h9 : _GEN_34034; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34036 = 10'h133 == _T_509[9:0] ? 4'h8 : _GEN_34035; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34037 = 10'h134 == _T_509[9:0] ? 4'h9 : _GEN_34036; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34038 = 10'h135 == _T_509[9:0] ? 4'h8 : _GEN_34037; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34039 = 10'h136 == _T_509[9:0] ? 4'h7 : _GEN_34038; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34040 = 10'h137 == _T_509[9:0] ? 4'h6 : _GEN_34039; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34041 = 10'h138 == _T_509[9:0] ? 4'h8 : _GEN_34040; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34042 = 10'h139 == _T_509[9:0] ? 4'h3 : _GEN_34041; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34043 = 10'h13a == _T_509[9:0] ? 4'h3 : _GEN_34042; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34044 = 10'h13b == _T_509[9:0] ? 4'h4 : _GEN_34043; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34045 = 10'h13c == _T_509[9:0] ? 4'h4 : _GEN_34044; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34046 = 10'h13d == _T_509[9:0] ? 4'h3 : _GEN_34045; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34047 = 10'h13e == _T_509[9:0] ? 4'h5 : _GEN_34046; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34048 = 10'h13f == _T_509[9:0] ? 4'h9 : _GEN_34047; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34049 = 10'h140 == _T_509[9:0] ? 4'ha : _GEN_34048; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34050 = 10'h141 == _T_509[9:0] ? 4'ha : _GEN_34049; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34051 = 10'h142 == _T_509[9:0] ? 4'ha : _GEN_34050; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34052 = 10'h143 == _T_509[9:0] ? 4'h5 : _GEN_34051; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34053 = 10'h144 == _T_509[9:0] ? 4'h3 : _GEN_34052; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34054 = 10'h145 == _T_509[9:0] ? 4'h3 : _GEN_34053; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34055 = 10'h146 == _T_509[9:0] ? 4'h3 : _GEN_34054; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34056 = 10'h147 == _T_509[9:0] ? 4'h4 : _GEN_34055; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34057 = 10'h148 == _T_509[9:0] ? 4'h3 : _GEN_34056; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34058 = 10'h149 == _T_509[9:0] ? 4'h3 : _GEN_34057; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34059 = 10'h14a == _T_509[9:0] ? 4'h3 : _GEN_34058; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34060 = 10'h14b == _T_509[9:0] ? 4'h6 : _GEN_34059; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34061 = 10'h14c == _T_509[9:0] ? 4'h8 : _GEN_34060; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34062 = 10'h14d == _T_509[9:0] ? 4'h5 : _GEN_34061; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34063 = 10'h14e == _T_509[9:0] ? 4'h4 : _GEN_34062; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34064 = 10'h14f == _T_509[9:0] ? 4'h3 : _GEN_34063; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34065 = 10'h150 == _T_509[9:0] ? 4'h3 : _GEN_34064; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34066 = 10'h151 == _T_509[9:0] ? 4'h3 : _GEN_34065; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34067 = 10'h152 == _T_509[9:0] ? 4'h3 : _GEN_34066; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34068 = 10'h153 == _T_509[9:0] ? 4'h3 : _GEN_34067; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34069 = 10'h154 == _T_509[9:0] ? 4'h3 : _GEN_34068; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34070 = 10'h155 == _T_509[9:0] ? 4'h4 : _GEN_34069; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34071 = 10'h156 == _T_509[9:0] ? 4'h9 : _GEN_34070; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34072 = 10'h157 == _T_509[9:0] ? 4'h8 : _GEN_34071; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34073 = 10'h158 == _T_509[9:0] ? 4'h8 : _GEN_34072; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34074 = 10'h159 == _T_509[9:0] ? 4'h8 : _GEN_34073; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34075 = 10'h15a == _T_509[9:0] ? 4'h8 : _GEN_34074; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34076 = 10'h15b == _T_509[9:0] ? 4'h8 : _GEN_34075; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34077 = 10'h15c == _T_509[9:0] ? 4'h7 : _GEN_34076; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34078 = 10'h15d == _T_509[9:0] ? 4'h7 : _GEN_34077; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34079 = 10'h15e == _T_509[9:0] ? 4'h8 : _GEN_34078; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34080 = 10'h15f == _T_509[9:0] ? 4'h3 : _GEN_34079; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34081 = 10'h160 == _T_509[9:0] ? 4'h4 : _GEN_34080; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34082 = 10'h161 == _T_509[9:0] ? 4'h4 : _GEN_34081; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34083 = 10'h162 == _T_509[9:0] ? 4'h4 : _GEN_34082; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34084 = 10'h163 == _T_509[9:0] ? 4'h4 : _GEN_34083; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34085 = 10'h164 == _T_509[9:0] ? 4'h5 : _GEN_34084; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34086 = 10'h165 == _T_509[9:0] ? 4'ha : _GEN_34085; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34087 = 10'h166 == _T_509[9:0] ? 4'h9 : _GEN_34086; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34088 = 10'h167 == _T_509[9:0] ? 4'ha : _GEN_34087; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34089 = 10'h168 == _T_509[9:0] ? 4'ha : _GEN_34088; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34090 = 10'h169 == _T_509[9:0] ? 4'h6 : _GEN_34089; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34091 = 10'h16a == _T_509[9:0] ? 4'h3 : _GEN_34090; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34092 = 10'h16b == _T_509[9:0] ? 4'h3 : _GEN_34091; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34093 = 10'h16c == _T_509[9:0] ? 4'h3 : _GEN_34092; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34094 = 10'h16d == _T_509[9:0] ? 4'h4 : _GEN_34093; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34095 = 10'h16e == _T_509[9:0] ? 4'h3 : _GEN_34094; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34096 = 10'h16f == _T_509[9:0] ? 4'h3 : _GEN_34095; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34097 = 10'h170 == _T_509[9:0] ? 4'h3 : _GEN_34096; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34098 = 10'h171 == _T_509[9:0] ? 4'h7 : _GEN_34097; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34099 = 10'h172 == _T_509[9:0] ? 4'ha : _GEN_34098; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34100 = 10'h173 == _T_509[9:0] ? 4'h5 : _GEN_34099; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34101 = 10'h174 == _T_509[9:0] ? 4'h3 : _GEN_34100; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34102 = 10'h175 == _T_509[9:0] ? 4'h4 : _GEN_34101; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34103 = 10'h176 == _T_509[9:0] ? 4'h4 : _GEN_34102; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34104 = 10'h177 == _T_509[9:0] ? 4'h4 : _GEN_34103; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34105 = 10'h178 == _T_509[9:0] ? 4'h4 : _GEN_34104; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34106 = 10'h179 == _T_509[9:0] ? 4'h3 : _GEN_34105; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34107 = 10'h17a == _T_509[9:0] ? 4'h3 : _GEN_34106; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34108 = 10'h17b == _T_509[9:0] ? 4'h3 : _GEN_34107; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34109 = 10'h17c == _T_509[9:0] ? 4'h8 : _GEN_34108; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34110 = 10'h17d == _T_509[9:0] ? 4'h8 : _GEN_34109; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34111 = 10'h17e == _T_509[9:0] ? 4'h8 : _GEN_34110; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34112 = 10'h17f == _T_509[9:0] ? 4'h8 : _GEN_34111; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34113 = 10'h180 == _T_509[9:0] ? 4'h8 : _GEN_34112; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34114 = 10'h181 == _T_509[9:0] ? 4'h8 : _GEN_34113; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34115 = 10'h182 == _T_509[9:0] ? 4'h8 : _GEN_34114; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34116 = 10'h183 == _T_509[9:0] ? 4'h8 : _GEN_34115; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34117 = 10'h184 == _T_509[9:0] ? 4'h8 : _GEN_34116; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34118 = 10'h185 == _T_509[9:0] ? 4'h5 : _GEN_34117; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34119 = 10'h186 == _T_509[9:0] ? 4'h3 : _GEN_34118; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34120 = 10'h187 == _T_509[9:0] ? 4'h4 : _GEN_34119; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34121 = 10'h188 == _T_509[9:0] ? 4'h4 : _GEN_34120; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34122 = 10'h189 == _T_509[9:0] ? 4'h4 : _GEN_34121; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34123 = 10'h18a == _T_509[9:0] ? 4'h5 : _GEN_34122; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34124 = 10'h18b == _T_509[9:0] ? 4'ha : _GEN_34123; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34125 = 10'h18c == _T_509[9:0] ? 4'ha : _GEN_34124; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34126 = 10'h18d == _T_509[9:0] ? 4'h9 : _GEN_34125; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34127 = 10'h18e == _T_509[9:0] ? 4'ha : _GEN_34126; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34128 = 10'h18f == _T_509[9:0] ? 4'h4 : _GEN_34127; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34129 = 10'h190 == _T_509[9:0] ? 4'h3 : _GEN_34128; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34130 = 10'h191 == _T_509[9:0] ? 4'h3 : _GEN_34129; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34131 = 10'h192 == _T_509[9:0] ? 4'h5 : _GEN_34130; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34132 = 10'h193 == _T_509[9:0] ? 4'h6 : _GEN_34131; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34133 = 10'h194 == _T_509[9:0] ? 4'h5 : _GEN_34132; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34134 = 10'h195 == _T_509[9:0] ? 4'h3 : _GEN_34133; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34135 = 10'h196 == _T_509[9:0] ? 4'h3 : _GEN_34134; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34136 = 10'h197 == _T_509[9:0] ? 4'h5 : _GEN_34135; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34137 = 10'h198 == _T_509[9:0] ? 4'ha : _GEN_34136; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34138 = 10'h199 == _T_509[9:0] ? 4'h3 : _GEN_34137; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34139 = 10'h19a == _T_509[9:0] ? 4'h1 : _GEN_34138; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34140 = 10'h19b == _T_509[9:0] ? 4'h2 : _GEN_34139; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34141 = 10'h19c == _T_509[9:0] ? 4'h4 : _GEN_34140; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34142 = 10'h19d == _T_509[9:0] ? 4'h3 : _GEN_34141; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34143 = 10'h19e == _T_509[9:0] ? 4'h1 : _GEN_34142; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34144 = 10'h19f == _T_509[9:0] ? 4'h2 : _GEN_34143; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34145 = 10'h1a0 == _T_509[9:0] ? 4'h3 : _GEN_34144; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34146 = 10'h1a1 == _T_509[9:0] ? 4'h4 : _GEN_34145; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34147 = 10'h1a2 == _T_509[9:0] ? 4'h8 : _GEN_34146; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34148 = 10'h1a3 == _T_509[9:0] ? 4'h8 : _GEN_34147; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34149 = 10'h1a4 == _T_509[9:0] ? 4'h8 : _GEN_34148; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34150 = 10'h1a5 == _T_509[9:0] ? 4'h8 : _GEN_34149; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34151 = 10'h1a6 == _T_509[9:0] ? 4'h7 : _GEN_34150; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34152 = 10'h1a7 == _T_509[9:0] ? 4'h8 : _GEN_34151; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34153 = 10'h1a8 == _T_509[9:0] ? 4'h8 : _GEN_34152; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34154 = 10'h1a9 == _T_509[9:0] ? 4'h8 : _GEN_34153; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34155 = 10'h1aa == _T_509[9:0] ? 4'h7 : _GEN_34154; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34156 = 10'h1ab == _T_509[9:0] ? 4'h4 : _GEN_34155; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34157 = 10'h1ac == _T_509[9:0] ? 4'h4 : _GEN_34156; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34158 = 10'h1ad == _T_509[9:0] ? 4'h3 : _GEN_34157; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34159 = 10'h1ae == _T_509[9:0] ? 4'h3 : _GEN_34158; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34160 = 10'h1af == _T_509[9:0] ? 4'h4 : _GEN_34159; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34161 = 10'h1b0 == _T_509[9:0] ? 4'h6 : _GEN_34160; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34162 = 10'h1b1 == _T_509[9:0] ? 4'ha : _GEN_34161; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34163 = 10'h1b2 == _T_509[9:0] ? 4'ha : _GEN_34162; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34164 = 10'h1b3 == _T_509[9:0] ? 4'h9 : _GEN_34163; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34165 = 10'h1b4 == _T_509[9:0] ? 4'h9 : _GEN_34164; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34166 = 10'h1b5 == _T_509[9:0] ? 4'h3 : _GEN_34165; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34167 = 10'h1b6 == _T_509[9:0] ? 4'h3 : _GEN_34166; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34168 = 10'h1b7 == _T_509[9:0] ? 4'h4 : _GEN_34167; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34169 = 10'h1b8 == _T_509[9:0] ? 4'h5 : _GEN_34168; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34170 = 10'h1b9 == _T_509[9:0] ? 4'h6 : _GEN_34169; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34171 = 10'h1ba == _T_509[9:0] ? 4'h4 : _GEN_34170; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34172 = 10'h1bb == _T_509[9:0] ? 4'h3 : _GEN_34171; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34173 = 10'h1bc == _T_509[9:0] ? 4'h3 : _GEN_34172; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34174 = 10'h1bd == _T_509[9:0] ? 4'h4 : _GEN_34173; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34175 = 10'h1be == _T_509[9:0] ? 4'ha : _GEN_34174; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34176 = 10'h1bf == _T_509[9:0] ? 4'h4 : _GEN_34175; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34177 = 10'h1c0 == _T_509[9:0] ? 4'h5 : _GEN_34176; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34178 = 10'h1c1 == _T_509[9:0] ? 4'h5 : _GEN_34177; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34179 = 10'h1c2 == _T_509[9:0] ? 4'h4 : _GEN_34178; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34180 = 10'h1c3 == _T_509[9:0] ? 4'h5 : _GEN_34179; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34181 = 10'h1c4 == _T_509[9:0] ? 4'h4 : _GEN_34180; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34182 = 10'h1c5 == _T_509[9:0] ? 4'h3 : _GEN_34181; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34183 = 10'h1c6 == _T_509[9:0] ? 4'h4 : _GEN_34182; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34184 = 10'h1c7 == _T_509[9:0] ? 4'h3 : _GEN_34183; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34185 = 10'h1c8 == _T_509[9:0] ? 4'h8 : _GEN_34184; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34186 = 10'h1c9 == _T_509[9:0] ? 4'h8 : _GEN_34185; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34187 = 10'h1ca == _T_509[9:0] ? 4'h8 : _GEN_34186; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34188 = 10'h1cb == _T_509[9:0] ? 4'h8 : _GEN_34187; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34189 = 10'h1cc == _T_509[9:0] ? 4'h8 : _GEN_34188; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34190 = 10'h1cd == _T_509[9:0] ? 4'h8 : _GEN_34189; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34191 = 10'h1ce == _T_509[9:0] ? 4'h8 : _GEN_34190; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34192 = 10'h1cf == _T_509[9:0] ? 4'h8 : _GEN_34191; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34193 = 10'h1d0 == _T_509[9:0] ? 4'h5 : _GEN_34192; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34194 = 10'h1d1 == _T_509[9:0] ? 4'h4 : _GEN_34193; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34195 = 10'h1d2 == _T_509[9:0] ? 4'h6 : _GEN_34194; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34196 = 10'h1d3 == _T_509[9:0] ? 4'h6 : _GEN_34195; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34197 = 10'h1d4 == _T_509[9:0] ? 4'h6 : _GEN_34196; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34198 = 10'h1d5 == _T_509[9:0] ? 4'h5 : _GEN_34197; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34199 = 10'h1d6 == _T_509[9:0] ? 4'h8 : _GEN_34198; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34200 = 10'h1d7 == _T_509[9:0] ? 4'ha : _GEN_34199; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34201 = 10'h1d8 == _T_509[9:0] ? 4'ha : _GEN_34200; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34202 = 10'h1d9 == _T_509[9:0] ? 4'ha : _GEN_34201; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34203 = 10'h1da == _T_509[9:0] ? 4'h6 : _GEN_34202; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34204 = 10'h1db == _T_509[9:0] ? 4'h3 : _GEN_34203; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34205 = 10'h1dc == _T_509[9:0] ? 4'h5 : _GEN_34204; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34206 = 10'h1dd == _T_509[9:0] ? 4'h2 : _GEN_34205; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34207 = 10'h1de == _T_509[9:0] ? 4'h5 : _GEN_34206; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34208 = 10'h1df == _T_509[9:0] ? 4'h5 : _GEN_34207; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34209 = 10'h1e0 == _T_509[9:0] ? 4'h5 : _GEN_34208; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34210 = 10'h1e1 == _T_509[9:0] ? 4'h3 : _GEN_34209; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34211 = 10'h1e2 == _T_509[9:0] ? 4'h3 : _GEN_34210; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34212 = 10'h1e3 == _T_509[9:0] ? 4'h3 : _GEN_34211; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34213 = 10'h1e4 == _T_509[9:0] ? 4'h9 : _GEN_34212; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34214 = 10'h1e5 == _T_509[9:0] ? 4'h4 : _GEN_34213; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34215 = 10'h1e6 == _T_509[9:0] ? 4'h4 : _GEN_34214; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34216 = 10'h1e7 == _T_509[9:0] ? 4'h4 : _GEN_34215; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34217 = 10'h1e8 == _T_509[9:0] ? 4'h4 : _GEN_34216; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34218 = 10'h1e9 == _T_509[9:0] ? 4'h4 : _GEN_34217; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34219 = 10'h1ea == _T_509[9:0] ? 4'h4 : _GEN_34218; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34220 = 10'h1eb == _T_509[9:0] ? 4'h4 : _GEN_34219; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34221 = 10'h1ec == _T_509[9:0] ? 4'h4 : _GEN_34220; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34222 = 10'h1ed == _T_509[9:0] ? 4'h4 : _GEN_34221; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34223 = 10'h1ee == _T_509[9:0] ? 4'h8 : _GEN_34222; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34224 = 10'h1ef == _T_509[9:0] ? 4'h8 : _GEN_34223; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34225 = 10'h1f0 == _T_509[9:0] ? 4'h8 : _GEN_34224; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34226 = 10'h1f1 == _T_509[9:0] ? 4'h8 : _GEN_34225; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34227 = 10'h1f2 == _T_509[9:0] ? 4'h8 : _GEN_34226; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34228 = 10'h1f3 == _T_509[9:0] ? 4'h8 : _GEN_34227; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34229 = 10'h1f4 == _T_509[9:0] ? 4'h9 : _GEN_34228; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34230 = 10'h1f5 == _T_509[9:0] ? 4'h9 : _GEN_34229; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34231 = 10'h1f6 == _T_509[9:0] ? 4'ha : _GEN_34230; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34232 = 10'h1f7 == _T_509[9:0] ? 4'h5 : _GEN_34231; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34233 = 10'h1f8 == _T_509[9:0] ? 4'h5 : _GEN_34232; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34234 = 10'h1f9 == _T_509[9:0] ? 4'h7 : _GEN_34233; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34235 = 10'h1fa == _T_509[9:0] ? 4'h7 : _GEN_34234; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34236 = 10'h1fb == _T_509[9:0] ? 4'h5 : _GEN_34235; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34237 = 10'h1fc == _T_509[9:0] ? 4'ha : _GEN_34236; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34238 = 10'h1fd == _T_509[9:0] ? 4'hb : _GEN_34237; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34239 = 10'h1fe == _T_509[9:0] ? 4'hb : _GEN_34238; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34240 = 10'h1ff == _T_509[9:0] ? 4'ha : _GEN_34239; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34241 = 10'h200 == _T_509[9:0] ? 4'h4 : _GEN_34240; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34242 = 10'h201 == _T_509[9:0] ? 4'h3 : _GEN_34241; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34243 = 10'h202 == _T_509[9:0] ? 4'h2 : _GEN_34242; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34244 = 10'h203 == _T_509[9:0] ? 4'h2 : _GEN_34243; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34245 = 10'h204 == _T_509[9:0] ? 4'h2 : _GEN_34244; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34246 = 10'h205 == _T_509[9:0] ? 4'h2 : _GEN_34245; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34247 = 10'h206 == _T_509[9:0] ? 4'h2 : _GEN_34246; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34248 = 10'h207 == _T_509[9:0] ? 4'h2 : _GEN_34247; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34249 = 10'h208 == _T_509[9:0] ? 4'h3 : _GEN_34248; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34250 = 10'h209 == _T_509[9:0] ? 4'h3 : _GEN_34249; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34251 = 10'h20a == _T_509[9:0] ? 4'h8 : _GEN_34250; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34252 = 10'h20b == _T_509[9:0] ? 4'h4 : _GEN_34251; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34253 = 10'h20c == _T_509[9:0] ? 4'h4 : _GEN_34252; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34254 = 10'h20d == _T_509[9:0] ? 4'h4 : _GEN_34253; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34255 = 10'h20e == _T_509[9:0] ? 4'h4 : _GEN_34254; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34256 = 10'h20f == _T_509[9:0] ? 4'h4 : _GEN_34255; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34257 = 10'h210 == _T_509[9:0] ? 4'h4 : _GEN_34256; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34258 = 10'h211 == _T_509[9:0] ? 4'h4 : _GEN_34257; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34259 = 10'h212 == _T_509[9:0] ? 4'h4 : _GEN_34258; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34260 = 10'h213 == _T_509[9:0] ? 4'h6 : _GEN_34259; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34261 = 10'h214 == _T_509[9:0] ? 4'h7 : _GEN_34260; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34262 = 10'h215 == _T_509[9:0] ? 4'h8 : _GEN_34261; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34263 = 10'h216 == _T_509[9:0] ? 4'h8 : _GEN_34262; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34264 = 10'h217 == _T_509[9:0] ? 4'h8 : _GEN_34263; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34265 = 10'h218 == _T_509[9:0] ? 4'h8 : _GEN_34264; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34266 = 10'h219 == _T_509[9:0] ? 4'h8 : _GEN_34265; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34267 = 10'h21a == _T_509[9:0] ? 4'h8 : _GEN_34266; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34268 = 10'h21b == _T_509[9:0] ? 4'h8 : _GEN_34267; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34269 = 10'h21c == _T_509[9:0] ? 4'ha : _GEN_34268; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34270 = 10'h21d == _T_509[9:0] ? 4'h9 : _GEN_34269; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34271 = 10'h21e == _T_509[9:0] ? 4'h6 : _GEN_34270; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34272 = 10'h21f == _T_509[9:0] ? 4'h4 : _GEN_34271; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34273 = 10'h220 == _T_509[9:0] ? 4'h4 : _GEN_34272; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34274 = 10'h221 == _T_509[9:0] ? 4'h5 : _GEN_34273; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34275 = 10'h222 == _T_509[9:0] ? 4'ha : _GEN_34274; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34276 = 10'h223 == _T_509[9:0] ? 4'ha : _GEN_34275; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34277 = 10'h224 == _T_509[9:0] ? 4'ha : _GEN_34276; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34278 = 10'h225 == _T_509[9:0] ? 4'h8 : _GEN_34277; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34279 = 10'h226 == _T_509[9:0] ? 4'h4 : _GEN_34278; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34280 = 10'h227 == _T_509[9:0] ? 4'h2 : _GEN_34279; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34281 = 10'h228 == _T_509[9:0] ? 4'h2 : _GEN_34280; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34282 = 10'h229 == _T_509[9:0] ? 4'h2 : _GEN_34281; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34283 = 10'h22a == _T_509[9:0] ? 4'h2 : _GEN_34282; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34284 = 10'h22b == _T_509[9:0] ? 4'h2 : _GEN_34283; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34285 = 10'h22c == _T_509[9:0] ? 4'h2 : _GEN_34284; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34286 = 10'h22d == _T_509[9:0] ? 4'h2 : _GEN_34285; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34287 = 10'h22e == _T_509[9:0] ? 4'h2 : _GEN_34286; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34288 = 10'h22f == _T_509[9:0] ? 4'h3 : _GEN_34287; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34289 = 10'h230 == _T_509[9:0] ? 4'h3 : _GEN_34288; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34290 = 10'h231 == _T_509[9:0] ? 4'h3 : _GEN_34289; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34291 = 10'h232 == _T_509[9:0] ? 4'h4 : _GEN_34290; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34292 = 10'h233 == _T_509[9:0] ? 4'h6 : _GEN_34291; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34293 = 10'h234 == _T_509[9:0] ? 4'h6 : _GEN_34292; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34294 = 10'h235 == _T_509[9:0] ? 4'h4 : _GEN_34293; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34295 = 10'h236 == _T_509[9:0] ? 4'h4 : _GEN_34294; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34296 = 10'h237 == _T_509[9:0] ? 4'h4 : _GEN_34295; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34297 = 10'h238 == _T_509[9:0] ? 4'h4 : _GEN_34296; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34298 = 10'h239 == _T_509[9:0] ? 4'h3 : _GEN_34297; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34299 = 10'h23a == _T_509[9:0] ? 4'h7 : _GEN_34298; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34300 = 10'h23b == _T_509[9:0] ? 4'h7 : _GEN_34299; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34301 = 10'h23c == _T_509[9:0] ? 4'h7 : _GEN_34300; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34302 = 10'h23d == _T_509[9:0] ? 4'h7 : _GEN_34301; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34303 = 10'h23e == _T_509[9:0] ? 4'h7 : _GEN_34302; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34304 = 10'h23f == _T_509[9:0] ? 4'h7 : _GEN_34303; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34305 = 10'h240 == _T_509[9:0] ? 4'h7 : _GEN_34304; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34306 = 10'h241 == _T_509[9:0] ? 4'h8 : _GEN_34305; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34307 = 10'h242 == _T_509[9:0] ? 4'ha : _GEN_34306; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34308 = 10'h243 == _T_509[9:0] ? 4'ha : _GEN_34307; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34309 = 10'h244 == _T_509[9:0] ? 4'ha : _GEN_34308; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34310 = 10'h245 == _T_509[9:0] ? 4'h8 : _GEN_34309; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34311 = 10'h246 == _T_509[9:0] ? 4'h7 : _GEN_34310; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34312 = 10'h247 == _T_509[9:0] ? 4'h8 : _GEN_34311; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34313 = 10'h248 == _T_509[9:0] ? 4'ha : _GEN_34312; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34314 = 10'h249 == _T_509[9:0] ? 4'ha : _GEN_34313; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34315 = 10'h24a == _T_509[9:0] ? 4'ha : _GEN_34314; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34316 = 10'h24b == _T_509[9:0] ? 4'h4 : _GEN_34315; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34317 = 10'h24c == _T_509[9:0] ? 4'h4 : _GEN_34316; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34318 = 10'h24d == _T_509[9:0] ? 4'h2 : _GEN_34317; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34319 = 10'h24e == _T_509[9:0] ? 4'h2 : _GEN_34318; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34320 = 10'h24f == _T_509[9:0] ? 4'h2 : _GEN_34319; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34321 = 10'h250 == _T_509[9:0] ? 4'h2 : _GEN_34320; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34322 = 10'h251 == _T_509[9:0] ? 4'h2 : _GEN_34321; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34323 = 10'h252 == _T_509[9:0] ? 4'h2 : _GEN_34322; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34324 = 10'h253 == _T_509[9:0] ? 4'h2 : _GEN_34323; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34325 = 10'h254 == _T_509[9:0] ? 4'h2 : _GEN_34324; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34326 = 10'h255 == _T_509[9:0] ? 4'h3 : _GEN_34325; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34327 = 10'h256 == _T_509[9:0] ? 4'h4 : _GEN_34326; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34328 = 10'h257 == _T_509[9:0] ? 4'h3 : _GEN_34327; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34329 = 10'h258 == _T_509[9:0] ? 4'h4 : _GEN_34328; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34330 = 10'h259 == _T_509[9:0] ? 4'h4 : _GEN_34329; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34331 = 10'h25a == _T_509[9:0] ? 4'h4 : _GEN_34330; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34332 = 10'h25b == _T_509[9:0] ? 4'h3 : _GEN_34331; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34333 = 10'h25c == _T_509[9:0] ? 4'h4 : _GEN_34332; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34334 = 10'h25d == _T_509[9:0] ? 4'h4 : _GEN_34333; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34335 = 10'h25e == _T_509[9:0] ? 4'h3 : _GEN_34334; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34336 = 10'h25f == _T_509[9:0] ? 4'h3 : _GEN_34335; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34337 = 10'h260 == _T_509[9:0] ? 4'h8 : _GEN_34336; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34338 = 10'h261 == _T_509[9:0] ? 4'h7 : _GEN_34337; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34339 = 10'h262 == _T_509[9:0] ? 4'h6 : _GEN_34338; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34340 = 10'h263 == _T_509[9:0] ? 4'h5 : _GEN_34339; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34341 = 10'h264 == _T_509[9:0] ? 4'h6 : _GEN_34340; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34342 = 10'h265 == _T_509[9:0] ? 4'h5 : _GEN_34341; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34343 = 10'h266 == _T_509[9:0] ? 4'h5 : _GEN_34342; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34344 = 10'h267 == _T_509[9:0] ? 4'h7 : _GEN_34343; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34345 = 10'h268 == _T_509[9:0] ? 4'ha : _GEN_34344; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34346 = 10'h269 == _T_509[9:0] ? 4'ha : _GEN_34345; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34347 = 10'h26a == _T_509[9:0] ? 4'ha : _GEN_34346; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34348 = 10'h26b == _T_509[9:0] ? 4'ha : _GEN_34347; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34349 = 10'h26c == _T_509[9:0] ? 4'ha : _GEN_34348; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34350 = 10'h26d == _T_509[9:0] ? 4'ha : _GEN_34349; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34351 = 10'h26e == _T_509[9:0] ? 4'ha : _GEN_34350; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34352 = 10'h26f == _T_509[9:0] ? 4'ha : _GEN_34351; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34353 = 10'h270 == _T_509[9:0] ? 4'h5 : _GEN_34352; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34354 = 10'h271 == _T_509[9:0] ? 4'h4 : _GEN_34353; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34355 = 10'h272 == _T_509[9:0] ? 4'h3 : _GEN_34354; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34356 = 10'h273 == _T_509[9:0] ? 4'h2 : _GEN_34355; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34357 = 10'h274 == _T_509[9:0] ? 4'h2 : _GEN_34356; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34358 = 10'h275 == _T_509[9:0] ? 4'h2 : _GEN_34357; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34359 = 10'h276 == _T_509[9:0] ? 4'h2 : _GEN_34358; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34360 = 10'h277 == _T_509[9:0] ? 4'h2 : _GEN_34359; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34361 = 10'h278 == _T_509[9:0] ? 4'h2 : _GEN_34360; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34362 = 10'h279 == _T_509[9:0] ? 4'h2 : _GEN_34361; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34363 = 10'h27a == _T_509[9:0] ? 4'h2 : _GEN_34362; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34364 = 10'h27b == _T_509[9:0] ? 4'h4 : _GEN_34363; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34365 = 10'h27c == _T_509[9:0] ? 4'h3 : _GEN_34364; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34366 = 10'h27d == _T_509[9:0] ? 4'h4 : _GEN_34365; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34367 = 10'h27e == _T_509[9:0] ? 4'h5 : _GEN_34366; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34368 = 10'h27f == _T_509[9:0] ? 4'h4 : _GEN_34367; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34369 = 10'h280 == _T_509[9:0] ? 4'h4 : _GEN_34368; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34370 = 10'h281 == _T_509[9:0] ? 4'h4 : _GEN_34369; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34371 = 10'h282 == _T_509[9:0] ? 4'h4 : _GEN_34370; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34372 = 10'h283 == _T_509[9:0] ? 4'h3 : _GEN_34371; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34373 = 10'h284 == _T_509[9:0] ? 4'h3 : _GEN_34372; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34374 = 10'h285 == _T_509[9:0] ? 4'h3 : _GEN_34373; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34375 = 10'h286 == _T_509[9:0] ? 4'h8 : _GEN_34374; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34376 = 10'h287 == _T_509[9:0] ? 4'h6 : _GEN_34375; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34377 = 10'h288 == _T_509[9:0] ? 4'h6 : _GEN_34376; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34378 = 10'h289 == _T_509[9:0] ? 4'h6 : _GEN_34377; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34379 = 10'h28a == _T_509[9:0] ? 4'h7 : _GEN_34378; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34380 = 10'h28b == _T_509[9:0] ? 4'h7 : _GEN_34379; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34381 = 10'h28c == _T_509[9:0] ? 4'h6 : _GEN_34380; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34382 = 10'h28d == _T_509[9:0] ? 4'h6 : _GEN_34381; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34383 = 10'h28e == _T_509[9:0] ? 4'h4 : _GEN_34382; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34384 = 10'h28f == _T_509[9:0] ? 4'h7 : _GEN_34383; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34385 = 10'h290 == _T_509[9:0] ? 4'h9 : _GEN_34384; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34386 = 10'h291 == _T_509[9:0] ? 4'ha : _GEN_34385; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34387 = 10'h292 == _T_509[9:0] ? 4'ha : _GEN_34386; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34388 = 10'h293 == _T_509[9:0] ? 4'ha : _GEN_34387; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34389 = 10'h294 == _T_509[9:0] ? 4'h9 : _GEN_34388; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34390 = 10'h295 == _T_509[9:0] ? 4'h5 : _GEN_34389; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34391 = 10'h296 == _T_509[9:0] ? 4'h4 : _GEN_34390; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34392 = 10'h297 == _T_509[9:0] ? 4'h4 : _GEN_34391; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34393 = 10'h298 == _T_509[9:0] ? 4'h3 : _GEN_34392; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34394 = 10'h299 == _T_509[9:0] ? 4'h3 : _GEN_34393; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34395 = 10'h29a == _T_509[9:0] ? 4'h2 : _GEN_34394; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34396 = 10'h29b == _T_509[9:0] ? 4'h2 : _GEN_34395; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34397 = 10'h29c == _T_509[9:0] ? 4'h2 : _GEN_34396; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34398 = 10'h29d == _T_509[9:0] ? 4'h2 : _GEN_34397; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34399 = 10'h29e == _T_509[9:0] ? 4'h2 : _GEN_34398; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34400 = 10'h29f == _T_509[9:0] ? 4'h2 : _GEN_34399; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34401 = 10'h2a0 == _T_509[9:0] ? 4'h2 : _GEN_34400; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34402 = 10'h2a1 == _T_509[9:0] ? 4'h4 : _GEN_34401; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34403 = 10'h2a2 == _T_509[9:0] ? 4'h3 : _GEN_34402; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34404 = 10'h2a3 == _T_509[9:0] ? 4'h4 : _GEN_34403; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34405 = 10'h2a4 == _T_509[9:0] ? 4'h5 : _GEN_34404; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34406 = 10'h2a5 == _T_509[9:0] ? 4'h4 : _GEN_34405; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34407 = 10'h2a6 == _T_509[9:0] ? 4'h4 : _GEN_34406; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34408 = 10'h2a7 == _T_509[9:0] ? 4'h4 : _GEN_34407; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34409 = 10'h2a8 == _T_509[9:0] ? 4'h3 : _GEN_34408; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34410 = 10'h2a9 == _T_509[9:0] ? 4'h3 : _GEN_34409; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34411 = 10'h2aa == _T_509[9:0] ? 4'h3 : _GEN_34410; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34412 = 10'h2ab == _T_509[9:0] ? 4'h3 : _GEN_34411; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34413 = 10'h2ac == _T_509[9:0] ? 4'h8 : _GEN_34412; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34414 = 10'h2ad == _T_509[9:0] ? 4'h7 : _GEN_34413; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34415 = 10'h2ae == _T_509[9:0] ? 4'h5 : _GEN_34414; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34416 = 10'h2af == _T_509[9:0] ? 4'h6 : _GEN_34415; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34417 = 10'h2b0 == _T_509[9:0] ? 4'h7 : _GEN_34416; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34418 = 10'h2b1 == _T_509[9:0] ? 4'h6 : _GEN_34417; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34419 = 10'h2b2 == _T_509[9:0] ? 4'h6 : _GEN_34418; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34420 = 10'h2b3 == _T_509[9:0] ? 4'h6 : _GEN_34419; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34421 = 10'h2b4 == _T_509[9:0] ? 4'h3 : _GEN_34420; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34422 = 10'h2b5 == _T_509[9:0] ? 4'h3 : _GEN_34421; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34423 = 10'h2b6 == _T_509[9:0] ? 4'h3 : _GEN_34422; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34424 = 10'h2b7 == _T_509[9:0] ? 4'h4 : _GEN_34423; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34425 = 10'h2b8 == _T_509[9:0] ? 4'h6 : _GEN_34424; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34426 = 10'h2b9 == _T_509[9:0] ? 4'h9 : _GEN_34425; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34427 = 10'h2ba == _T_509[9:0] ? 4'h4 : _GEN_34426; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34428 = 10'h2bb == _T_509[9:0] ? 4'h3 : _GEN_34427; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34429 = 10'h2bc == _T_509[9:0] ? 4'h4 : _GEN_34428; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34430 = 10'h2bd == _T_509[9:0] ? 4'h3 : _GEN_34429; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34431 = 10'h2be == _T_509[9:0] ? 4'h3 : _GEN_34430; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34432 = 10'h2bf == _T_509[9:0] ? 4'h3 : _GEN_34431; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34433 = 10'h2c0 == _T_509[9:0] ? 4'h2 : _GEN_34432; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34434 = 10'h2c1 == _T_509[9:0] ? 4'h2 : _GEN_34433; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34435 = 10'h2c2 == _T_509[9:0] ? 4'h2 : _GEN_34434; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34436 = 10'h2c3 == _T_509[9:0] ? 4'h2 : _GEN_34435; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34437 = 10'h2c4 == _T_509[9:0] ? 4'h2 : _GEN_34436; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34438 = 10'h2c5 == _T_509[9:0] ? 4'h2 : _GEN_34437; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34439 = 10'h2c6 == _T_509[9:0] ? 4'h2 : _GEN_34438; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34440 = 10'h2c7 == _T_509[9:0] ? 4'h4 : _GEN_34439; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34441 = 10'h2c8 == _T_509[9:0] ? 4'h3 : _GEN_34440; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34442 = 10'h2c9 == _T_509[9:0] ? 4'h4 : _GEN_34441; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34443 = 10'h2ca == _T_509[9:0] ? 4'h5 : _GEN_34442; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34444 = 10'h2cb == _T_509[9:0] ? 4'h3 : _GEN_34443; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34445 = 10'h2cc == _T_509[9:0] ? 4'h3 : _GEN_34444; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34446 = 10'h2cd == _T_509[9:0] ? 4'h3 : _GEN_34445; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34447 = 10'h2ce == _T_509[9:0] ? 4'h3 : _GEN_34446; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34448 = 10'h2cf == _T_509[9:0] ? 4'h3 : _GEN_34447; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34449 = 10'h2d0 == _T_509[9:0] ? 4'h3 : _GEN_34448; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34450 = 10'h2d1 == _T_509[9:0] ? 4'h3 : _GEN_34449; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34451 = 10'h2d2 == _T_509[9:0] ? 4'h8 : _GEN_34450; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34452 = 10'h2d3 == _T_509[9:0] ? 4'h6 : _GEN_34451; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34453 = 10'h2d4 == _T_509[9:0] ? 4'h6 : _GEN_34452; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34454 = 10'h2d5 == _T_509[9:0] ? 4'h7 : _GEN_34453; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34455 = 10'h2d6 == _T_509[9:0] ? 4'h7 : _GEN_34454; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34456 = 10'h2d7 == _T_509[9:0] ? 4'h7 : _GEN_34455; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34457 = 10'h2d8 == _T_509[9:0] ? 4'h6 : _GEN_34456; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34458 = 10'h2d9 == _T_509[9:0] ? 4'h7 : _GEN_34457; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34459 = 10'h2da == _T_509[9:0] ? 4'h5 : _GEN_34458; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34460 = 10'h2db == _T_509[9:0] ? 4'h3 : _GEN_34459; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34461 = 10'h2dc == _T_509[9:0] ? 4'h3 : _GEN_34460; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34462 = 10'h2dd == _T_509[9:0] ? 4'h3 : _GEN_34461; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34463 = 10'h2de == _T_509[9:0] ? 4'h3 : _GEN_34462; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34464 = 10'h2df == _T_509[9:0] ? 4'h4 : _GEN_34463; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34465 = 10'h2e0 == _T_509[9:0] ? 4'h3 : _GEN_34464; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34466 = 10'h2e1 == _T_509[9:0] ? 4'h3 : _GEN_34465; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34467 = 10'h2e2 == _T_509[9:0] ? 4'h3 : _GEN_34466; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34468 = 10'h2e3 == _T_509[9:0] ? 4'h3 : _GEN_34467; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34469 = 10'h2e4 == _T_509[9:0] ? 4'h3 : _GEN_34468; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34470 = 10'h2e5 == _T_509[9:0] ? 4'h3 : _GEN_34469; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34471 = 10'h2e6 == _T_509[9:0] ? 4'h2 : _GEN_34470; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34472 = 10'h2e7 == _T_509[9:0] ? 4'h2 : _GEN_34471; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34473 = 10'h2e8 == _T_509[9:0] ? 4'h2 : _GEN_34472; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34474 = 10'h2e9 == _T_509[9:0] ? 4'h2 : _GEN_34473; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34475 = 10'h2ea == _T_509[9:0] ? 4'h2 : _GEN_34474; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34476 = 10'h2eb == _T_509[9:0] ? 4'h2 : _GEN_34475; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34477 = 10'h2ec == _T_509[9:0] ? 4'h3 : _GEN_34476; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34478 = 10'h2ed == _T_509[9:0] ? 4'h4 : _GEN_34477; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34479 = 10'h2ee == _T_509[9:0] ? 4'h3 : _GEN_34478; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34480 = 10'h2ef == _T_509[9:0] ? 4'h3 : _GEN_34479; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34481 = 10'h2f0 == _T_509[9:0] ? 4'h6 : _GEN_34480; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34482 = 10'h2f1 == _T_509[9:0] ? 4'h3 : _GEN_34481; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34483 = 10'h2f2 == _T_509[9:0] ? 4'h3 : _GEN_34482; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34484 = 10'h2f3 == _T_509[9:0] ? 4'h3 : _GEN_34483; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34485 = 10'h2f4 == _T_509[9:0] ? 4'h3 : _GEN_34484; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34486 = 10'h2f5 == _T_509[9:0] ? 4'h3 : _GEN_34485; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34487 = 10'h2f6 == _T_509[9:0] ? 4'h3 : _GEN_34486; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34488 = 10'h2f7 == _T_509[9:0] ? 4'h3 : _GEN_34487; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34489 = 10'h2f8 == _T_509[9:0] ? 4'h8 : _GEN_34488; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34490 = 10'h2f9 == _T_509[9:0] ? 4'h6 : _GEN_34489; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34491 = 10'h2fa == _T_509[9:0] ? 4'h7 : _GEN_34490; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34492 = 10'h2fb == _T_509[9:0] ? 4'h7 : _GEN_34491; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34493 = 10'h2fc == _T_509[9:0] ? 4'h6 : _GEN_34492; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34494 = 10'h2fd == _T_509[9:0] ? 4'h6 : _GEN_34493; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34495 = 10'h2fe == _T_509[9:0] ? 4'h6 : _GEN_34494; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34496 = 10'h2ff == _T_509[9:0] ? 4'h8 : _GEN_34495; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34497 = 10'h300 == _T_509[9:0] ? 4'h9 : _GEN_34496; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34498 = 10'h301 == _T_509[9:0] ? 4'h7 : _GEN_34497; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34499 = 10'h302 == _T_509[9:0] ? 4'h4 : _GEN_34498; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34500 = 10'h303 == _T_509[9:0] ? 4'h4 : _GEN_34499; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34501 = 10'h304 == _T_509[9:0] ? 4'h3 : _GEN_34500; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34502 = 10'h305 == _T_509[9:0] ? 4'h3 : _GEN_34501; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34503 = 10'h306 == _T_509[9:0] ? 4'h3 : _GEN_34502; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34504 = 10'h307 == _T_509[9:0] ? 4'h3 : _GEN_34503; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34505 = 10'h308 == _T_509[9:0] ? 4'h3 : _GEN_34504; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34506 = 10'h309 == _T_509[9:0] ? 4'h3 : _GEN_34505; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34507 = 10'h30a == _T_509[9:0] ? 4'h3 : _GEN_34506; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34508 = 10'h30b == _T_509[9:0] ? 4'h3 : _GEN_34507; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34509 = 10'h30c == _T_509[9:0] ? 4'h2 : _GEN_34508; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34510 = 10'h30d == _T_509[9:0] ? 4'h2 : _GEN_34509; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34511 = 10'h30e == _T_509[9:0] ? 4'h2 : _GEN_34510; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34512 = 10'h30f == _T_509[9:0] ? 4'h2 : _GEN_34511; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34513 = 10'h310 == _T_509[9:0] ? 4'h2 : _GEN_34512; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34514 = 10'h311 == _T_509[9:0] ? 4'h2 : _GEN_34513; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34515 = 10'h312 == _T_509[9:0] ? 4'h3 : _GEN_34514; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34516 = 10'h313 == _T_509[9:0] ? 4'h4 : _GEN_34515; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34517 = 10'h314 == _T_509[9:0] ? 4'h3 : _GEN_34516; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34518 = 10'h315 == _T_509[9:0] ? 4'h3 : _GEN_34517; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34519 = 10'h316 == _T_509[9:0] ? 4'h5 : _GEN_34518; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34520 = 10'h317 == _T_509[9:0] ? 4'h5 : _GEN_34519; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34521 = 10'h318 == _T_509[9:0] ? 4'h3 : _GEN_34520; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34522 = 10'h319 == _T_509[9:0] ? 4'h3 : _GEN_34521; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34523 = 10'h31a == _T_509[9:0] ? 4'h3 : _GEN_34522; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34524 = 10'h31b == _T_509[9:0] ? 4'h3 : _GEN_34523; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34525 = 10'h31c == _T_509[9:0] ? 4'h3 : _GEN_34524; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34526 = 10'h31d == _T_509[9:0] ? 4'h3 : _GEN_34525; // @[Filter.scala 230:62]
  wire [4:0] _GEN_39038 = {{1'd0}, _GEN_34526}; // @[Filter.scala 230:62]
  wire [8:0] _T_511 = _GEN_39038 * 5'h14; // @[Filter.scala 230:62]
  wire [3:0] _GEN_34550 = 10'h17 == _T_509[9:0] ? 4'hb : 4'he; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34551 = 10'h18 == _T_509[9:0] ? 4'hc : _GEN_34550; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34552 = 10'h19 == _T_509[9:0] ? 4'he : _GEN_34551; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34553 = 10'h1a == _T_509[9:0] ? 4'he : _GEN_34552; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34554 = 10'h1b == _T_509[9:0] ? 4'he : _GEN_34553; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34555 = 10'h1c == _T_509[9:0] ? 4'he : _GEN_34554; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34556 = 10'h1d == _T_509[9:0] ? 4'he : _GEN_34555; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34557 = 10'h1e == _T_509[9:0] ? 4'he : _GEN_34556; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34558 = 10'h1f == _T_509[9:0] ? 4'he : _GEN_34557; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34559 = 10'h20 == _T_509[9:0] ? 4'he : _GEN_34558; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34560 = 10'h21 == _T_509[9:0] ? 4'he : _GEN_34559; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34561 = 10'h22 == _T_509[9:0] ? 4'he : _GEN_34560; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34562 = 10'h23 == _T_509[9:0] ? 4'he : _GEN_34561; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34563 = 10'h24 == _T_509[9:0] ? 4'he : _GEN_34562; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34564 = 10'h25 == _T_509[9:0] ? 4'he : _GEN_34563; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34565 = 10'h26 == _T_509[9:0] ? 4'he : _GEN_34564; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34566 = 10'h27 == _T_509[9:0] ? 4'he : _GEN_34565; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34567 = 10'h28 == _T_509[9:0] ? 4'he : _GEN_34566; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34568 = 10'h29 == _T_509[9:0] ? 4'he : _GEN_34567; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34569 = 10'h2a == _T_509[9:0] ? 4'he : _GEN_34568; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34570 = 10'h2b == _T_509[9:0] ? 4'he : _GEN_34569; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34571 = 10'h2c == _T_509[9:0] ? 4'he : _GEN_34570; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34572 = 10'h2d == _T_509[9:0] ? 4'he : _GEN_34571; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34573 = 10'h2e == _T_509[9:0] ? 4'he : _GEN_34572; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34574 = 10'h2f == _T_509[9:0] ? 4'he : _GEN_34573; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34575 = 10'h30 == _T_509[9:0] ? 4'he : _GEN_34574; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34576 = 10'h31 == _T_509[9:0] ? 4'he : _GEN_34575; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34577 = 10'h32 == _T_509[9:0] ? 4'he : _GEN_34576; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34578 = 10'h33 == _T_509[9:0] ? 4'he : _GEN_34577; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34579 = 10'h34 == _T_509[9:0] ? 4'he : _GEN_34578; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34580 = 10'h35 == _T_509[9:0] ? 4'he : _GEN_34579; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34581 = 10'h36 == _T_509[9:0] ? 4'he : _GEN_34580; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34582 = 10'h37 == _T_509[9:0] ? 4'he : _GEN_34581; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34583 = 10'h38 == _T_509[9:0] ? 4'he : _GEN_34582; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34584 = 10'h39 == _T_509[9:0] ? 4'he : _GEN_34583; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34585 = 10'h3a == _T_509[9:0] ? 4'he : _GEN_34584; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34586 = 10'h3b == _T_509[9:0] ? 4'he : _GEN_34585; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34587 = 10'h3c == _T_509[9:0] ? 4'ha : _GEN_34586; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34588 = 10'h3d == _T_509[9:0] ? 4'hc : _GEN_34587; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34589 = 10'h3e == _T_509[9:0] ? 4'hb : _GEN_34588; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34590 = 10'h3f == _T_509[9:0] ? 4'he : _GEN_34589; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34591 = 10'h40 == _T_509[9:0] ? 4'he : _GEN_34590; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34592 = 10'h41 == _T_509[9:0] ? 4'he : _GEN_34591; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34593 = 10'h42 == _T_509[9:0] ? 4'he : _GEN_34592; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34594 = 10'h43 == _T_509[9:0] ? 4'he : _GEN_34593; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34595 = 10'h44 == _T_509[9:0] ? 4'he : _GEN_34594; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34596 = 10'h45 == _T_509[9:0] ? 4'he : _GEN_34595; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34597 = 10'h46 == _T_509[9:0] ? 4'he : _GEN_34596; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34598 = 10'h47 == _T_509[9:0] ? 4'he : _GEN_34597; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34599 = 10'h48 == _T_509[9:0] ? 4'he : _GEN_34598; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34600 = 10'h49 == _T_509[9:0] ? 4'he : _GEN_34599; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34601 = 10'h4a == _T_509[9:0] ? 4'he : _GEN_34600; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34602 = 10'h4b == _T_509[9:0] ? 4'he : _GEN_34601; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34603 = 10'h4c == _T_509[9:0] ? 4'he : _GEN_34602; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34604 = 10'h4d == _T_509[9:0] ? 4'he : _GEN_34603; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34605 = 10'h4e == _T_509[9:0] ? 4'he : _GEN_34604; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34606 = 10'h4f == _T_509[9:0] ? 4'he : _GEN_34605; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34607 = 10'h50 == _T_509[9:0] ? 4'he : _GEN_34606; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34608 = 10'h51 == _T_509[9:0] ? 4'he : _GEN_34607; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34609 = 10'h52 == _T_509[9:0] ? 4'he : _GEN_34608; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34610 = 10'h53 == _T_509[9:0] ? 4'he : _GEN_34609; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34611 = 10'h54 == _T_509[9:0] ? 4'he : _GEN_34610; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34612 = 10'h55 == _T_509[9:0] ? 4'he : _GEN_34611; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34613 = 10'h56 == _T_509[9:0] ? 4'he : _GEN_34612; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34614 = 10'h57 == _T_509[9:0] ? 4'he : _GEN_34613; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34615 = 10'h58 == _T_509[9:0] ? 4'he : _GEN_34614; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34616 = 10'h59 == _T_509[9:0] ? 4'he : _GEN_34615; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34617 = 10'h5a == _T_509[9:0] ? 4'hc : _GEN_34616; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34618 = 10'h5b == _T_509[9:0] ? 4'hd : _GEN_34617; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34619 = 10'h5c == _T_509[9:0] ? 4'he : _GEN_34618; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34620 = 10'h5d == _T_509[9:0] ? 4'he : _GEN_34619; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34621 = 10'h5e == _T_509[9:0] ? 4'he : _GEN_34620; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34622 = 10'h5f == _T_509[9:0] ? 4'he : _GEN_34621; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34623 = 10'h60 == _T_509[9:0] ? 4'he : _GEN_34622; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34624 = 10'h61 == _T_509[9:0] ? 4'hd : _GEN_34623; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34625 = 10'h62 == _T_509[9:0] ? 4'hb : _GEN_34624; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34626 = 10'h63 == _T_509[9:0] ? 4'hc : _GEN_34625; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34627 = 10'h64 == _T_509[9:0] ? 4'ha : _GEN_34626; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34628 = 10'h65 == _T_509[9:0] ? 4'hd : _GEN_34627; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34629 = 10'h66 == _T_509[9:0] ? 4'he : _GEN_34628; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34630 = 10'h67 == _T_509[9:0] ? 4'he : _GEN_34629; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34631 = 10'h68 == _T_509[9:0] ? 4'he : _GEN_34630; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34632 = 10'h69 == _T_509[9:0] ? 4'he : _GEN_34631; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34633 = 10'h6a == _T_509[9:0] ? 4'he : _GEN_34632; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34634 = 10'h6b == _T_509[9:0] ? 4'hd : _GEN_34633; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34635 = 10'h6c == _T_509[9:0] ? 4'hc : _GEN_34634; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34636 = 10'h6d == _T_509[9:0] ? 4'hc : _GEN_34635; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34637 = 10'h6e == _T_509[9:0] ? 4'he : _GEN_34636; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34638 = 10'h6f == _T_509[9:0] ? 4'he : _GEN_34637; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34639 = 10'h70 == _T_509[9:0] ? 4'he : _GEN_34638; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34640 = 10'h71 == _T_509[9:0] ? 4'he : _GEN_34639; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34641 = 10'h72 == _T_509[9:0] ? 4'he : _GEN_34640; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34642 = 10'h73 == _T_509[9:0] ? 4'he : _GEN_34641; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34643 = 10'h74 == _T_509[9:0] ? 4'he : _GEN_34642; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34644 = 10'h75 == _T_509[9:0] ? 4'he : _GEN_34643; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34645 = 10'h76 == _T_509[9:0] ? 4'he : _GEN_34644; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34646 = 10'h77 == _T_509[9:0] ? 4'he : _GEN_34645; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34647 = 10'h78 == _T_509[9:0] ? 4'he : _GEN_34646; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34648 = 10'h79 == _T_509[9:0] ? 4'he : _GEN_34647; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34649 = 10'h7a == _T_509[9:0] ? 4'he : _GEN_34648; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34650 = 10'h7b == _T_509[9:0] ? 4'he : _GEN_34649; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34651 = 10'h7c == _T_509[9:0] ? 4'he : _GEN_34650; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34652 = 10'h7d == _T_509[9:0] ? 4'he : _GEN_34651; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34653 = 10'h7e == _T_509[9:0] ? 4'he : _GEN_34652; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34654 = 10'h7f == _T_509[9:0] ? 4'he : _GEN_34653; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34655 = 10'h80 == _T_509[9:0] ? 4'he : _GEN_34654; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34656 = 10'h81 == _T_509[9:0] ? 4'hb : _GEN_34655; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34657 = 10'h82 == _T_509[9:0] ? 4'hc : _GEN_34656; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34658 = 10'h83 == _T_509[9:0] ? 4'hc : _GEN_34657; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34659 = 10'h84 == _T_509[9:0] ? 4'he : _GEN_34658; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34660 = 10'h85 == _T_509[9:0] ? 4'he : _GEN_34659; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34661 = 10'h86 == _T_509[9:0] ? 4'he : _GEN_34660; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34662 = 10'h87 == _T_509[9:0] ? 4'ha : _GEN_34661; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34663 = 10'h88 == _T_509[9:0] ? 4'hd : _GEN_34662; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34664 = 10'h89 == _T_509[9:0] ? 4'hd : _GEN_34663; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34665 = 10'h8a == _T_509[9:0] ? 4'hc : _GEN_34664; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34666 = 10'h8b == _T_509[9:0] ? 4'he : _GEN_34665; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34667 = 10'h8c == _T_509[9:0] ? 4'he : _GEN_34666; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34668 = 10'h8d == _T_509[9:0] ? 4'he : _GEN_34667; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34669 = 10'h8e == _T_509[9:0] ? 4'he : _GEN_34668; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34670 = 10'h8f == _T_509[9:0] ? 4'hb : _GEN_34669; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34671 = 10'h90 == _T_509[9:0] ? 4'hc : _GEN_34670; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34672 = 10'h91 == _T_509[9:0] ? 4'hc : _GEN_34671; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34673 = 10'h92 == _T_509[9:0] ? 4'hd : _GEN_34672; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34674 = 10'h93 == _T_509[9:0] ? 4'he : _GEN_34673; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34675 = 10'h94 == _T_509[9:0] ? 4'he : _GEN_34674; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34676 = 10'h95 == _T_509[9:0] ? 4'he : _GEN_34675; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34677 = 10'h96 == _T_509[9:0] ? 4'he : _GEN_34676; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34678 = 10'h97 == _T_509[9:0] ? 4'he : _GEN_34677; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34679 = 10'h98 == _T_509[9:0] ? 4'he : _GEN_34678; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34680 = 10'h99 == _T_509[9:0] ? 4'he : _GEN_34679; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34681 = 10'h9a == _T_509[9:0] ? 4'he : _GEN_34680; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34682 = 10'h9b == _T_509[9:0] ? 4'he : _GEN_34681; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34683 = 10'h9c == _T_509[9:0] ? 4'he : _GEN_34682; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34684 = 10'h9d == _T_509[9:0] ? 4'he : _GEN_34683; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34685 = 10'h9e == _T_509[9:0] ? 4'he : _GEN_34684; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34686 = 10'h9f == _T_509[9:0] ? 4'he : _GEN_34685; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34687 = 10'ha0 == _T_509[9:0] ? 4'he : _GEN_34686; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34688 = 10'ha1 == _T_509[9:0] ? 4'he : _GEN_34687; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34689 = 10'ha2 == _T_509[9:0] ? 4'he : _GEN_34688; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34690 = 10'ha3 == _T_509[9:0] ? 4'he : _GEN_34689; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34691 = 10'ha4 == _T_509[9:0] ? 4'he : _GEN_34690; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34692 = 10'ha5 == _T_509[9:0] ? 4'he : _GEN_34691; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34693 = 10'ha6 == _T_509[9:0] ? 4'he : _GEN_34692; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34694 = 10'ha7 == _T_509[9:0] ? 4'he : _GEN_34693; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34695 = 10'ha8 == _T_509[9:0] ? 4'hb : _GEN_34694; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34696 = 10'ha9 == _T_509[9:0] ? 4'hc : _GEN_34695; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34697 = 10'haa == _T_509[9:0] ? 4'hb : _GEN_34696; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34698 = 10'hab == _T_509[9:0] ? 4'hc : _GEN_34697; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34699 = 10'hac == _T_509[9:0] ? 4'hd : _GEN_34698; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34700 = 10'had == _T_509[9:0] ? 4'ha : _GEN_34699; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34701 = 10'hae == _T_509[9:0] ? 4'hd : _GEN_34700; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34702 = 10'haf == _T_509[9:0] ? 4'hd : _GEN_34701; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34703 = 10'hb0 == _T_509[9:0] ? 4'hb : _GEN_34702; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34704 = 10'hb1 == _T_509[9:0] ? 4'hc : _GEN_34703; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34705 = 10'hb2 == _T_509[9:0] ? 4'he : _GEN_34704; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34706 = 10'hb3 == _T_509[9:0] ? 4'hb : _GEN_34705; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34707 = 10'hb4 == _T_509[9:0] ? 4'hc : _GEN_34706; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34708 = 10'hb5 == _T_509[9:0] ? 4'hd : _GEN_34707; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34709 = 10'hb6 == _T_509[9:0] ? 4'hd : _GEN_34708; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34710 = 10'hb7 == _T_509[9:0] ? 4'hc : _GEN_34709; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34711 = 10'hb8 == _T_509[9:0] ? 4'he : _GEN_34710; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34712 = 10'hb9 == _T_509[9:0] ? 4'he : _GEN_34711; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34713 = 10'hba == _T_509[9:0] ? 4'he : _GEN_34712; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34714 = 10'hbb == _T_509[9:0] ? 4'he : _GEN_34713; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34715 = 10'hbc == _T_509[9:0] ? 4'he : _GEN_34714; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34716 = 10'hbd == _T_509[9:0] ? 4'he : _GEN_34715; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34717 = 10'hbe == _T_509[9:0] ? 4'he : _GEN_34716; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34718 = 10'hbf == _T_509[9:0] ? 4'he : _GEN_34717; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34719 = 10'hc0 == _T_509[9:0] ? 4'he : _GEN_34718; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34720 = 10'hc1 == _T_509[9:0] ? 4'he : _GEN_34719; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34721 = 10'hc2 == _T_509[9:0] ? 4'he : _GEN_34720; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34722 = 10'hc3 == _T_509[9:0] ? 4'he : _GEN_34721; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34723 = 10'hc4 == _T_509[9:0] ? 4'he : _GEN_34722; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34724 = 10'hc5 == _T_509[9:0] ? 4'he : _GEN_34723; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34725 = 10'hc6 == _T_509[9:0] ? 4'he : _GEN_34724; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34726 = 10'hc7 == _T_509[9:0] ? 4'hd : _GEN_34725; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34727 = 10'hc8 == _T_509[9:0] ? 4'hb : _GEN_34726; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34728 = 10'hc9 == _T_509[9:0] ? 4'hc : _GEN_34727; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34729 = 10'hca == _T_509[9:0] ? 4'he : _GEN_34728; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34730 = 10'hcb == _T_509[9:0] ? 4'he : _GEN_34729; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34731 = 10'hcc == _T_509[9:0] ? 4'he : _GEN_34730; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34732 = 10'hcd == _T_509[9:0] ? 4'he : _GEN_34731; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34733 = 10'hce == _T_509[9:0] ? 4'hd : _GEN_34732; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34734 = 10'hcf == _T_509[9:0] ? 4'hb : _GEN_34733; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34735 = 10'hd0 == _T_509[9:0] ? 4'hc : _GEN_34734; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34736 = 10'hd1 == _T_509[9:0] ? 4'hc : _GEN_34735; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34737 = 10'hd2 == _T_509[9:0] ? 4'hb : _GEN_34736; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34738 = 10'hd3 == _T_509[9:0] ? 4'hd : _GEN_34737; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34739 = 10'hd4 == _T_509[9:0] ? 4'hd : _GEN_34738; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34740 = 10'hd5 == _T_509[9:0] ? 4'hd : _GEN_34739; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34741 = 10'hd6 == _T_509[9:0] ? 4'hd : _GEN_34740; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34742 = 10'hd7 == _T_509[9:0] ? 4'hc : _GEN_34741; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34743 = 10'hd8 == _T_509[9:0] ? 4'hc : _GEN_34742; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34744 = 10'hd9 == _T_509[9:0] ? 4'hc : _GEN_34743; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34745 = 10'hda == _T_509[9:0] ? 4'hd : _GEN_34744; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34746 = 10'hdb == _T_509[9:0] ? 4'hc : _GEN_34745; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34747 = 10'hdc == _T_509[9:0] ? 4'h9 : _GEN_34746; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34748 = 10'hdd == _T_509[9:0] ? 4'he : _GEN_34747; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34749 = 10'hde == _T_509[9:0] ? 4'he : _GEN_34748; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34750 = 10'hdf == _T_509[9:0] ? 4'he : _GEN_34749; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34751 = 10'he0 == _T_509[9:0] ? 4'he : _GEN_34750; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34752 = 10'he1 == _T_509[9:0] ? 4'he : _GEN_34751; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34753 = 10'he2 == _T_509[9:0] ? 4'he : _GEN_34752; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34754 = 10'he3 == _T_509[9:0] ? 4'h9 : _GEN_34753; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34755 = 10'he4 == _T_509[9:0] ? 4'he : _GEN_34754; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34756 = 10'he5 == _T_509[9:0] ? 4'he : _GEN_34755; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34757 = 10'he6 == _T_509[9:0] ? 4'he : _GEN_34756; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34758 = 10'he7 == _T_509[9:0] ? 4'he : _GEN_34757; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34759 = 10'he8 == _T_509[9:0] ? 4'he : _GEN_34758; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34760 = 10'he9 == _T_509[9:0] ? 4'he : _GEN_34759; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34761 = 10'hea == _T_509[9:0] ? 4'he : _GEN_34760; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34762 = 10'heb == _T_509[9:0] ? 4'hc : _GEN_34761; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34763 = 10'hec == _T_509[9:0] ? 4'h7 : _GEN_34762; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34764 = 10'hed == _T_509[9:0] ? 4'h1 : _GEN_34763; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34765 = 10'hee == _T_509[9:0] ? 4'h0 : _GEN_34764; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34766 = 10'hef == _T_509[9:0] ? 4'h0 : _GEN_34765; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34767 = 10'hf0 == _T_509[9:0] ? 4'h2 : _GEN_34766; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34768 = 10'hf1 == _T_509[9:0] ? 4'h9 : _GEN_34767; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34769 = 10'hf2 == _T_509[9:0] ? 4'he : _GEN_34768; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34770 = 10'hf3 == _T_509[9:0] ? 4'he : _GEN_34769; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34771 = 10'hf4 == _T_509[9:0] ? 4'he : _GEN_34770; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34772 = 10'hf5 == _T_509[9:0] ? 4'hc : _GEN_34771; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34773 = 10'hf6 == _T_509[9:0] ? 4'hc : _GEN_34772; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34774 = 10'hf7 == _T_509[9:0] ? 4'hd : _GEN_34773; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34775 = 10'hf8 == _T_509[9:0] ? 4'hd : _GEN_34774; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34776 = 10'hf9 == _T_509[9:0] ? 4'hd : _GEN_34775; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34777 = 10'hfa == _T_509[9:0] ? 4'hd : _GEN_34776; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34778 = 10'hfb == _T_509[9:0] ? 4'hd : _GEN_34777; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34779 = 10'hfc == _T_509[9:0] ? 4'hd : _GEN_34778; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34780 = 10'hfd == _T_509[9:0] ? 4'hd : _GEN_34779; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34781 = 10'hfe == _T_509[9:0] ? 4'hd : _GEN_34780; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34782 = 10'hff == _T_509[9:0] ? 4'hd : _GEN_34781; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34783 = 10'h100 == _T_509[9:0] ? 4'hd : _GEN_34782; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34784 = 10'h101 == _T_509[9:0] ? 4'h9 : _GEN_34783; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34785 = 10'h102 == _T_509[9:0] ? 4'h9 : _GEN_34784; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34786 = 10'h103 == _T_509[9:0] ? 4'he : _GEN_34785; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34787 = 10'h104 == _T_509[9:0] ? 4'he : _GEN_34786; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34788 = 10'h105 == _T_509[9:0] ? 4'he : _GEN_34787; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34789 = 10'h106 == _T_509[9:0] ? 4'he : _GEN_34788; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34790 = 10'h107 == _T_509[9:0] ? 4'he : _GEN_34789; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34791 = 10'h108 == _T_509[9:0] ? 4'he : _GEN_34790; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34792 = 10'h109 == _T_509[9:0] ? 4'h6 : _GEN_34791; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34793 = 10'h10a == _T_509[9:0] ? 4'he : _GEN_34792; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34794 = 10'h10b == _T_509[9:0] ? 4'he : _GEN_34793; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34795 = 10'h10c == _T_509[9:0] ? 4'he : _GEN_34794; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34796 = 10'h10d == _T_509[9:0] ? 4'he : _GEN_34795; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34797 = 10'h10e == _T_509[9:0] ? 4'he : _GEN_34796; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34798 = 10'h10f == _T_509[9:0] ? 4'ha : _GEN_34797; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34799 = 10'h110 == _T_509[9:0] ? 4'hd : _GEN_34798; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34800 = 10'h111 == _T_509[9:0] ? 4'h4 : _GEN_34799; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34801 = 10'h112 == _T_509[9:0] ? 4'h7 : _GEN_34800; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34802 = 10'h113 == _T_509[9:0] ? 4'h0 : _GEN_34801; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34803 = 10'h114 == _T_509[9:0] ? 4'h0 : _GEN_34802; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34804 = 10'h115 == _T_509[9:0] ? 4'h0 : _GEN_34803; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34805 = 10'h116 == _T_509[9:0] ? 4'h0 : _GEN_34804; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34806 = 10'h117 == _T_509[9:0] ? 4'h0 : _GEN_34805; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34807 = 10'h118 == _T_509[9:0] ? 4'ha : _GEN_34806; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34808 = 10'h119 == _T_509[9:0] ? 4'he : _GEN_34807; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34809 = 10'h11a == _T_509[9:0] ? 4'he : _GEN_34808; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34810 = 10'h11b == _T_509[9:0] ? 4'he : _GEN_34809; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34811 = 10'h11c == _T_509[9:0] ? 4'hb : _GEN_34810; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34812 = 10'h11d == _T_509[9:0] ? 4'hc : _GEN_34811; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34813 = 10'h11e == _T_509[9:0] ? 4'hd : _GEN_34812; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34814 = 10'h11f == _T_509[9:0] ? 4'hb : _GEN_34813; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34815 = 10'h120 == _T_509[9:0] ? 4'ha : _GEN_34814; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34816 = 10'h121 == _T_509[9:0] ? 4'hc : _GEN_34815; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34817 = 10'h122 == _T_509[9:0] ? 4'ha : _GEN_34816; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34818 = 10'h123 == _T_509[9:0] ? 4'ha : _GEN_34817; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34819 = 10'h124 == _T_509[9:0] ? 4'hd : _GEN_34818; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34820 = 10'h125 == _T_509[9:0] ? 4'hd : _GEN_34819; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34821 = 10'h126 == _T_509[9:0] ? 4'hb : _GEN_34820; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34822 = 10'h127 == _T_509[9:0] ? 4'h9 : _GEN_34821; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34823 = 10'h128 == _T_509[9:0] ? 4'h7 : _GEN_34822; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34824 = 10'h129 == _T_509[9:0] ? 4'hd : _GEN_34823; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34825 = 10'h12a == _T_509[9:0] ? 4'hc : _GEN_34824; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34826 = 10'h12b == _T_509[9:0] ? 4'hb : _GEN_34825; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34827 = 10'h12c == _T_509[9:0] ? 4'hc : _GEN_34826; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34828 = 10'h12d == _T_509[9:0] ? 4'hb : _GEN_34827; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34829 = 10'h12e == _T_509[9:0] ? 4'ha : _GEN_34828; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34830 = 10'h12f == _T_509[9:0] ? 4'h6 : _GEN_34829; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34831 = 10'h130 == _T_509[9:0] ? 4'he : _GEN_34830; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34832 = 10'h131 == _T_509[9:0] ? 4'hc : _GEN_34831; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34833 = 10'h132 == _T_509[9:0] ? 4'ha : _GEN_34832; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34834 = 10'h133 == _T_509[9:0] ? 4'h9 : _GEN_34833; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34835 = 10'h134 == _T_509[9:0] ? 4'hb : _GEN_34834; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34836 = 10'h135 == _T_509[9:0] ? 4'h8 : _GEN_34835; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34837 = 10'h136 == _T_509[9:0] ? 4'h8 : _GEN_34836; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34838 = 10'h137 == _T_509[9:0] ? 4'h4 : _GEN_34837; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34839 = 10'h138 == _T_509[9:0] ? 4'h7 : _GEN_34838; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34840 = 10'h139 == _T_509[9:0] ? 4'h0 : _GEN_34839; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34841 = 10'h13a == _T_509[9:0] ? 4'h0 : _GEN_34840; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34842 = 10'h13b == _T_509[9:0] ? 4'h0 : _GEN_34841; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34843 = 10'h13c == _T_509[9:0] ? 4'h0 : _GEN_34842; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34844 = 10'h13d == _T_509[9:0] ? 4'h0 : _GEN_34843; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34845 = 10'h13e == _T_509[9:0] ? 4'h4 : _GEN_34844; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34846 = 10'h13f == _T_509[9:0] ? 4'hc : _GEN_34845; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34847 = 10'h140 == _T_509[9:0] ? 4'he : _GEN_34846; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34848 = 10'h141 == _T_509[9:0] ? 4'he : _GEN_34847; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34849 = 10'h142 == _T_509[9:0] ? 4'he : _GEN_34848; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34850 = 10'h143 == _T_509[9:0] ? 4'hc : _GEN_34849; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34851 = 10'h144 == _T_509[9:0] ? 4'hd : _GEN_34850; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34852 = 10'h145 == _T_509[9:0] ? 4'hb : _GEN_34851; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34853 = 10'h146 == _T_509[9:0] ? 4'hb : _GEN_34852; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34854 = 10'h147 == _T_509[9:0] ? 4'ha : _GEN_34853; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34855 = 10'h148 == _T_509[9:0] ? 4'ha : _GEN_34854; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34856 = 10'h149 == _T_509[9:0] ? 4'hc : _GEN_34855; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34857 = 10'h14a == _T_509[9:0] ? 4'hd : _GEN_34856; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34858 = 10'h14b == _T_509[9:0] ? 4'hc : _GEN_34857; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34859 = 10'h14c == _T_509[9:0] ? 4'hd : _GEN_34858; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34860 = 10'h14d == _T_509[9:0] ? 4'h9 : _GEN_34859; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34861 = 10'h14e == _T_509[9:0] ? 4'h7 : _GEN_34860; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34862 = 10'h14f == _T_509[9:0] ? 4'ha : _GEN_34861; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34863 = 10'h150 == _T_509[9:0] ? 4'ha : _GEN_34862; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34864 = 10'h151 == _T_509[9:0] ? 4'hb : _GEN_34863; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34865 = 10'h152 == _T_509[9:0] ? 4'hb : _GEN_34864; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34866 = 10'h153 == _T_509[9:0] ? 4'hc : _GEN_34865; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34867 = 10'h154 == _T_509[9:0] ? 4'hb : _GEN_34866; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34868 = 10'h155 == _T_509[9:0] ? 4'h6 : _GEN_34867; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34869 = 10'h156 == _T_509[9:0] ? 4'hb : _GEN_34868; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34870 = 10'h157 == _T_509[9:0] ? 4'h7 : _GEN_34869; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34871 = 10'h158 == _T_509[9:0] ? 4'h7 : _GEN_34870; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34872 = 10'h159 == _T_509[9:0] ? 4'h7 : _GEN_34871; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34873 = 10'h15a == _T_509[9:0] ? 4'h7 : _GEN_34872; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34874 = 10'h15b == _T_509[9:0] ? 4'h7 : _GEN_34873; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34875 = 10'h15c == _T_509[9:0] ? 4'h7 : _GEN_34874; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34876 = 10'h15d == _T_509[9:0] ? 4'h6 : _GEN_34875; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34877 = 10'h15e == _T_509[9:0] ? 4'h7 : _GEN_34876; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34878 = 10'h15f == _T_509[9:0] ? 4'h0 : _GEN_34877; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34879 = 10'h160 == _T_509[9:0] ? 4'h0 : _GEN_34878; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34880 = 10'h161 == _T_509[9:0] ? 4'h0 : _GEN_34879; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34881 = 10'h162 == _T_509[9:0] ? 4'h0 : _GEN_34880; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34882 = 10'h163 == _T_509[9:0] ? 4'h2 : _GEN_34881; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34883 = 10'h164 == _T_509[9:0] ? 4'h4 : _GEN_34882; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34884 = 10'h165 == _T_509[9:0] ? 4'hb : _GEN_34883; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34885 = 10'h166 == _T_509[9:0] ? 4'hb : _GEN_34884; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34886 = 10'h167 == _T_509[9:0] ? 4'he : _GEN_34885; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34887 = 10'h168 == _T_509[9:0] ? 4'he : _GEN_34886; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34888 = 10'h169 == _T_509[9:0] ? 4'hc : _GEN_34887; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34889 = 10'h16a == _T_509[9:0] ? 4'hd : _GEN_34888; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34890 = 10'h16b == _T_509[9:0] ? 4'hd : _GEN_34889; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34891 = 10'h16c == _T_509[9:0] ? 4'ha : _GEN_34890; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34892 = 10'h16d == _T_509[9:0] ? 4'ha : _GEN_34891; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34893 = 10'h16e == _T_509[9:0] ? 4'ha : _GEN_34892; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34894 = 10'h16f == _T_509[9:0] ? 4'hd : _GEN_34893; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34895 = 10'h170 == _T_509[9:0] ? 4'hd : _GEN_34894; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34896 = 10'h171 == _T_509[9:0] ? 4'hd : _GEN_34895; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34897 = 10'h172 == _T_509[9:0] ? 4'he : _GEN_34896; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34898 = 10'h173 == _T_509[9:0] ? 4'h8 : _GEN_34897; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34899 = 10'h174 == _T_509[9:0] ? 4'h5 : _GEN_34898; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34900 = 10'h175 == _T_509[9:0] ? 4'h6 : _GEN_34899; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34901 = 10'h176 == _T_509[9:0] ? 4'h6 : _GEN_34900; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34902 = 10'h177 == _T_509[9:0] ? 4'h6 : _GEN_34901; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34903 = 10'h178 == _T_509[9:0] ? 4'h7 : _GEN_34902; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34904 = 10'h179 == _T_509[9:0] ? 4'h9 : _GEN_34903; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34905 = 10'h17a == _T_509[9:0] ? 4'h9 : _GEN_34904; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34906 = 10'h17b == _T_509[9:0] ? 4'h6 : _GEN_34905; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34907 = 10'h17c == _T_509[9:0] ? 4'h7 : _GEN_34906; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34908 = 10'h17d == _T_509[9:0] ? 4'h7 : _GEN_34907; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34909 = 10'h17e == _T_509[9:0] ? 4'h7 : _GEN_34908; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34910 = 10'h17f == _T_509[9:0] ? 4'h7 : _GEN_34909; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34911 = 10'h180 == _T_509[9:0] ? 4'h7 : _GEN_34910; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34912 = 10'h181 == _T_509[9:0] ? 4'h7 : _GEN_34911; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34913 = 10'h182 == _T_509[9:0] ? 4'h8 : _GEN_34912; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34914 = 10'h183 == _T_509[9:0] ? 4'h8 : _GEN_34913; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34915 = 10'h184 == _T_509[9:0] ? 4'h8 : _GEN_34914; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34916 = 10'h185 == _T_509[9:0] ? 4'h7 : _GEN_34915; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34917 = 10'h186 == _T_509[9:0] ? 4'h1 : _GEN_34916; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34918 = 10'h187 == _T_509[9:0] ? 4'h0 : _GEN_34917; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34919 = 10'h188 == _T_509[9:0] ? 4'h0 : _GEN_34918; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34920 = 10'h189 == _T_509[9:0] ? 4'h4 : _GEN_34919; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34921 = 10'h18a == _T_509[9:0] ? 4'h4 : _GEN_34920; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34922 = 10'h18b == _T_509[9:0] ? 4'hb : _GEN_34921; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34923 = 10'h18c == _T_509[9:0] ? 4'hb : _GEN_34922; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34924 = 10'h18d == _T_509[9:0] ? 4'hc : _GEN_34923; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34925 = 10'h18e == _T_509[9:0] ? 4'he : _GEN_34924; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34926 = 10'h18f == _T_509[9:0] ? 4'hb : _GEN_34925; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34927 = 10'h190 == _T_509[9:0] ? 4'hd : _GEN_34926; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34928 = 10'h191 == _T_509[9:0] ? 4'hc : _GEN_34927; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34929 = 10'h192 == _T_509[9:0] ? 4'h9 : _GEN_34928; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34930 = 10'h193 == _T_509[9:0] ? 4'ha : _GEN_34929; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34931 = 10'h194 == _T_509[9:0] ? 4'h9 : _GEN_34930; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34932 = 10'h195 == _T_509[9:0] ? 4'hd : _GEN_34931; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34933 = 10'h196 == _T_509[9:0] ? 4'hd : _GEN_34932; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34934 = 10'h197 == _T_509[9:0] ? 4'hb : _GEN_34933; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34935 = 10'h198 == _T_509[9:0] ? 4'he : _GEN_34934; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34936 = 10'h199 == _T_509[9:0] ? 4'h5 : _GEN_34935; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34937 = 10'h19a == _T_509[9:0] ? 4'h1 : _GEN_34936; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34938 = 10'h19b == _T_509[9:0] ? 4'h3 : _GEN_34937; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34939 = 10'h19c == _T_509[9:0] ? 4'h6 : _GEN_34938; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34940 = 10'h19d == _T_509[9:0] ? 4'h4 : _GEN_34939; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34941 = 10'h19e == _T_509[9:0] ? 4'h1 : _GEN_34940; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34942 = 10'h19f == _T_509[9:0] ? 4'h3 : _GEN_34941; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34943 = 10'h1a0 == _T_509[9:0] ? 4'h6 : _GEN_34942; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34944 = 10'h1a1 == _T_509[9:0] ? 4'h6 : _GEN_34943; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34945 = 10'h1a2 == _T_509[9:0] ? 4'h7 : _GEN_34944; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34946 = 10'h1a3 == _T_509[9:0] ? 4'h7 : _GEN_34945; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34947 = 10'h1a4 == _T_509[9:0] ? 4'h7 : _GEN_34946; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34948 = 10'h1a5 == _T_509[9:0] ? 4'h7 : _GEN_34947; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34949 = 10'h1a6 == _T_509[9:0] ? 4'h7 : _GEN_34948; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34950 = 10'h1a7 == _T_509[9:0] ? 4'h7 : _GEN_34949; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34951 = 10'h1a8 == _T_509[9:0] ? 4'h8 : _GEN_34950; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34952 = 10'h1a9 == _T_509[9:0] ? 4'h8 : _GEN_34951; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34953 = 10'h1aa == _T_509[9:0] ? 4'h7 : _GEN_34952; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34954 = 10'h1ab == _T_509[9:0] ? 4'h8 : _GEN_34953; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34955 = 10'h1ac == _T_509[9:0] ? 4'h8 : _GEN_34954; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34956 = 10'h1ad == _T_509[9:0] ? 4'h3 : _GEN_34955; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34957 = 10'h1ae == _T_509[9:0] ? 4'h2 : _GEN_34956; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34958 = 10'h1af == _T_509[9:0] ? 4'h8 : _GEN_34957; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34959 = 10'h1b0 == _T_509[9:0] ? 4'h6 : _GEN_34958; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34960 = 10'h1b1 == _T_509[9:0] ? 4'hb : _GEN_34959; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34961 = 10'h1b2 == _T_509[9:0] ? 4'hb : _GEN_34960; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34962 = 10'h1b3 == _T_509[9:0] ? 4'ha : _GEN_34961; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34963 = 10'h1b4 == _T_509[9:0] ? 4'he : _GEN_34962; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34964 = 10'h1b5 == _T_509[9:0] ? 4'hb : _GEN_34963; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34965 = 10'h1b6 == _T_509[9:0] ? 4'hc : _GEN_34964; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34966 = 10'h1b7 == _T_509[9:0] ? 4'ha : _GEN_34965; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34967 = 10'h1b8 == _T_509[9:0] ? 4'h9 : _GEN_34966; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34968 = 10'h1b9 == _T_509[9:0] ? 4'h9 : _GEN_34967; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34969 = 10'h1ba == _T_509[9:0] ? 4'h9 : _GEN_34968; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34970 = 10'h1bb == _T_509[9:0] ? 4'hb : _GEN_34969; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34971 = 10'h1bc == _T_509[9:0] ? 4'hd : _GEN_34970; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34972 = 10'h1bd == _T_509[9:0] ? 4'hd : _GEN_34971; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34973 = 10'h1be == _T_509[9:0] ? 4'he : _GEN_34972; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34974 = 10'h1bf == _T_509[9:0] ? 4'h7 : _GEN_34973; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34975 = 10'h1c0 == _T_509[9:0] ? 4'h6 : _GEN_34974; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34976 = 10'h1c1 == _T_509[9:0] ? 4'h6 : _GEN_34975; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34977 = 10'h1c2 == _T_509[9:0] ? 4'h5 : _GEN_34976; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34978 = 10'h1c3 == _T_509[9:0] ? 4'h5 : _GEN_34977; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34979 = 10'h1c4 == _T_509[9:0] ? 4'h4 : _GEN_34978; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34980 = 10'h1c5 == _T_509[9:0] ? 4'h5 : _GEN_34979; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34981 = 10'h1c6 == _T_509[9:0] ? 4'h6 : _GEN_34980; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34982 = 10'h1c7 == _T_509[9:0] ? 4'h6 : _GEN_34981; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34983 = 10'h1c8 == _T_509[9:0] ? 4'h7 : _GEN_34982; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34984 = 10'h1c9 == _T_509[9:0] ? 4'h7 : _GEN_34983; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34985 = 10'h1ca == _T_509[9:0] ? 4'h7 : _GEN_34984; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34986 = 10'h1cb == _T_509[9:0] ? 4'h7 : _GEN_34985; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34987 = 10'h1cc == _T_509[9:0] ? 4'h7 : _GEN_34986; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34988 = 10'h1cd == _T_509[9:0] ? 4'h8 : _GEN_34987; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34989 = 10'h1ce == _T_509[9:0] ? 4'h8 : _GEN_34988; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34990 = 10'h1cf == _T_509[9:0] ? 4'h8 : _GEN_34989; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34991 = 10'h1d0 == _T_509[9:0] ? 4'h5 : _GEN_34990; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34992 = 10'h1d1 == _T_509[9:0] ? 4'h8 : _GEN_34991; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34993 = 10'h1d2 == _T_509[9:0] ? 4'h8 : _GEN_34992; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34994 = 10'h1d3 == _T_509[9:0] ? 4'h8 : _GEN_34993; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34995 = 10'h1d4 == _T_509[9:0] ? 4'h8 : _GEN_34994; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34996 = 10'h1d5 == _T_509[9:0] ? 4'h7 : _GEN_34995; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34997 = 10'h1d6 == _T_509[9:0] ? 4'h9 : _GEN_34996; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34998 = 10'h1d7 == _T_509[9:0] ? 4'hb : _GEN_34997; // @[Filter.scala 230:102]
  wire [3:0] _GEN_34999 = 10'h1d8 == _T_509[9:0] ? 4'hb : _GEN_34998; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35000 = 10'h1d9 == _T_509[9:0] ? 4'hb : _GEN_34999; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35001 = 10'h1da == _T_509[9:0] ? 4'ha : _GEN_35000; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35002 = 10'h1db == _T_509[9:0] ? 4'hc : _GEN_35001; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35003 = 10'h1dc == _T_509[9:0] ? 4'hb : _GEN_35002; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35004 = 10'h1dd == _T_509[9:0] ? 4'h5 : _GEN_35003; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35005 = 10'h1de == _T_509[9:0] ? 4'h9 : _GEN_35004; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35006 = 10'h1df == _T_509[9:0] ? 4'h9 : _GEN_35005; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35007 = 10'h1e0 == _T_509[9:0] ? 4'h9 : _GEN_35006; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35008 = 10'h1e1 == _T_509[9:0] ? 4'h7 : _GEN_35007; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35009 = 10'h1e2 == _T_509[9:0] ? 4'hc : _GEN_35008; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35010 = 10'h1e3 == _T_509[9:0] ? 4'hc : _GEN_35009; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35011 = 10'h1e4 == _T_509[9:0] ? 4'hd : _GEN_35010; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35012 = 10'h1e5 == _T_509[9:0] ? 4'h7 : _GEN_35011; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35013 = 10'h1e6 == _T_509[9:0] ? 4'h6 : _GEN_35012; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35014 = 10'h1e7 == _T_509[9:0] ? 4'h6 : _GEN_35013; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35015 = 10'h1e8 == _T_509[9:0] ? 4'h6 : _GEN_35014; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35016 = 10'h1e9 == _T_509[9:0] ? 4'h6 : _GEN_35015; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35017 = 10'h1ea == _T_509[9:0] ? 4'h6 : _GEN_35016; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35018 = 10'h1eb == _T_509[9:0] ? 4'h6 : _GEN_35017; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35019 = 10'h1ec == _T_509[9:0] ? 4'h6 : _GEN_35018; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35020 = 10'h1ed == _T_509[9:0] ? 4'h8 : _GEN_35019; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35021 = 10'h1ee == _T_509[9:0] ? 4'h7 : _GEN_35020; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35022 = 10'h1ef == _T_509[9:0] ? 4'h7 : _GEN_35021; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35023 = 10'h1f0 == _T_509[9:0] ? 4'h7 : _GEN_35022; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35024 = 10'h1f1 == _T_509[9:0] ? 4'h7 : _GEN_35023; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35025 = 10'h1f2 == _T_509[9:0] ? 4'h7 : _GEN_35024; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35026 = 10'h1f3 == _T_509[9:0] ? 4'h8 : _GEN_35025; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35027 = 10'h1f4 == _T_509[9:0] ? 4'h8 : _GEN_35026; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35028 = 10'h1f5 == _T_509[9:0] ? 4'h8 : _GEN_35027; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35029 = 10'h1f6 == _T_509[9:0] ? 4'ha : _GEN_35028; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35030 = 10'h1f7 == _T_509[9:0] ? 4'h8 : _GEN_35029; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35031 = 10'h1f8 == _T_509[9:0] ? 4'h8 : _GEN_35030; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35032 = 10'h1f9 == _T_509[9:0] ? 4'h9 : _GEN_35031; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35033 = 10'h1fa == _T_509[9:0] ? 4'h9 : _GEN_35032; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35034 = 10'h1fb == _T_509[9:0] ? 4'h8 : _GEN_35033; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35035 = 10'h1fc == _T_509[9:0] ? 4'hb : _GEN_35034; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35036 = 10'h1fd == _T_509[9:0] ? 4'hb : _GEN_35035; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35037 = 10'h1fe == _T_509[9:0] ? 4'hb : _GEN_35036; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35038 = 10'h1ff == _T_509[9:0] ? 4'ha : _GEN_35037; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35039 = 10'h200 == _T_509[9:0] ? 4'h3 : _GEN_35038; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35040 = 10'h201 == _T_509[9:0] ? 4'h9 : _GEN_35039; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35041 = 10'h202 == _T_509[9:0] ? 4'h5 : _GEN_35040; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35042 = 10'h203 == _T_509[9:0] ? 4'h3 : _GEN_35041; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35043 = 10'h204 == _T_509[9:0] ? 4'h4 : _GEN_35042; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35044 = 10'h205 == _T_509[9:0] ? 4'h4 : _GEN_35043; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35045 = 10'h206 == _T_509[9:0] ? 4'h4 : _GEN_35044; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35046 = 10'h207 == _T_509[9:0] ? 4'h4 : _GEN_35045; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35047 = 10'h208 == _T_509[9:0] ? 4'h8 : _GEN_35046; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35048 = 10'h209 == _T_509[9:0] ? 4'hc : _GEN_35047; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35049 = 10'h20a == _T_509[9:0] ? 4'hd : _GEN_35048; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35050 = 10'h20b == _T_509[9:0] ? 4'h7 : _GEN_35049; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35051 = 10'h20c == _T_509[9:0] ? 4'h6 : _GEN_35050; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35052 = 10'h20d == _T_509[9:0] ? 4'h6 : _GEN_35051; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35053 = 10'h20e == _T_509[9:0] ? 4'h6 : _GEN_35052; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35054 = 10'h20f == _T_509[9:0] ? 4'h5 : _GEN_35053; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35055 = 10'h210 == _T_509[9:0] ? 4'h6 : _GEN_35054; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35056 = 10'h211 == _T_509[9:0] ? 4'h6 : _GEN_35055; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35057 = 10'h212 == _T_509[9:0] ? 4'h7 : _GEN_35056; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35058 = 10'h213 == _T_509[9:0] ? 4'ha : _GEN_35057; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35059 = 10'h214 == _T_509[9:0] ? 4'h6 : _GEN_35058; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35060 = 10'h215 == _T_509[9:0] ? 4'h7 : _GEN_35059; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35061 = 10'h216 == _T_509[9:0] ? 4'h7 : _GEN_35060; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35062 = 10'h217 == _T_509[9:0] ? 4'h7 : _GEN_35061; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35063 = 10'h218 == _T_509[9:0] ? 4'h7 : _GEN_35062; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35064 = 10'h219 == _T_509[9:0] ? 4'h8 : _GEN_35063; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35065 = 10'h21a == _T_509[9:0] ? 4'h7 : _GEN_35064; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35066 = 10'h21b == _T_509[9:0] ? 4'h8 : _GEN_35065; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35067 = 10'h21c == _T_509[9:0] ? 4'hb : _GEN_35066; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35068 = 10'h21d == _T_509[9:0] ? 4'ha : _GEN_35067; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35069 = 10'h21e == _T_509[9:0] ? 4'h9 : _GEN_35068; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35070 = 10'h21f == _T_509[9:0] ? 4'h9 : _GEN_35069; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35071 = 10'h220 == _T_509[9:0] ? 4'h8 : _GEN_35070; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35072 = 10'h221 == _T_509[9:0] ? 4'h9 : _GEN_35071; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35073 = 10'h222 == _T_509[9:0] ? 4'hb : _GEN_35072; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35074 = 10'h223 == _T_509[9:0] ? 4'hb : _GEN_35073; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35075 = 10'h224 == _T_509[9:0] ? 4'hb : _GEN_35074; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35076 = 10'h225 == _T_509[9:0] ? 4'h8 : _GEN_35075; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35077 = 10'h226 == _T_509[9:0] ? 4'h1 : _GEN_35076; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35078 = 10'h227 == _T_509[9:0] ? 4'h3 : _GEN_35077; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35079 = 10'h228 == _T_509[9:0] ? 4'h3 : _GEN_35078; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35080 = 10'h229 == _T_509[9:0] ? 4'h3 : _GEN_35079; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35081 = 10'h22a == _T_509[9:0] ? 4'h3 : _GEN_35080; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35082 = 10'h22b == _T_509[9:0] ? 4'h3 : _GEN_35081; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35083 = 10'h22c == _T_509[9:0] ? 4'h3 : _GEN_35082; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35084 = 10'h22d == _T_509[9:0] ? 4'h3 : _GEN_35083; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35085 = 10'h22e == _T_509[9:0] ? 4'h3 : _GEN_35084; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35086 = 10'h22f == _T_509[9:0] ? 4'h9 : _GEN_35085; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35087 = 10'h230 == _T_509[9:0] ? 4'h6 : _GEN_35086; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35088 = 10'h231 == _T_509[9:0] ? 4'h7 : _GEN_35087; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35089 = 10'h232 == _T_509[9:0] ? 4'h6 : _GEN_35088; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35090 = 10'h233 == _T_509[9:0] ? 4'h7 : _GEN_35089; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35091 = 10'h234 == _T_509[9:0] ? 4'h7 : _GEN_35090; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35092 = 10'h235 == _T_509[9:0] ? 4'h6 : _GEN_35091; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35093 = 10'h236 == _T_509[9:0] ? 4'h6 : _GEN_35092; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35094 = 10'h237 == _T_509[9:0] ? 4'h6 : _GEN_35093; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35095 = 10'h238 == _T_509[9:0] ? 4'h6 : _GEN_35094; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35096 = 10'h239 == _T_509[9:0] ? 4'h8 : _GEN_35095; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35097 = 10'h23a == _T_509[9:0] ? 4'h6 : _GEN_35096; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35098 = 10'h23b == _T_509[9:0] ? 4'h7 : _GEN_35097; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35099 = 10'h23c == _T_509[9:0] ? 4'h7 : _GEN_35098; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35100 = 10'h23d == _T_509[9:0] ? 4'h7 : _GEN_35099; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35101 = 10'h23e == _T_509[9:0] ? 4'h7 : _GEN_35100; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35102 = 10'h23f == _T_509[9:0] ? 4'h7 : _GEN_35101; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35103 = 10'h240 == _T_509[9:0] ? 4'h7 : _GEN_35102; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35104 = 10'h241 == _T_509[9:0] ? 4'h8 : _GEN_35103; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35105 = 10'h242 == _T_509[9:0] ? 4'hb : _GEN_35104; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35106 = 10'h243 == _T_509[9:0] ? 4'hb : _GEN_35105; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35107 = 10'h244 == _T_509[9:0] ? 4'hb : _GEN_35106; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35108 = 10'h245 == _T_509[9:0] ? 4'ha : _GEN_35107; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35109 = 10'h246 == _T_509[9:0] ? 4'h9 : _GEN_35108; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35110 = 10'h247 == _T_509[9:0] ? 4'ha : _GEN_35109; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35111 = 10'h248 == _T_509[9:0] ? 4'hb : _GEN_35110; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35112 = 10'h249 == _T_509[9:0] ? 4'hb : _GEN_35111; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35113 = 10'h24a == _T_509[9:0] ? 4'ha : _GEN_35112; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35114 = 10'h24b == _T_509[9:0] ? 4'h2 : _GEN_35113; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35115 = 10'h24c == _T_509[9:0] ? 4'h0 : _GEN_35114; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35116 = 10'h24d == _T_509[9:0] ? 4'h2 : _GEN_35115; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35117 = 10'h24e == _T_509[9:0] ? 4'h3 : _GEN_35116; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35118 = 10'h24f == _T_509[9:0] ? 4'h3 : _GEN_35117; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35119 = 10'h250 == _T_509[9:0] ? 4'h3 : _GEN_35118; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35120 = 10'h251 == _T_509[9:0] ? 4'h3 : _GEN_35119; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35121 = 10'h252 == _T_509[9:0] ? 4'h3 : _GEN_35120; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35122 = 10'h253 == _T_509[9:0] ? 4'h3 : _GEN_35121; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35123 = 10'h254 == _T_509[9:0] ? 4'h3 : _GEN_35122; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35124 = 10'h255 == _T_509[9:0] ? 4'h5 : _GEN_35123; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35125 = 10'h256 == _T_509[9:0] ? 4'h6 : _GEN_35124; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35126 = 10'h257 == _T_509[9:0] ? 4'h8 : _GEN_35125; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35127 = 10'h258 == _T_509[9:0] ? 4'h5 : _GEN_35126; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35128 = 10'h259 == _T_509[9:0] ? 4'h6 : _GEN_35127; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35129 = 10'h25a == _T_509[9:0] ? 4'h6 : _GEN_35128; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35130 = 10'h25b == _T_509[9:0] ? 4'h5 : _GEN_35129; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35131 = 10'h25c == _T_509[9:0] ? 4'h6 : _GEN_35130; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35132 = 10'h25d == _T_509[9:0] ? 4'h6 : _GEN_35131; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35133 = 10'h25e == _T_509[9:0] ? 4'h9 : _GEN_35132; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35134 = 10'h25f == _T_509[9:0] ? 4'hc : _GEN_35133; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35135 = 10'h260 == _T_509[9:0] ? 4'h7 : _GEN_35134; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35136 = 10'h261 == _T_509[9:0] ? 4'h9 : _GEN_35135; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35137 = 10'h262 == _T_509[9:0] ? 4'ha : _GEN_35136; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35138 = 10'h263 == _T_509[9:0] ? 4'h8 : _GEN_35137; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35139 = 10'h264 == _T_509[9:0] ? 4'ha : _GEN_35138; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35140 = 10'h265 == _T_509[9:0] ? 4'h9 : _GEN_35139; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35141 = 10'h266 == _T_509[9:0] ? 4'h8 : _GEN_35140; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35142 = 10'h267 == _T_509[9:0] ? 4'h8 : _GEN_35141; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35143 = 10'h268 == _T_509[9:0] ? 4'ha : _GEN_35142; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35144 = 10'h269 == _T_509[9:0] ? 4'ha : _GEN_35143; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35145 = 10'h26a == _T_509[9:0] ? 4'hb : _GEN_35144; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35146 = 10'h26b == _T_509[9:0] ? 4'hb : _GEN_35145; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35147 = 10'h26c == _T_509[9:0] ? 4'hb : _GEN_35146; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35148 = 10'h26d == _T_509[9:0] ? 4'hb : _GEN_35147; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35149 = 10'h26e == _T_509[9:0] ? 4'hb : _GEN_35148; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35150 = 10'h26f == _T_509[9:0] ? 4'ha : _GEN_35149; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35151 = 10'h270 == _T_509[9:0] ? 4'h3 : _GEN_35150; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35152 = 10'h271 == _T_509[9:0] ? 4'h0 : _GEN_35151; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35153 = 10'h272 == _T_509[9:0] ? 4'h0 : _GEN_35152; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35154 = 10'h273 == _T_509[9:0] ? 4'h2 : _GEN_35153; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35155 = 10'h274 == _T_509[9:0] ? 4'h3 : _GEN_35154; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35156 = 10'h275 == _T_509[9:0] ? 4'h3 : _GEN_35155; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35157 = 10'h276 == _T_509[9:0] ? 4'h3 : _GEN_35156; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35158 = 10'h277 == _T_509[9:0] ? 4'h3 : _GEN_35157; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35159 = 10'h278 == _T_509[9:0] ? 4'h3 : _GEN_35158; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35160 = 10'h279 == _T_509[9:0] ? 4'h3 : _GEN_35159; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35161 = 10'h27a == _T_509[9:0] ? 4'h3 : _GEN_35160; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35162 = 10'h27b == _T_509[9:0] ? 4'h6 : _GEN_35161; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35163 = 10'h27c == _T_509[9:0] ? 4'h7 : _GEN_35162; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35164 = 10'h27d == _T_509[9:0] ? 4'h7 : _GEN_35163; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35165 = 10'h27e == _T_509[9:0] ? 4'h4 : _GEN_35164; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35166 = 10'h27f == _T_509[9:0] ? 4'h6 : _GEN_35165; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35167 = 10'h280 == _T_509[9:0] ? 4'h6 : _GEN_35166; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35168 = 10'h281 == _T_509[9:0] ? 4'h6 : _GEN_35167; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35169 = 10'h282 == _T_509[9:0] ? 4'h6 : _GEN_35168; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35170 = 10'h283 == _T_509[9:0] ? 4'ha : _GEN_35169; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35171 = 10'h284 == _T_509[9:0] ? 4'hc : _GEN_35170; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35172 = 10'h285 == _T_509[9:0] ? 4'hc : _GEN_35171; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35173 = 10'h286 == _T_509[9:0] ? 4'h8 : _GEN_35172; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35174 = 10'h287 == _T_509[9:0] ? 4'ha : _GEN_35173; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35175 = 10'h288 == _T_509[9:0] ? 4'ha : _GEN_35174; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35176 = 10'h289 == _T_509[9:0] ? 4'ha : _GEN_35175; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35177 = 10'h28a == _T_509[9:0] ? 4'hc : _GEN_35176; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35178 = 10'h28b == _T_509[9:0] ? 4'hb : _GEN_35177; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35179 = 10'h28c == _T_509[9:0] ? 4'ha : _GEN_35178; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35180 = 10'h28d == _T_509[9:0] ? 4'h7 : _GEN_35179; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35181 = 10'h28e == _T_509[9:0] ? 4'h2 : _GEN_35180; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35182 = 10'h28f == _T_509[9:0] ? 4'h5 : _GEN_35181; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35183 = 10'h290 == _T_509[9:0] ? 4'h8 : _GEN_35182; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35184 = 10'h291 == _T_509[9:0] ? 4'ha : _GEN_35183; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35185 = 10'h292 == _T_509[9:0] ? 4'ha : _GEN_35184; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35186 = 10'h293 == _T_509[9:0] ? 4'ha : _GEN_35185; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35187 = 10'h294 == _T_509[9:0] ? 4'h9 : _GEN_35186; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35188 = 10'h295 == _T_509[9:0] ? 4'h3 : _GEN_35187; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35189 = 10'h296 == _T_509[9:0] ? 4'h0 : _GEN_35188; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35190 = 10'h297 == _T_509[9:0] ? 4'h0 : _GEN_35189; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35191 = 10'h298 == _T_509[9:0] ? 4'h0 : _GEN_35190; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35192 = 10'h299 == _T_509[9:0] ? 4'h1 : _GEN_35191; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35193 = 10'h29a == _T_509[9:0] ? 4'h3 : _GEN_35192; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35194 = 10'h29b == _T_509[9:0] ? 4'h3 : _GEN_35193; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35195 = 10'h29c == _T_509[9:0] ? 4'h3 : _GEN_35194; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35196 = 10'h29d == _T_509[9:0] ? 4'h3 : _GEN_35195; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35197 = 10'h29e == _T_509[9:0] ? 4'h3 : _GEN_35196; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35198 = 10'h29f == _T_509[9:0] ? 4'h3 : _GEN_35197; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35199 = 10'h2a0 == _T_509[9:0] ? 4'h4 : _GEN_35198; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35200 = 10'h2a1 == _T_509[9:0] ? 4'h6 : _GEN_35199; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35201 = 10'h2a2 == _T_509[9:0] ? 4'h7 : _GEN_35200; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35202 = 10'h2a3 == _T_509[9:0] ? 4'h6 : _GEN_35201; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35203 = 10'h2a4 == _T_509[9:0] ? 4'h4 : _GEN_35202; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35204 = 10'h2a5 == _T_509[9:0] ? 4'h6 : _GEN_35203; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35205 = 10'h2a6 == _T_509[9:0] ? 4'h6 : _GEN_35204; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35206 = 10'h2a7 == _T_509[9:0] ? 4'h7 : _GEN_35205; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35207 = 10'h2a8 == _T_509[9:0] ? 4'ha : _GEN_35206; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35208 = 10'h2a9 == _T_509[9:0] ? 4'hb : _GEN_35207; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35209 = 10'h2aa == _T_509[9:0] ? 4'hb : _GEN_35208; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35210 = 10'h2ab == _T_509[9:0] ? 4'hb : _GEN_35209; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35211 = 10'h2ac == _T_509[9:0] ? 4'h8 : _GEN_35210; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35212 = 10'h2ad == _T_509[9:0] ? 4'hb : _GEN_35211; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35213 = 10'h2ae == _T_509[9:0] ? 4'ha : _GEN_35212; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35214 = 10'h2af == _T_509[9:0] ? 4'hb : _GEN_35213; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35215 = 10'h2b0 == _T_509[9:0] ? 4'hc : _GEN_35214; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35216 = 10'h2b1 == _T_509[9:0] ? 4'hb : _GEN_35215; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35217 = 10'h2b2 == _T_509[9:0] ? 4'ha : _GEN_35216; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35218 = 10'h2b3 == _T_509[9:0] ? 4'h6 : _GEN_35217; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35219 = 10'h2b4 == _T_509[9:0] ? 4'h0 : _GEN_35218; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35220 = 10'h2b5 == _T_509[9:0] ? 4'h0 : _GEN_35219; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35221 = 10'h2b6 == _T_509[9:0] ? 4'h0 : _GEN_35220; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35222 = 10'h2b7 == _T_509[9:0] ? 4'h1 : _GEN_35221; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35223 = 10'h2b8 == _T_509[9:0] ? 4'h5 : _GEN_35222; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35224 = 10'h2b9 == _T_509[9:0] ? 4'h9 : _GEN_35223; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35225 = 10'h2ba == _T_509[9:0] ? 4'h1 : _GEN_35224; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35226 = 10'h2bb == _T_509[9:0] ? 4'h0 : _GEN_35225; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35227 = 10'h2bc == _T_509[9:0] ? 4'h0 : _GEN_35226; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35228 = 10'h2bd == _T_509[9:0] ? 4'h0 : _GEN_35227; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35229 = 10'h2be == _T_509[9:0] ? 4'h0 : _GEN_35228; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35230 = 10'h2bf == _T_509[9:0] ? 4'h0 : _GEN_35229; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35231 = 10'h2c0 == _T_509[9:0] ? 4'h3 : _GEN_35230; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35232 = 10'h2c1 == _T_509[9:0] ? 4'h3 : _GEN_35231; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35233 = 10'h2c2 == _T_509[9:0] ? 4'h3 : _GEN_35232; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35234 = 10'h2c3 == _T_509[9:0] ? 4'h3 : _GEN_35233; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35235 = 10'h2c4 == _T_509[9:0] ? 4'h3 : _GEN_35234; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35236 = 10'h2c5 == _T_509[9:0] ? 4'h3 : _GEN_35235; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35237 = 10'h2c6 == _T_509[9:0] ? 4'h4 : _GEN_35236; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35238 = 10'h2c7 == _T_509[9:0] ? 4'h5 : _GEN_35237; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35239 = 10'h2c8 == _T_509[9:0] ? 4'h7 : _GEN_35238; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35240 = 10'h2c9 == _T_509[9:0] ? 4'h7 : _GEN_35239; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35241 = 10'h2ca == _T_509[9:0] ? 4'h4 : _GEN_35240; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35242 = 10'h2cb == _T_509[9:0] ? 4'h9 : _GEN_35241; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35243 = 10'h2cc == _T_509[9:0] ? 4'h9 : _GEN_35242; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35244 = 10'h2cd == _T_509[9:0] ? 4'hb : _GEN_35243; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35245 = 10'h2ce == _T_509[9:0] ? 4'hb : _GEN_35244; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35246 = 10'h2cf == _T_509[9:0] ? 4'hb : _GEN_35245; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35247 = 10'h2d0 == _T_509[9:0] ? 4'hb : _GEN_35246; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35248 = 10'h2d1 == _T_509[9:0] ? 4'hb : _GEN_35247; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35249 = 10'h2d2 == _T_509[9:0] ? 4'h8 : _GEN_35248; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35250 = 10'h2d3 == _T_509[9:0] ? 4'ha : _GEN_35249; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35251 = 10'h2d4 == _T_509[9:0] ? 4'hb : _GEN_35250; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35252 = 10'h2d5 == _T_509[9:0] ? 4'ha : _GEN_35251; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35253 = 10'h2d6 == _T_509[9:0] ? 4'ha : _GEN_35252; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35254 = 10'h2d7 == _T_509[9:0] ? 4'ha : _GEN_35253; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35255 = 10'h2d8 == _T_509[9:0] ? 4'ha : _GEN_35254; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35256 = 10'h2d9 == _T_509[9:0] ? 4'h7 : _GEN_35255; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35257 = 10'h2da == _T_509[9:0] ? 4'h2 : _GEN_35256; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35258 = 10'h2db == _T_509[9:0] ? 4'h0 : _GEN_35257; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35259 = 10'h2dc == _T_509[9:0] ? 4'h0 : _GEN_35258; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35260 = 10'h2dd == _T_509[9:0] ? 4'h0 : _GEN_35259; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35261 = 10'h2de == _T_509[9:0] ? 4'h0 : _GEN_35260; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35262 = 10'h2df == _T_509[9:0] ? 4'h2 : _GEN_35261; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35263 = 10'h2e0 == _T_509[9:0] ? 4'h0 : _GEN_35262; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35264 = 10'h2e1 == _T_509[9:0] ? 4'h0 : _GEN_35263; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35265 = 10'h2e2 == _T_509[9:0] ? 4'h0 : _GEN_35264; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35266 = 10'h2e3 == _T_509[9:0] ? 4'h0 : _GEN_35265; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35267 = 10'h2e4 == _T_509[9:0] ? 4'h0 : _GEN_35266; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35268 = 10'h2e5 == _T_509[9:0] ? 4'h0 : _GEN_35267; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35269 = 10'h2e6 == _T_509[9:0] ? 4'h2 : _GEN_35268; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35270 = 10'h2e7 == _T_509[9:0] ? 4'h3 : _GEN_35269; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35271 = 10'h2e8 == _T_509[9:0] ? 4'h3 : _GEN_35270; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35272 = 10'h2e9 == _T_509[9:0] ? 4'h3 : _GEN_35271; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35273 = 10'h2ea == _T_509[9:0] ? 4'h3 : _GEN_35272; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35274 = 10'h2eb == _T_509[9:0] ? 4'h3 : _GEN_35273; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35275 = 10'h2ec == _T_509[9:0] ? 4'h4 : _GEN_35274; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35276 = 10'h2ed == _T_509[9:0] ? 4'h5 : _GEN_35275; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35277 = 10'h2ee == _T_509[9:0] ? 4'h6 : _GEN_35276; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35278 = 10'h2ef == _T_509[9:0] ? 4'h8 : _GEN_35277; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35279 = 10'h2f0 == _T_509[9:0] ? 4'h4 : _GEN_35278; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35280 = 10'h2f1 == _T_509[9:0] ? 4'h9 : _GEN_35279; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35281 = 10'h2f2 == _T_509[9:0] ? 4'hb : _GEN_35280; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35282 = 10'h2f3 == _T_509[9:0] ? 4'hb : _GEN_35281; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35283 = 10'h2f4 == _T_509[9:0] ? 4'hb : _GEN_35282; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35284 = 10'h2f5 == _T_509[9:0] ? 4'hb : _GEN_35283; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35285 = 10'h2f6 == _T_509[9:0] ? 4'hb : _GEN_35284; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35286 = 10'h2f7 == _T_509[9:0] ? 4'hb : _GEN_35285; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35287 = 10'h2f8 == _T_509[9:0] ? 4'h8 : _GEN_35286; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35288 = 10'h2f9 == _T_509[9:0] ? 4'h9 : _GEN_35287; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35289 = 10'h2fa == _T_509[9:0] ? 4'hb : _GEN_35288; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35290 = 10'h2fb == _T_509[9:0] ? 4'hb : _GEN_35289; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35291 = 10'h2fc == _T_509[9:0] ? 4'ha : _GEN_35290; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35292 = 10'h2fd == _T_509[9:0] ? 4'ha : _GEN_35291; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35293 = 10'h2fe == _T_509[9:0] ? 4'h9 : _GEN_35292; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35294 = 10'h2ff == _T_509[9:0] ? 4'h8 : _GEN_35293; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35295 = 10'h300 == _T_509[9:0] ? 4'h8 : _GEN_35294; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35296 = 10'h301 == _T_509[9:0] ? 4'h6 : _GEN_35295; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35297 = 10'h302 == _T_509[9:0] ? 4'h1 : _GEN_35296; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35298 = 10'h303 == _T_509[9:0] ? 4'h0 : _GEN_35297; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35299 = 10'h304 == _T_509[9:0] ? 4'h0 : _GEN_35298; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35300 = 10'h305 == _T_509[9:0] ? 4'h0 : _GEN_35299; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35301 = 10'h306 == _T_509[9:0] ? 4'h0 : _GEN_35300; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35302 = 10'h307 == _T_509[9:0] ? 4'h0 : _GEN_35301; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35303 = 10'h308 == _T_509[9:0] ? 4'h0 : _GEN_35302; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35304 = 10'h309 == _T_509[9:0] ? 4'h0 : _GEN_35303; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35305 = 10'h30a == _T_509[9:0] ? 4'h0 : _GEN_35304; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35306 = 10'h30b == _T_509[9:0] ? 4'h0 : _GEN_35305; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35307 = 10'h30c == _T_509[9:0] ? 4'h2 : _GEN_35306; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35308 = 10'h30d == _T_509[9:0] ? 4'h3 : _GEN_35307; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35309 = 10'h30e == _T_509[9:0] ? 4'h3 : _GEN_35308; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35310 = 10'h30f == _T_509[9:0] ? 4'h3 : _GEN_35309; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35311 = 10'h310 == _T_509[9:0] ? 4'h3 : _GEN_35310; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35312 = 10'h311 == _T_509[9:0] ? 4'h3 : _GEN_35311; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35313 = 10'h312 == _T_509[9:0] ? 4'h4 : _GEN_35312; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35314 = 10'h313 == _T_509[9:0] ? 4'h5 : _GEN_35313; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35315 = 10'h314 == _T_509[9:0] ? 4'h5 : _GEN_35314; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35316 = 10'h315 == _T_509[9:0] ? 4'h8 : _GEN_35315; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35317 = 10'h316 == _T_509[9:0] ? 4'h4 : _GEN_35316; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35318 = 10'h317 == _T_509[9:0] ? 4'h6 : _GEN_35317; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35319 = 10'h318 == _T_509[9:0] ? 4'hb : _GEN_35318; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35320 = 10'h319 == _T_509[9:0] ? 4'hb : _GEN_35319; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35321 = 10'h31a == _T_509[9:0] ? 4'hb : _GEN_35320; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35322 = 10'h31b == _T_509[9:0] ? 4'hb : _GEN_35321; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35323 = 10'h31c == _T_509[9:0] ? 4'hb : _GEN_35322; // @[Filter.scala 230:102]
  wire [3:0] _GEN_35324 = 10'h31d == _T_509[9:0] ? 4'hb : _GEN_35323; // @[Filter.scala 230:102]
  wire [6:0] _GEN_39040 = {{3'd0}, _GEN_35324}; // @[Filter.scala 230:102]
  wire [10:0] _T_516 = _GEN_39040 * 7'h46; // @[Filter.scala 230:102]
  wire [10:0] _GEN_39041 = {{2'd0}, _T_511}; // @[Filter.scala 230:69]
  wire [10:0] _T_518 = _GEN_39041 + _T_516; // @[Filter.scala 230:69]
  wire [3:0] _GEN_35347 = 10'h16 == _T_509[9:0] ? 4'hb : 4'hc; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35348 = 10'h17 == _T_509[9:0] ? 4'h8 : _GEN_35347; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35349 = 10'h18 == _T_509[9:0] ? 4'ha : _GEN_35348; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35350 = 10'h19 == _T_509[9:0] ? 4'hc : _GEN_35349; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35351 = 10'h1a == _T_509[9:0] ? 4'hc : _GEN_35350; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35352 = 10'h1b == _T_509[9:0] ? 4'hc : _GEN_35351; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35353 = 10'h1c == _T_509[9:0] ? 4'hc : _GEN_35352; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35354 = 10'h1d == _T_509[9:0] ? 4'hc : _GEN_35353; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35355 = 10'h1e == _T_509[9:0] ? 4'hc : _GEN_35354; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35356 = 10'h1f == _T_509[9:0] ? 4'hc : _GEN_35355; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35357 = 10'h20 == _T_509[9:0] ? 4'hc : _GEN_35356; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35358 = 10'h21 == _T_509[9:0] ? 4'hc : _GEN_35357; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35359 = 10'h22 == _T_509[9:0] ? 4'hc : _GEN_35358; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35360 = 10'h23 == _T_509[9:0] ? 4'hc : _GEN_35359; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35361 = 10'h24 == _T_509[9:0] ? 4'hc : _GEN_35360; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35362 = 10'h25 == _T_509[9:0] ? 4'hc : _GEN_35361; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35363 = 10'h26 == _T_509[9:0] ? 4'hc : _GEN_35362; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35364 = 10'h27 == _T_509[9:0] ? 4'hc : _GEN_35363; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35365 = 10'h28 == _T_509[9:0] ? 4'hc : _GEN_35364; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35366 = 10'h29 == _T_509[9:0] ? 4'hc : _GEN_35365; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35367 = 10'h2a == _T_509[9:0] ? 4'hc : _GEN_35366; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35368 = 10'h2b == _T_509[9:0] ? 4'hc : _GEN_35367; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35369 = 10'h2c == _T_509[9:0] ? 4'hc : _GEN_35368; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35370 = 10'h2d == _T_509[9:0] ? 4'hc : _GEN_35369; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35371 = 10'h2e == _T_509[9:0] ? 4'hc : _GEN_35370; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35372 = 10'h2f == _T_509[9:0] ? 4'hc : _GEN_35371; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35373 = 10'h30 == _T_509[9:0] ? 4'hc : _GEN_35372; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35374 = 10'h31 == _T_509[9:0] ? 4'hc : _GEN_35373; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35375 = 10'h32 == _T_509[9:0] ? 4'hc : _GEN_35374; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35376 = 10'h33 == _T_509[9:0] ? 4'hc : _GEN_35375; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35377 = 10'h34 == _T_509[9:0] ? 4'hc : _GEN_35376; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35378 = 10'h35 == _T_509[9:0] ? 4'hc : _GEN_35377; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35379 = 10'h36 == _T_509[9:0] ? 4'hc : _GEN_35378; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35380 = 10'h37 == _T_509[9:0] ? 4'hc : _GEN_35379; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35381 = 10'h38 == _T_509[9:0] ? 4'hc : _GEN_35380; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35382 = 10'h39 == _T_509[9:0] ? 4'hc : _GEN_35381; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35383 = 10'h3a == _T_509[9:0] ? 4'hc : _GEN_35382; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35384 = 10'h3b == _T_509[9:0] ? 4'hc : _GEN_35383; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35385 = 10'h3c == _T_509[9:0] ? 4'h7 : _GEN_35384; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35386 = 10'h3d == _T_509[9:0] ? 4'h9 : _GEN_35385; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35387 = 10'h3e == _T_509[9:0] ? 4'h8 : _GEN_35386; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35388 = 10'h3f == _T_509[9:0] ? 4'hc : _GEN_35387; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35389 = 10'h40 == _T_509[9:0] ? 4'hc : _GEN_35388; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35390 = 10'h41 == _T_509[9:0] ? 4'hc : _GEN_35389; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35391 = 10'h42 == _T_509[9:0] ? 4'hc : _GEN_35390; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35392 = 10'h43 == _T_509[9:0] ? 4'hc : _GEN_35391; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35393 = 10'h44 == _T_509[9:0] ? 4'hc : _GEN_35392; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35394 = 10'h45 == _T_509[9:0] ? 4'hc : _GEN_35393; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35395 = 10'h46 == _T_509[9:0] ? 4'hc : _GEN_35394; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35396 = 10'h47 == _T_509[9:0] ? 4'hc : _GEN_35395; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35397 = 10'h48 == _T_509[9:0] ? 4'hc : _GEN_35396; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35398 = 10'h49 == _T_509[9:0] ? 4'hc : _GEN_35397; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35399 = 10'h4a == _T_509[9:0] ? 4'hc : _GEN_35398; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35400 = 10'h4b == _T_509[9:0] ? 4'hc : _GEN_35399; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35401 = 10'h4c == _T_509[9:0] ? 4'hc : _GEN_35400; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35402 = 10'h4d == _T_509[9:0] ? 4'hc : _GEN_35401; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35403 = 10'h4e == _T_509[9:0] ? 4'hc : _GEN_35402; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35404 = 10'h4f == _T_509[9:0] ? 4'hc : _GEN_35403; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35405 = 10'h50 == _T_509[9:0] ? 4'hc : _GEN_35404; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35406 = 10'h51 == _T_509[9:0] ? 4'hc : _GEN_35405; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35407 = 10'h52 == _T_509[9:0] ? 4'hc : _GEN_35406; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35408 = 10'h53 == _T_509[9:0] ? 4'hc : _GEN_35407; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35409 = 10'h54 == _T_509[9:0] ? 4'hc : _GEN_35408; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35410 = 10'h55 == _T_509[9:0] ? 4'hc : _GEN_35409; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35411 = 10'h56 == _T_509[9:0] ? 4'hc : _GEN_35410; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35412 = 10'h57 == _T_509[9:0] ? 4'hc : _GEN_35411; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35413 = 10'h58 == _T_509[9:0] ? 4'hc : _GEN_35412; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35414 = 10'h59 == _T_509[9:0] ? 4'hc : _GEN_35413; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35415 = 10'h5a == _T_509[9:0] ? 4'h9 : _GEN_35414; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35416 = 10'h5b == _T_509[9:0] ? 4'ha : _GEN_35415; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35417 = 10'h5c == _T_509[9:0] ? 4'hc : _GEN_35416; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35418 = 10'h5d == _T_509[9:0] ? 4'hc : _GEN_35417; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35419 = 10'h5e == _T_509[9:0] ? 4'hc : _GEN_35418; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35420 = 10'h5f == _T_509[9:0] ? 4'hc : _GEN_35419; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35421 = 10'h60 == _T_509[9:0] ? 4'hc : _GEN_35420; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35422 = 10'h61 == _T_509[9:0] ? 4'hb : _GEN_35421; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35423 = 10'h62 == _T_509[9:0] ? 4'h8 : _GEN_35422; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35424 = 10'h63 == _T_509[9:0] ? 4'h9 : _GEN_35423; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35425 = 10'h64 == _T_509[9:0] ? 4'h7 : _GEN_35424; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35426 = 10'h65 == _T_509[9:0] ? 4'hb : _GEN_35425; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35427 = 10'h66 == _T_509[9:0] ? 4'hc : _GEN_35426; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35428 = 10'h67 == _T_509[9:0] ? 4'hc : _GEN_35427; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35429 = 10'h68 == _T_509[9:0] ? 4'hc : _GEN_35428; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35430 = 10'h69 == _T_509[9:0] ? 4'hc : _GEN_35429; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35431 = 10'h6a == _T_509[9:0] ? 4'hc : _GEN_35430; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35432 = 10'h6b == _T_509[9:0] ? 4'hb : _GEN_35431; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35433 = 10'h6c == _T_509[9:0] ? 4'h9 : _GEN_35432; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35434 = 10'h6d == _T_509[9:0] ? 4'ha : _GEN_35433; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35435 = 10'h6e == _T_509[9:0] ? 4'hc : _GEN_35434; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35436 = 10'h6f == _T_509[9:0] ? 4'hc : _GEN_35435; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35437 = 10'h70 == _T_509[9:0] ? 4'hc : _GEN_35436; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35438 = 10'h71 == _T_509[9:0] ? 4'hc : _GEN_35437; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35439 = 10'h72 == _T_509[9:0] ? 4'hc : _GEN_35438; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35440 = 10'h73 == _T_509[9:0] ? 4'hc : _GEN_35439; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35441 = 10'h74 == _T_509[9:0] ? 4'hc : _GEN_35440; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35442 = 10'h75 == _T_509[9:0] ? 4'hc : _GEN_35441; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35443 = 10'h76 == _T_509[9:0] ? 4'hc : _GEN_35442; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35444 = 10'h77 == _T_509[9:0] ? 4'hc : _GEN_35443; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35445 = 10'h78 == _T_509[9:0] ? 4'hc : _GEN_35444; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35446 = 10'h79 == _T_509[9:0] ? 4'hc : _GEN_35445; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35447 = 10'h7a == _T_509[9:0] ? 4'hc : _GEN_35446; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35448 = 10'h7b == _T_509[9:0] ? 4'hc : _GEN_35447; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35449 = 10'h7c == _T_509[9:0] ? 4'hc : _GEN_35448; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35450 = 10'h7d == _T_509[9:0] ? 4'hc : _GEN_35449; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35451 = 10'h7e == _T_509[9:0] ? 4'hc : _GEN_35450; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35452 = 10'h7f == _T_509[9:0] ? 4'hc : _GEN_35451; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35453 = 10'h80 == _T_509[9:0] ? 4'hc : _GEN_35452; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35454 = 10'h81 == _T_509[9:0] ? 4'h9 : _GEN_35453; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35455 = 10'h82 == _T_509[9:0] ? 4'h9 : _GEN_35454; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35456 = 10'h83 == _T_509[9:0] ? 4'h9 : _GEN_35455; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35457 = 10'h84 == _T_509[9:0] ? 4'hc : _GEN_35456; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35458 = 10'h85 == _T_509[9:0] ? 4'hc : _GEN_35457; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35459 = 10'h86 == _T_509[9:0] ? 4'hc : _GEN_35458; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35460 = 10'h87 == _T_509[9:0] ? 4'h8 : _GEN_35459; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35461 = 10'h88 == _T_509[9:0] ? 4'h9 : _GEN_35460; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35462 = 10'h89 == _T_509[9:0] ? 4'h9 : _GEN_35461; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35463 = 10'h8a == _T_509[9:0] ? 4'h9 : _GEN_35462; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35464 = 10'h8b == _T_509[9:0] ? 4'hc : _GEN_35463; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35465 = 10'h8c == _T_509[9:0] ? 4'hc : _GEN_35464; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35466 = 10'h8d == _T_509[9:0] ? 4'hc : _GEN_35465; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35467 = 10'h8e == _T_509[9:0] ? 4'hc : _GEN_35466; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35468 = 10'h8f == _T_509[9:0] ? 4'h9 : _GEN_35467; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35469 = 10'h90 == _T_509[9:0] ? 4'h9 : _GEN_35468; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35470 = 10'h91 == _T_509[9:0] ? 4'h9 : _GEN_35469; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35471 = 10'h92 == _T_509[9:0] ? 4'ha : _GEN_35470; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35472 = 10'h93 == _T_509[9:0] ? 4'hc : _GEN_35471; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35473 = 10'h94 == _T_509[9:0] ? 4'hc : _GEN_35472; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35474 = 10'h95 == _T_509[9:0] ? 4'hc : _GEN_35473; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35475 = 10'h96 == _T_509[9:0] ? 4'hc : _GEN_35474; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35476 = 10'h97 == _T_509[9:0] ? 4'hc : _GEN_35475; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35477 = 10'h98 == _T_509[9:0] ? 4'hc : _GEN_35476; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35478 = 10'h99 == _T_509[9:0] ? 4'hc : _GEN_35477; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35479 = 10'h9a == _T_509[9:0] ? 4'hc : _GEN_35478; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35480 = 10'h9b == _T_509[9:0] ? 4'hc : _GEN_35479; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35481 = 10'h9c == _T_509[9:0] ? 4'hc : _GEN_35480; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35482 = 10'h9d == _T_509[9:0] ? 4'hc : _GEN_35481; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35483 = 10'h9e == _T_509[9:0] ? 4'hc : _GEN_35482; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35484 = 10'h9f == _T_509[9:0] ? 4'hc : _GEN_35483; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35485 = 10'ha0 == _T_509[9:0] ? 4'hc : _GEN_35484; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35486 = 10'ha1 == _T_509[9:0] ? 4'hc : _GEN_35485; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35487 = 10'ha2 == _T_509[9:0] ? 4'hc : _GEN_35486; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35488 = 10'ha3 == _T_509[9:0] ? 4'hc : _GEN_35487; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35489 = 10'ha4 == _T_509[9:0] ? 4'hc : _GEN_35488; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35490 = 10'ha5 == _T_509[9:0] ? 4'hc : _GEN_35489; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35491 = 10'ha6 == _T_509[9:0] ? 4'hc : _GEN_35490; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35492 = 10'ha7 == _T_509[9:0] ? 4'hc : _GEN_35491; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35493 = 10'ha8 == _T_509[9:0] ? 4'h9 : _GEN_35492; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35494 = 10'ha9 == _T_509[9:0] ? 4'h8 : _GEN_35493; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35495 = 10'haa == _T_509[9:0] ? 4'h8 : _GEN_35494; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35496 = 10'hab == _T_509[9:0] ? 4'ha : _GEN_35495; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35497 = 10'hac == _T_509[9:0] ? 4'hb : _GEN_35496; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35498 = 10'had == _T_509[9:0] ? 4'h7 : _GEN_35497; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35499 = 10'hae == _T_509[9:0] ? 4'h9 : _GEN_35498; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35500 = 10'haf == _T_509[9:0] ? 4'h9 : _GEN_35499; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35501 = 10'hb0 == _T_509[9:0] ? 4'h8 : _GEN_35500; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35502 = 10'hb1 == _T_509[9:0] ? 4'h9 : _GEN_35501; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35503 = 10'hb2 == _T_509[9:0] ? 4'hc : _GEN_35502; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35504 = 10'hb3 == _T_509[9:0] ? 4'h9 : _GEN_35503; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35505 = 10'hb4 == _T_509[9:0] ? 4'h9 : _GEN_35504; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35506 = 10'hb5 == _T_509[9:0] ? 4'h9 : _GEN_35505; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35507 = 10'hb6 == _T_509[9:0] ? 4'h9 : _GEN_35506; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35508 = 10'hb7 == _T_509[9:0] ? 4'ha : _GEN_35507; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35509 = 10'hb8 == _T_509[9:0] ? 4'hc : _GEN_35508; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35510 = 10'hb9 == _T_509[9:0] ? 4'hc : _GEN_35509; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35511 = 10'hba == _T_509[9:0] ? 4'hc : _GEN_35510; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35512 = 10'hbb == _T_509[9:0] ? 4'hc : _GEN_35511; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35513 = 10'hbc == _T_509[9:0] ? 4'hc : _GEN_35512; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35514 = 10'hbd == _T_509[9:0] ? 4'hb : _GEN_35513; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35515 = 10'hbe == _T_509[9:0] ? 4'hc : _GEN_35514; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35516 = 10'hbf == _T_509[9:0] ? 4'hc : _GEN_35515; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35517 = 10'hc0 == _T_509[9:0] ? 4'hc : _GEN_35516; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35518 = 10'hc1 == _T_509[9:0] ? 4'hc : _GEN_35517; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35519 = 10'hc2 == _T_509[9:0] ? 4'hc : _GEN_35518; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35520 = 10'hc3 == _T_509[9:0] ? 4'hc : _GEN_35519; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35521 = 10'hc4 == _T_509[9:0] ? 4'hc : _GEN_35520; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35522 = 10'hc5 == _T_509[9:0] ? 4'hc : _GEN_35521; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35523 = 10'hc6 == _T_509[9:0] ? 4'hb : _GEN_35522; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35524 = 10'hc7 == _T_509[9:0] ? 4'hb : _GEN_35523; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35525 = 10'hc8 == _T_509[9:0] ? 4'ha : _GEN_35524; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35526 = 10'hc9 == _T_509[9:0] ? 4'ha : _GEN_35525; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35527 = 10'hca == _T_509[9:0] ? 4'hb : _GEN_35526; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35528 = 10'hcb == _T_509[9:0] ? 4'hc : _GEN_35527; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35529 = 10'hcc == _T_509[9:0] ? 4'hc : _GEN_35528; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35530 = 10'hcd == _T_509[9:0] ? 4'hc : _GEN_35529; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35531 = 10'hce == _T_509[9:0] ? 4'ha : _GEN_35530; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35532 = 10'hcf == _T_509[9:0] ? 4'h8 : _GEN_35531; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35533 = 10'hd0 == _T_509[9:0] ? 4'h9 : _GEN_35532; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35534 = 10'hd1 == _T_509[9:0] ? 4'h8 : _GEN_35533; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35535 = 10'hd2 == _T_509[9:0] ? 4'h9 : _GEN_35534; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35536 = 10'hd3 == _T_509[9:0] ? 4'h9 : _GEN_35535; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35537 = 10'hd4 == _T_509[9:0] ? 4'h9 : _GEN_35536; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35538 = 10'hd5 == _T_509[9:0] ? 4'h9 : _GEN_35537; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35539 = 10'hd6 == _T_509[9:0] ? 4'ha : _GEN_35538; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35540 = 10'hd7 == _T_509[9:0] ? 4'h9 : _GEN_35539; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35541 = 10'hd8 == _T_509[9:0] ? 4'h9 : _GEN_35540; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35542 = 10'hd9 == _T_509[9:0] ? 4'h9 : _GEN_35541; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35543 = 10'hda == _T_509[9:0] ? 4'ha : _GEN_35542; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35544 = 10'hdb == _T_509[9:0] ? 4'h9 : _GEN_35543; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35545 = 10'hdc == _T_509[9:0] ? 4'h7 : _GEN_35544; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35546 = 10'hdd == _T_509[9:0] ? 4'hc : _GEN_35545; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35547 = 10'hde == _T_509[9:0] ? 4'hc : _GEN_35546; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35548 = 10'hdf == _T_509[9:0] ? 4'hc : _GEN_35547; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35549 = 10'he0 == _T_509[9:0] ? 4'hc : _GEN_35548; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35550 = 10'he1 == _T_509[9:0] ? 4'hc : _GEN_35549; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35551 = 10'he2 == _T_509[9:0] ? 4'hc : _GEN_35550; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35552 = 10'he3 == _T_509[9:0] ? 4'h8 : _GEN_35551; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35553 = 10'he4 == _T_509[9:0] ? 4'hc : _GEN_35552; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35554 = 10'he5 == _T_509[9:0] ? 4'hc : _GEN_35553; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35555 = 10'he6 == _T_509[9:0] ? 4'hc : _GEN_35554; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35556 = 10'he7 == _T_509[9:0] ? 4'hc : _GEN_35555; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35557 = 10'he8 == _T_509[9:0] ? 4'hc : _GEN_35556; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35558 = 10'he9 == _T_509[9:0] ? 4'hc : _GEN_35557; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35559 = 10'hea == _T_509[9:0] ? 4'hc : _GEN_35558; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35560 = 10'heb == _T_509[9:0] ? 4'ha : _GEN_35559; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35561 = 10'hec == _T_509[9:0] ? 4'h7 : _GEN_35560; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35562 = 10'hed == _T_509[9:0] ? 4'h3 : _GEN_35561; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35563 = 10'hee == _T_509[9:0] ? 4'h3 : _GEN_35562; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35564 = 10'hef == _T_509[9:0] ? 4'h3 : _GEN_35563; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35565 = 10'hf0 == _T_509[9:0] ? 4'h3 : _GEN_35564; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35566 = 10'hf1 == _T_509[9:0] ? 4'h8 : _GEN_35565; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35567 = 10'hf2 == _T_509[9:0] ? 4'hc : _GEN_35566; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35568 = 10'hf3 == _T_509[9:0] ? 4'hc : _GEN_35567; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35569 = 10'hf4 == _T_509[9:0] ? 4'hc : _GEN_35568; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35570 = 10'hf5 == _T_509[9:0] ? 4'h9 : _GEN_35569; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35571 = 10'hf6 == _T_509[9:0] ? 4'h9 : _GEN_35570; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35572 = 10'hf7 == _T_509[9:0] ? 4'h9 : _GEN_35571; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35573 = 10'hf8 == _T_509[9:0] ? 4'h9 : _GEN_35572; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35574 = 10'hf9 == _T_509[9:0] ? 4'ha : _GEN_35573; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35575 = 10'hfa == _T_509[9:0] ? 4'h9 : _GEN_35574; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35576 = 10'hfb == _T_509[9:0] ? 4'h9 : _GEN_35575; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35577 = 10'hfc == _T_509[9:0] ? 4'h9 : _GEN_35576; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35578 = 10'hfd == _T_509[9:0] ? 4'h9 : _GEN_35577; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35579 = 10'hfe == _T_509[9:0] ? 4'h9 : _GEN_35578; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35580 = 10'hff == _T_509[9:0] ? 4'ha : _GEN_35579; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35581 = 10'h100 == _T_509[9:0] ? 4'ha : _GEN_35580; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35582 = 10'h101 == _T_509[9:0] ? 4'h7 : _GEN_35581; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35583 = 10'h102 == _T_509[9:0] ? 4'h9 : _GEN_35582; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35584 = 10'h103 == _T_509[9:0] ? 4'hc : _GEN_35583; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35585 = 10'h104 == _T_509[9:0] ? 4'hc : _GEN_35584; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35586 = 10'h105 == _T_509[9:0] ? 4'hb : _GEN_35585; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35587 = 10'h106 == _T_509[9:0] ? 4'hb : _GEN_35586; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35588 = 10'h107 == _T_509[9:0] ? 4'hb : _GEN_35587; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35589 = 10'h108 == _T_509[9:0] ? 4'hb : _GEN_35588; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35590 = 10'h109 == _T_509[9:0] ? 4'h7 : _GEN_35589; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35591 = 10'h10a == _T_509[9:0] ? 4'hc : _GEN_35590; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35592 = 10'h10b == _T_509[9:0] ? 4'hc : _GEN_35591; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35593 = 10'h10c == _T_509[9:0] ? 4'hc : _GEN_35592; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35594 = 10'h10d == _T_509[9:0] ? 4'hc : _GEN_35593; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35595 = 10'h10e == _T_509[9:0] ? 4'hc : _GEN_35594; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35596 = 10'h10f == _T_509[9:0] ? 4'h9 : _GEN_35595; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35597 = 10'h110 == _T_509[9:0] ? 4'hb : _GEN_35596; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35598 = 10'h111 == _T_509[9:0] ? 4'h4 : _GEN_35597; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35599 = 10'h112 == _T_509[9:0] ? 4'h7 : _GEN_35598; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35600 = 10'h113 == _T_509[9:0] ? 4'h3 : _GEN_35599; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35601 = 10'h114 == _T_509[9:0] ? 4'h3 : _GEN_35600; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35602 = 10'h115 == _T_509[9:0] ? 4'h3 : _GEN_35601; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35603 = 10'h116 == _T_509[9:0] ? 4'h3 : _GEN_35602; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35604 = 10'h117 == _T_509[9:0] ? 4'h2 : _GEN_35603; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35605 = 10'h118 == _T_509[9:0] ? 4'h9 : _GEN_35604; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35606 = 10'h119 == _T_509[9:0] ? 4'hc : _GEN_35605; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35607 = 10'h11a == _T_509[9:0] ? 4'hc : _GEN_35606; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35608 = 10'h11b == _T_509[9:0] ? 4'hc : _GEN_35607; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35609 = 10'h11c == _T_509[9:0] ? 4'h9 : _GEN_35608; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35610 = 10'h11d == _T_509[9:0] ? 4'h9 : _GEN_35609; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35611 = 10'h11e == _T_509[9:0] ? 4'h9 : _GEN_35610; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35612 = 10'h11f == _T_509[9:0] ? 4'h8 : _GEN_35611; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35613 = 10'h120 == _T_509[9:0] ? 4'h7 : _GEN_35612; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35614 = 10'h121 == _T_509[9:0] ? 4'h9 : _GEN_35613; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35615 = 10'h122 == _T_509[9:0] ? 4'h7 : _GEN_35614; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35616 = 10'h123 == _T_509[9:0] ? 4'h7 : _GEN_35615; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35617 = 10'h124 == _T_509[9:0] ? 4'h9 : _GEN_35616; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35618 = 10'h125 == _T_509[9:0] ? 4'h9 : _GEN_35617; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35619 = 10'h126 == _T_509[9:0] ? 4'h8 : _GEN_35618; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35620 = 10'h127 == _T_509[9:0] ? 4'h9 : _GEN_35619; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35621 = 10'h128 == _T_509[9:0] ? 4'h8 : _GEN_35620; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35622 = 10'h129 == _T_509[9:0] ? 4'ha : _GEN_35621; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35623 = 10'h12a == _T_509[9:0] ? 4'h5 : _GEN_35622; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35624 = 10'h12b == _T_509[9:0] ? 4'h3 : _GEN_35623; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35625 = 10'h12c == _T_509[9:0] ? 4'h3 : _GEN_35624; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35626 = 10'h12d == _T_509[9:0] ? 4'h3 : _GEN_35625; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35627 = 10'h12e == _T_509[9:0] ? 4'h5 : _GEN_35626; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35628 = 10'h12f == _T_509[9:0] ? 4'h8 : _GEN_35627; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35629 = 10'h130 == _T_509[9:0] ? 4'hc : _GEN_35628; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35630 = 10'h131 == _T_509[9:0] ? 4'hb : _GEN_35629; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35631 = 10'h132 == _T_509[9:0] ? 4'h9 : _GEN_35630; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35632 = 10'h133 == _T_509[9:0] ? 4'h8 : _GEN_35631; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35633 = 10'h134 == _T_509[9:0] ? 4'h9 : _GEN_35632; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35634 = 10'h135 == _T_509[9:0] ? 4'h7 : _GEN_35633; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35635 = 10'h136 == _T_509[9:0] ? 4'h7 : _GEN_35634; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35636 = 10'h137 == _T_509[9:0] ? 4'h5 : _GEN_35635; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35637 = 10'h138 == _T_509[9:0] ? 4'h7 : _GEN_35636; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35638 = 10'h139 == _T_509[9:0] ? 4'h3 : _GEN_35637; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35639 = 10'h13a == _T_509[9:0] ? 4'h3 : _GEN_35638; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35640 = 10'h13b == _T_509[9:0] ? 4'h3 : _GEN_35639; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35641 = 10'h13c == _T_509[9:0] ? 4'h3 : _GEN_35640; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35642 = 10'h13d == _T_509[9:0] ? 4'h3 : _GEN_35641; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35643 = 10'h13e == _T_509[9:0] ? 4'h5 : _GEN_35642; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35644 = 10'h13f == _T_509[9:0] ? 4'ha : _GEN_35643; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35645 = 10'h140 == _T_509[9:0] ? 4'hc : _GEN_35644; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35646 = 10'h141 == _T_509[9:0] ? 4'hc : _GEN_35645; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35647 = 10'h142 == _T_509[9:0] ? 4'hc : _GEN_35646; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35648 = 10'h143 == _T_509[9:0] ? 4'h9 : _GEN_35647; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35649 = 10'h144 == _T_509[9:0] ? 4'h9 : _GEN_35648; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35650 = 10'h145 == _T_509[9:0] ? 4'h8 : _GEN_35649; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35651 = 10'h146 == _T_509[9:0] ? 4'h8 : _GEN_35650; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35652 = 10'h147 == _T_509[9:0] ? 4'h7 : _GEN_35651; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35653 = 10'h148 == _T_509[9:0] ? 4'h8 : _GEN_35652; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35654 = 10'h149 == _T_509[9:0] ? 4'h9 : _GEN_35653; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35655 = 10'h14a == _T_509[9:0] ? 4'ha : _GEN_35654; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35656 = 10'h14b == _T_509[9:0] ? 4'h9 : _GEN_35655; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35657 = 10'h14c == _T_509[9:0] ? 4'ha : _GEN_35656; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35658 = 10'h14d == _T_509[9:0] ? 4'h9 : _GEN_35657; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35659 = 10'h14e == _T_509[9:0] ? 4'h7 : _GEN_35658; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35660 = 10'h14f == _T_509[9:0] ? 4'h3 : _GEN_35659; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35661 = 10'h150 == _T_509[9:0] ? 4'h3 : _GEN_35660; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35662 = 10'h151 == _T_509[9:0] ? 4'h3 : _GEN_35661; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35663 = 10'h152 == _T_509[9:0] ? 4'h3 : _GEN_35662; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35664 = 10'h153 == _T_509[9:0] ? 4'h3 : _GEN_35663; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35665 = 10'h154 == _T_509[9:0] ? 4'h3 : _GEN_35664; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35666 = 10'h155 == _T_509[9:0] ? 4'h8 : _GEN_35665; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35667 = 10'h156 == _T_509[9:0] ? 4'ha : _GEN_35666; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35668 = 10'h157 == _T_509[9:0] ? 4'h7 : _GEN_35667; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35669 = 10'h158 == _T_509[9:0] ? 4'h7 : _GEN_35668; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35670 = 10'h159 == _T_509[9:0] ? 4'h7 : _GEN_35669; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35671 = 10'h15a == _T_509[9:0] ? 4'h7 : _GEN_35670; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35672 = 10'h15b == _T_509[9:0] ? 4'h7 : _GEN_35671; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35673 = 10'h15c == _T_509[9:0] ? 4'h7 : _GEN_35672; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35674 = 10'h15d == _T_509[9:0] ? 4'h7 : _GEN_35673; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35675 = 10'h15e == _T_509[9:0] ? 4'h7 : _GEN_35674; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35676 = 10'h15f == _T_509[9:0] ? 4'h3 : _GEN_35675; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35677 = 10'h160 == _T_509[9:0] ? 4'h3 : _GEN_35676; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35678 = 10'h161 == _T_509[9:0] ? 4'h3 : _GEN_35677; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35679 = 10'h162 == _T_509[9:0] ? 4'h3 : _GEN_35678; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35680 = 10'h163 == _T_509[9:0] ? 4'h3 : _GEN_35679; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35681 = 10'h164 == _T_509[9:0] ? 4'h4 : _GEN_35680; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35682 = 10'h165 == _T_509[9:0] ? 4'ha : _GEN_35681; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35683 = 10'h166 == _T_509[9:0] ? 4'ha : _GEN_35682; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35684 = 10'h167 == _T_509[9:0] ? 4'hc : _GEN_35683; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35685 = 10'h168 == _T_509[9:0] ? 4'hc : _GEN_35684; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35686 = 10'h169 == _T_509[9:0] ? 4'h9 : _GEN_35685; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35687 = 10'h16a == _T_509[9:0] ? 4'h9 : _GEN_35686; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35688 = 10'h16b == _T_509[9:0] ? 4'ha : _GEN_35687; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35689 = 10'h16c == _T_509[9:0] ? 4'h7 : _GEN_35688; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35690 = 10'h16d == _T_509[9:0] ? 4'h7 : _GEN_35689; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35691 = 10'h16e == _T_509[9:0] ? 4'h7 : _GEN_35690; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35692 = 10'h16f == _T_509[9:0] ? 4'ha : _GEN_35691; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35693 = 10'h170 == _T_509[9:0] ? 4'ha : _GEN_35692; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35694 = 10'h171 == _T_509[9:0] ? 4'ha : _GEN_35693; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35695 = 10'h172 == _T_509[9:0] ? 4'hc : _GEN_35694; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35696 = 10'h173 == _T_509[9:0] ? 4'h8 : _GEN_35695; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35697 = 10'h174 == _T_509[9:0] ? 4'h5 : _GEN_35696; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35698 = 10'h175 == _T_509[9:0] ? 4'h8 : _GEN_35697; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35699 = 10'h176 == _T_509[9:0] ? 4'h7 : _GEN_35698; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35700 = 10'h177 == _T_509[9:0] ? 4'h8 : _GEN_35699; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35701 = 10'h178 == _T_509[9:0] ? 4'h7 : _GEN_35700; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35702 = 10'h179 == _T_509[9:0] ? 4'h5 : _GEN_35701; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35703 = 10'h17a == _T_509[9:0] ? 4'h5 : _GEN_35702; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35704 = 10'h17b == _T_509[9:0] ? 4'h7 : _GEN_35703; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35705 = 10'h17c == _T_509[9:0] ? 4'h7 : _GEN_35704; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35706 = 10'h17d == _T_509[9:0] ? 4'h7 : _GEN_35705; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35707 = 10'h17e == _T_509[9:0] ? 4'h7 : _GEN_35706; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35708 = 10'h17f == _T_509[9:0] ? 4'h7 : _GEN_35707; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35709 = 10'h180 == _T_509[9:0] ? 4'h7 : _GEN_35708; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35710 = 10'h181 == _T_509[9:0] ? 4'h7 : _GEN_35709; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35711 = 10'h182 == _T_509[9:0] ? 4'h7 : _GEN_35710; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35712 = 10'h183 == _T_509[9:0] ? 4'h7 : _GEN_35711; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35713 = 10'h184 == _T_509[9:0] ? 4'h7 : _GEN_35712; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35714 = 10'h185 == _T_509[9:0] ? 4'h5 : _GEN_35713; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35715 = 10'h186 == _T_509[9:0] ? 4'h3 : _GEN_35714; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35716 = 10'h187 == _T_509[9:0] ? 4'h3 : _GEN_35715; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35717 = 10'h188 == _T_509[9:0] ? 4'h3 : _GEN_35716; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35718 = 10'h189 == _T_509[9:0] ? 4'h4 : _GEN_35717; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35719 = 10'h18a == _T_509[9:0] ? 4'h5 : _GEN_35718; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35720 = 10'h18b == _T_509[9:0] ? 4'ha : _GEN_35719; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35721 = 10'h18c == _T_509[9:0] ? 4'ha : _GEN_35720; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35722 = 10'h18d == _T_509[9:0] ? 4'ha : _GEN_35721; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35723 = 10'h18e == _T_509[9:0] ? 4'hc : _GEN_35722; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35724 = 10'h18f == _T_509[9:0] ? 4'h8 : _GEN_35723; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35725 = 10'h190 == _T_509[9:0] ? 4'h9 : _GEN_35724; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35726 = 10'h191 == _T_509[9:0] ? 4'h8 : _GEN_35725; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35727 = 10'h192 == _T_509[9:0] ? 4'h7 : _GEN_35726; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35728 = 10'h193 == _T_509[9:0] ? 4'h7 : _GEN_35727; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35729 = 10'h194 == _T_509[9:0] ? 4'h7 : _GEN_35728; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35730 = 10'h195 == _T_509[9:0] ? 4'h9 : _GEN_35729; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35731 = 10'h196 == _T_509[9:0] ? 4'ha : _GEN_35730; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35732 = 10'h197 == _T_509[9:0] ? 4'h8 : _GEN_35731; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35733 = 10'h198 == _T_509[9:0] ? 4'hc : _GEN_35732; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35734 = 10'h199 == _T_509[9:0] ? 4'h5 : _GEN_35733; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35735 = 10'h19a == _T_509[9:0] ? 4'h1 : _GEN_35734; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35736 = 10'h19b == _T_509[9:0] ? 4'h4 : _GEN_35735; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35737 = 10'h19c == _T_509[9:0] ? 4'h7 : _GEN_35736; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35738 = 10'h19d == _T_509[9:0] ? 4'h5 : _GEN_35737; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35739 = 10'h19e == _T_509[9:0] ? 4'h2 : _GEN_35738; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35740 = 10'h19f == _T_509[9:0] ? 4'h3 : _GEN_35739; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35741 = 10'h1a0 == _T_509[9:0] ? 4'h7 : _GEN_35740; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35742 = 10'h1a1 == _T_509[9:0] ? 4'h7 : _GEN_35741; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35743 = 10'h1a2 == _T_509[9:0] ? 4'h7 : _GEN_35742; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35744 = 10'h1a3 == _T_509[9:0] ? 4'h7 : _GEN_35743; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35745 = 10'h1a4 == _T_509[9:0] ? 4'h7 : _GEN_35744; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35746 = 10'h1a5 == _T_509[9:0] ? 4'h7 : _GEN_35745; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35747 = 10'h1a6 == _T_509[9:0] ? 4'h7 : _GEN_35746; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35748 = 10'h1a7 == _T_509[9:0] ? 4'h7 : _GEN_35747; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35749 = 10'h1a8 == _T_509[9:0] ? 4'h8 : _GEN_35748; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35750 = 10'h1a9 == _T_509[9:0] ? 4'h8 : _GEN_35749; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35751 = 10'h1aa == _T_509[9:0] ? 4'h6 : _GEN_35750; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35752 = 10'h1ab == _T_509[9:0] ? 4'h6 : _GEN_35751; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35753 = 10'h1ac == _T_509[9:0] ? 4'h5 : _GEN_35752; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35754 = 10'h1ad == _T_509[9:0] ? 4'h4 : _GEN_35753; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35755 = 10'h1ae == _T_509[9:0] ? 4'h3 : _GEN_35754; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35756 = 10'h1af == _T_509[9:0] ? 4'h6 : _GEN_35755; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35757 = 10'h1b0 == _T_509[9:0] ? 4'h6 : _GEN_35756; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35758 = 10'h1b1 == _T_509[9:0] ? 4'ha : _GEN_35757; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35759 = 10'h1b2 == _T_509[9:0] ? 4'ha : _GEN_35758; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35760 = 10'h1b3 == _T_509[9:0] ? 4'h9 : _GEN_35759; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35761 = 10'h1b4 == _T_509[9:0] ? 4'hb : _GEN_35760; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35762 = 10'h1b5 == _T_509[9:0] ? 4'h8 : _GEN_35761; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35763 = 10'h1b6 == _T_509[9:0] ? 4'h8 : _GEN_35762; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35764 = 10'h1b7 == _T_509[9:0] ? 4'h7 : _GEN_35763; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35765 = 10'h1b8 == _T_509[9:0] ? 4'h6 : _GEN_35764; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35766 = 10'h1b9 == _T_509[9:0] ? 4'h7 : _GEN_35765; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35767 = 10'h1ba == _T_509[9:0] ? 4'h6 : _GEN_35766; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35768 = 10'h1bb == _T_509[9:0] ? 4'h8 : _GEN_35767; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35769 = 10'h1bc == _T_509[9:0] ? 4'ha : _GEN_35768; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35770 = 10'h1bd == _T_509[9:0] ? 4'h9 : _GEN_35769; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35771 = 10'h1be == _T_509[9:0] ? 4'hc : _GEN_35770; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35772 = 10'h1bf == _T_509[9:0] ? 4'h7 : _GEN_35771; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35773 = 10'h1c0 == _T_509[9:0] ? 4'h6 : _GEN_35772; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35774 = 10'h1c1 == _T_509[9:0] ? 4'h7 : _GEN_35773; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35775 = 10'h1c2 == _T_509[9:0] ? 4'h7 : _GEN_35774; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35776 = 10'h1c3 == _T_509[9:0] ? 4'h6 : _GEN_35775; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35777 = 10'h1c4 == _T_509[9:0] ? 4'h5 : _GEN_35776; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35778 = 10'h1c5 == _T_509[9:0] ? 4'h6 : _GEN_35777; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35779 = 10'h1c6 == _T_509[9:0] ? 4'h8 : _GEN_35778; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35780 = 10'h1c7 == _T_509[9:0] ? 4'h7 : _GEN_35779; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35781 = 10'h1c8 == _T_509[9:0] ? 4'h7 : _GEN_35780; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35782 = 10'h1c9 == _T_509[9:0] ? 4'h7 : _GEN_35781; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35783 = 10'h1ca == _T_509[9:0] ? 4'h7 : _GEN_35782; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35784 = 10'h1cb == _T_509[9:0] ? 4'h7 : _GEN_35783; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35785 = 10'h1cc == _T_509[9:0] ? 4'h7 : _GEN_35784; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35786 = 10'h1cd == _T_509[9:0] ? 4'h8 : _GEN_35785; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35787 = 10'h1ce == _T_509[9:0] ? 4'h8 : _GEN_35786; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35788 = 10'h1cf == _T_509[9:0] ? 4'h8 : _GEN_35787; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35789 = 10'h1d0 == _T_509[9:0] ? 4'h5 : _GEN_35788; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35790 = 10'h1d1 == _T_509[9:0] ? 4'h6 : _GEN_35789; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35791 = 10'h1d2 == _T_509[9:0] ? 4'h7 : _GEN_35790; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35792 = 10'h1d3 == _T_509[9:0] ? 4'h7 : _GEN_35791; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35793 = 10'h1d4 == _T_509[9:0] ? 4'h7 : _GEN_35792; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35794 = 10'h1d5 == _T_509[9:0] ? 4'h6 : _GEN_35793; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35795 = 10'h1d6 == _T_509[9:0] ? 4'h8 : _GEN_35794; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35796 = 10'h1d7 == _T_509[9:0] ? 4'ha : _GEN_35795; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35797 = 10'h1d8 == _T_509[9:0] ? 4'ha : _GEN_35796; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35798 = 10'h1d9 == _T_509[9:0] ? 4'ha : _GEN_35797; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35799 = 10'h1da == _T_509[9:0] ? 4'h8 : _GEN_35798; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35800 = 10'h1db == _T_509[9:0] ? 4'h9 : _GEN_35799; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35801 = 10'h1dc == _T_509[9:0] ? 4'h9 : _GEN_35800; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35802 = 10'h1dd == _T_509[9:0] ? 4'h5 : _GEN_35801; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35803 = 10'h1de == _T_509[9:0] ? 4'h7 : _GEN_35802; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35804 = 10'h1df == _T_509[9:0] ? 4'h7 : _GEN_35803; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35805 = 10'h1e0 == _T_509[9:0] ? 4'h7 : _GEN_35804; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35806 = 10'h1e1 == _T_509[9:0] ? 4'h6 : _GEN_35805; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35807 = 10'h1e2 == _T_509[9:0] ? 4'h9 : _GEN_35806; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35808 = 10'h1e3 == _T_509[9:0] ? 4'h9 : _GEN_35807; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35809 = 10'h1e4 == _T_509[9:0] ? 4'hb : _GEN_35808; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35810 = 10'h1e5 == _T_509[9:0] ? 4'h8 : _GEN_35809; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35811 = 10'h1e6 == _T_509[9:0] ? 4'h7 : _GEN_35810; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35812 = 10'h1e7 == _T_509[9:0] ? 4'h8 : _GEN_35811; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35813 = 10'h1e8 == _T_509[9:0] ? 4'h8 : _GEN_35812; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35814 = 10'h1e9 == _T_509[9:0] ? 4'h8 : _GEN_35813; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35815 = 10'h1ea == _T_509[9:0] ? 4'h8 : _GEN_35814; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35816 = 10'h1eb == _T_509[9:0] ? 4'h8 : _GEN_35815; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35817 = 10'h1ec == _T_509[9:0] ? 4'h8 : _GEN_35816; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35818 = 10'h1ed == _T_509[9:0] ? 4'h6 : _GEN_35817; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35819 = 10'h1ee == _T_509[9:0] ? 4'h7 : _GEN_35818; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35820 = 10'h1ef == _T_509[9:0] ? 4'h7 : _GEN_35819; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35821 = 10'h1f0 == _T_509[9:0] ? 4'h7 : _GEN_35820; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35822 = 10'h1f1 == _T_509[9:0] ? 4'h7 : _GEN_35821; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35823 = 10'h1f2 == _T_509[9:0] ? 4'h7 : _GEN_35822; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35824 = 10'h1f3 == _T_509[9:0] ? 4'h8 : _GEN_35823; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35825 = 10'h1f4 == _T_509[9:0] ? 4'h8 : _GEN_35824; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35826 = 10'h1f5 == _T_509[9:0] ? 4'h8 : _GEN_35825; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35827 = 10'h1f6 == _T_509[9:0] ? 4'ha : _GEN_35826; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35828 = 10'h1f7 == _T_509[9:0] ? 4'h6 : _GEN_35827; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35829 = 10'h1f8 == _T_509[9:0] ? 4'h6 : _GEN_35828; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35830 = 10'h1f9 == _T_509[9:0] ? 4'h8 : _GEN_35829; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35831 = 10'h1fa == _T_509[9:0] ? 4'h8 : _GEN_35830; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35832 = 10'h1fb == _T_509[9:0] ? 4'h6 : _GEN_35831; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35833 = 10'h1fc == _T_509[9:0] ? 4'ha : _GEN_35832; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35834 = 10'h1fd == _T_509[9:0] ? 4'hb : _GEN_35833; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35835 = 10'h1fe == _T_509[9:0] ? 4'ha : _GEN_35834; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35836 = 10'h1ff == _T_509[9:0] ? 4'ha : _GEN_35835; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35837 = 10'h200 == _T_509[9:0] ? 4'h4 : _GEN_35836; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35838 = 10'h201 == _T_509[9:0] ? 4'h7 : _GEN_35837; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35839 = 10'h202 == _T_509[9:0] ? 4'h6 : _GEN_35838; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35840 = 10'h203 == _T_509[9:0] ? 4'h6 : _GEN_35839; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35841 = 10'h204 == _T_509[9:0] ? 4'h5 : _GEN_35840; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35842 = 10'h205 == _T_509[9:0] ? 4'h6 : _GEN_35841; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35843 = 10'h206 == _T_509[9:0] ? 4'h6 : _GEN_35842; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35844 = 10'h207 == _T_509[9:0] ? 4'h5 : _GEN_35843; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35845 = 10'h208 == _T_509[9:0] ? 4'h7 : _GEN_35844; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35846 = 10'h209 == _T_509[9:0] ? 4'h9 : _GEN_35845; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35847 = 10'h20a == _T_509[9:0] ? 4'hb : _GEN_35846; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35848 = 10'h20b == _T_509[9:0] ? 4'h7 : _GEN_35847; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35849 = 10'h20c == _T_509[9:0] ? 4'h7 : _GEN_35848; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35850 = 10'h20d == _T_509[9:0] ? 4'h7 : _GEN_35849; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35851 = 10'h20e == _T_509[9:0] ? 4'h7 : _GEN_35850; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35852 = 10'h20f == _T_509[9:0] ? 4'h7 : _GEN_35851; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35853 = 10'h210 == _T_509[9:0] ? 4'h7 : _GEN_35852; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35854 = 10'h211 == _T_509[9:0] ? 4'h8 : _GEN_35853; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35855 = 10'h212 == _T_509[9:0] ? 4'h8 : _GEN_35854; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35856 = 10'h213 == _T_509[9:0] ? 4'h9 : _GEN_35855; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35857 = 10'h214 == _T_509[9:0] ? 4'h6 : _GEN_35856; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35858 = 10'h215 == _T_509[9:0] ? 4'h7 : _GEN_35857; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35859 = 10'h216 == _T_509[9:0] ? 4'h7 : _GEN_35858; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35860 = 10'h217 == _T_509[9:0] ? 4'h7 : _GEN_35859; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35861 = 10'h218 == _T_509[9:0] ? 4'h7 : _GEN_35860; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35862 = 10'h219 == _T_509[9:0] ? 4'h8 : _GEN_35861; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35863 = 10'h21a == _T_509[9:0] ? 4'h7 : _GEN_35862; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35864 = 10'h21b == _T_509[9:0] ? 4'h8 : _GEN_35863; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35865 = 10'h21c == _T_509[9:0] ? 4'ha : _GEN_35864; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35866 = 10'h21d == _T_509[9:0] ? 4'ha : _GEN_35865; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35867 = 10'h21e == _T_509[9:0] ? 4'h7 : _GEN_35866; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35868 = 10'h21f == _T_509[9:0] ? 4'h6 : _GEN_35867; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35869 = 10'h220 == _T_509[9:0] ? 4'h6 : _GEN_35868; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35870 = 10'h221 == _T_509[9:0] ? 4'h7 : _GEN_35869; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35871 = 10'h222 == _T_509[9:0] ? 4'ha : _GEN_35870; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35872 = 10'h223 == _T_509[9:0] ? 4'ha : _GEN_35871; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35873 = 10'h224 == _T_509[9:0] ? 4'ha : _GEN_35872; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35874 = 10'h225 == _T_509[9:0] ? 4'h8 : _GEN_35873; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35875 = 10'h226 == _T_509[9:0] ? 4'h3 : _GEN_35874; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35876 = 10'h227 == _T_509[9:0] ? 4'h4 : _GEN_35875; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35877 = 10'h228 == _T_509[9:0] ? 4'h6 : _GEN_35876; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35878 = 10'h229 == _T_509[9:0] ? 4'h6 : _GEN_35877; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35879 = 10'h22a == _T_509[9:0] ? 4'h6 : _GEN_35878; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35880 = 10'h22b == _T_509[9:0] ? 4'h6 : _GEN_35879; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35881 = 10'h22c == _T_509[9:0] ? 4'h5 : _GEN_35880; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35882 = 10'h22d == _T_509[9:0] ? 4'h6 : _GEN_35881; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35883 = 10'h22e == _T_509[9:0] ? 4'h6 : _GEN_35882; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35884 = 10'h22f == _T_509[9:0] ? 4'h8 : _GEN_35883; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35885 = 10'h230 == _T_509[9:0] ? 4'h7 : _GEN_35884; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35886 = 10'h231 == _T_509[9:0] ? 4'h5 : _GEN_35885; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35887 = 10'h232 == _T_509[9:0] ? 4'h6 : _GEN_35886; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35888 = 10'h233 == _T_509[9:0] ? 4'h8 : _GEN_35887; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35889 = 10'h234 == _T_509[9:0] ? 4'h8 : _GEN_35888; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35890 = 10'h235 == _T_509[9:0] ? 4'h8 : _GEN_35889; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35891 = 10'h236 == _T_509[9:0] ? 4'h8 : _GEN_35890; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35892 = 10'h237 == _T_509[9:0] ? 4'h8 : _GEN_35891; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35893 = 10'h238 == _T_509[9:0] ? 4'h8 : _GEN_35892; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35894 = 10'h239 == _T_509[9:0] ? 4'h6 : _GEN_35893; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35895 = 10'h23a == _T_509[9:0] ? 4'h6 : _GEN_35894; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35896 = 10'h23b == _T_509[9:0] ? 4'h7 : _GEN_35895; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35897 = 10'h23c == _T_509[9:0] ? 4'h6 : _GEN_35896; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35898 = 10'h23d == _T_509[9:0] ? 4'h7 : _GEN_35897; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35899 = 10'h23e == _T_509[9:0] ? 4'h7 : _GEN_35898; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35900 = 10'h23f == _T_509[9:0] ? 4'h6 : _GEN_35899; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35901 = 10'h240 == _T_509[9:0] ? 4'h6 : _GEN_35900; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35902 = 10'h241 == _T_509[9:0] ? 4'h8 : _GEN_35901; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35903 = 10'h242 == _T_509[9:0] ? 4'ha : _GEN_35902; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35904 = 10'h243 == _T_509[9:0] ? 4'ha : _GEN_35903; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35905 = 10'h244 == _T_509[9:0] ? 4'ha : _GEN_35904; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35906 = 10'h245 == _T_509[9:0] ? 4'h8 : _GEN_35905; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35907 = 10'h246 == _T_509[9:0] ? 4'h8 : _GEN_35906; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35908 = 10'h247 == _T_509[9:0] ? 4'h9 : _GEN_35907; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35909 = 10'h248 == _T_509[9:0] ? 4'ha : _GEN_35908; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35910 = 10'h249 == _T_509[9:0] ? 4'ha : _GEN_35909; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35911 = 10'h24a == _T_509[9:0] ? 4'ha : _GEN_35910; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35912 = 10'h24b == _T_509[9:0] ? 4'h4 : _GEN_35911; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35913 = 10'h24c == _T_509[9:0] ? 4'h3 : _GEN_35912; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35914 = 10'h24d == _T_509[9:0] ? 4'h4 : _GEN_35913; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35915 = 10'h24e == _T_509[9:0] ? 4'h5 : _GEN_35914; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35916 = 10'h24f == _T_509[9:0] ? 4'h5 : _GEN_35915; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35917 = 10'h250 == _T_509[9:0] ? 4'h5 : _GEN_35916; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35918 = 10'h251 == _T_509[9:0] ? 4'h5 : _GEN_35917; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35919 = 10'h252 == _T_509[9:0] ? 4'h5 : _GEN_35918; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35920 = 10'h253 == _T_509[9:0] ? 4'h5 : _GEN_35919; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35921 = 10'h254 == _T_509[9:0] ? 4'h5 : _GEN_35920; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35922 = 10'h255 == _T_509[9:0] ? 4'h6 : _GEN_35921; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35923 = 10'h256 == _T_509[9:0] ? 4'h7 : _GEN_35922; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35924 = 10'h257 == _T_509[9:0] ? 4'h3 : _GEN_35923; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35925 = 10'h258 == _T_509[9:0] ? 4'h6 : _GEN_35924; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35926 = 10'h259 == _T_509[9:0] ? 4'h7 : _GEN_35925; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35927 = 10'h25a == _T_509[9:0] ? 4'h7 : _GEN_35926; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35928 = 10'h25b == _T_509[9:0] ? 4'h7 : _GEN_35927; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35929 = 10'h25c == _T_509[9:0] ? 4'h8 : _GEN_35928; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35930 = 10'h25d == _T_509[9:0] ? 4'h8 : _GEN_35929; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35931 = 10'h25e == _T_509[9:0] ? 4'h4 : _GEN_35930; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35932 = 10'h25f == _T_509[9:0] ? 4'h3 : _GEN_35931; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35933 = 10'h260 == _T_509[9:0] ? 4'h7 : _GEN_35932; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35934 = 10'h261 == _T_509[9:0] ? 4'h7 : _GEN_35933; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35935 = 10'h262 == _T_509[9:0] ? 4'h7 : _GEN_35934; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35936 = 10'h263 == _T_509[9:0] ? 4'h6 : _GEN_35935; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35937 = 10'h264 == _T_509[9:0] ? 4'h7 : _GEN_35936; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35938 = 10'h265 == _T_509[9:0] ? 4'h6 : _GEN_35937; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35939 = 10'h266 == _T_509[9:0] ? 4'h5 : _GEN_35938; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35940 = 10'h267 == _T_509[9:0] ? 4'h7 : _GEN_35939; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35941 = 10'h268 == _T_509[9:0] ? 4'ha : _GEN_35940; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35942 = 10'h269 == _T_509[9:0] ? 4'ha : _GEN_35941; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35943 = 10'h26a == _T_509[9:0] ? 4'ha : _GEN_35942; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35944 = 10'h26b == _T_509[9:0] ? 4'ha : _GEN_35943; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35945 = 10'h26c == _T_509[9:0] ? 4'ha : _GEN_35944; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35946 = 10'h26d == _T_509[9:0] ? 4'ha : _GEN_35945; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35947 = 10'h26e == _T_509[9:0] ? 4'ha : _GEN_35946; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35948 = 10'h26f == _T_509[9:0] ? 4'ha : _GEN_35947; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35949 = 10'h270 == _T_509[9:0] ? 4'h5 : _GEN_35948; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35950 = 10'h271 == _T_509[9:0] ? 4'h3 : _GEN_35949; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35951 = 10'h272 == _T_509[9:0] ? 4'h3 : _GEN_35950; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35952 = 10'h273 == _T_509[9:0] ? 4'h4 : _GEN_35951; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35953 = 10'h274 == _T_509[9:0] ? 4'h6 : _GEN_35952; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35954 = 10'h275 == _T_509[9:0] ? 4'h5 : _GEN_35953; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35955 = 10'h276 == _T_509[9:0] ? 4'h6 : _GEN_35954; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35956 = 10'h277 == _T_509[9:0] ? 4'h5 : _GEN_35955; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35957 = 10'h278 == _T_509[9:0] ? 4'h6 : _GEN_35956; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35958 = 10'h279 == _T_509[9:0] ? 4'h6 : _GEN_35957; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35959 = 10'h27a == _T_509[9:0] ? 4'h6 : _GEN_35958; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35960 = 10'h27b == _T_509[9:0] ? 4'h8 : _GEN_35959; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35961 = 10'h27c == _T_509[9:0] ? 4'h6 : _GEN_35960; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35962 = 10'h27d == _T_509[9:0] ? 4'h2 : _GEN_35961; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35963 = 10'h27e == _T_509[9:0] ? 4'h5 : _GEN_35962; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35964 = 10'h27f == _T_509[9:0] ? 4'h7 : _GEN_35963; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35965 = 10'h280 == _T_509[9:0] ? 4'h7 : _GEN_35964; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35966 = 10'h281 == _T_509[9:0] ? 4'h8 : _GEN_35965; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35967 = 10'h282 == _T_509[9:0] ? 4'h7 : _GEN_35966; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35968 = 10'h283 == _T_509[9:0] ? 4'h3 : _GEN_35967; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35969 = 10'h284 == _T_509[9:0] ? 4'h3 : _GEN_35968; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35970 = 10'h285 == _T_509[9:0] ? 4'h3 : _GEN_35969; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35971 = 10'h286 == _T_509[9:0] ? 4'h7 : _GEN_35970; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35972 = 10'h287 == _T_509[9:0] ? 4'h7 : _GEN_35971; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35973 = 10'h288 == _T_509[9:0] ? 4'h7 : _GEN_35972; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35974 = 10'h289 == _T_509[9:0] ? 4'h7 : _GEN_35973; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35975 = 10'h28a == _T_509[9:0] ? 4'h8 : _GEN_35974; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35976 = 10'h28b == _T_509[9:0] ? 4'h8 : _GEN_35975; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35977 = 10'h28c == _T_509[9:0] ? 4'h7 : _GEN_35976; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35978 = 10'h28d == _T_509[9:0] ? 4'h6 : _GEN_35977; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35979 = 10'h28e == _T_509[9:0] ? 4'h3 : _GEN_35978; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35980 = 10'h28f == _T_509[9:0] ? 4'h6 : _GEN_35979; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35981 = 10'h290 == _T_509[9:0] ? 4'h8 : _GEN_35980; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35982 = 10'h291 == _T_509[9:0] ? 4'ha : _GEN_35981; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35983 = 10'h292 == _T_509[9:0] ? 4'ha : _GEN_35982; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35984 = 10'h293 == _T_509[9:0] ? 4'ha : _GEN_35983; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35985 = 10'h294 == _T_509[9:0] ? 4'h9 : _GEN_35984; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35986 = 10'h295 == _T_509[9:0] ? 4'h4 : _GEN_35985; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35987 = 10'h296 == _T_509[9:0] ? 4'h3 : _GEN_35986; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35988 = 10'h297 == _T_509[9:0] ? 4'h3 : _GEN_35987; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35989 = 10'h298 == _T_509[9:0] ? 4'h3 : _GEN_35988; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35990 = 10'h299 == _T_509[9:0] ? 4'h4 : _GEN_35989; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35991 = 10'h29a == _T_509[9:0] ? 4'h5 : _GEN_35990; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35992 = 10'h29b == _T_509[9:0] ? 4'h5 : _GEN_35991; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35993 = 10'h29c == _T_509[9:0] ? 4'h5 : _GEN_35992; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35994 = 10'h29d == _T_509[9:0] ? 4'h5 : _GEN_35993; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35995 = 10'h29e == _T_509[9:0] ? 4'h5 : _GEN_35994; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35996 = 10'h29f == _T_509[9:0] ? 4'h5 : _GEN_35995; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35997 = 10'h2a0 == _T_509[9:0] ? 4'h6 : _GEN_35996; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35998 = 10'h2a1 == _T_509[9:0] ? 4'h7 : _GEN_35997; // @[Filter.scala 230:142]
  wire [3:0] _GEN_35999 = 10'h2a2 == _T_509[9:0] ? 4'h5 : _GEN_35998; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36000 = 10'h2a3 == _T_509[9:0] ? 4'h2 : _GEN_35999; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36001 = 10'h2a4 == _T_509[9:0] ? 4'h3 : _GEN_36000; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36002 = 10'h2a5 == _T_509[9:0] ? 4'h7 : _GEN_36001; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36003 = 10'h2a6 == _T_509[9:0] ? 4'h8 : _GEN_36002; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36004 = 10'h2a7 == _T_509[9:0] ? 4'h7 : _GEN_36003; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36005 = 10'h2a8 == _T_509[9:0] ? 4'h3 : _GEN_36004; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36006 = 10'h2a9 == _T_509[9:0] ? 4'h2 : _GEN_36005; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36007 = 10'h2aa == _T_509[9:0] ? 4'h3 : _GEN_36006; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36008 = 10'h2ab == _T_509[9:0] ? 4'h3 : _GEN_36007; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36009 = 10'h2ac == _T_509[9:0] ? 4'h7 : _GEN_36008; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36010 = 10'h2ad == _T_509[9:0] ? 4'h8 : _GEN_36009; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36011 = 10'h2ae == _T_509[9:0] ? 4'h7 : _GEN_36010; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36012 = 10'h2af == _T_509[9:0] ? 4'h8 : _GEN_36011; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36013 = 10'h2b0 == _T_509[9:0] ? 4'h8 : _GEN_36012; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36014 = 10'h2b1 == _T_509[9:0] ? 4'h8 : _GEN_36013; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36015 = 10'h2b2 == _T_509[9:0] ? 4'h7 : _GEN_36014; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36016 = 10'h2b3 == _T_509[9:0] ? 4'h6 : _GEN_36015; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36017 = 10'h2b4 == _T_509[9:0] ? 4'h2 : _GEN_36016; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36018 = 10'h2b5 == _T_509[9:0] ? 4'h2 : _GEN_36017; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36019 = 10'h2b6 == _T_509[9:0] ? 4'h3 : _GEN_36018; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36020 = 10'h2b7 == _T_509[9:0] ? 4'h3 : _GEN_36019; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36021 = 10'h2b8 == _T_509[9:0] ? 4'h6 : _GEN_36020; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36022 = 10'h2b9 == _T_509[9:0] ? 4'h9 : _GEN_36021; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36023 = 10'h2ba == _T_509[9:0] ? 4'h3 : _GEN_36022; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36024 = 10'h2bb == _T_509[9:0] ? 4'h3 : _GEN_36023; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36025 = 10'h2bc == _T_509[9:0] ? 4'h3 : _GEN_36024; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36026 = 10'h2bd == _T_509[9:0] ? 4'h2 : _GEN_36025; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36027 = 10'h2be == _T_509[9:0] ? 4'h3 : _GEN_36026; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36028 = 10'h2bf == _T_509[9:0] ? 4'h3 : _GEN_36027; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36029 = 10'h2c0 == _T_509[9:0] ? 4'h5 : _GEN_36028; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36030 = 10'h2c1 == _T_509[9:0] ? 4'h5 : _GEN_36029; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36031 = 10'h2c2 == _T_509[9:0] ? 4'h5 : _GEN_36030; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36032 = 10'h2c3 == _T_509[9:0] ? 4'h5 : _GEN_36031; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36033 = 10'h2c4 == _T_509[9:0] ? 4'h5 : _GEN_36032; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36034 = 10'h2c5 == _T_509[9:0] ? 4'h5 : _GEN_36033; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36035 = 10'h2c6 == _T_509[9:0] ? 4'h6 : _GEN_36034; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36036 = 10'h2c7 == _T_509[9:0] ? 4'h7 : _GEN_36035; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36037 = 10'h2c8 == _T_509[9:0] ? 4'h5 : _GEN_36036; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36038 = 10'h2c9 == _T_509[9:0] ? 4'h2 : _GEN_36037; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36039 = 10'h2ca == _T_509[9:0] ? 4'h2 : _GEN_36038; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36040 = 10'h2cb == _T_509[9:0] ? 4'h3 : _GEN_36039; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36041 = 10'h2cc == _T_509[9:0] ? 4'h3 : _GEN_36040; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36042 = 10'h2cd == _T_509[9:0] ? 4'h2 : _GEN_36041; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36043 = 10'h2ce == _T_509[9:0] ? 4'h2 : _GEN_36042; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36044 = 10'h2cf == _T_509[9:0] ? 4'h2 : _GEN_36043; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36045 = 10'h2d0 == _T_509[9:0] ? 4'h2 : _GEN_36044; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36046 = 10'h2d1 == _T_509[9:0] ? 4'h2 : _GEN_36045; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36047 = 10'h2d2 == _T_509[9:0] ? 4'h7 : _GEN_36046; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36048 = 10'h2d3 == _T_509[9:0] ? 4'h7 : _GEN_36047; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36049 = 10'h2d4 == _T_509[9:0] ? 4'h8 : _GEN_36048; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36050 = 10'h2d5 == _T_509[9:0] ? 4'h8 : _GEN_36049; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36051 = 10'h2d6 == _T_509[9:0] ? 4'h8 : _GEN_36050; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36052 = 10'h2d7 == _T_509[9:0] ? 4'h8 : _GEN_36051; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36053 = 10'h2d8 == _T_509[9:0] ? 4'h7 : _GEN_36052; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36054 = 10'h2d9 == _T_509[9:0] ? 4'h6 : _GEN_36053; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36055 = 10'h2da == _T_509[9:0] ? 4'h4 : _GEN_36054; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36056 = 10'h2db == _T_509[9:0] ? 4'h2 : _GEN_36055; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36057 = 10'h2dc == _T_509[9:0] ? 4'h2 : _GEN_36056; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36058 = 10'h2dd == _T_509[9:0] ? 4'h3 : _GEN_36057; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36059 = 10'h2de == _T_509[9:0] ? 4'h3 : _GEN_36058; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36060 = 10'h2df == _T_509[9:0] ? 4'h3 : _GEN_36059; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36061 = 10'h2e0 == _T_509[9:0] ? 4'h3 : _GEN_36060; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36062 = 10'h2e1 == _T_509[9:0] ? 4'h3 : _GEN_36061; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36063 = 10'h2e2 == _T_509[9:0] ? 4'h3 : _GEN_36062; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36064 = 10'h2e3 == _T_509[9:0] ? 4'h2 : _GEN_36063; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36065 = 10'h2e4 == _T_509[9:0] ? 4'h3 : _GEN_36064; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36066 = 10'h2e5 == _T_509[9:0] ? 4'h2 : _GEN_36065; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36067 = 10'h2e6 == _T_509[9:0] ? 4'h5 : _GEN_36066; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36068 = 10'h2e7 == _T_509[9:0] ? 4'h5 : _GEN_36067; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36069 = 10'h2e8 == _T_509[9:0] ? 4'h5 : _GEN_36068; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36070 = 10'h2e9 == _T_509[9:0] ? 4'h5 : _GEN_36069; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36071 = 10'h2ea == _T_509[9:0] ? 4'h5 : _GEN_36070; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36072 = 10'h2eb == _T_509[9:0] ? 4'h5 : _GEN_36071; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36073 = 10'h2ec == _T_509[9:0] ? 4'h6 : _GEN_36072; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36074 = 10'h2ed == _T_509[9:0] ? 4'h7 : _GEN_36073; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36075 = 10'h2ee == _T_509[9:0] ? 4'h6 : _GEN_36074; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36076 = 10'h2ef == _T_509[9:0] ? 4'h2 : _GEN_36075; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36077 = 10'h2f0 == _T_509[9:0] ? 4'h2 : _GEN_36076; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36078 = 10'h2f1 == _T_509[9:0] ? 4'h2 : _GEN_36077; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36079 = 10'h2f2 == _T_509[9:0] ? 4'h2 : _GEN_36078; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36080 = 10'h2f3 == _T_509[9:0] ? 4'h2 : _GEN_36079; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36081 = 10'h2f4 == _T_509[9:0] ? 4'h2 : _GEN_36080; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36082 = 10'h2f5 == _T_509[9:0] ? 4'h2 : _GEN_36081; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36083 = 10'h2f6 == _T_509[9:0] ? 4'h2 : _GEN_36082; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36084 = 10'h2f7 == _T_509[9:0] ? 4'h2 : _GEN_36083; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36085 = 10'h2f8 == _T_509[9:0] ? 4'h7 : _GEN_36084; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36086 = 10'h2f9 == _T_509[9:0] ? 4'h7 : _GEN_36085; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36087 = 10'h2fa == _T_509[9:0] ? 4'h8 : _GEN_36086; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36088 = 10'h2fb == _T_509[9:0] ? 4'h8 : _GEN_36087; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36089 = 10'h2fc == _T_509[9:0] ? 4'h7 : _GEN_36088; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36090 = 10'h2fd == _T_509[9:0] ? 4'h7 : _GEN_36089; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36091 = 10'h2fe == _T_509[9:0] ? 4'h7 : _GEN_36090; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36092 = 10'h2ff == _T_509[9:0] ? 4'h7 : _GEN_36091; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36093 = 10'h300 == _T_509[9:0] ? 4'h8 : _GEN_36092; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36094 = 10'h301 == _T_509[9:0] ? 4'h7 : _GEN_36093; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36095 = 10'h302 == _T_509[9:0] ? 4'h3 : _GEN_36094; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36096 = 10'h303 == _T_509[9:0] ? 4'h3 : _GEN_36095; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36097 = 10'h304 == _T_509[9:0] ? 4'h2 : _GEN_36096; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36098 = 10'h305 == _T_509[9:0] ? 4'h2 : _GEN_36097; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36099 = 10'h306 == _T_509[9:0] ? 4'h2 : _GEN_36098; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36100 = 10'h307 == _T_509[9:0] ? 4'h2 : _GEN_36099; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36101 = 10'h308 == _T_509[9:0] ? 4'h2 : _GEN_36100; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36102 = 10'h309 == _T_509[9:0] ? 4'h2 : _GEN_36101; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36103 = 10'h30a == _T_509[9:0] ? 4'h2 : _GEN_36102; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36104 = 10'h30b == _T_509[9:0] ? 4'h3 : _GEN_36103; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36105 = 10'h30c == _T_509[9:0] ? 4'h4 : _GEN_36104; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36106 = 10'h30d == _T_509[9:0] ? 4'h5 : _GEN_36105; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36107 = 10'h30e == _T_509[9:0] ? 4'h5 : _GEN_36106; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36108 = 10'h30f == _T_509[9:0] ? 4'h5 : _GEN_36107; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36109 = 10'h310 == _T_509[9:0] ? 4'h5 : _GEN_36108; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36110 = 10'h311 == _T_509[9:0] ? 4'h5 : _GEN_36109; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36111 = 10'h312 == _T_509[9:0] ? 4'h6 : _GEN_36110; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36112 = 10'h313 == _T_509[9:0] ? 4'h7 : _GEN_36111; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36113 = 10'h314 == _T_509[9:0] ? 4'h7 : _GEN_36112; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36114 = 10'h315 == _T_509[9:0] ? 4'h3 : _GEN_36113; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36115 = 10'h316 == _T_509[9:0] ? 4'h2 : _GEN_36114; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36116 = 10'h317 == _T_509[9:0] ? 4'h2 : _GEN_36115; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36117 = 10'h318 == _T_509[9:0] ? 4'h2 : _GEN_36116; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36118 = 10'h319 == _T_509[9:0] ? 4'h2 : _GEN_36117; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36119 = 10'h31a == _T_509[9:0] ? 4'h2 : _GEN_36118; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36120 = 10'h31b == _T_509[9:0] ? 4'h2 : _GEN_36119; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36121 = 10'h31c == _T_509[9:0] ? 4'h2 : _GEN_36120; // @[Filter.scala 230:142]
  wire [3:0] _GEN_36122 = 10'h31d == _T_509[9:0] ? 4'h2 : _GEN_36121; // @[Filter.scala 230:142]
  wire [7:0] _T_523 = _GEN_36122 * 4'ha; // @[Filter.scala 230:142]
  wire [10:0] _GEN_39043 = {{3'd0}, _T_523}; // @[Filter.scala 230:109]
  wire [10:0] _T_525 = _T_518 + _GEN_39043; // @[Filter.scala 230:109]
  wire [10:0] _T_526 = _T_525 / 11'h64; // @[Filter.scala 230:150]
  wire  _T_528 = _T_499 >= 6'h20; // @[Filter.scala 233:31]
  wire  _T_532 = _T_506 >= 32'h12; // @[Filter.scala 233:63]
  wire  _T_533 = _T_528 | _T_532; // @[Filter.scala 233:58]
  wire [10:0] _GEN_36921 = io_SPI_distort ? _T_526 : {{7'd0}, _GEN_34526}; // @[Filter.scala 235:35]
  wire [10:0] _GEN_36922 = _T_533 ? 11'h0 : _GEN_36921; // @[Filter.scala 233:80]
  wire [10:0] _GEN_37721 = io_SPI_distort ? _T_526 : {{7'd0}, _GEN_35324}; // @[Filter.scala 235:35]
  wire [10:0] _GEN_37722 = _T_533 ? 11'h0 : _GEN_37721; // @[Filter.scala 233:80]
  wire [10:0] _GEN_38521 = io_SPI_distort ? _T_526 : {{7'd0}, _GEN_36122}; // @[Filter.scala 235:35]
  wire [10:0] _GEN_38522 = _T_533 ? 11'h0 : _GEN_38521; // @[Filter.scala 233:80]
  reg [8:0] pixOut_0_0; // @[Filter.scala 244:32]
  reg [8:0] pixOut_0_1; // @[Filter.scala 244:32]
  reg [8:0] pixOut_0_2; // @[Filter.scala 244:32]
  reg [8:0] pixOut_0_3; // @[Filter.scala 244:32]
  reg [8:0] pixOut_0_4; // @[Filter.scala 244:32]
  reg [8:0] pixOut_0_5; // @[Filter.scala 244:32]
  reg [8:0] pixOut_0_6; // @[Filter.scala 244:32]
  reg [8:0] pixOut_0_7; // @[Filter.scala 244:32]
  reg [8:0] pixOut_1_0; // @[Filter.scala 244:87]
  reg [8:0] pixOut_1_1; // @[Filter.scala 244:87]
  reg [8:0] pixOut_1_2; // @[Filter.scala 244:87]
  reg [8:0] pixOut_1_3; // @[Filter.scala 244:87]
  reg [8:0] pixOut_1_4; // @[Filter.scala 244:87]
  reg [8:0] pixOut_1_5; // @[Filter.scala 244:87]
  reg [8:0] pixOut_1_6; // @[Filter.scala 244:87]
  reg [8:0] pixOut_1_7; // @[Filter.scala 244:87]
  reg [8:0] pixOut_2_0; // @[Filter.scala 244:142]
  reg [8:0] pixOut_2_1; // @[Filter.scala 244:142]
  reg [8:0] pixOut_2_2; // @[Filter.scala 244:142]
  reg [8:0] pixOut_2_3; // @[Filter.scala 244:142]
  reg [8:0] pixOut_2_4; // @[Filter.scala 244:142]
  reg [8:0] pixOut_2_5; // @[Filter.scala 244:142]
  reg [8:0] pixOut_2_6; // @[Filter.scala 244:142]
  reg [8:0] pixOut_2_7; // @[Filter.scala 244:142]
  reg  validOut; // @[Filter.scala 245:29]
  wire [7:0] _GEN_38524 = 3'h1 == io_SPI_filterIndex[2:0] ? $signed(8'sh9) : $signed(8'sh1); // @[Filter.scala 249:64]
  wire [7:0] _GEN_38525 = 3'h2 == io_SPI_filterIndex[2:0] ? $signed(8'sh10) : $signed(_GEN_38524); // @[Filter.scala 249:64]
  wire [7:0] _GEN_38526 = 3'h3 == io_SPI_filterIndex[2:0] ? $signed(8'sh1) : $signed(_GEN_38525); // @[Filter.scala 249:64]
  wire [7:0] _GEN_38527 = 3'h4 == io_SPI_filterIndex[2:0] ? $signed(8'sh1) : $signed(_GEN_38526); // @[Filter.scala 249:64]
  wire [7:0] _GEN_38528 = 3'h5 == io_SPI_filterIndex[2:0] ? $signed(8'sh1) : $signed(_GEN_38527); // @[Filter.scala 249:64]
  wire [8:0] _GEN_39047 = {{1{_GEN_38528[7]}},_GEN_38528}; // @[Filter.scala 249:64]
  wire [9:0] _T_564 = $signed(KernelConvolution_io_pixelVal_out_0) / $signed(_GEN_39047); // @[Filter.scala 249:64]
  wire  _T_565 = $signed(pixOut_0_0) < 9'sh0; // @[Filter.scala 251:30]
  wire  _T_568 = $signed(pixOut_0_0) > 9'shf; // @[Filter.scala 256:36]
  wire [8:0] _GEN_38530 = _T_568 ? 9'hf : pixOut_0_0; // @[Filter.scala 258:44]
  wire [8:0] _GEN_38532 = _T_565 ? 9'h0 : _GEN_38530; // @[Filter.scala 253:43]
  wire [9:0] _T_575 = $signed(KernelConvolution_io_pixelVal_out_1) / $signed(_GEN_39047); // @[Filter.scala 249:64]
  wire  _T_576 = $signed(pixOut_0_1) < 9'sh0; // @[Filter.scala 251:30]
  wire  _T_579 = $signed(pixOut_0_1) > 9'shf; // @[Filter.scala 256:36]
  wire [8:0] _GEN_38535 = _T_579 ? 9'hf : pixOut_0_1; // @[Filter.scala 258:44]
  wire [8:0] _GEN_38537 = _T_576 ? 9'h0 : _GEN_38535; // @[Filter.scala 253:43]
  wire [9:0] _T_586 = $signed(KernelConvolution_io_pixelVal_out_2) / $signed(_GEN_39047); // @[Filter.scala 249:64]
  wire  _T_587 = $signed(pixOut_0_2) < 9'sh0; // @[Filter.scala 251:30]
  wire  _T_590 = $signed(pixOut_0_2) > 9'shf; // @[Filter.scala 256:36]
  wire [8:0] _GEN_38540 = _T_590 ? 9'hf : pixOut_0_2; // @[Filter.scala 258:44]
  wire [8:0] _GEN_38542 = _T_587 ? 9'h0 : _GEN_38540; // @[Filter.scala 253:43]
  wire [9:0] _T_597 = $signed(KernelConvolution_io_pixelVal_out_3) / $signed(_GEN_39047); // @[Filter.scala 249:64]
  wire  _T_598 = $signed(pixOut_0_3) < 9'sh0; // @[Filter.scala 251:30]
  wire  _T_601 = $signed(pixOut_0_3) > 9'shf; // @[Filter.scala 256:36]
  wire [8:0] _GEN_38545 = _T_601 ? 9'hf : pixOut_0_3; // @[Filter.scala 258:44]
  wire [8:0] _GEN_38547 = _T_598 ? 9'h0 : _GEN_38545; // @[Filter.scala 253:43]
  wire [9:0] _T_608 = $signed(KernelConvolution_io_pixelVal_out_4) / $signed(_GEN_39047); // @[Filter.scala 249:64]
  wire  _T_609 = $signed(pixOut_0_4) < 9'sh0; // @[Filter.scala 251:30]
  wire  _T_612 = $signed(pixOut_0_4) > 9'shf; // @[Filter.scala 256:36]
  wire [8:0] _GEN_38550 = _T_612 ? 9'hf : pixOut_0_4; // @[Filter.scala 258:44]
  wire [8:0] _GEN_38552 = _T_609 ? 9'h0 : _GEN_38550; // @[Filter.scala 253:43]
  wire [9:0] _T_619 = $signed(KernelConvolution_io_pixelVal_out_5) / $signed(_GEN_39047); // @[Filter.scala 249:64]
  wire  _T_620 = $signed(pixOut_0_5) < 9'sh0; // @[Filter.scala 251:30]
  wire  _T_623 = $signed(pixOut_0_5) > 9'shf; // @[Filter.scala 256:36]
  wire [8:0] _GEN_38555 = _T_623 ? 9'hf : pixOut_0_5; // @[Filter.scala 258:44]
  wire [8:0] _GEN_38557 = _T_620 ? 9'h0 : _GEN_38555; // @[Filter.scala 253:43]
  wire [9:0] _T_630 = $signed(KernelConvolution_io_pixelVal_out_6) / $signed(_GEN_39047); // @[Filter.scala 249:64]
  wire  _T_631 = $signed(pixOut_0_6) < 9'sh0; // @[Filter.scala 251:30]
  wire  _T_634 = $signed(pixOut_0_6) > 9'shf; // @[Filter.scala 256:36]
  wire [8:0] _GEN_38560 = _T_634 ? 9'hf : pixOut_0_6; // @[Filter.scala 258:44]
  wire [8:0] _GEN_38562 = _T_631 ? 9'h0 : _GEN_38560; // @[Filter.scala 253:43]
  wire [9:0] _T_641 = $signed(KernelConvolution_io_pixelVal_out_7) / $signed(_GEN_39047); // @[Filter.scala 249:64]
  wire  _T_642 = $signed(pixOut_0_7) < 9'sh0; // @[Filter.scala 251:30]
  wire  _T_645 = $signed(pixOut_0_7) > 9'shf; // @[Filter.scala 256:36]
  wire [8:0] _GEN_38565 = _T_645 ? 9'hf : pixOut_0_7; // @[Filter.scala 258:44]
  wire [8:0] _GEN_38567 = _T_642 ? 9'h0 : _GEN_38565; // @[Filter.scala 253:43]
  wire [9:0] _T_652 = $signed(KernelConvolution_1_io_pixelVal_out_0) / $signed(_GEN_39047); // @[Filter.scala 249:64]
  wire  _T_653 = $signed(pixOut_1_0) < 9'sh0; // @[Filter.scala 251:30]
  wire  _T_656 = $signed(pixOut_1_0) > 9'shf; // @[Filter.scala 256:36]
  wire [8:0] _GEN_38570 = _T_656 ? 9'hf : pixOut_1_0; // @[Filter.scala 258:44]
  wire [8:0] _GEN_38572 = _T_653 ? 9'h0 : _GEN_38570; // @[Filter.scala 253:43]
  wire [9:0] _T_663 = $signed(KernelConvolution_1_io_pixelVal_out_1) / $signed(_GEN_39047); // @[Filter.scala 249:64]
  wire  _T_664 = $signed(pixOut_1_1) < 9'sh0; // @[Filter.scala 251:30]
  wire  _T_667 = $signed(pixOut_1_1) > 9'shf; // @[Filter.scala 256:36]
  wire [8:0] _GEN_38575 = _T_667 ? 9'hf : pixOut_1_1; // @[Filter.scala 258:44]
  wire [8:0] _GEN_38577 = _T_664 ? 9'h0 : _GEN_38575; // @[Filter.scala 253:43]
  wire [9:0] _T_674 = $signed(KernelConvolution_1_io_pixelVal_out_2) / $signed(_GEN_39047); // @[Filter.scala 249:64]
  wire  _T_675 = $signed(pixOut_1_2) < 9'sh0; // @[Filter.scala 251:30]
  wire  _T_678 = $signed(pixOut_1_2) > 9'shf; // @[Filter.scala 256:36]
  wire [8:0] _GEN_38580 = _T_678 ? 9'hf : pixOut_1_2; // @[Filter.scala 258:44]
  wire [8:0] _GEN_38582 = _T_675 ? 9'h0 : _GEN_38580; // @[Filter.scala 253:43]
  wire [9:0] _T_685 = $signed(KernelConvolution_1_io_pixelVal_out_3) / $signed(_GEN_39047); // @[Filter.scala 249:64]
  wire  _T_686 = $signed(pixOut_1_3) < 9'sh0; // @[Filter.scala 251:30]
  wire  _T_689 = $signed(pixOut_1_3) > 9'shf; // @[Filter.scala 256:36]
  wire [8:0] _GEN_38585 = _T_689 ? 9'hf : pixOut_1_3; // @[Filter.scala 258:44]
  wire [8:0] _GEN_38587 = _T_686 ? 9'h0 : _GEN_38585; // @[Filter.scala 253:43]
  wire [9:0] _T_696 = $signed(KernelConvolution_1_io_pixelVal_out_4) / $signed(_GEN_39047); // @[Filter.scala 249:64]
  wire  _T_697 = $signed(pixOut_1_4) < 9'sh0; // @[Filter.scala 251:30]
  wire  _T_700 = $signed(pixOut_1_4) > 9'shf; // @[Filter.scala 256:36]
  wire [8:0] _GEN_38590 = _T_700 ? 9'hf : pixOut_1_4; // @[Filter.scala 258:44]
  wire [8:0] _GEN_38592 = _T_697 ? 9'h0 : _GEN_38590; // @[Filter.scala 253:43]
  wire [9:0] _T_707 = $signed(KernelConvolution_1_io_pixelVal_out_5) / $signed(_GEN_39047); // @[Filter.scala 249:64]
  wire  _T_708 = $signed(pixOut_1_5) < 9'sh0; // @[Filter.scala 251:30]
  wire  _T_711 = $signed(pixOut_1_5) > 9'shf; // @[Filter.scala 256:36]
  wire [8:0] _GEN_38595 = _T_711 ? 9'hf : pixOut_1_5; // @[Filter.scala 258:44]
  wire [8:0] _GEN_38597 = _T_708 ? 9'h0 : _GEN_38595; // @[Filter.scala 253:43]
  wire [9:0] _T_718 = $signed(KernelConvolution_1_io_pixelVal_out_6) / $signed(_GEN_39047); // @[Filter.scala 249:64]
  wire  _T_719 = $signed(pixOut_1_6) < 9'sh0; // @[Filter.scala 251:30]
  wire  _T_722 = $signed(pixOut_1_6) > 9'shf; // @[Filter.scala 256:36]
  wire [8:0] _GEN_38600 = _T_722 ? 9'hf : pixOut_1_6; // @[Filter.scala 258:44]
  wire [8:0] _GEN_38602 = _T_719 ? 9'h0 : _GEN_38600; // @[Filter.scala 253:43]
  wire [9:0] _T_729 = $signed(KernelConvolution_1_io_pixelVal_out_7) / $signed(_GEN_39047); // @[Filter.scala 249:64]
  wire  _T_730 = $signed(pixOut_1_7) < 9'sh0; // @[Filter.scala 251:30]
  wire  _T_733 = $signed(pixOut_1_7) > 9'shf; // @[Filter.scala 256:36]
  wire [8:0] _GEN_38605 = _T_733 ? 9'hf : pixOut_1_7; // @[Filter.scala 258:44]
  wire [8:0] _GEN_38607 = _T_730 ? 9'h0 : _GEN_38605; // @[Filter.scala 253:43]
  wire [9:0] _T_740 = $signed(KernelConvolution_2_io_pixelVal_out_0) / $signed(_GEN_39047); // @[Filter.scala 249:64]
  wire  _T_741 = $signed(pixOut_2_0) < 9'sh0; // @[Filter.scala 251:30]
  wire  _T_744 = $signed(pixOut_2_0) > 9'shf; // @[Filter.scala 256:36]
  wire [8:0] _GEN_38610 = _T_744 ? 9'hf : pixOut_2_0; // @[Filter.scala 258:44]
  wire [8:0] _GEN_38612 = _T_741 ? 9'h0 : _GEN_38610; // @[Filter.scala 253:43]
  wire [9:0] _T_751 = $signed(KernelConvolution_2_io_pixelVal_out_1) / $signed(_GEN_39047); // @[Filter.scala 249:64]
  wire  _T_752 = $signed(pixOut_2_1) < 9'sh0; // @[Filter.scala 251:30]
  wire  _T_755 = $signed(pixOut_2_1) > 9'shf; // @[Filter.scala 256:36]
  wire [8:0] _GEN_38615 = _T_755 ? 9'hf : pixOut_2_1; // @[Filter.scala 258:44]
  wire [8:0] _GEN_38617 = _T_752 ? 9'h0 : _GEN_38615; // @[Filter.scala 253:43]
  wire [9:0] _T_762 = $signed(KernelConvolution_2_io_pixelVal_out_2) / $signed(_GEN_39047); // @[Filter.scala 249:64]
  wire  _T_763 = $signed(pixOut_2_2) < 9'sh0; // @[Filter.scala 251:30]
  wire  _T_766 = $signed(pixOut_2_2) > 9'shf; // @[Filter.scala 256:36]
  wire [8:0] _GEN_38620 = _T_766 ? 9'hf : pixOut_2_2; // @[Filter.scala 258:44]
  wire [8:0] _GEN_38622 = _T_763 ? 9'h0 : _GEN_38620; // @[Filter.scala 253:43]
  wire [9:0] _T_773 = $signed(KernelConvolution_2_io_pixelVal_out_3) / $signed(_GEN_39047); // @[Filter.scala 249:64]
  wire  _T_774 = $signed(pixOut_2_3) < 9'sh0; // @[Filter.scala 251:30]
  wire  _T_777 = $signed(pixOut_2_3) > 9'shf; // @[Filter.scala 256:36]
  wire [8:0] _GEN_38625 = _T_777 ? 9'hf : pixOut_2_3; // @[Filter.scala 258:44]
  wire [8:0] _GEN_38627 = _T_774 ? 9'h0 : _GEN_38625; // @[Filter.scala 253:43]
  wire [9:0] _T_784 = $signed(KernelConvolution_2_io_pixelVal_out_4) / $signed(_GEN_39047); // @[Filter.scala 249:64]
  wire  _T_785 = $signed(pixOut_2_4) < 9'sh0; // @[Filter.scala 251:30]
  wire  _T_788 = $signed(pixOut_2_4) > 9'shf; // @[Filter.scala 256:36]
  wire [8:0] _GEN_38630 = _T_788 ? 9'hf : pixOut_2_4; // @[Filter.scala 258:44]
  wire [8:0] _GEN_38632 = _T_785 ? 9'h0 : _GEN_38630; // @[Filter.scala 253:43]
  wire [9:0] _T_795 = $signed(KernelConvolution_2_io_pixelVal_out_5) / $signed(_GEN_39047); // @[Filter.scala 249:64]
  wire  _T_796 = $signed(pixOut_2_5) < 9'sh0; // @[Filter.scala 251:30]
  wire  _T_799 = $signed(pixOut_2_5) > 9'shf; // @[Filter.scala 256:36]
  wire [8:0] _GEN_38635 = _T_799 ? 9'hf : pixOut_2_5; // @[Filter.scala 258:44]
  wire [8:0] _GEN_38637 = _T_796 ? 9'h0 : _GEN_38635; // @[Filter.scala 253:43]
  wire [9:0] _T_806 = $signed(KernelConvolution_2_io_pixelVal_out_6) / $signed(_GEN_39047); // @[Filter.scala 249:64]
  wire  _T_807 = $signed(pixOut_2_6) < 9'sh0; // @[Filter.scala 251:30]
  wire  _T_810 = $signed(pixOut_2_6) > 9'shf; // @[Filter.scala 256:36]
  wire [8:0] _GEN_38640 = _T_810 ? 9'hf : pixOut_2_6; // @[Filter.scala 258:44]
  wire [8:0] _GEN_38642 = _T_807 ? 9'h0 : _GEN_38640; // @[Filter.scala 253:43]
  wire [9:0] _T_817 = $signed(KernelConvolution_2_io_pixelVal_out_7) / $signed(_GEN_39047); // @[Filter.scala 249:64]
  wire  _T_818 = $signed(pixOut_2_7) < 9'sh0; // @[Filter.scala 251:30]
  wire  _T_821 = $signed(pixOut_2_7) > 9'shf; // @[Filter.scala 256:36]
  wire [8:0] _GEN_38645 = _T_821 ? 9'hf : pixOut_2_7; // @[Filter.scala 258:44]
  wire [8:0] _GEN_38647 = _T_818 ? 9'h0 : _GEN_38645; // @[Filter.scala 253:43]
  wire [31:0] _T_829 = pixelIndex + 32'h8; // @[Filter.scala 273:34]
  wire [10:0] _T_830 = 6'h20 * 6'h12; // @[Filter.scala 274:42]
  wire [31:0] _GEN_39071 = {{21'd0}, _T_830}; // @[Filter.scala 274:25]
  wire  _T_831 = pixelIndex == _GEN_39071; // @[Filter.scala 274:25]
  KernelConvolution KernelConvolution ( // @[Filter.scala 212:36]
    .clock(KernelConvolution_clock),
    .reset(KernelConvolution_reset),
    .io_kernelVal_in(KernelConvolution_io_kernelVal_in),
    .io_pixelVal_in_0(KernelConvolution_io_pixelVal_in_0),
    .io_pixelVal_in_1(KernelConvolution_io_pixelVal_in_1),
    .io_pixelVal_in_2(KernelConvolution_io_pixelVal_in_2),
    .io_pixelVal_in_3(KernelConvolution_io_pixelVal_in_3),
    .io_pixelVal_in_4(KernelConvolution_io_pixelVal_in_4),
    .io_pixelVal_in_5(KernelConvolution_io_pixelVal_in_5),
    .io_pixelVal_in_6(KernelConvolution_io_pixelVal_in_6),
    .io_pixelVal_in_7(KernelConvolution_io_pixelVal_in_7),
    .io_pixelVal_out_0(KernelConvolution_io_pixelVal_out_0),
    .io_pixelVal_out_1(KernelConvolution_io_pixelVal_out_1),
    .io_pixelVal_out_2(KernelConvolution_io_pixelVal_out_2),
    .io_pixelVal_out_3(KernelConvolution_io_pixelVal_out_3),
    .io_pixelVal_out_4(KernelConvolution_io_pixelVal_out_4),
    .io_pixelVal_out_5(KernelConvolution_io_pixelVal_out_5),
    .io_pixelVal_out_6(KernelConvolution_io_pixelVal_out_6),
    .io_pixelVal_out_7(KernelConvolution_io_pixelVal_out_7),
    .io_valid_out(KernelConvolution_io_valid_out)
  );
  KernelConvolution KernelConvolution_1 ( // @[Filter.scala 213:36]
    .clock(KernelConvolution_1_clock),
    .reset(KernelConvolution_1_reset),
    .io_kernelVal_in(KernelConvolution_1_io_kernelVal_in),
    .io_pixelVal_in_0(KernelConvolution_1_io_pixelVal_in_0),
    .io_pixelVal_in_1(KernelConvolution_1_io_pixelVal_in_1),
    .io_pixelVal_in_2(KernelConvolution_1_io_pixelVal_in_2),
    .io_pixelVal_in_3(KernelConvolution_1_io_pixelVal_in_3),
    .io_pixelVal_in_4(KernelConvolution_1_io_pixelVal_in_4),
    .io_pixelVal_in_5(KernelConvolution_1_io_pixelVal_in_5),
    .io_pixelVal_in_6(KernelConvolution_1_io_pixelVal_in_6),
    .io_pixelVal_in_7(KernelConvolution_1_io_pixelVal_in_7),
    .io_pixelVal_out_0(KernelConvolution_1_io_pixelVal_out_0),
    .io_pixelVal_out_1(KernelConvolution_1_io_pixelVal_out_1),
    .io_pixelVal_out_2(KernelConvolution_1_io_pixelVal_out_2),
    .io_pixelVal_out_3(KernelConvolution_1_io_pixelVal_out_3),
    .io_pixelVal_out_4(KernelConvolution_1_io_pixelVal_out_4),
    .io_pixelVal_out_5(KernelConvolution_1_io_pixelVal_out_5),
    .io_pixelVal_out_6(KernelConvolution_1_io_pixelVal_out_6),
    .io_pixelVal_out_7(KernelConvolution_1_io_pixelVal_out_7),
    .io_valid_out(KernelConvolution_1_io_valid_out)
  );
  KernelConvolution KernelConvolution_2 ( // @[Filter.scala 214:36]
    .clock(KernelConvolution_2_clock),
    .reset(KernelConvolution_2_reset),
    .io_kernelVal_in(KernelConvolution_2_io_kernelVal_in),
    .io_pixelVal_in_0(KernelConvolution_2_io_pixelVal_in_0),
    .io_pixelVal_in_1(KernelConvolution_2_io_pixelVal_in_1),
    .io_pixelVal_in_2(KernelConvolution_2_io_pixelVal_in_2),
    .io_pixelVal_in_3(KernelConvolution_2_io_pixelVal_in_3),
    .io_pixelVal_in_4(KernelConvolution_2_io_pixelVal_in_4),
    .io_pixelVal_in_5(KernelConvolution_2_io_pixelVal_in_5),
    .io_pixelVal_in_6(KernelConvolution_2_io_pixelVal_in_6),
    .io_pixelVal_in_7(KernelConvolution_2_io_pixelVal_in_7),
    .io_pixelVal_out_0(KernelConvolution_2_io_pixelVal_out_0),
    .io_pixelVal_out_1(KernelConvolution_2_io_pixelVal_out_1),
    .io_pixelVal_out_2(KernelConvolution_2_io_pixelVal_out_2),
    .io_pixelVal_out_3(KernelConvolution_2_io_pixelVal_out_3),
    .io_pixelVal_out_4(KernelConvolution_2_io_pixelVal_out_4),
    .io_pixelVal_out_5(KernelConvolution_2_io_pixelVal_out_5),
    .io_pixelVal_out_6(KernelConvolution_2_io_pixelVal_out_6),
    .io_pixelVal_out_7(KernelConvolution_2_io_pixelVal_out_7),
    .io_valid_out(KernelConvolution_2_io_valid_out)
  );
  assign io_pixelVal_out_0_0 = _GEN_38532[3:0]; // @[Filter.scala 252:35 Filter.scala 254:37 Filter.scala 257:35 Filter.scala 259:35 Filter.scala 261:35 Filter.scala 263:35]
  assign io_pixelVal_out_0_1 = _GEN_38537[3:0]; // @[Filter.scala 252:35 Filter.scala 254:37 Filter.scala 257:35 Filter.scala 259:35 Filter.scala 261:35 Filter.scala 263:35]
  assign io_pixelVal_out_0_2 = _GEN_38542[3:0]; // @[Filter.scala 252:35 Filter.scala 254:37 Filter.scala 257:35 Filter.scala 259:35 Filter.scala 261:35 Filter.scala 263:35]
  assign io_pixelVal_out_0_3 = _GEN_38547[3:0]; // @[Filter.scala 252:35 Filter.scala 254:37 Filter.scala 257:35 Filter.scala 259:35 Filter.scala 261:35 Filter.scala 263:35]
  assign io_pixelVal_out_0_4 = _GEN_38552[3:0]; // @[Filter.scala 252:35 Filter.scala 254:37 Filter.scala 257:35 Filter.scala 259:35 Filter.scala 261:35 Filter.scala 263:35]
  assign io_pixelVal_out_0_5 = _GEN_38557[3:0]; // @[Filter.scala 252:35 Filter.scala 254:37 Filter.scala 257:35 Filter.scala 259:35 Filter.scala 261:35 Filter.scala 263:35]
  assign io_pixelVal_out_0_6 = _GEN_38562[3:0]; // @[Filter.scala 252:35 Filter.scala 254:37 Filter.scala 257:35 Filter.scala 259:35 Filter.scala 261:35 Filter.scala 263:35]
  assign io_pixelVal_out_0_7 = _GEN_38567[3:0]; // @[Filter.scala 252:35 Filter.scala 254:37 Filter.scala 257:35 Filter.scala 259:35 Filter.scala 261:35 Filter.scala 263:35]
  assign io_pixelVal_out_1_0 = _GEN_38572[3:0]; // @[Filter.scala 252:35 Filter.scala 254:37 Filter.scala 257:35 Filter.scala 259:35 Filter.scala 261:35 Filter.scala 263:35]
  assign io_pixelVal_out_1_1 = _GEN_38577[3:0]; // @[Filter.scala 252:35 Filter.scala 254:37 Filter.scala 257:35 Filter.scala 259:35 Filter.scala 261:35 Filter.scala 263:35]
  assign io_pixelVal_out_1_2 = _GEN_38582[3:0]; // @[Filter.scala 252:35 Filter.scala 254:37 Filter.scala 257:35 Filter.scala 259:35 Filter.scala 261:35 Filter.scala 263:35]
  assign io_pixelVal_out_1_3 = _GEN_38587[3:0]; // @[Filter.scala 252:35 Filter.scala 254:37 Filter.scala 257:35 Filter.scala 259:35 Filter.scala 261:35 Filter.scala 263:35]
  assign io_pixelVal_out_1_4 = _GEN_38592[3:0]; // @[Filter.scala 252:35 Filter.scala 254:37 Filter.scala 257:35 Filter.scala 259:35 Filter.scala 261:35 Filter.scala 263:35]
  assign io_pixelVal_out_1_5 = _GEN_38597[3:0]; // @[Filter.scala 252:35 Filter.scala 254:37 Filter.scala 257:35 Filter.scala 259:35 Filter.scala 261:35 Filter.scala 263:35]
  assign io_pixelVal_out_1_6 = _GEN_38602[3:0]; // @[Filter.scala 252:35 Filter.scala 254:37 Filter.scala 257:35 Filter.scala 259:35 Filter.scala 261:35 Filter.scala 263:35]
  assign io_pixelVal_out_1_7 = _GEN_38607[3:0]; // @[Filter.scala 252:35 Filter.scala 254:37 Filter.scala 257:35 Filter.scala 259:35 Filter.scala 261:35 Filter.scala 263:35]
  assign io_pixelVal_out_2_0 = _GEN_38612[3:0]; // @[Filter.scala 252:35 Filter.scala 254:37 Filter.scala 257:35 Filter.scala 259:35 Filter.scala 261:35 Filter.scala 263:35]
  assign io_pixelVal_out_2_1 = _GEN_38617[3:0]; // @[Filter.scala 252:35 Filter.scala 254:37 Filter.scala 257:35 Filter.scala 259:35 Filter.scala 261:35 Filter.scala 263:35]
  assign io_pixelVal_out_2_2 = _GEN_38622[3:0]; // @[Filter.scala 252:35 Filter.scala 254:37 Filter.scala 257:35 Filter.scala 259:35 Filter.scala 261:35 Filter.scala 263:35]
  assign io_pixelVal_out_2_3 = _GEN_38627[3:0]; // @[Filter.scala 252:35 Filter.scala 254:37 Filter.scala 257:35 Filter.scala 259:35 Filter.scala 261:35 Filter.scala 263:35]
  assign io_pixelVal_out_2_4 = _GEN_38632[3:0]; // @[Filter.scala 252:35 Filter.scala 254:37 Filter.scala 257:35 Filter.scala 259:35 Filter.scala 261:35 Filter.scala 263:35]
  assign io_pixelVal_out_2_5 = _GEN_38637[3:0]; // @[Filter.scala 252:35 Filter.scala 254:37 Filter.scala 257:35 Filter.scala 259:35 Filter.scala 261:35 Filter.scala 263:35]
  assign io_pixelVal_out_2_6 = _GEN_38642[3:0]; // @[Filter.scala 252:35 Filter.scala 254:37 Filter.scala 257:35 Filter.scala 259:35 Filter.scala 261:35 Filter.scala 263:35]
  assign io_pixelVal_out_2_7 = _GEN_38647[3:0]; // @[Filter.scala 252:35 Filter.scala 254:37 Filter.scala 257:35 Filter.scala 259:35 Filter.scala 261:35 Filter.scala 263:35]
  assign io_valid_out = validOut; // @[Filter.scala 270:18]
  assign KernelConvolution_clock = clock;
  assign KernelConvolution_reset = reset;
  assign KernelConvolution_io_kernelVal_in = _GEN_38733 & _GEN_38660 ? $signed(5'sh0) : $signed(_GEN_55); // @[Filter.scala 220:41]
  assign KernelConvolution_io_pixelVal_in_0 = _GEN_3364[3:0]; // @[Filter.scala 234:53 Filter.scala 236:51 Filter.scala 238:51]
  assign KernelConvolution_io_pixelVal_in_1 = _GEN_8158[3:0]; // @[Filter.scala 234:53 Filter.scala 236:51 Filter.scala 238:51]
  assign KernelConvolution_io_pixelVal_in_2 = _GEN_12952[3:0]; // @[Filter.scala 234:53 Filter.scala 236:51 Filter.scala 238:51]
  assign KernelConvolution_io_pixelVal_in_3 = _GEN_17746[3:0]; // @[Filter.scala 234:53 Filter.scala 236:51 Filter.scala 238:51]
  assign KernelConvolution_io_pixelVal_in_4 = _GEN_22540[3:0]; // @[Filter.scala 234:53 Filter.scala 236:51 Filter.scala 238:51]
  assign KernelConvolution_io_pixelVal_in_5 = _GEN_27334[3:0]; // @[Filter.scala 234:53 Filter.scala 236:51 Filter.scala 238:51]
  assign KernelConvolution_io_pixelVal_in_6 = _GEN_32128[3:0]; // @[Filter.scala 234:53 Filter.scala 236:51 Filter.scala 238:51]
  assign KernelConvolution_io_pixelVal_in_7 = _GEN_36922[3:0]; // @[Filter.scala 234:53 Filter.scala 236:51 Filter.scala 238:51]
  assign KernelConvolution_1_clock = clock;
  assign KernelConvolution_1_reset = reset;
  assign KernelConvolution_1_io_kernelVal_in = _GEN_38733 & _GEN_38660 ? $signed(5'sh0) : $signed(_GEN_55); // @[Filter.scala 220:41]
  assign KernelConvolution_1_io_pixelVal_in_0 = _GEN_4164[3:0]; // @[Filter.scala 234:53 Filter.scala 236:51 Filter.scala 238:51]
  assign KernelConvolution_1_io_pixelVal_in_1 = _GEN_8958[3:0]; // @[Filter.scala 234:53 Filter.scala 236:51 Filter.scala 238:51]
  assign KernelConvolution_1_io_pixelVal_in_2 = _GEN_13752[3:0]; // @[Filter.scala 234:53 Filter.scala 236:51 Filter.scala 238:51]
  assign KernelConvolution_1_io_pixelVal_in_3 = _GEN_18546[3:0]; // @[Filter.scala 234:53 Filter.scala 236:51 Filter.scala 238:51]
  assign KernelConvolution_1_io_pixelVal_in_4 = _GEN_23340[3:0]; // @[Filter.scala 234:53 Filter.scala 236:51 Filter.scala 238:51]
  assign KernelConvolution_1_io_pixelVal_in_5 = _GEN_28134[3:0]; // @[Filter.scala 234:53 Filter.scala 236:51 Filter.scala 238:51]
  assign KernelConvolution_1_io_pixelVal_in_6 = _GEN_32928[3:0]; // @[Filter.scala 234:53 Filter.scala 236:51 Filter.scala 238:51]
  assign KernelConvolution_1_io_pixelVal_in_7 = _GEN_37722[3:0]; // @[Filter.scala 234:53 Filter.scala 236:51 Filter.scala 238:51]
  assign KernelConvolution_2_clock = clock;
  assign KernelConvolution_2_reset = reset;
  assign KernelConvolution_2_io_kernelVal_in = _GEN_38733 & _GEN_38660 ? $signed(5'sh0) : $signed(_GEN_55); // @[Filter.scala 220:41]
  assign KernelConvolution_2_io_pixelVal_in_0 = _GEN_4964[3:0]; // @[Filter.scala 234:53 Filter.scala 236:51 Filter.scala 238:51]
  assign KernelConvolution_2_io_pixelVal_in_1 = _GEN_9758[3:0]; // @[Filter.scala 234:53 Filter.scala 236:51 Filter.scala 238:51]
  assign KernelConvolution_2_io_pixelVal_in_2 = _GEN_14552[3:0]; // @[Filter.scala 234:53 Filter.scala 236:51 Filter.scala 238:51]
  assign KernelConvolution_2_io_pixelVal_in_3 = _GEN_19346[3:0]; // @[Filter.scala 234:53 Filter.scala 236:51 Filter.scala 238:51]
  assign KernelConvolution_2_io_pixelVal_in_4 = _GEN_24140[3:0]; // @[Filter.scala 234:53 Filter.scala 236:51 Filter.scala 238:51]
  assign KernelConvolution_2_io_pixelVal_in_5 = _GEN_28934[3:0]; // @[Filter.scala 234:53 Filter.scala 236:51 Filter.scala 238:51]
  assign KernelConvolution_2_io_pixelVal_in_6 = _GEN_33728[3:0]; // @[Filter.scala 234:53 Filter.scala 236:51 Filter.scala 238:51]
  assign KernelConvolution_2_io_pixelVal_in_7 = _GEN_38522[3:0]; // @[Filter.scala 234:53 Filter.scala 236:51 Filter.scala 238:51]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  kernelCounter = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  imageCounterX = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  imageCounterY = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  pixelIndex = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  pixOut_0_0 = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  pixOut_0_1 = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  pixOut_0_2 = _RAND_6[8:0];
  _RAND_7 = {1{`RANDOM}};
  pixOut_0_3 = _RAND_7[8:0];
  _RAND_8 = {1{`RANDOM}};
  pixOut_0_4 = _RAND_8[8:0];
  _RAND_9 = {1{`RANDOM}};
  pixOut_0_5 = _RAND_9[8:0];
  _RAND_10 = {1{`RANDOM}};
  pixOut_0_6 = _RAND_10[8:0];
  _RAND_11 = {1{`RANDOM}};
  pixOut_0_7 = _RAND_11[8:0];
  _RAND_12 = {1{`RANDOM}};
  pixOut_1_0 = _RAND_12[8:0];
  _RAND_13 = {1{`RANDOM}};
  pixOut_1_1 = _RAND_13[8:0];
  _RAND_14 = {1{`RANDOM}};
  pixOut_1_2 = _RAND_14[8:0];
  _RAND_15 = {1{`RANDOM}};
  pixOut_1_3 = _RAND_15[8:0];
  _RAND_16 = {1{`RANDOM}};
  pixOut_1_4 = _RAND_16[8:0];
  _RAND_17 = {1{`RANDOM}};
  pixOut_1_5 = _RAND_17[8:0];
  _RAND_18 = {1{`RANDOM}};
  pixOut_1_6 = _RAND_18[8:0];
  _RAND_19 = {1{`RANDOM}};
  pixOut_1_7 = _RAND_19[8:0];
  _RAND_20 = {1{`RANDOM}};
  pixOut_2_0 = _RAND_20[8:0];
  _RAND_21 = {1{`RANDOM}};
  pixOut_2_1 = _RAND_21[8:0];
  _RAND_22 = {1{`RANDOM}};
  pixOut_2_2 = _RAND_22[8:0];
  _RAND_23 = {1{`RANDOM}};
  pixOut_2_3 = _RAND_23[8:0];
  _RAND_24 = {1{`RANDOM}};
  pixOut_2_4 = _RAND_24[8:0];
  _RAND_25 = {1{`RANDOM}};
  pixOut_2_5 = _RAND_25[8:0];
  _RAND_26 = {1{`RANDOM}};
  pixOut_2_6 = _RAND_26[8:0];
  _RAND_27 = {1{`RANDOM}};
  pixOut_2_7 = _RAND_27[8:0];
  _RAND_28 = {1{`RANDOM}};
  validOut = _RAND_28[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      kernelCounter <= 4'h0;
    end else if (kernelCountReset) begin
      kernelCounter <= 4'h0;
    end else begin
      kernelCounter <= _T_14;
    end
    if (reset) begin
      imageCounterX <= 2'h0;
    end else if (imageCounterXReset) begin
      imageCounterX <= 2'h0;
    end else begin
      imageCounterX <= _T_20;
    end
    if (reset) begin
      imageCounterY <= 2'h0;
    end else if (imageCounterXReset) begin
      if (_T_21) begin
        imageCounterY <= 2'h0;
      end else begin
        imageCounterY <= _T_23;
      end
    end
    if (reset) begin
      pixelIndex <= 32'h0;
    end else if (kernelCountReset) begin
      if (_T_831) begin
        pixelIndex <= 32'h0;
      end else begin
        pixelIndex <= _T_829;
      end
    end
    if (reset) begin
      pixOut_0_0 <= 9'sh0;
    end else begin
      pixOut_0_0 <= _T_564[8:0];
    end
    if (reset) begin
      pixOut_0_1 <= 9'sh0;
    end else begin
      pixOut_0_1 <= _T_575[8:0];
    end
    if (reset) begin
      pixOut_0_2 <= 9'sh0;
    end else begin
      pixOut_0_2 <= _T_586[8:0];
    end
    if (reset) begin
      pixOut_0_3 <= 9'sh0;
    end else begin
      pixOut_0_3 <= _T_597[8:0];
    end
    if (reset) begin
      pixOut_0_4 <= 9'sh0;
    end else begin
      pixOut_0_4 <= _T_608[8:0];
    end
    if (reset) begin
      pixOut_0_5 <= 9'sh0;
    end else begin
      pixOut_0_5 <= _T_619[8:0];
    end
    if (reset) begin
      pixOut_0_6 <= 9'sh0;
    end else begin
      pixOut_0_6 <= _T_630[8:0];
    end
    if (reset) begin
      pixOut_0_7 <= 9'sh0;
    end else begin
      pixOut_0_7 <= _T_641[8:0];
    end
    if (reset) begin
      pixOut_1_0 <= 9'sh0;
    end else begin
      pixOut_1_0 <= _T_652[8:0];
    end
    if (reset) begin
      pixOut_1_1 <= 9'sh0;
    end else begin
      pixOut_1_1 <= _T_663[8:0];
    end
    if (reset) begin
      pixOut_1_2 <= 9'sh0;
    end else begin
      pixOut_1_2 <= _T_674[8:0];
    end
    if (reset) begin
      pixOut_1_3 <= 9'sh0;
    end else begin
      pixOut_1_3 <= _T_685[8:0];
    end
    if (reset) begin
      pixOut_1_4 <= 9'sh0;
    end else begin
      pixOut_1_4 <= _T_696[8:0];
    end
    if (reset) begin
      pixOut_1_5 <= 9'sh0;
    end else begin
      pixOut_1_5 <= _T_707[8:0];
    end
    if (reset) begin
      pixOut_1_6 <= 9'sh0;
    end else begin
      pixOut_1_6 <= _T_718[8:0];
    end
    if (reset) begin
      pixOut_1_7 <= 9'sh0;
    end else begin
      pixOut_1_7 <= _T_729[8:0];
    end
    if (reset) begin
      pixOut_2_0 <= 9'sh0;
    end else begin
      pixOut_2_0 <= _T_740[8:0];
    end
    if (reset) begin
      pixOut_2_1 <= 9'sh0;
    end else begin
      pixOut_2_1 <= _T_751[8:0];
    end
    if (reset) begin
      pixOut_2_2 <= 9'sh0;
    end else begin
      pixOut_2_2 <= _T_762[8:0];
    end
    if (reset) begin
      pixOut_2_3 <= 9'sh0;
    end else begin
      pixOut_2_3 <= _T_773[8:0];
    end
    if (reset) begin
      pixOut_2_4 <= 9'sh0;
    end else begin
      pixOut_2_4 <= _T_784[8:0];
    end
    if (reset) begin
      pixOut_2_5 <= 9'sh0;
    end else begin
      pixOut_2_5 <= _T_795[8:0];
    end
    if (reset) begin
      pixOut_2_6 <= 9'sh0;
    end else begin
      pixOut_2_6 <= _T_806[8:0];
    end
    if (reset) begin
      pixOut_2_7 <= 9'sh0;
    end else begin
      pixOut_2_7 <= _T_817[8:0];
    end
    if (reset) begin
      validOut <= 1'h0;
    end else begin
      validOut <= KernelConvolution_io_valid_out;
    end
  end
endmodule
module VideoBuffer(
  input         clock,
  input         reset,
  input  [3:0]  io_pixelVal_in_0_0,
  input  [3:0]  io_pixelVal_in_0_1,
  input  [3:0]  io_pixelVal_in_0_2,
  input  [3:0]  io_pixelVal_in_0_3,
  input  [3:0]  io_pixelVal_in_0_4,
  input  [3:0]  io_pixelVal_in_0_5,
  input  [3:0]  io_pixelVal_in_0_6,
  input  [3:0]  io_pixelVal_in_0_7,
  input  [3:0]  io_pixelVal_in_1_0,
  input  [3:0]  io_pixelVal_in_1_1,
  input  [3:0]  io_pixelVal_in_1_2,
  input  [3:0]  io_pixelVal_in_1_3,
  input  [3:0]  io_pixelVal_in_1_4,
  input  [3:0]  io_pixelVal_in_1_5,
  input  [3:0]  io_pixelVal_in_1_6,
  input  [3:0]  io_pixelVal_in_1_7,
  input  [3:0]  io_pixelVal_in_2_0,
  input  [3:0]  io_pixelVal_in_2_1,
  input  [3:0]  io_pixelVal_in_2_2,
  input  [3:0]  io_pixelVal_in_2_3,
  input  [3:0]  io_pixelVal_in_2_4,
  input  [3:0]  io_pixelVal_in_2_5,
  input  [3:0]  io_pixelVal_in_2_6,
  input  [3:0]  io_pixelVal_in_2_7,
  input         io_valid_in,
  input  [10:0] io_rowIndex,
  input  [10:0] io_colIndex,
  output [3:0]  io_pixelVal_out_0,
  output [3:0]  io_pixelVal_out_1,
  output [3:0]  io_pixelVal_out_2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [31:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1285;
  reg [31:0] _RAND_1286;
  reg [31:0] _RAND_1287;
  reg [31:0] _RAND_1288;
  reg [31:0] _RAND_1289;
  reg [31:0] _RAND_1290;
  reg [31:0] _RAND_1291;
  reg [31:0] _RAND_1292;
  reg [31:0] _RAND_1293;
  reg [31:0] _RAND_1294;
  reg [31:0] _RAND_1295;
  reg [31:0] _RAND_1296;
  reg [31:0] _RAND_1297;
  reg [31:0] _RAND_1298;
  reg [31:0] _RAND_1299;
  reg [31:0] _RAND_1300;
  reg [31:0] _RAND_1301;
  reg [31:0] _RAND_1302;
  reg [31:0] _RAND_1303;
  reg [31:0] _RAND_1304;
  reg [31:0] _RAND_1305;
  reg [31:0] _RAND_1306;
  reg [31:0] _RAND_1307;
  reg [31:0] _RAND_1308;
  reg [31:0] _RAND_1309;
  reg [31:0] _RAND_1310;
  reg [31:0] _RAND_1311;
  reg [31:0] _RAND_1312;
  reg [31:0] _RAND_1313;
  reg [31:0] _RAND_1314;
  reg [31:0] _RAND_1315;
  reg [31:0] _RAND_1316;
  reg [31:0] _RAND_1317;
  reg [31:0] _RAND_1318;
  reg [31:0] _RAND_1319;
  reg [31:0] _RAND_1320;
  reg [31:0] _RAND_1321;
  reg [31:0] _RAND_1322;
  reg [31:0] _RAND_1323;
  reg [31:0] _RAND_1324;
  reg [31:0] _RAND_1325;
  reg [31:0] _RAND_1326;
  reg [31:0] _RAND_1327;
  reg [31:0] _RAND_1328;
  reg [31:0] _RAND_1329;
  reg [31:0] _RAND_1330;
  reg [31:0] _RAND_1331;
  reg [31:0] _RAND_1332;
  reg [31:0] _RAND_1333;
  reg [31:0] _RAND_1334;
  reg [31:0] _RAND_1335;
  reg [31:0] _RAND_1336;
  reg [31:0] _RAND_1337;
  reg [31:0] _RAND_1338;
  reg [31:0] _RAND_1339;
  reg [31:0] _RAND_1340;
  reg [31:0] _RAND_1341;
  reg [31:0] _RAND_1342;
  reg [31:0] _RAND_1343;
  reg [31:0] _RAND_1344;
  reg [31:0] _RAND_1345;
  reg [31:0] _RAND_1346;
  reg [31:0] _RAND_1347;
  reg [31:0] _RAND_1348;
  reg [31:0] _RAND_1349;
  reg [31:0] _RAND_1350;
  reg [31:0] _RAND_1351;
  reg [31:0] _RAND_1352;
  reg [31:0] _RAND_1353;
  reg [31:0] _RAND_1354;
  reg [31:0] _RAND_1355;
  reg [31:0] _RAND_1356;
  reg [31:0] _RAND_1357;
  reg [31:0] _RAND_1358;
  reg [31:0] _RAND_1359;
  reg [31:0] _RAND_1360;
  reg [31:0] _RAND_1361;
  reg [31:0] _RAND_1362;
  reg [31:0] _RAND_1363;
  reg [31:0] _RAND_1364;
  reg [31:0] _RAND_1365;
  reg [31:0] _RAND_1366;
  reg [31:0] _RAND_1367;
  reg [31:0] _RAND_1368;
  reg [31:0] _RAND_1369;
  reg [31:0] _RAND_1370;
  reg [31:0] _RAND_1371;
  reg [31:0] _RAND_1372;
  reg [31:0] _RAND_1373;
  reg [31:0] _RAND_1374;
  reg [31:0] _RAND_1375;
  reg [31:0] _RAND_1376;
  reg [31:0] _RAND_1377;
  reg [31:0] _RAND_1378;
  reg [31:0] _RAND_1379;
  reg [31:0] _RAND_1380;
  reg [31:0] _RAND_1381;
  reg [31:0] _RAND_1382;
  reg [31:0] _RAND_1383;
  reg [31:0] _RAND_1384;
  reg [31:0] _RAND_1385;
  reg [31:0] _RAND_1386;
  reg [31:0] _RAND_1387;
  reg [31:0] _RAND_1388;
  reg [31:0] _RAND_1389;
  reg [31:0] _RAND_1390;
  reg [31:0] _RAND_1391;
  reg [31:0] _RAND_1392;
  reg [31:0] _RAND_1393;
  reg [31:0] _RAND_1394;
  reg [31:0] _RAND_1395;
  reg [31:0] _RAND_1396;
  reg [31:0] _RAND_1397;
  reg [31:0] _RAND_1398;
  reg [31:0] _RAND_1399;
  reg [31:0] _RAND_1400;
  reg [31:0] _RAND_1401;
  reg [31:0] _RAND_1402;
  reg [31:0] _RAND_1403;
  reg [31:0] _RAND_1404;
  reg [31:0] _RAND_1405;
  reg [31:0] _RAND_1406;
  reg [31:0] _RAND_1407;
  reg [31:0] _RAND_1408;
  reg [31:0] _RAND_1409;
  reg [31:0] _RAND_1410;
  reg [31:0] _RAND_1411;
  reg [31:0] _RAND_1412;
  reg [31:0] _RAND_1413;
  reg [31:0] _RAND_1414;
  reg [31:0] _RAND_1415;
  reg [31:0] _RAND_1416;
  reg [31:0] _RAND_1417;
  reg [31:0] _RAND_1418;
  reg [31:0] _RAND_1419;
  reg [31:0] _RAND_1420;
  reg [31:0] _RAND_1421;
  reg [31:0] _RAND_1422;
  reg [31:0] _RAND_1423;
  reg [31:0] _RAND_1424;
  reg [31:0] _RAND_1425;
  reg [31:0] _RAND_1426;
  reg [31:0] _RAND_1427;
  reg [31:0] _RAND_1428;
  reg [31:0] _RAND_1429;
  reg [31:0] _RAND_1430;
  reg [31:0] _RAND_1431;
  reg [31:0] _RAND_1432;
  reg [31:0] _RAND_1433;
  reg [31:0] _RAND_1434;
  reg [31:0] _RAND_1435;
  reg [31:0] _RAND_1436;
  reg [31:0] _RAND_1437;
  reg [31:0] _RAND_1438;
  reg [31:0] _RAND_1439;
  reg [31:0] _RAND_1440;
  reg [31:0] _RAND_1441;
  reg [31:0] _RAND_1442;
  reg [31:0] _RAND_1443;
  reg [31:0] _RAND_1444;
  reg [31:0] _RAND_1445;
  reg [31:0] _RAND_1446;
  reg [31:0] _RAND_1447;
  reg [31:0] _RAND_1448;
  reg [31:0] _RAND_1449;
  reg [31:0] _RAND_1450;
  reg [31:0] _RAND_1451;
  reg [31:0] _RAND_1452;
  reg [31:0] _RAND_1453;
  reg [31:0] _RAND_1454;
  reg [31:0] _RAND_1455;
  reg [31:0] _RAND_1456;
  reg [31:0] _RAND_1457;
  reg [31:0] _RAND_1458;
  reg [31:0] _RAND_1459;
  reg [31:0] _RAND_1460;
  reg [31:0] _RAND_1461;
  reg [31:0] _RAND_1462;
  reg [31:0] _RAND_1463;
  reg [31:0] _RAND_1464;
  reg [31:0] _RAND_1465;
  reg [31:0] _RAND_1466;
  reg [31:0] _RAND_1467;
  reg [31:0] _RAND_1468;
  reg [31:0] _RAND_1469;
  reg [31:0] _RAND_1470;
  reg [31:0] _RAND_1471;
  reg [31:0] _RAND_1472;
  reg [31:0] _RAND_1473;
  reg [31:0] _RAND_1474;
  reg [31:0] _RAND_1475;
  reg [31:0] _RAND_1476;
  reg [31:0] _RAND_1477;
  reg [31:0] _RAND_1478;
  reg [31:0] _RAND_1479;
  reg [31:0] _RAND_1480;
  reg [31:0] _RAND_1481;
  reg [31:0] _RAND_1482;
  reg [31:0] _RAND_1483;
  reg [31:0] _RAND_1484;
  reg [31:0] _RAND_1485;
  reg [31:0] _RAND_1486;
  reg [31:0] _RAND_1487;
  reg [31:0] _RAND_1488;
  reg [31:0] _RAND_1489;
  reg [31:0] _RAND_1490;
  reg [31:0] _RAND_1491;
  reg [31:0] _RAND_1492;
  reg [31:0] _RAND_1493;
  reg [31:0] _RAND_1494;
  reg [31:0] _RAND_1495;
  reg [31:0] _RAND_1496;
  reg [31:0] _RAND_1497;
  reg [31:0] _RAND_1498;
  reg [31:0] _RAND_1499;
  reg [31:0] _RAND_1500;
  reg [31:0] _RAND_1501;
  reg [31:0] _RAND_1502;
  reg [31:0] _RAND_1503;
  reg [31:0] _RAND_1504;
  reg [31:0] _RAND_1505;
  reg [31:0] _RAND_1506;
  reg [31:0] _RAND_1507;
  reg [31:0] _RAND_1508;
  reg [31:0] _RAND_1509;
  reg [31:0] _RAND_1510;
  reg [31:0] _RAND_1511;
  reg [31:0] _RAND_1512;
  reg [31:0] _RAND_1513;
  reg [31:0] _RAND_1514;
  reg [31:0] _RAND_1515;
  reg [31:0] _RAND_1516;
  reg [31:0] _RAND_1517;
  reg [31:0] _RAND_1518;
  reg [31:0] _RAND_1519;
  reg [31:0] _RAND_1520;
  reg [31:0] _RAND_1521;
  reg [31:0] _RAND_1522;
  reg [31:0] _RAND_1523;
  reg [31:0] _RAND_1524;
  reg [31:0] _RAND_1525;
  reg [31:0] _RAND_1526;
  reg [31:0] _RAND_1527;
  reg [31:0] _RAND_1528;
  reg [31:0] _RAND_1529;
  reg [31:0] _RAND_1530;
  reg [31:0] _RAND_1531;
  reg [31:0] _RAND_1532;
  reg [31:0] _RAND_1533;
  reg [31:0] _RAND_1534;
  reg [31:0] _RAND_1535;
  reg [31:0] _RAND_1536;
  reg [31:0] _RAND_1537;
  reg [31:0] _RAND_1538;
  reg [31:0] _RAND_1539;
  reg [31:0] _RAND_1540;
  reg [31:0] _RAND_1541;
  reg [31:0] _RAND_1542;
  reg [31:0] _RAND_1543;
  reg [31:0] _RAND_1544;
  reg [31:0] _RAND_1545;
  reg [31:0] _RAND_1546;
  reg [31:0] _RAND_1547;
  reg [31:0] _RAND_1548;
  reg [31:0] _RAND_1549;
  reg [31:0] _RAND_1550;
  reg [31:0] _RAND_1551;
  reg [31:0] _RAND_1552;
  reg [31:0] _RAND_1553;
  reg [31:0] _RAND_1554;
  reg [31:0] _RAND_1555;
  reg [31:0] _RAND_1556;
  reg [31:0] _RAND_1557;
  reg [31:0] _RAND_1558;
  reg [31:0] _RAND_1559;
  reg [31:0] _RAND_1560;
  reg [31:0] _RAND_1561;
  reg [31:0] _RAND_1562;
  reg [31:0] _RAND_1563;
  reg [31:0] _RAND_1564;
  reg [31:0] _RAND_1565;
  reg [31:0] _RAND_1566;
  reg [31:0] _RAND_1567;
  reg [31:0] _RAND_1568;
  reg [31:0] _RAND_1569;
  reg [31:0] _RAND_1570;
  reg [31:0] _RAND_1571;
  reg [31:0] _RAND_1572;
  reg [31:0] _RAND_1573;
  reg [31:0] _RAND_1574;
  reg [31:0] _RAND_1575;
  reg [31:0] _RAND_1576;
  reg [31:0] _RAND_1577;
  reg [31:0] _RAND_1578;
  reg [31:0] _RAND_1579;
  reg [31:0] _RAND_1580;
  reg [31:0] _RAND_1581;
  reg [31:0] _RAND_1582;
  reg [31:0] _RAND_1583;
  reg [31:0] _RAND_1584;
  reg [31:0] _RAND_1585;
  reg [31:0] _RAND_1586;
  reg [31:0] _RAND_1587;
  reg [31:0] _RAND_1588;
  reg [31:0] _RAND_1589;
  reg [31:0] _RAND_1590;
  reg [31:0] _RAND_1591;
  reg [31:0] _RAND_1592;
  reg [31:0] _RAND_1593;
  reg [31:0] _RAND_1594;
  reg [31:0] _RAND_1595;
  reg [31:0] _RAND_1596;
  reg [31:0] _RAND_1597;
  reg [31:0] _RAND_1598;
  reg [31:0] _RAND_1599;
  reg [31:0] _RAND_1600;
  reg [31:0] _RAND_1601;
  reg [31:0] _RAND_1602;
  reg [31:0] _RAND_1603;
  reg [31:0] _RAND_1604;
  reg [31:0] _RAND_1605;
  reg [31:0] _RAND_1606;
  reg [31:0] _RAND_1607;
  reg [31:0] _RAND_1608;
  reg [31:0] _RAND_1609;
  reg [31:0] _RAND_1610;
  reg [31:0] _RAND_1611;
  reg [31:0] _RAND_1612;
  reg [31:0] _RAND_1613;
  reg [31:0] _RAND_1614;
  reg [31:0] _RAND_1615;
  reg [31:0] _RAND_1616;
  reg [31:0] _RAND_1617;
  reg [31:0] _RAND_1618;
  reg [31:0] _RAND_1619;
  reg [31:0] _RAND_1620;
  reg [31:0] _RAND_1621;
  reg [31:0] _RAND_1622;
  reg [31:0] _RAND_1623;
  reg [31:0] _RAND_1624;
  reg [31:0] _RAND_1625;
  reg [31:0] _RAND_1626;
  reg [31:0] _RAND_1627;
  reg [31:0] _RAND_1628;
  reg [31:0] _RAND_1629;
  reg [31:0] _RAND_1630;
  reg [31:0] _RAND_1631;
  reg [31:0] _RAND_1632;
  reg [31:0] _RAND_1633;
  reg [31:0] _RAND_1634;
  reg [31:0] _RAND_1635;
  reg [31:0] _RAND_1636;
  reg [31:0] _RAND_1637;
  reg [31:0] _RAND_1638;
  reg [31:0] _RAND_1639;
  reg [31:0] _RAND_1640;
  reg [31:0] _RAND_1641;
  reg [31:0] _RAND_1642;
  reg [31:0] _RAND_1643;
  reg [31:0] _RAND_1644;
  reg [31:0] _RAND_1645;
  reg [31:0] _RAND_1646;
  reg [31:0] _RAND_1647;
  reg [31:0] _RAND_1648;
  reg [31:0] _RAND_1649;
  reg [31:0] _RAND_1650;
  reg [31:0] _RAND_1651;
  reg [31:0] _RAND_1652;
  reg [31:0] _RAND_1653;
  reg [31:0] _RAND_1654;
  reg [31:0] _RAND_1655;
  reg [31:0] _RAND_1656;
  reg [31:0] _RAND_1657;
  reg [31:0] _RAND_1658;
  reg [31:0] _RAND_1659;
  reg [31:0] _RAND_1660;
  reg [31:0] _RAND_1661;
  reg [31:0] _RAND_1662;
  reg [31:0] _RAND_1663;
  reg [31:0] _RAND_1664;
  reg [31:0] _RAND_1665;
  reg [31:0] _RAND_1666;
  reg [31:0] _RAND_1667;
  reg [31:0] _RAND_1668;
  reg [31:0] _RAND_1669;
  reg [31:0] _RAND_1670;
  reg [31:0] _RAND_1671;
  reg [31:0] _RAND_1672;
  reg [31:0] _RAND_1673;
  reg [31:0] _RAND_1674;
  reg [31:0] _RAND_1675;
  reg [31:0] _RAND_1676;
  reg [31:0] _RAND_1677;
  reg [31:0] _RAND_1678;
  reg [31:0] _RAND_1679;
  reg [31:0] _RAND_1680;
  reg [31:0] _RAND_1681;
  reg [31:0] _RAND_1682;
  reg [31:0] _RAND_1683;
  reg [31:0] _RAND_1684;
  reg [31:0] _RAND_1685;
  reg [31:0] _RAND_1686;
  reg [31:0] _RAND_1687;
  reg [31:0] _RAND_1688;
  reg [31:0] _RAND_1689;
  reg [31:0] _RAND_1690;
  reg [31:0] _RAND_1691;
  reg [31:0] _RAND_1692;
  reg [31:0] _RAND_1693;
  reg [31:0] _RAND_1694;
  reg [31:0] _RAND_1695;
  reg [31:0] _RAND_1696;
  reg [31:0] _RAND_1697;
  reg [31:0] _RAND_1698;
  reg [31:0] _RAND_1699;
  reg [31:0] _RAND_1700;
  reg [31:0] _RAND_1701;
  reg [31:0] _RAND_1702;
  reg [31:0] _RAND_1703;
  reg [31:0] _RAND_1704;
  reg [31:0] _RAND_1705;
  reg [31:0] _RAND_1706;
  reg [31:0] _RAND_1707;
  reg [31:0] _RAND_1708;
  reg [31:0] _RAND_1709;
  reg [31:0] _RAND_1710;
  reg [31:0] _RAND_1711;
  reg [31:0] _RAND_1712;
  reg [31:0] _RAND_1713;
  reg [31:0] _RAND_1714;
  reg [31:0] _RAND_1715;
  reg [31:0] _RAND_1716;
  reg [31:0] _RAND_1717;
  reg [31:0] _RAND_1718;
  reg [31:0] _RAND_1719;
  reg [31:0] _RAND_1720;
  reg [31:0] _RAND_1721;
  reg [31:0] _RAND_1722;
  reg [31:0] _RAND_1723;
  reg [31:0] _RAND_1724;
  reg [31:0] _RAND_1725;
  reg [31:0] _RAND_1726;
  reg [31:0] _RAND_1727;
  reg [31:0] _RAND_1728;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] image_0_0; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_1; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_2; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_3; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_4; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_5; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_6; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_7; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_8; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_9; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_10; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_11; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_12; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_13; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_14; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_15; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_16; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_17; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_18; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_19; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_20; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_21; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_22; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_23; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_24; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_25; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_26; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_27; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_28; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_29; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_30; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_31; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_32; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_33; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_34; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_35; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_36; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_37; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_38; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_39; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_40; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_41; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_42; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_43; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_44; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_45; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_46; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_47; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_48; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_49; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_50; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_51; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_52; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_53; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_54; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_55; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_56; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_57; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_58; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_59; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_60; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_61; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_62; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_63; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_64; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_65; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_66; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_67; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_68; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_69; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_70; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_71; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_72; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_73; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_74; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_75; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_76; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_77; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_78; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_79; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_80; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_81; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_82; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_83; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_84; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_85; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_86; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_87; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_88; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_89; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_90; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_91; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_92; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_93; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_94; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_95; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_96; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_97; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_98; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_99; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_100; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_101; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_102; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_103; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_104; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_105; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_106; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_107; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_108; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_109; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_110; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_111; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_112; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_113; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_114; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_115; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_116; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_117; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_118; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_119; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_120; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_121; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_122; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_123; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_124; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_125; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_126; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_127; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_128; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_129; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_130; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_131; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_132; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_133; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_134; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_135; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_136; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_137; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_138; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_139; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_140; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_141; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_142; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_143; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_144; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_145; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_146; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_147; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_148; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_149; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_150; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_151; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_152; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_153; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_154; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_155; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_156; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_157; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_158; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_159; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_160; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_161; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_162; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_163; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_164; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_165; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_166; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_167; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_168; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_169; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_170; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_171; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_172; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_173; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_174; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_175; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_176; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_177; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_178; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_179; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_180; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_181; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_182; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_183; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_184; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_185; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_186; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_187; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_188; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_189; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_190; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_191; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_192; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_193; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_194; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_195; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_196; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_197; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_198; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_199; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_200; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_201; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_202; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_203; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_204; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_205; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_206; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_207; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_208; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_209; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_210; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_211; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_212; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_213; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_214; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_215; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_216; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_217; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_218; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_219; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_220; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_221; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_222; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_223; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_224; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_225; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_226; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_227; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_228; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_229; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_230; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_231; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_232; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_233; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_234; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_235; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_236; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_237; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_238; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_239; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_240; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_241; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_242; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_243; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_244; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_245; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_246; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_247; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_248; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_249; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_250; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_251; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_252; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_253; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_254; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_255; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_256; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_257; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_258; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_259; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_260; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_261; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_262; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_263; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_264; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_265; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_266; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_267; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_268; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_269; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_270; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_271; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_272; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_273; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_274; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_275; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_276; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_277; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_278; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_279; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_280; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_281; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_282; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_283; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_284; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_285; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_286; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_287; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_288; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_289; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_290; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_291; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_292; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_293; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_294; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_295; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_296; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_297; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_298; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_299; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_300; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_301; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_302; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_303; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_304; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_305; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_306; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_307; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_308; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_309; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_310; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_311; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_312; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_313; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_314; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_315; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_316; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_317; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_318; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_319; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_320; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_321; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_322; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_323; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_324; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_325; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_326; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_327; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_328; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_329; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_330; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_331; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_332; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_333; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_334; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_335; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_336; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_337; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_338; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_339; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_340; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_341; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_342; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_343; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_344; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_345; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_346; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_347; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_348; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_349; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_350; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_351; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_352; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_353; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_354; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_355; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_356; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_357; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_358; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_359; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_360; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_361; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_362; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_363; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_364; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_365; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_366; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_367; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_368; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_369; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_370; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_371; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_372; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_373; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_374; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_375; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_376; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_377; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_378; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_379; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_380; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_381; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_382; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_383; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_384; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_385; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_386; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_387; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_388; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_389; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_390; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_391; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_392; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_393; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_394; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_395; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_396; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_397; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_398; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_399; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_400; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_401; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_402; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_403; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_404; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_405; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_406; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_407; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_408; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_409; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_410; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_411; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_412; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_413; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_414; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_415; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_416; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_417; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_418; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_419; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_420; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_421; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_422; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_423; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_424; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_425; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_426; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_427; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_428; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_429; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_430; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_431; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_432; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_433; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_434; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_435; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_436; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_437; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_438; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_439; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_440; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_441; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_442; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_443; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_444; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_445; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_446; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_447; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_448; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_449; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_450; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_451; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_452; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_453; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_454; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_455; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_456; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_457; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_458; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_459; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_460; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_461; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_462; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_463; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_464; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_465; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_466; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_467; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_468; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_469; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_470; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_471; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_472; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_473; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_474; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_475; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_476; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_477; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_478; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_479; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_480; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_481; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_482; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_483; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_484; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_485; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_486; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_487; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_488; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_489; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_490; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_491; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_492; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_493; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_494; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_495; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_496; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_497; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_498; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_499; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_500; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_501; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_502; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_503; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_504; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_505; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_506; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_507; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_508; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_509; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_510; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_511; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_512; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_513; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_514; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_515; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_516; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_517; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_518; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_519; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_520; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_521; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_522; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_523; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_524; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_525; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_526; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_527; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_528; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_529; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_530; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_531; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_532; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_533; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_534; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_535; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_536; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_537; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_538; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_539; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_540; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_541; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_542; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_543; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_544; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_545; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_546; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_547; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_548; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_549; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_550; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_551; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_552; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_553; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_554; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_555; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_556; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_557; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_558; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_559; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_560; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_561; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_562; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_563; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_564; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_565; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_566; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_567; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_568; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_569; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_570; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_571; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_572; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_573; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_574; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_575; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_1_0; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_1; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_2; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_3; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_4; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_5; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_6; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_7; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_8; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_9; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_10; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_11; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_12; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_13; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_14; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_15; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_16; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_17; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_18; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_19; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_20; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_21; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_22; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_23; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_24; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_25; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_26; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_27; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_28; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_29; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_30; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_31; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_32; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_33; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_34; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_35; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_36; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_37; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_38; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_39; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_40; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_41; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_42; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_43; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_44; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_45; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_46; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_47; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_48; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_49; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_50; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_51; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_52; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_53; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_54; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_55; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_56; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_57; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_58; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_59; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_60; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_61; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_62; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_63; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_64; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_65; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_66; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_67; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_68; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_69; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_70; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_71; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_72; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_73; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_74; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_75; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_76; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_77; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_78; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_79; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_80; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_81; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_82; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_83; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_84; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_85; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_86; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_87; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_88; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_89; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_90; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_91; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_92; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_93; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_94; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_95; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_96; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_97; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_98; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_99; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_100; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_101; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_102; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_103; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_104; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_105; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_106; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_107; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_108; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_109; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_110; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_111; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_112; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_113; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_114; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_115; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_116; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_117; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_118; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_119; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_120; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_121; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_122; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_123; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_124; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_125; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_126; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_127; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_128; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_129; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_130; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_131; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_132; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_133; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_134; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_135; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_136; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_137; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_138; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_139; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_140; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_141; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_142; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_143; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_144; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_145; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_146; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_147; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_148; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_149; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_150; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_151; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_152; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_153; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_154; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_155; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_156; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_157; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_158; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_159; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_160; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_161; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_162; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_163; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_164; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_165; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_166; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_167; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_168; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_169; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_170; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_171; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_172; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_173; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_174; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_175; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_176; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_177; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_178; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_179; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_180; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_181; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_182; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_183; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_184; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_185; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_186; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_187; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_188; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_189; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_190; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_191; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_192; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_193; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_194; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_195; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_196; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_197; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_198; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_199; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_200; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_201; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_202; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_203; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_204; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_205; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_206; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_207; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_208; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_209; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_210; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_211; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_212; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_213; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_214; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_215; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_216; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_217; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_218; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_219; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_220; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_221; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_222; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_223; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_224; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_225; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_226; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_227; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_228; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_229; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_230; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_231; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_232; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_233; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_234; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_235; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_236; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_237; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_238; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_239; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_240; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_241; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_242; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_243; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_244; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_245; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_246; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_247; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_248; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_249; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_250; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_251; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_252; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_253; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_254; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_255; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_256; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_257; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_258; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_259; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_260; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_261; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_262; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_263; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_264; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_265; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_266; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_267; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_268; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_269; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_270; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_271; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_272; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_273; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_274; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_275; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_276; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_277; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_278; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_279; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_280; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_281; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_282; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_283; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_284; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_285; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_286; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_287; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_288; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_289; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_290; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_291; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_292; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_293; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_294; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_295; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_296; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_297; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_298; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_299; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_300; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_301; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_302; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_303; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_304; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_305; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_306; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_307; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_308; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_309; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_310; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_311; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_312; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_313; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_314; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_315; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_316; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_317; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_318; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_319; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_320; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_321; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_322; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_323; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_324; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_325; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_326; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_327; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_328; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_329; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_330; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_331; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_332; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_333; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_334; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_335; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_336; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_337; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_338; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_339; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_340; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_341; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_342; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_343; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_344; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_345; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_346; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_347; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_348; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_349; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_350; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_351; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_352; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_353; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_354; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_355; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_356; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_357; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_358; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_359; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_360; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_361; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_362; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_363; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_364; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_365; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_366; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_367; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_368; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_369; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_370; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_371; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_372; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_373; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_374; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_375; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_376; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_377; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_378; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_379; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_380; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_381; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_382; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_383; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_384; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_385; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_386; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_387; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_388; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_389; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_390; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_391; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_392; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_393; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_394; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_395; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_396; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_397; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_398; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_399; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_400; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_401; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_402; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_403; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_404; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_405; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_406; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_407; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_408; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_409; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_410; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_411; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_412; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_413; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_414; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_415; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_416; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_417; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_418; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_419; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_420; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_421; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_422; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_423; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_424; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_425; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_426; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_427; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_428; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_429; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_430; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_431; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_432; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_433; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_434; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_435; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_436; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_437; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_438; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_439; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_440; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_441; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_442; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_443; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_444; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_445; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_446; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_447; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_448; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_449; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_450; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_451; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_452; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_453; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_454; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_455; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_456; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_457; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_458; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_459; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_460; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_461; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_462; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_463; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_464; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_465; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_466; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_467; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_468; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_469; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_470; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_471; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_472; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_473; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_474; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_475; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_476; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_477; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_478; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_479; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_480; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_481; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_482; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_483; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_484; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_485; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_486; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_487; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_488; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_489; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_490; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_491; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_492; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_493; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_494; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_495; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_496; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_497; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_498; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_499; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_500; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_501; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_502; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_503; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_504; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_505; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_506; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_507; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_508; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_509; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_510; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_511; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_512; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_513; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_514; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_515; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_516; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_517; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_518; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_519; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_520; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_521; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_522; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_523; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_524; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_525; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_526; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_527; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_528; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_529; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_530; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_531; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_532; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_533; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_534; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_535; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_536; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_537; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_538; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_539; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_540; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_541; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_542; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_543; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_544; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_545; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_546; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_547; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_548; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_549; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_550; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_551; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_552; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_553; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_554; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_555; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_556; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_557; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_558; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_559; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_560; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_561; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_562; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_563; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_564; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_565; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_566; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_567; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_568; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_569; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_570; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_571; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_572; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_573; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_574; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_575; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_2_0; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_1; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_2; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_3; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_4; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_5; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_6; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_7; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_8; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_9; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_10; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_11; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_12; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_13; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_14; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_15; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_16; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_17; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_18; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_19; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_20; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_21; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_22; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_23; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_24; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_25; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_26; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_27; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_28; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_29; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_30; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_31; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_32; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_33; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_34; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_35; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_36; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_37; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_38; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_39; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_40; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_41; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_42; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_43; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_44; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_45; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_46; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_47; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_48; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_49; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_50; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_51; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_52; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_53; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_54; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_55; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_56; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_57; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_58; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_59; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_60; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_61; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_62; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_63; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_64; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_65; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_66; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_67; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_68; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_69; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_70; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_71; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_72; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_73; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_74; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_75; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_76; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_77; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_78; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_79; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_80; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_81; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_82; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_83; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_84; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_85; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_86; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_87; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_88; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_89; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_90; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_91; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_92; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_93; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_94; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_95; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_96; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_97; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_98; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_99; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_100; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_101; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_102; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_103; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_104; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_105; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_106; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_107; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_108; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_109; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_110; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_111; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_112; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_113; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_114; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_115; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_116; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_117; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_118; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_119; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_120; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_121; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_122; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_123; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_124; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_125; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_126; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_127; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_128; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_129; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_130; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_131; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_132; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_133; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_134; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_135; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_136; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_137; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_138; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_139; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_140; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_141; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_142; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_143; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_144; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_145; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_146; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_147; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_148; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_149; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_150; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_151; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_152; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_153; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_154; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_155; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_156; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_157; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_158; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_159; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_160; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_161; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_162; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_163; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_164; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_165; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_166; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_167; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_168; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_169; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_170; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_171; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_172; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_173; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_174; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_175; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_176; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_177; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_178; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_179; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_180; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_181; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_182; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_183; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_184; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_185; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_186; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_187; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_188; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_189; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_190; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_191; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_192; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_193; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_194; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_195; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_196; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_197; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_198; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_199; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_200; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_201; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_202; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_203; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_204; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_205; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_206; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_207; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_208; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_209; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_210; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_211; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_212; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_213; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_214; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_215; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_216; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_217; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_218; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_219; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_220; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_221; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_222; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_223; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_224; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_225; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_226; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_227; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_228; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_229; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_230; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_231; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_232; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_233; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_234; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_235; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_236; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_237; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_238; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_239; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_240; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_241; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_242; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_243; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_244; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_245; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_246; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_247; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_248; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_249; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_250; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_251; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_252; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_253; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_254; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_255; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_256; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_257; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_258; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_259; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_260; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_261; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_262; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_263; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_264; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_265; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_266; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_267; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_268; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_269; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_270; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_271; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_272; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_273; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_274; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_275; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_276; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_277; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_278; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_279; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_280; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_281; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_282; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_283; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_284; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_285; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_286; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_287; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_288; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_289; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_290; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_291; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_292; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_293; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_294; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_295; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_296; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_297; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_298; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_299; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_300; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_301; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_302; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_303; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_304; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_305; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_306; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_307; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_308; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_309; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_310; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_311; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_312; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_313; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_314; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_315; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_316; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_317; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_318; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_319; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_320; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_321; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_322; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_323; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_324; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_325; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_326; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_327; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_328; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_329; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_330; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_331; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_332; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_333; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_334; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_335; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_336; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_337; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_338; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_339; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_340; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_341; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_342; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_343; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_344; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_345; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_346; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_347; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_348; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_349; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_350; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_351; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_352; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_353; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_354; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_355; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_356; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_357; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_358; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_359; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_360; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_361; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_362; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_363; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_364; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_365; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_366; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_367; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_368; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_369; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_370; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_371; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_372; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_373; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_374; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_375; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_376; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_377; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_378; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_379; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_380; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_381; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_382; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_383; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_384; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_385; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_386; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_387; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_388; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_389; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_390; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_391; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_392; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_393; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_394; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_395; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_396; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_397; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_398; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_399; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_400; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_401; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_402; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_403; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_404; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_405; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_406; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_407; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_408; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_409; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_410; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_411; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_412; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_413; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_414; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_415; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_416; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_417; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_418; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_419; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_420; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_421; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_422; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_423; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_424; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_425; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_426; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_427; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_428; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_429; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_430; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_431; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_432; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_433; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_434; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_435; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_436; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_437; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_438; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_439; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_440; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_441; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_442; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_443; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_444; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_445; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_446; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_447; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_448; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_449; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_450; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_451; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_452; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_453; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_454; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_455; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_456; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_457; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_458; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_459; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_460; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_461; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_462; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_463; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_464; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_465; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_466; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_467; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_468; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_469; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_470; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_471; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_472; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_473; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_474; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_475; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_476; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_477; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_478; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_479; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_480; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_481; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_482; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_483; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_484; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_485; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_486; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_487; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_488; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_489; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_490; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_491; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_492; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_493; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_494; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_495; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_496; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_497; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_498; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_499; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_500; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_501; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_502; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_503; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_504; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_505; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_506; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_507; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_508; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_509; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_510; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_511; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_512; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_513; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_514; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_515; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_516; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_517; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_518; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_519; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_520; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_521; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_522; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_523; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_524; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_525; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_526; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_527; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_528; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_529; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_530; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_531; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_532; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_533; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_534; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_535; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_536; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_537; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_538; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_539; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_540; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_541; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_542; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_543; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_544; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_545; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_546; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_547; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_548; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_549; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_550; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_551; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_552; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_553; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_554; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_555; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_556; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_557; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_558; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_559; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_560; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_561; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_562; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_563; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_564; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_565; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_566; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_567; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_568; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_569; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_570; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_571; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_572; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_573; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_574; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_575; // @[VideoBuffer.scala 21:25]
  reg [31:0] pixelIndex; // @[VideoBuffer.scala 24:33]
  wire [16:0] _T_3 = io_rowIndex * 11'h20; // @[VideoBuffer.scala 27:54]
  wire [16:0] _GEN_17282 = {{6'd0}, io_colIndex}; // @[VideoBuffer.scala 27:69]
  wire [16:0] _T_5 = _T_3 + _GEN_17282; // @[VideoBuffer.scala 27:69]
  wire [3:0] _GEN_1 = 10'h1 == _T_5[9:0] ? image_0_1 : image_0_0; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2 = 10'h2 == _T_5[9:0] ? image_0_2 : _GEN_1; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3 = 10'h3 == _T_5[9:0] ? image_0_3 : _GEN_2; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4 = 10'h4 == _T_5[9:0] ? image_0_4 : _GEN_3; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_5 = 10'h5 == _T_5[9:0] ? image_0_5 : _GEN_4; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_6 = 10'h6 == _T_5[9:0] ? image_0_6 : _GEN_5; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_7 = 10'h7 == _T_5[9:0] ? image_0_7 : _GEN_6; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_8 = 10'h8 == _T_5[9:0] ? image_0_8 : _GEN_7; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_9 = 10'h9 == _T_5[9:0] ? image_0_9 : _GEN_8; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_10 = 10'ha == _T_5[9:0] ? image_0_10 : _GEN_9; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_11 = 10'hb == _T_5[9:0] ? image_0_11 : _GEN_10; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_12 = 10'hc == _T_5[9:0] ? image_0_12 : _GEN_11; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_13 = 10'hd == _T_5[9:0] ? image_0_13 : _GEN_12; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_14 = 10'he == _T_5[9:0] ? image_0_14 : _GEN_13; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_15 = 10'hf == _T_5[9:0] ? image_0_15 : _GEN_14; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_16 = 10'h10 == _T_5[9:0] ? image_0_16 : _GEN_15; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_17 = 10'h11 == _T_5[9:0] ? image_0_17 : _GEN_16; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_18 = 10'h12 == _T_5[9:0] ? image_0_18 : _GEN_17; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_19 = 10'h13 == _T_5[9:0] ? image_0_19 : _GEN_18; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_20 = 10'h14 == _T_5[9:0] ? image_0_20 : _GEN_19; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_21 = 10'h15 == _T_5[9:0] ? image_0_21 : _GEN_20; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_22 = 10'h16 == _T_5[9:0] ? image_0_22 : _GEN_21; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_23 = 10'h17 == _T_5[9:0] ? image_0_23 : _GEN_22; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_24 = 10'h18 == _T_5[9:0] ? image_0_24 : _GEN_23; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_25 = 10'h19 == _T_5[9:0] ? image_0_25 : _GEN_24; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_26 = 10'h1a == _T_5[9:0] ? image_0_26 : _GEN_25; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_27 = 10'h1b == _T_5[9:0] ? image_0_27 : _GEN_26; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_28 = 10'h1c == _T_5[9:0] ? image_0_28 : _GEN_27; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_29 = 10'h1d == _T_5[9:0] ? image_0_29 : _GEN_28; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_30 = 10'h1e == _T_5[9:0] ? image_0_30 : _GEN_29; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_31 = 10'h1f == _T_5[9:0] ? image_0_31 : _GEN_30; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_32 = 10'h20 == _T_5[9:0] ? image_0_32 : _GEN_31; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_33 = 10'h21 == _T_5[9:0] ? image_0_33 : _GEN_32; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_34 = 10'h22 == _T_5[9:0] ? image_0_34 : _GEN_33; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_35 = 10'h23 == _T_5[9:0] ? image_0_35 : _GEN_34; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_36 = 10'h24 == _T_5[9:0] ? image_0_36 : _GEN_35; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_37 = 10'h25 == _T_5[9:0] ? image_0_37 : _GEN_36; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_38 = 10'h26 == _T_5[9:0] ? image_0_38 : _GEN_37; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_39 = 10'h27 == _T_5[9:0] ? image_0_39 : _GEN_38; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_40 = 10'h28 == _T_5[9:0] ? image_0_40 : _GEN_39; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_41 = 10'h29 == _T_5[9:0] ? image_0_41 : _GEN_40; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_42 = 10'h2a == _T_5[9:0] ? image_0_42 : _GEN_41; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_43 = 10'h2b == _T_5[9:0] ? image_0_43 : _GEN_42; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_44 = 10'h2c == _T_5[9:0] ? image_0_44 : _GEN_43; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_45 = 10'h2d == _T_5[9:0] ? image_0_45 : _GEN_44; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_46 = 10'h2e == _T_5[9:0] ? image_0_46 : _GEN_45; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_47 = 10'h2f == _T_5[9:0] ? image_0_47 : _GEN_46; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_48 = 10'h30 == _T_5[9:0] ? image_0_48 : _GEN_47; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_49 = 10'h31 == _T_5[9:0] ? image_0_49 : _GEN_48; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_50 = 10'h32 == _T_5[9:0] ? image_0_50 : _GEN_49; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_51 = 10'h33 == _T_5[9:0] ? image_0_51 : _GEN_50; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_52 = 10'h34 == _T_5[9:0] ? image_0_52 : _GEN_51; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_53 = 10'h35 == _T_5[9:0] ? image_0_53 : _GEN_52; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_54 = 10'h36 == _T_5[9:0] ? image_0_54 : _GEN_53; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_55 = 10'h37 == _T_5[9:0] ? image_0_55 : _GEN_54; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_56 = 10'h38 == _T_5[9:0] ? image_0_56 : _GEN_55; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_57 = 10'h39 == _T_5[9:0] ? image_0_57 : _GEN_56; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_58 = 10'h3a == _T_5[9:0] ? image_0_58 : _GEN_57; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_59 = 10'h3b == _T_5[9:0] ? image_0_59 : _GEN_58; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_60 = 10'h3c == _T_5[9:0] ? image_0_60 : _GEN_59; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_61 = 10'h3d == _T_5[9:0] ? image_0_61 : _GEN_60; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_62 = 10'h3e == _T_5[9:0] ? image_0_62 : _GEN_61; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_63 = 10'h3f == _T_5[9:0] ? image_0_63 : _GEN_62; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_64 = 10'h40 == _T_5[9:0] ? image_0_64 : _GEN_63; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_65 = 10'h41 == _T_5[9:0] ? image_0_65 : _GEN_64; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_66 = 10'h42 == _T_5[9:0] ? image_0_66 : _GEN_65; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_67 = 10'h43 == _T_5[9:0] ? image_0_67 : _GEN_66; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_68 = 10'h44 == _T_5[9:0] ? image_0_68 : _GEN_67; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_69 = 10'h45 == _T_5[9:0] ? image_0_69 : _GEN_68; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_70 = 10'h46 == _T_5[9:0] ? image_0_70 : _GEN_69; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_71 = 10'h47 == _T_5[9:0] ? image_0_71 : _GEN_70; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_72 = 10'h48 == _T_5[9:0] ? image_0_72 : _GEN_71; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_73 = 10'h49 == _T_5[9:0] ? image_0_73 : _GEN_72; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_74 = 10'h4a == _T_5[9:0] ? image_0_74 : _GEN_73; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_75 = 10'h4b == _T_5[9:0] ? image_0_75 : _GEN_74; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_76 = 10'h4c == _T_5[9:0] ? image_0_76 : _GEN_75; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_77 = 10'h4d == _T_5[9:0] ? image_0_77 : _GEN_76; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_78 = 10'h4e == _T_5[9:0] ? image_0_78 : _GEN_77; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_79 = 10'h4f == _T_5[9:0] ? image_0_79 : _GEN_78; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_80 = 10'h50 == _T_5[9:0] ? image_0_80 : _GEN_79; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_81 = 10'h51 == _T_5[9:0] ? image_0_81 : _GEN_80; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_82 = 10'h52 == _T_5[9:0] ? image_0_82 : _GEN_81; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_83 = 10'h53 == _T_5[9:0] ? image_0_83 : _GEN_82; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_84 = 10'h54 == _T_5[9:0] ? image_0_84 : _GEN_83; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_85 = 10'h55 == _T_5[9:0] ? image_0_85 : _GEN_84; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_86 = 10'h56 == _T_5[9:0] ? image_0_86 : _GEN_85; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_87 = 10'h57 == _T_5[9:0] ? image_0_87 : _GEN_86; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_88 = 10'h58 == _T_5[9:0] ? image_0_88 : _GEN_87; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_89 = 10'h59 == _T_5[9:0] ? image_0_89 : _GEN_88; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_90 = 10'h5a == _T_5[9:0] ? image_0_90 : _GEN_89; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_91 = 10'h5b == _T_5[9:0] ? image_0_91 : _GEN_90; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_92 = 10'h5c == _T_5[9:0] ? image_0_92 : _GEN_91; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_93 = 10'h5d == _T_5[9:0] ? image_0_93 : _GEN_92; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_94 = 10'h5e == _T_5[9:0] ? image_0_94 : _GEN_93; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_95 = 10'h5f == _T_5[9:0] ? image_0_95 : _GEN_94; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_96 = 10'h60 == _T_5[9:0] ? image_0_96 : _GEN_95; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_97 = 10'h61 == _T_5[9:0] ? image_0_97 : _GEN_96; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_98 = 10'h62 == _T_5[9:0] ? image_0_98 : _GEN_97; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_99 = 10'h63 == _T_5[9:0] ? image_0_99 : _GEN_98; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_100 = 10'h64 == _T_5[9:0] ? image_0_100 : _GEN_99; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_101 = 10'h65 == _T_5[9:0] ? image_0_101 : _GEN_100; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_102 = 10'h66 == _T_5[9:0] ? image_0_102 : _GEN_101; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_103 = 10'h67 == _T_5[9:0] ? image_0_103 : _GEN_102; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_104 = 10'h68 == _T_5[9:0] ? image_0_104 : _GEN_103; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_105 = 10'h69 == _T_5[9:0] ? image_0_105 : _GEN_104; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_106 = 10'h6a == _T_5[9:0] ? image_0_106 : _GEN_105; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_107 = 10'h6b == _T_5[9:0] ? image_0_107 : _GEN_106; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_108 = 10'h6c == _T_5[9:0] ? image_0_108 : _GEN_107; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_109 = 10'h6d == _T_5[9:0] ? image_0_109 : _GEN_108; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_110 = 10'h6e == _T_5[9:0] ? image_0_110 : _GEN_109; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_111 = 10'h6f == _T_5[9:0] ? image_0_111 : _GEN_110; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_112 = 10'h70 == _T_5[9:0] ? image_0_112 : _GEN_111; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_113 = 10'h71 == _T_5[9:0] ? image_0_113 : _GEN_112; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_114 = 10'h72 == _T_5[9:0] ? image_0_114 : _GEN_113; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_115 = 10'h73 == _T_5[9:0] ? image_0_115 : _GEN_114; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_116 = 10'h74 == _T_5[9:0] ? image_0_116 : _GEN_115; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_117 = 10'h75 == _T_5[9:0] ? image_0_117 : _GEN_116; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_118 = 10'h76 == _T_5[9:0] ? image_0_118 : _GEN_117; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_119 = 10'h77 == _T_5[9:0] ? image_0_119 : _GEN_118; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_120 = 10'h78 == _T_5[9:0] ? image_0_120 : _GEN_119; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_121 = 10'h79 == _T_5[9:0] ? image_0_121 : _GEN_120; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_122 = 10'h7a == _T_5[9:0] ? image_0_122 : _GEN_121; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_123 = 10'h7b == _T_5[9:0] ? image_0_123 : _GEN_122; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_124 = 10'h7c == _T_5[9:0] ? image_0_124 : _GEN_123; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_125 = 10'h7d == _T_5[9:0] ? image_0_125 : _GEN_124; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_126 = 10'h7e == _T_5[9:0] ? image_0_126 : _GEN_125; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_127 = 10'h7f == _T_5[9:0] ? image_0_127 : _GEN_126; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_128 = 10'h80 == _T_5[9:0] ? image_0_128 : _GEN_127; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_129 = 10'h81 == _T_5[9:0] ? image_0_129 : _GEN_128; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_130 = 10'h82 == _T_5[9:0] ? image_0_130 : _GEN_129; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_131 = 10'h83 == _T_5[9:0] ? image_0_131 : _GEN_130; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_132 = 10'h84 == _T_5[9:0] ? image_0_132 : _GEN_131; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_133 = 10'h85 == _T_5[9:0] ? image_0_133 : _GEN_132; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_134 = 10'h86 == _T_5[9:0] ? image_0_134 : _GEN_133; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_135 = 10'h87 == _T_5[9:0] ? image_0_135 : _GEN_134; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_136 = 10'h88 == _T_5[9:0] ? image_0_136 : _GEN_135; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_137 = 10'h89 == _T_5[9:0] ? image_0_137 : _GEN_136; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_138 = 10'h8a == _T_5[9:0] ? image_0_138 : _GEN_137; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_139 = 10'h8b == _T_5[9:0] ? image_0_139 : _GEN_138; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_140 = 10'h8c == _T_5[9:0] ? image_0_140 : _GEN_139; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_141 = 10'h8d == _T_5[9:0] ? image_0_141 : _GEN_140; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_142 = 10'h8e == _T_5[9:0] ? image_0_142 : _GEN_141; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_143 = 10'h8f == _T_5[9:0] ? image_0_143 : _GEN_142; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_144 = 10'h90 == _T_5[9:0] ? image_0_144 : _GEN_143; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_145 = 10'h91 == _T_5[9:0] ? image_0_145 : _GEN_144; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_146 = 10'h92 == _T_5[9:0] ? image_0_146 : _GEN_145; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_147 = 10'h93 == _T_5[9:0] ? image_0_147 : _GEN_146; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_148 = 10'h94 == _T_5[9:0] ? image_0_148 : _GEN_147; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_149 = 10'h95 == _T_5[9:0] ? image_0_149 : _GEN_148; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_150 = 10'h96 == _T_5[9:0] ? image_0_150 : _GEN_149; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_151 = 10'h97 == _T_5[9:0] ? image_0_151 : _GEN_150; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_152 = 10'h98 == _T_5[9:0] ? image_0_152 : _GEN_151; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_153 = 10'h99 == _T_5[9:0] ? image_0_153 : _GEN_152; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_154 = 10'h9a == _T_5[9:0] ? image_0_154 : _GEN_153; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_155 = 10'h9b == _T_5[9:0] ? image_0_155 : _GEN_154; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_156 = 10'h9c == _T_5[9:0] ? image_0_156 : _GEN_155; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_157 = 10'h9d == _T_5[9:0] ? image_0_157 : _GEN_156; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_158 = 10'h9e == _T_5[9:0] ? image_0_158 : _GEN_157; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_159 = 10'h9f == _T_5[9:0] ? image_0_159 : _GEN_158; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_160 = 10'ha0 == _T_5[9:0] ? image_0_160 : _GEN_159; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_161 = 10'ha1 == _T_5[9:0] ? image_0_161 : _GEN_160; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_162 = 10'ha2 == _T_5[9:0] ? image_0_162 : _GEN_161; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_163 = 10'ha3 == _T_5[9:0] ? image_0_163 : _GEN_162; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_164 = 10'ha4 == _T_5[9:0] ? image_0_164 : _GEN_163; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_165 = 10'ha5 == _T_5[9:0] ? image_0_165 : _GEN_164; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_166 = 10'ha6 == _T_5[9:0] ? image_0_166 : _GEN_165; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_167 = 10'ha7 == _T_5[9:0] ? image_0_167 : _GEN_166; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_168 = 10'ha8 == _T_5[9:0] ? image_0_168 : _GEN_167; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_169 = 10'ha9 == _T_5[9:0] ? image_0_169 : _GEN_168; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_170 = 10'haa == _T_5[9:0] ? image_0_170 : _GEN_169; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_171 = 10'hab == _T_5[9:0] ? image_0_171 : _GEN_170; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_172 = 10'hac == _T_5[9:0] ? image_0_172 : _GEN_171; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_173 = 10'had == _T_5[9:0] ? image_0_173 : _GEN_172; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_174 = 10'hae == _T_5[9:0] ? image_0_174 : _GEN_173; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_175 = 10'haf == _T_5[9:0] ? image_0_175 : _GEN_174; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_176 = 10'hb0 == _T_5[9:0] ? image_0_176 : _GEN_175; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_177 = 10'hb1 == _T_5[9:0] ? image_0_177 : _GEN_176; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_178 = 10'hb2 == _T_5[9:0] ? image_0_178 : _GEN_177; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_179 = 10'hb3 == _T_5[9:0] ? image_0_179 : _GEN_178; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_180 = 10'hb4 == _T_5[9:0] ? image_0_180 : _GEN_179; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_181 = 10'hb5 == _T_5[9:0] ? image_0_181 : _GEN_180; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_182 = 10'hb6 == _T_5[9:0] ? image_0_182 : _GEN_181; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_183 = 10'hb7 == _T_5[9:0] ? image_0_183 : _GEN_182; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_184 = 10'hb8 == _T_5[9:0] ? image_0_184 : _GEN_183; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_185 = 10'hb9 == _T_5[9:0] ? image_0_185 : _GEN_184; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_186 = 10'hba == _T_5[9:0] ? image_0_186 : _GEN_185; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_187 = 10'hbb == _T_5[9:0] ? image_0_187 : _GEN_186; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_188 = 10'hbc == _T_5[9:0] ? image_0_188 : _GEN_187; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_189 = 10'hbd == _T_5[9:0] ? image_0_189 : _GEN_188; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_190 = 10'hbe == _T_5[9:0] ? image_0_190 : _GEN_189; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_191 = 10'hbf == _T_5[9:0] ? image_0_191 : _GEN_190; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_192 = 10'hc0 == _T_5[9:0] ? image_0_192 : _GEN_191; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_193 = 10'hc1 == _T_5[9:0] ? image_0_193 : _GEN_192; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_194 = 10'hc2 == _T_5[9:0] ? image_0_194 : _GEN_193; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_195 = 10'hc3 == _T_5[9:0] ? image_0_195 : _GEN_194; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_196 = 10'hc4 == _T_5[9:0] ? image_0_196 : _GEN_195; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_197 = 10'hc5 == _T_5[9:0] ? image_0_197 : _GEN_196; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_198 = 10'hc6 == _T_5[9:0] ? image_0_198 : _GEN_197; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_199 = 10'hc7 == _T_5[9:0] ? image_0_199 : _GEN_198; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_200 = 10'hc8 == _T_5[9:0] ? image_0_200 : _GEN_199; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_201 = 10'hc9 == _T_5[9:0] ? image_0_201 : _GEN_200; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_202 = 10'hca == _T_5[9:0] ? image_0_202 : _GEN_201; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_203 = 10'hcb == _T_5[9:0] ? image_0_203 : _GEN_202; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_204 = 10'hcc == _T_5[9:0] ? image_0_204 : _GEN_203; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_205 = 10'hcd == _T_5[9:0] ? image_0_205 : _GEN_204; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_206 = 10'hce == _T_5[9:0] ? image_0_206 : _GEN_205; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_207 = 10'hcf == _T_5[9:0] ? image_0_207 : _GEN_206; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_208 = 10'hd0 == _T_5[9:0] ? image_0_208 : _GEN_207; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_209 = 10'hd1 == _T_5[9:0] ? image_0_209 : _GEN_208; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_210 = 10'hd2 == _T_5[9:0] ? image_0_210 : _GEN_209; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_211 = 10'hd3 == _T_5[9:0] ? image_0_211 : _GEN_210; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_212 = 10'hd4 == _T_5[9:0] ? image_0_212 : _GEN_211; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_213 = 10'hd5 == _T_5[9:0] ? image_0_213 : _GEN_212; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_214 = 10'hd6 == _T_5[9:0] ? image_0_214 : _GEN_213; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_215 = 10'hd7 == _T_5[9:0] ? image_0_215 : _GEN_214; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_216 = 10'hd8 == _T_5[9:0] ? image_0_216 : _GEN_215; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_217 = 10'hd9 == _T_5[9:0] ? image_0_217 : _GEN_216; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_218 = 10'hda == _T_5[9:0] ? image_0_218 : _GEN_217; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_219 = 10'hdb == _T_5[9:0] ? image_0_219 : _GEN_218; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_220 = 10'hdc == _T_5[9:0] ? image_0_220 : _GEN_219; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_221 = 10'hdd == _T_5[9:0] ? image_0_221 : _GEN_220; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_222 = 10'hde == _T_5[9:0] ? image_0_222 : _GEN_221; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_223 = 10'hdf == _T_5[9:0] ? image_0_223 : _GEN_222; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_224 = 10'he0 == _T_5[9:0] ? image_0_224 : _GEN_223; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_225 = 10'he1 == _T_5[9:0] ? image_0_225 : _GEN_224; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_226 = 10'he2 == _T_5[9:0] ? image_0_226 : _GEN_225; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_227 = 10'he3 == _T_5[9:0] ? image_0_227 : _GEN_226; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_228 = 10'he4 == _T_5[9:0] ? image_0_228 : _GEN_227; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_229 = 10'he5 == _T_5[9:0] ? image_0_229 : _GEN_228; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_230 = 10'he6 == _T_5[9:0] ? image_0_230 : _GEN_229; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_231 = 10'he7 == _T_5[9:0] ? image_0_231 : _GEN_230; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_232 = 10'he8 == _T_5[9:0] ? image_0_232 : _GEN_231; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_233 = 10'he9 == _T_5[9:0] ? image_0_233 : _GEN_232; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_234 = 10'hea == _T_5[9:0] ? image_0_234 : _GEN_233; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_235 = 10'heb == _T_5[9:0] ? image_0_235 : _GEN_234; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_236 = 10'hec == _T_5[9:0] ? image_0_236 : _GEN_235; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_237 = 10'hed == _T_5[9:0] ? image_0_237 : _GEN_236; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_238 = 10'hee == _T_5[9:0] ? image_0_238 : _GEN_237; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_239 = 10'hef == _T_5[9:0] ? image_0_239 : _GEN_238; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_240 = 10'hf0 == _T_5[9:0] ? image_0_240 : _GEN_239; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_241 = 10'hf1 == _T_5[9:0] ? image_0_241 : _GEN_240; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_242 = 10'hf2 == _T_5[9:0] ? image_0_242 : _GEN_241; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_243 = 10'hf3 == _T_5[9:0] ? image_0_243 : _GEN_242; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_244 = 10'hf4 == _T_5[9:0] ? image_0_244 : _GEN_243; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_245 = 10'hf5 == _T_5[9:0] ? image_0_245 : _GEN_244; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_246 = 10'hf6 == _T_5[9:0] ? image_0_246 : _GEN_245; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_247 = 10'hf7 == _T_5[9:0] ? image_0_247 : _GEN_246; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_248 = 10'hf8 == _T_5[9:0] ? image_0_248 : _GEN_247; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_249 = 10'hf9 == _T_5[9:0] ? image_0_249 : _GEN_248; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_250 = 10'hfa == _T_5[9:0] ? image_0_250 : _GEN_249; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_251 = 10'hfb == _T_5[9:0] ? image_0_251 : _GEN_250; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_252 = 10'hfc == _T_5[9:0] ? image_0_252 : _GEN_251; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_253 = 10'hfd == _T_5[9:0] ? image_0_253 : _GEN_252; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_254 = 10'hfe == _T_5[9:0] ? image_0_254 : _GEN_253; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_255 = 10'hff == _T_5[9:0] ? image_0_255 : _GEN_254; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_256 = 10'h100 == _T_5[9:0] ? image_0_256 : _GEN_255; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_257 = 10'h101 == _T_5[9:0] ? image_0_257 : _GEN_256; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_258 = 10'h102 == _T_5[9:0] ? image_0_258 : _GEN_257; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_259 = 10'h103 == _T_5[9:0] ? image_0_259 : _GEN_258; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_260 = 10'h104 == _T_5[9:0] ? image_0_260 : _GEN_259; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_261 = 10'h105 == _T_5[9:0] ? image_0_261 : _GEN_260; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_262 = 10'h106 == _T_5[9:0] ? image_0_262 : _GEN_261; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_263 = 10'h107 == _T_5[9:0] ? image_0_263 : _GEN_262; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_264 = 10'h108 == _T_5[9:0] ? image_0_264 : _GEN_263; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_265 = 10'h109 == _T_5[9:0] ? image_0_265 : _GEN_264; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_266 = 10'h10a == _T_5[9:0] ? image_0_266 : _GEN_265; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_267 = 10'h10b == _T_5[9:0] ? image_0_267 : _GEN_266; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_268 = 10'h10c == _T_5[9:0] ? image_0_268 : _GEN_267; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_269 = 10'h10d == _T_5[9:0] ? image_0_269 : _GEN_268; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_270 = 10'h10e == _T_5[9:0] ? image_0_270 : _GEN_269; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_271 = 10'h10f == _T_5[9:0] ? image_0_271 : _GEN_270; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_272 = 10'h110 == _T_5[9:0] ? image_0_272 : _GEN_271; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_273 = 10'h111 == _T_5[9:0] ? image_0_273 : _GEN_272; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_274 = 10'h112 == _T_5[9:0] ? image_0_274 : _GEN_273; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_275 = 10'h113 == _T_5[9:0] ? image_0_275 : _GEN_274; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_276 = 10'h114 == _T_5[9:0] ? image_0_276 : _GEN_275; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_277 = 10'h115 == _T_5[9:0] ? image_0_277 : _GEN_276; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_278 = 10'h116 == _T_5[9:0] ? image_0_278 : _GEN_277; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_279 = 10'h117 == _T_5[9:0] ? image_0_279 : _GEN_278; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_280 = 10'h118 == _T_5[9:0] ? image_0_280 : _GEN_279; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_281 = 10'h119 == _T_5[9:0] ? image_0_281 : _GEN_280; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_282 = 10'h11a == _T_5[9:0] ? image_0_282 : _GEN_281; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_283 = 10'h11b == _T_5[9:0] ? image_0_283 : _GEN_282; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_284 = 10'h11c == _T_5[9:0] ? image_0_284 : _GEN_283; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_285 = 10'h11d == _T_5[9:0] ? image_0_285 : _GEN_284; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_286 = 10'h11e == _T_5[9:0] ? image_0_286 : _GEN_285; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_287 = 10'h11f == _T_5[9:0] ? image_0_287 : _GEN_286; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_288 = 10'h120 == _T_5[9:0] ? image_0_288 : _GEN_287; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_289 = 10'h121 == _T_5[9:0] ? image_0_289 : _GEN_288; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_290 = 10'h122 == _T_5[9:0] ? image_0_290 : _GEN_289; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_291 = 10'h123 == _T_5[9:0] ? image_0_291 : _GEN_290; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_292 = 10'h124 == _T_5[9:0] ? image_0_292 : _GEN_291; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_293 = 10'h125 == _T_5[9:0] ? image_0_293 : _GEN_292; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_294 = 10'h126 == _T_5[9:0] ? image_0_294 : _GEN_293; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_295 = 10'h127 == _T_5[9:0] ? image_0_295 : _GEN_294; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_296 = 10'h128 == _T_5[9:0] ? image_0_296 : _GEN_295; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_297 = 10'h129 == _T_5[9:0] ? image_0_297 : _GEN_296; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_298 = 10'h12a == _T_5[9:0] ? image_0_298 : _GEN_297; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_299 = 10'h12b == _T_5[9:0] ? image_0_299 : _GEN_298; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_300 = 10'h12c == _T_5[9:0] ? image_0_300 : _GEN_299; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_301 = 10'h12d == _T_5[9:0] ? image_0_301 : _GEN_300; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_302 = 10'h12e == _T_5[9:0] ? image_0_302 : _GEN_301; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_303 = 10'h12f == _T_5[9:0] ? image_0_303 : _GEN_302; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_304 = 10'h130 == _T_5[9:0] ? image_0_304 : _GEN_303; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_305 = 10'h131 == _T_5[9:0] ? image_0_305 : _GEN_304; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_306 = 10'h132 == _T_5[9:0] ? image_0_306 : _GEN_305; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_307 = 10'h133 == _T_5[9:0] ? image_0_307 : _GEN_306; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_308 = 10'h134 == _T_5[9:0] ? image_0_308 : _GEN_307; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_309 = 10'h135 == _T_5[9:0] ? image_0_309 : _GEN_308; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_310 = 10'h136 == _T_5[9:0] ? image_0_310 : _GEN_309; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_311 = 10'h137 == _T_5[9:0] ? image_0_311 : _GEN_310; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_312 = 10'h138 == _T_5[9:0] ? image_0_312 : _GEN_311; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_313 = 10'h139 == _T_5[9:0] ? image_0_313 : _GEN_312; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_314 = 10'h13a == _T_5[9:0] ? image_0_314 : _GEN_313; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_315 = 10'h13b == _T_5[9:0] ? image_0_315 : _GEN_314; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_316 = 10'h13c == _T_5[9:0] ? image_0_316 : _GEN_315; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_317 = 10'h13d == _T_5[9:0] ? image_0_317 : _GEN_316; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_318 = 10'h13e == _T_5[9:0] ? image_0_318 : _GEN_317; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_319 = 10'h13f == _T_5[9:0] ? image_0_319 : _GEN_318; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_320 = 10'h140 == _T_5[9:0] ? image_0_320 : _GEN_319; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_321 = 10'h141 == _T_5[9:0] ? image_0_321 : _GEN_320; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_322 = 10'h142 == _T_5[9:0] ? image_0_322 : _GEN_321; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_323 = 10'h143 == _T_5[9:0] ? image_0_323 : _GEN_322; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_324 = 10'h144 == _T_5[9:0] ? image_0_324 : _GEN_323; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_325 = 10'h145 == _T_5[9:0] ? image_0_325 : _GEN_324; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_326 = 10'h146 == _T_5[9:0] ? image_0_326 : _GEN_325; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_327 = 10'h147 == _T_5[9:0] ? image_0_327 : _GEN_326; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_328 = 10'h148 == _T_5[9:0] ? image_0_328 : _GEN_327; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_329 = 10'h149 == _T_5[9:0] ? image_0_329 : _GEN_328; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_330 = 10'h14a == _T_5[9:0] ? image_0_330 : _GEN_329; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_331 = 10'h14b == _T_5[9:0] ? image_0_331 : _GEN_330; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_332 = 10'h14c == _T_5[9:0] ? image_0_332 : _GEN_331; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_333 = 10'h14d == _T_5[9:0] ? image_0_333 : _GEN_332; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_334 = 10'h14e == _T_5[9:0] ? image_0_334 : _GEN_333; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_335 = 10'h14f == _T_5[9:0] ? image_0_335 : _GEN_334; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_336 = 10'h150 == _T_5[9:0] ? image_0_336 : _GEN_335; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_337 = 10'h151 == _T_5[9:0] ? image_0_337 : _GEN_336; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_338 = 10'h152 == _T_5[9:0] ? image_0_338 : _GEN_337; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_339 = 10'h153 == _T_5[9:0] ? image_0_339 : _GEN_338; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_340 = 10'h154 == _T_5[9:0] ? image_0_340 : _GEN_339; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_341 = 10'h155 == _T_5[9:0] ? image_0_341 : _GEN_340; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_342 = 10'h156 == _T_5[9:0] ? image_0_342 : _GEN_341; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_343 = 10'h157 == _T_5[9:0] ? image_0_343 : _GEN_342; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_344 = 10'h158 == _T_5[9:0] ? image_0_344 : _GEN_343; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_345 = 10'h159 == _T_5[9:0] ? image_0_345 : _GEN_344; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_346 = 10'h15a == _T_5[9:0] ? image_0_346 : _GEN_345; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_347 = 10'h15b == _T_5[9:0] ? image_0_347 : _GEN_346; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_348 = 10'h15c == _T_5[9:0] ? image_0_348 : _GEN_347; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_349 = 10'h15d == _T_5[9:0] ? image_0_349 : _GEN_348; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_350 = 10'h15e == _T_5[9:0] ? image_0_350 : _GEN_349; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_351 = 10'h15f == _T_5[9:0] ? image_0_351 : _GEN_350; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_352 = 10'h160 == _T_5[9:0] ? image_0_352 : _GEN_351; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_353 = 10'h161 == _T_5[9:0] ? image_0_353 : _GEN_352; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_354 = 10'h162 == _T_5[9:0] ? image_0_354 : _GEN_353; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_355 = 10'h163 == _T_5[9:0] ? image_0_355 : _GEN_354; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_356 = 10'h164 == _T_5[9:0] ? image_0_356 : _GEN_355; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_357 = 10'h165 == _T_5[9:0] ? image_0_357 : _GEN_356; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_358 = 10'h166 == _T_5[9:0] ? image_0_358 : _GEN_357; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_359 = 10'h167 == _T_5[9:0] ? image_0_359 : _GEN_358; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_360 = 10'h168 == _T_5[9:0] ? image_0_360 : _GEN_359; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_361 = 10'h169 == _T_5[9:0] ? image_0_361 : _GEN_360; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_362 = 10'h16a == _T_5[9:0] ? image_0_362 : _GEN_361; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_363 = 10'h16b == _T_5[9:0] ? image_0_363 : _GEN_362; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_364 = 10'h16c == _T_5[9:0] ? image_0_364 : _GEN_363; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_365 = 10'h16d == _T_5[9:0] ? image_0_365 : _GEN_364; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_366 = 10'h16e == _T_5[9:0] ? image_0_366 : _GEN_365; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_367 = 10'h16f == _T_5[9:0] ? image_0_367 : _GEN_366; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_368 = 10'h170 == _T_5[9:0] ? image_0_368 : _GEN_367; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_369 = 10'h171 == _T_5[9:0] ? image_0_369 : _GEN_368; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_370 = 10'h172 == _T_5[9:0] ? image_0_370 : _GEN_369; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_371 = 10'h173 == _T_5[9:0] ? image_0_371 : _GEN_370; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_372 = 10'h174 == _T_5[9:0] ? image_0_372 : _GEN_371; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_373 = 10'h175 == _T_5[9:0] ? image_0_373 : _GEN_372; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_374 = 10'h176 == _T_5[9:0] ? image_0_374 : _GEN_373; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_375 = 10'h177 == _T_5[9:0] ? image_0_375 : _GEN_374; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_376 = 10'h178 == _T_5[9:0] ? image_0_376 : _GEN_375; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_377 = 10'h179 == _T_5[9:0] ? image_0_377 : _GEN_376; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_378 = 10'h17a == _T_5[9:0] ? image_0_378 : _GEN_377; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_379 = 10'h17b == _T_5[9:0] ? image_0_379 : _GEN_378; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_380 = 10'h17c == _T_5[9:0] ? image_0_380 : _GEN_379; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_381 = 10'h17d == _T_5[9:0] ? image_0_381 : _GEN_380; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_382 = 10'h17e == _T_5[9:0] ? image_0_382 : _GEN_381; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_383 = 10'h17f == _T_5[9:0] ? image_0_383 : _GEN_382; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_384 = 10'h180 == _T_5[9:0] ? image_0_384 : _GEN_383; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_385 = 10'h181 == _T_5[9:0] ? image_0_385 : _GEN_384; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_386 = 10'h182 == _T_5[9:0] ? image_0_386 : _GEN_385; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_387 = 10'h183 == _T_5[9:0] ? image_0_387 : _GEN_386; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_388 = 10'h184 == _T_5[9:0] ? image_0_388 : _GEN_387; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_389 = 10'h185 == _T_5[9:0] ? image_0_389 : _GEN_388; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_390 = 10'h186 == _T_5[9:0] ? image_0_390 : _GEN_389; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_391 = 10'h187 == _T_5[9:0] ? image_0_391 : _GEN_390; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_392 = 10'h188 == _T_5[9:0] ? image_0_392 : _GEN_391; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_393 = 10'h189 == _T_5[9:0] ? image_0_393 : _GEN_392; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_394 = 10'h18a == _T_5[9:0] ? image_0_394 : _GEN_393; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_395 = 10'h18b == _T_5[9:0] ? image_0_395 : _GEN_394; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_396 = 10'h18c == _T_5[9:0] ? image_0_396 : _GEN_395; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_397 = 10'h18d == _T_5[9:0] ? image_0_397 : _GEN_396; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_398 = 10'h18e == _T_5[9:0] ? image_0_398 : _GEN_397; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_399 = 10'h18f == _T_5[9:0] ? image_0_399 : _GEN_398; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_400 = 10'h190 == _T_5[9:0] ? image_0_400 : _GEN_399; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_401 = 10'h191 == _T_5[9:0] ? image_0_401 : _GEN_400; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_402 = 10'h192 == _T_5[9:0] ? image_0_402 : _GEN_401; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_403 = 10'h193 == _T_5[9:0] ? image_0_403 : _GEN_402; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_404 = 10'h194 == _T_5[9:0] ? image_0_404 : _GEN_403; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_405 = 10'h195 == _T_5[9:0] ? image_0_405 : _GEN_404; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_406 = 10'h196 == _T_5[9:0] ? image_0_406 : _GEN_405; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_407 = 10'h197 == _T_5[9:0] ? image_0_407 : _GEN_406; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_408 = 10'h198 == _T_5[9:0] ? image_0_408 : _GEN_407; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_409 = 10'h199 == _T_5[9:0] ? image_0_409 : _GEN_408; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_410 = 10'h19a == _T_5[9:0] ? image_0_410 : _GEN_409; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_411 = 10'h19b == _T_5[9:0] ? image_0_411 : _GEN_410; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_412 = 10'h19c == _T_5[9:0] ? image_0_412 : _GEN_411; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_413 = 10'h19d == _T_5[9:0] ? image_0_413 : _GEN_412; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_414 = 10'h19e == _T_5[9:0] ? image_0_414 : _GEN_413; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_415 = 10'h19f == _T_5[9:0] ? image_0_415 : _GEN_414; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_416 = 10'h1a0 == _T_5[9:0] ? image_0_416 : _GEN_415; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_417 = 10'h1a1 == _T_5[9:0] ? image_0_417 : _GEN_416; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_418 = 10'h1a2 == _T_5[9:0] ? image_0_418 : _GEN_417; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_419 = 10'h1a3 == _T_5[9:0] ? image_0_419 : _GEN_418; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_420 = 10'h1a4 == _T_5[9:0] ? image_0_420 : _GEN_419; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_421 = 10'h1a5 == _T_5[9:0] ? image_0_421 : _GEN_420; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_422 = 10'h1a6 == _T_5[9:0] ? image_0_422 : _GEN_421; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_423 = 10'h1a7 == _T_5[9:0] ? image_0_423 : _GEN_422; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_424 = 10'h1a8 == _T_5[9:0] ? image_0_424 : _GEN_423; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_425 = 10'h1a9 == _T_5[9:0] ? image_0_425 : _GEN_424; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_426 = 10'h1aa == _T_5[9:0] ? image_0_426 : _GEN_425; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_427 = 10'h1ab == _T_5[9:0] ? image_0_427 : _GEN_426; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_428 = 10'h1ac == _T_5[9:0] ? image_0_428 : _GEN_427; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_429 = 10'h1ad == _T_5[9:0] ? image_0_429 : _GEN_428; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_430 = 10'h1ae == _T_5[9:0] ? image_0_430 : _GEN_429; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_431 = 10'h1af == _T_5[9:0] ? image_0_431 : _GEN_430; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_432 = 10'h1b0 == _T_5[9:0] ? image_0_432 : _GEN_431; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_433 = 10'h1b1 == _T_5[9:0] ? image_0_433 : _GEN_432; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_434 = 10'h1b2 == _T_5[9:0] ? image_0_434 : _GEN_433; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_435 = 10'h1b3 == _T_5[9:0] ? image_0_435 : _GEN_434; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_436 = 10'h1b4 == _T_5[9:0] ? image_0_436 : _GEN_435; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_437 = 10'h1b5 == _T_5[9:0] ? image_0_437 : _GEN_436; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_438 = 10'h1b6 == _T_5[9:0] ? image_0_438 : _GEN_437; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_439 = 10'h1b7 == _T_5[9:0] ? image_0_439 : _GEN_438; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_440 = 10'h1b8 == _T_5[9:0] ? image_0_440 : _GEN_439; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_441 = 10'h1b9 == _T_5[9:0] ? image_0_441 : _GEN_440; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_442 = 10'h1ba == _T_5[9:0] ? image_0_442 : _GEN_441; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_443 = 10'h1bb == _T_5[9:0] ? image_0_443 : _GEN_442; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_444 = 10'h1bc == _T_5[9:0] ? image_0_444 : _GEN_443; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_445 = 10'h1bd == _T_5[9:0] ? image_0_445 : _GEN_444; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_446 = 10'h1be == _T_5[9:0] ? image_0_446 : _GEN_445; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_447 = 10'h1bf == _T_5[9:0] ? image_0_447 : _GEN_446; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_448 = 10'h1c0 == _T_5[9:0] ? image_0_448 : _GEN_447; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_449 = 10'h1c1 == _T_5[9:0] ? image_0_449 : _GEN_448; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_450 = 10'h1c2 == _T_5[9:0] ? image_0_450 : _GEN_449; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_451 = 10'h1c3 == _T_5[9:0] ? image_0_451 : _GEN_450; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_452 = 10'h1c4 == _T_5[9:0] ? image_0_452 : _GEN_451; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_453 = 10'h1c5 == _T_5[9:0] ? image_0_453 : _GEN_452; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_454 = 10'h1c6 == _T_5[9:0] ? image_0_454 : _GEN_453; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_455 = 10'h1c7 == _T_5[9:0] ? image_0_455 : _GEN_454; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_456 = 10'h1c8 == _T_5[9:0] ? image_0_456 : _GEN_455; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_457 = 10'h1c9 == _T_5[9:0] ? image_0_457 : _GEN_456; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_458 = 10'h1ca == _T_5[9:0] ? image_0_458 : _GEN_457; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_459 = 10'h1cb == _T_5[9:0] ? image_0_459 : _GEN_458; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_460 = 10'h1cc == _T_5[9:0] ? image_0_460 : _GEN_459; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_461 = 10'h1cd == _T_5[9:0] ? image_0_461 : _GEN_460; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_462 = 10'h1ce == _T_5[9:0] ? image_0_462 : _GEN_461; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_463 = 10'h1cf == _T_5[9:0] ? image_0_463 : _GEN_462; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_464 = 10'h1d0 == _T_5[9:0] ? image_0_464 : _GEN_463; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_465 = 10'h1d1 == _T_5[9:0] ? image_0_465 : _GEN_464; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_466 = 10'h1d2 == _T_5[9:0] ? image_0_466 : _GEN_465; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_467 = 10'h1d3 == _T_5[9:0] ? image_0_467 : _GEN_466; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_468 = 10'h1d4 == _T_5[9:0] ? image_0_468 : _GEN_467; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_469 = 10'h1d5 == _T_5[9:0] ? image_0_469 : _GEN_468; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_470 = 10'h1d6 == _T_5[9:0] ? image_0_470 : _GEN_469; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_471 = 10'h1d7 == _T_5[9:0] ? image_0_471 : _GEN_470; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_472 = 10'h1d8 == _T_5[9:0] ? image_0_472 : _GEN_471; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_473 = 10'h1d9 == _T_5[9:0] ? image_0_473 : _GEN_472; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_474 = 10'h1da == _T_5[9:0] ? image_0_474 : _GEN_473; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_475 = 10'h1db == _T_5[9:0] ? image_0_475 : _GEN_474; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_476 = 10'h1dc == _T_5[9:0] ? image_0_476 : _GEN_475; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_477 = 10'h1dd == _T_5[9:0] ? image_0_477 : _GEN_476; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_478 = 10'h1de == _T_5[9:0] ? image_0_478 : _GEN_477; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_479 = 10'h1df == _T_5[9:0] ? image_0_479 : _GEN_478; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_480 = 10'h1e0 == _T_5[9:0] ? image_0_480 : _GEN_479; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_481 = 10'h1e1 == _T_5[9:0] ? image_0_481 : _GEN_480; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_482 = 10'h1e2 == _T_5[9:0] ? image_0_482 : _GEN_481; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_483 = 10'h1e3 == _T_5[9:0] ? image_0_483 : _GEN_482; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_484 = 10'h1e4 == _T_5[9:0] ? image_0_484 : _GEN_483; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_485 = 10'h1e5 == _T_5[9:0] ? image_0_485 : _GEN_484; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_486 = 10'h1e6 == _T_5[9:0] ? image_0_486 : _GEN_485; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_487 = 10'h1e7 == _T_5[9:0] ? image_0_487 : _GEN_486; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_488 = 10'h1e8 == _T_5[9:0] ? image_0_488 : _GEN_487; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_489 = 10'h1e9 == _T_5[9:0] ? image_0_489 : _GEN_488; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_490 = 10'h1ea == _T_5[9:0] ? image_0_490 : _GEN_489; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_491 = 10'h1eb == _T_5[9:0] ? image_0_491 : _GEN_490; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_492 = 10'h1ec == _T_5[9:0] ? image_0_492 : _GEN_491; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_493 = 10'h1ed == _T_5[9:0] ? image_0_493 : _GEN_492; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_494 = 10'h1ee == _T_5[9:0] ? image_0_494 : _GEN_493; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_495 = 10'h1ef == _T_5[9:0] ? image_0_495 : _GEN_494; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_496 = 10'h1f0 == _T_5[9:0] ? image_0_496 : _GEN_495; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_497 = 10'h1f1 == _T_5[9:0] ? image_0_497 : _GEN_496; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_498 = 10'h1f2 == _T_5[9:0] ? image_0_498 : _GEN_497; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_499 = 10'h1f3 == _T_5[9:0] ? image_0_499 : _GEN_498; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_500 = 10'h1f4 == _T_5[9:0] ? image_0_500 : _GEN_499; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_501 = 10'h1f5 == _T_5[9:0] ? image_0_501 : _GEN_500; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_502 = 10'h1f6 == _T_5[9:0] ? image_0_502 : _GEN_501; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_503 = 10'h1f7 == _T_5[9:0] ? image_0_503 : _GEN_502; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_504 = 10'h1f8 == _T_5[9:0] ? image_0_504 : _GEN_503; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_505 = 10'h1f9 == _T_5[9:0] ? image_0_505 : _GEN_504; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_506 = 10'h1fa == _T_5[9:0] ? image_0_506 : _GEN_505; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_507 = 10'h1fb == _T_5[9:0] ? image_0_507 : _GEN_506; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_508 = 10'h1fc == _T_5[9:0] ? image_0_508 : _GEN_507; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_509 = 10'h1fd == _T_5[9:0] ? image_0_509 : _GEN_508; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_510 = 10'h1fe == _T_5[9:0] ? image_0_510 : _GEN_509; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_511 = 10'h1ff == _T_5[9:0] ? image_0_511 : _GEN_510; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_512 = 10'h200 == _T_5[9:0] ? image_0_512 : _GEN_511; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_513 = 10'h201 == _T_5[9:0] ? image_0_513 : _GEN_512; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_514 = 10'h202 == _T_5[9:0] ? image_0_514 : _GEN_513; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_515 = 10'h203 == _T_5[9:0] ? image_0_515 : _GEN_514; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_516 = 10'h204 == _T_5[9:0] ? image_0_516 : _GEN_515; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_517 = 10'h205 == _T_5[9:0] ? image_0_517 : _GEN_516; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_518 = 10'h206 == _T_5[9:0] ? image_0_518 : _GEN_517; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_519 = 10'h207 == _T_5[9:0] ? image_0_519 : _GEN_518; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_520 = 10'h208 == _T_5[9:0] ? image_0_520 : _GEN_519; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_521 = 10'h209 == _T_5[9:0] ? image_0_521 : _GEN_520; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_522 = 10'h20a == _T_5[9:0] ? image_0_522 : _GEN_521; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_523 = 10'h20b == _T_5[9:0] ? image_0_523 : _GEN_522; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_524 = 10'h20c == _T_5[9:0] ? image_0_524 : _GEN_523; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_525 = 10'h20d == _T_5[9:0] ? image_0_525 : _GEN_524; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_526 = 10'h20e == _T_5[9:0] ? image_0_526 : _GEN_525; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_527 = 10'h20f == _T_5[9:0] ? image_0_527 : _GEN_526; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_528 = 10'h210 == _T_5[9:0] ? image_0_528 : _GEN_527; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_529 = 10'h211 == _T_5[9:0] ? image_0_529 : _GEN_528; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_530 = 10'h212 == _T_5[9:0] ? image_0_530 : _GEN_529; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_531 = 10'h213 == _T_5[9:0] ? image_0_531 : _GEN_530; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_532 = 10'h214 == _T_5[9:0] ? image_0_532 : _GEN_531; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_533 = 10'h215 == _T_5[9:0] ? image_0_533 : _GEN_532; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_534 = 10'h216 == _T_5[9:0] ? image_0_534 : _GEN_533; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_535 = 10'h217 == _T_5[9:0] ? image_0_535 : _GEN_534; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_536 = 10'h218 == _T_5[9:0] ? image_0_536 : _GEN_535; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_537 = 10'h219 == _T_5[9:0] ? image_0_537 : _GEN_536; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_538 = 10'h21a == _T_5[9:0] ? image_0_538 : _GEN_537; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_539 = 10'h21b == _T_5[9:0] ? image_0_539 : _GEN_538; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_540 = 10'h21c == _T_5[9:0] ? image_0_540 : _GEN_539; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_541 = 10'h21d == _T_5[9:0] ? image_0_541 : _GEN_540; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_542 = 10'h21e == _T_5[9:0] ? image_0_542 : _GEN_541; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_543 = 10'h21f == _T_5[9:0] ? image_0_543 : _GEN_542; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_544 = 10'h220 == _T_5[9:0] ? image_0_544 : _GEN_543; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_545 = 10'h221 == _T_5[9:0] ? image_0_545 : _GEN_544; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_546 = 10'h222 == _T_5[9:0] ? image_0_546 : _GEN_545; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_547 = 10'h223 == _T_5[9:0] ? image_0_547 : _GEN_546; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_548 = 10'h224 == _T_5[9:0] ? image_0_548 : _GEN_547; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_549 = 10'h225 == _T_5[9:0] ? image_0_549 : _GEN_548; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_550 = 10'h226 == _T_5[9:0] ? image_0_550 : _GEN_549; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_551 = 10'h227 == _T_5[9:0] ? image_0_551 : _GEN_550; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_552 = 10'h228 == _T_5[9:0] ? image_0_552 : _GEN_551; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_553 = 10'h229 == _T_5[9:0] ? image_0_553 : _GEN_552; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_554 = 10'h22a == _T_5[9:0] ? image_0_554 : _GEN_553; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_555 = 10'h22b == _T_5[9:0] ? image_0_555 : _GEN_554; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_556 = 10'h22c == _T_5[9:0] ? image_0_556 : _GEN_555; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_557 = 10'h22d == _T_5[9:0] ? image_0_557 : _GEN_556; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_558 = 10'h22e == _T_5[9:0] ? image_0_558 : _GEN_557; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_559 = 10'h22f == _T_5[9:0] ? image_0_559 : _GEN_558; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_560 = 10'h230 == _T_5[9:0] ? image_0_560 : _GEN_559; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_561 = 10'h231 == _T_5[9:0] ? image_0_561 : _GEN_560; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_562 = 10'h232 == _T_5[9:0] ? image_0_562 : _GEN_561; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_563 = 10'h233 == _T_5[9:0] ? image_0_563 : _GEN_562; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_564 = 10'h234 == _T_5[9:0] ? image_0_564 : _GEN_563; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_565 = 10'h235 == _T_5[9:0] ? image_0_565 : _GEN_564; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_566 = 10'h236 == _T_5[9:0] ? image_0_566 : _GEN_565; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_567 = 10'h237 == _T_5[9:0] ? image_0_567 : _GEN_566; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_568 = 10'h238 == _T_5[9:0] ? image_0_568 : _GEN_567; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_569 = 10'h239 == _T_5[9:0] ? image_0_569 : _GEN_568; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_570 = 10'h23a == _T_5[9:0] ? image_0_570 : _GEN_569; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_571 = 10'h23b == _T_5[9:0] ? image_0_571 : _GEN_570; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_572 = 10'h23c == _T_5[9:0] ? image_0_572 : _GEN_571; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_573 = 10'h23d == _T_5[9:0] ? image_0_573 : _GEN_572; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_574 = 10'h23e == _T_5[9:0] ? image_0_574 : _GEN_573; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_577 = 10'h1 == _T_5[9:0] ? image_1_1 : image_1_0; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_578 = 10'h2 == _T_5[9:0] ? image_1_2 : _GEN_577; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_579 = 10'h3 == _T_5[9:0] ? image_1_3 : _GEN_578; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_580 = 10'h4 == _T_5[9:0] ? image_1_4 : _GEN_579; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_581 = 10'h5 == _T_5[9:0] ? image_1_5 : _GEN_580; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_582 = 10'h6 == _T_5[9:0] ? image_1_6 : _GEN_581; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_583 = 10'h7 == _T_5[9:0] ? image_1_7 : _GEN_582; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_584 = 10'h8 == _T_5[9:0] ? image_1_8 : _GEN_583; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_585 = 10'h9 == _T_5[9:0] ? image_1_9 : _GEN_584; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_586 = 10'ha == _T_5[9:0] ? image_1_10 : _GEN_585; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_587 = 10'hb == _T_5[9:0] ? image_1_11 : _GEN_586; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_588 = 10'hc == _T_5[9:0] ? image_1_12 : _GEN_587; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_589 = 10'hd == _T_5[9:0] ? image_1_13 : _GEN_588; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_590 = 10'he == _T_5[9:0] ? image_1_14 : _GEN_589; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_591 = 10'hf == _T_5[9:0] ? image_1_15 : _GEN_590; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_592 = 10'h10 == _T_5[9:0] ? image_1_16 : _GEN_591; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_593 = 10'h11 == _T_5[9:0] ? image_1_17 : _GEN_592; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_594 = 10'h12 == _T_5[9:0] ? image_1_18 : _GEN_593; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_595 = 10'h13 == _T_5[9:0] ? image_1_19 : _GEN_594; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_596 = 10'h14 == _T_5[9:0] ? image_1_20 : _GEN_595; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_597 = 10'h15 == _T_5[9:0] ? image_1_21 : _GEN_596; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_598 = 10'h16 == _T_5[9:0] ? image_1_22 : _GEN_597; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_599 = 10'h17 == _T_5[9:0] ? image_1_23 : _GEN_598; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_600 = 10'h18 == _T_5[9:0] ? image_1_24 : _GEN_599; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_601 = 10'h19 == _T_5[9:0] ? image_1_25 : _GEN_600; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_602 = 10'h1a == _T_5[9:0] ? image_1_26 : _GEN_601; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_603 = 10'h1b == _T_5[9:0] ? image_1_27 : _GEN_602; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_604 = 10'h1c == _T_5[9:0] ? image_1_28 : _GEN_603; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_605 = 10'h1d == _T_5[9:0] ? image_1_29 : _GEN_604; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_606 = 10'h1e == _T_5[9:0] ? image_1_30 : _GEN_605; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_607 = 10'h1f == _T_5[9:0] ? image_1_31 : _GEN_606; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_608 = 10'h20 == _T_5[9:0] ? image_1_32 : _GEN_607; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_609 = 10'h21 == _T_5[9:0] ? image_1_33 : _GEN_608; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_610 = 10'h22 == _T_5[9:0] ? image_1_34 : _GEN_609; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_611 = 10'h23 == _T_5[9:0] ? image_1_35 : _GEN_610; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_612 = 10'h24 == _T_5[9:0] ? image_1_36 : _GEN_611; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_613 = 10'h25 == _T_5[9:0] ? image_1_37 : _GEN_612; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_614 = 10'h26 == _T_5[9:0] ? image_1_38 : _GEN_613; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_615 = 10'h27 == _T_5[9:0] ? image_1_39 : _GEN_614; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_616 = 10'h28 == _T_5[9:0] ? image_1_40 : _GEN_615; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_617 = 10'h29 == _T_5[9:0] ? image_1_41 : _GEN_616; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_618 = 10'h2a == _T_5[9:0] ? image_1_42 : _GEN_617; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_619 = 10'h2b == _T_5[9:0] ? image_1_43 : _GEN_618; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_620 = 10'h2c == _T_5[9:0] ? image_1_44 : _GEN_619; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_621 = 10'h2d == _T_5[9:0] ? image_1_45 : _GEN_620; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_622 = 10'h2e == _T_5[9:0] ? image_1_46 : _GEN_621; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_623 = 10'h2f == _T_5[9:0] ? image_1_47 : _GEN_622; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_624 = 10'h30 == _T_5[9:0] ? image_1_48 : _GEN_623; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_625 = 10'h31 == _T_5[9:0] ? image_1_49 : _GEN_624; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_626 = 10'h32 == _T_5[9:0] ? image_1_50 : _GEN_625; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_627 = 10'h33 == _T_5[9:0] ? image_1_51 : _GEN_626; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_628 = 10'h34 == _T_5[9:0] ? image_1_52 : _GEN_627; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_629 = 10'h35 == _T_5[9:0] ? image_1_53 : _GEN_628; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_630 = 10'h36 == _T_5[9:0] ? image_1_54 : _GEN_629; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_631 = 10'h37 == _T_5[9:0] ? image_1_55 : _GEN_630; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_632 = 10'h38 == _T_5[9:0] ? image_1_56 : _GEN_631; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_633 = 10'h39 == _T_5[9:0] ? image_1_57 : _GEN_632; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_634 = 10'h3a == _T_5[9:0] ? image_1_58 : _GEN_633; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_635 = 10'h3b == _T_5[9:0] ? image_1_59 : _GEN_634; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_636 = 10'h3c == _T_5[9:0] ? image_1_60 : _GEN_635; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_637 = 10'h3d == _T_5[9:0] ? image_1_61 : _GEN_636; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_638 = 10'h3e == _T_5[9:0] ? image_1_62 : _GEN_637; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_639 = 10'h3f == _T_5[9:0] ? image_1_63 : _GEN_638; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_640 = 10'h40 == _T_5[9:0] ? image_1_64 : _GEN_639; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_641 = 10'h41 == _T_5[9:0] ? image_1_65 : _GEN_640; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_642 = 10'h42 == _T_5[9:0] ? image_1_66 : _GEN_641; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_643 = 10'h43 == _T_5[9:0] ? image_1_67 : _GEN_642; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_644 = 10'h44 == _T_5[9:0] ? image_1_68 : _GEN_643; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_645 = 10'h45 == _T_5[9:0] ? image_1_69 : _GEN_644; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_646 = 10'h46 == _T_5[9:0] ? image_1_70 : _GEN_645; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_647 = 10'h47 == _T_5[9:0] ? image_1_71 : _GEN_646; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_648 = 10'h48 == _T_5[9:0] ? image_1_72 : _GEN_647; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_649 = 10'h49 == _T_5[9:0] ? image_1_73 : _GEN_648; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_650 = 10'h4a == _T_5[9:0] ? image_1_74 : _GEN_649; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_651 = 10'h4b == _T_5[9:0] ? image_1_75 : _GEN_650; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_652 = 10'h4c == _T_5[9:0] ? image_1_76 : _GEN_651; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_653 = 10'h4d == _T_5[9:0] ? image_1_77 : _GEN_652; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_654 = 10'h4e == _T_5[9:0] ? image_1_78 : _GEN_653; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_655 = 10'h4f == _T_5[9:0] ? image_1_79 : _GEN_654; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_656 = 10'h50 == _T_5[9:0] ? image_1_80 : _GEN_655; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_657 = 10'h51 == _T_5[9:0] ? image_1_81 : _GEN_656; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_658 = 10'h52 == _T_5[9:0] ? image_1_82 : _GEN_657; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_659 = 10'h53 == _T_5[9:0] ? image_1_83 : _GEN_658; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_660 = 10'h54 == _T_5[9:0] ? image_1_84 : _GEN_659; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_661 = 10'h55 == _T_5[9:0] ? image_1_85 : _GEN_660; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_662 = 10'h56 == _T_5[9:0] ? image_1_86 : _GEN_661; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_663 = 10'h57 == _T_5[9:0] ? image_1_87 : _GEN_662; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_664 = 10'h58 == _T_5[9:0] ? image_1_88 : _GEN_663; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_665 = 10'h59 == _T_5[9:0] ? image_1_89 : _GEN_664; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_666 = 10'h5a == _T_5[9:0] ? image_1_90 : _GEN_665; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_667 = 10'h5b == _T_5[9:0] ? image_1_91 : _GEN_666; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_668 = 10'h5c == _T_5[9:0] ? image_1_92 : _GEN_667; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_669 = 10'h5d == _T_5[9:0] ? image_1_93 : _GEN_668; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_670 = 10'h5e == _T_5[9:0] ? image_1_94 : _GEN_669; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_671 = 10'h5f == _T_5[9:0] ? image_1_95 : _GEN_670; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_672 = 10'h60 == _T_5[9:0] ? image_1_96 : _GEN_671; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_673 = 10'h61 == _T_5[9:0] ? image_1_97 : _GEN_672; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_674 = 10'h62 == _T_5[9:0] ? image_1_98 : _GEN_673; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_675 = 10'h63 == _T_5[9:0] ? image_1_99 : _GEN_674; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_676 = 10'h64 == _T_5[9:0] ? image_1_100 : _GEN_675; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_677 = 10'h65 == _T_5[9:0] ? image_1_101 : _GEN_676; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_678 = 10'h66 == _T_5[9:0] ? image_1_102 : _GEN_677; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_679 = 10'h67 == _T_5[9:0] ? image_1_103 : _GEN_678; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_680 = 10'h68 == _T_5[9:0] ? image_1_104 : _GEN_679; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_681 = 10'h69 == _T_5[9:0] ? image_1_105 : _GEN_680; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_682 = 10'h6a == _T_5[9:0] ? image_1_106 : _GEN_681; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_683 = 10'h6b == _T_5[9:0] ? image_1_107 : _GEN_682; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_684 = 10'h6c == _T_5[9:0] ? image_1_108 : _GEN_683; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_685 = 10'h6d == _T_5[9:0] ? image_1_109 : _GEN_684; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_686 = 10'h6e == _T_5[9:0] ? image_1_110 : _GEN_685; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_687 = 10'h6f == _T_5[9:0] ? image_1_111 : _GEN_686; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_688 = 10'h70 == _T_5[9:0] ? image_1_112 : _GEN_687; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_689 = 10'h71 == _T_5[9:0] ? image_1_113 : _GEN_688; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_690 = 10'h72 == _T_5[9:0] ? image_1_114 : _GEN_689; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_691 = 10'h73 == _T_5[9:0] ? image_1_115 : _GEN_690; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_692 = 10'h74 == _T_5[9:0] ? image_1_116 : _GEN_691; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_693 = 10'h75 == _T_5[9:0] ? image_1_117 : _GEN_692; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_694 = 10'h76 == _T_5[9:0] ? image_1_118 : _GEN_693; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_695 = 10'h77 == _T_5[9:0] ? image_1_119 : _GEN_694; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_696 = 10'h78 == _T_5[9:0] ? image_1_120 : _GEN_695; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_697 = 10'h79 == _T_5[9:0] ? image_1_121 : _GEN_696; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_698 = 10'h7a == _T_5[9:0] ? image_1_122 : _GEN_697; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_699 = 10'h7b == _T_5[9:0] ? image_1_123 : _GEN_698; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_700 = 10'h7c == _T_5[9:0] ? image_1_124 : _GEN_699; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_701 = 10'h7d == _T_5[9:0] ? image_1_125 : _GEN_700; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_702 = 10'h7e == _T_5[9:0] ? image_1_126 : _GEN_701; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_703 = 10'h7f == _T_5[9:0] ? image_1_127 : _GEN_702; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_704 = 10'h80 == _T_5[9:0] ? image_1_128 : _GEN_703; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_705 = 10'h81 == _T_5[9:0] ? image_1_129 : _GEN_704; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_706 = 10'h82 == _T_5[9:0] ? image_1_130 : _GEN_705; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_707 = 10'h83 == _T_5[9:0] ? image_1_131 : _GEN_706; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_708 = 10'h84 == _T_5[9:0] ? image_1_132 : _GEN_707; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_709 = 10'h85 == _T_5[9:0] ? image_1_133 : _GEN_708; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_710 = 10'h86 == _T_5[9:0] ? image_1_134 : _GEN_709; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_711 = 10'h87 == _T_5[9:0] ? image_1_135 : _GEN_710; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_712 = 10'h88 == _T_5[9:0] ? image_1_136 : _GEN_711; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_713 = 10'h89 == _T_5[9:0] ? image_1_137 : _GEN_712; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_714 = 10'h8a == _T_5[9:0] ? image_1_138 : _GEN_713; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_715 = 10'h8b == _T_5[9:0] ? image_1_139 : _GEN_714; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_716 = 10'h8c == _T_5[9:0] ? image_1_140 : _GEN_715; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_717 = 10'h8d == _T_5[9:0] ? image_1_141 : _GEN_716; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_718 = 10'h8e == _T_5[9:0] ? image_1_142 : _GEN_717; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_719 = 10'h8f == _T_5[9:0] ? image_1_143 : _GEN_718; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_720 = 10'h90 == _T_5[9:0] ? image_1_144 : _GEN_719; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_721 = 10'h91 == _T_5[9:0] ? image_1_145 : _GEN_720; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_722 = 10'h92 == _T_5[9:0] ? image_1_146 : _GEN_721; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_723 = 10'h93 == _T_5[9:0] ? image_1_147 : _GEN_722; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_724 = 10'h94 == _T_5[9:0] ? image_1_148 : _GEN_723; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_725 = 10'h95 == _T_5[9:0] ? image_1_149 : _GEN_724; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_726 = 10'h96 == _T_5[9:0] ? image_1_150 : _GEN_725; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_727 = 10'h97 == _T_5[9:0] ? image_1_151 : _GEN_726; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_728 = 10'h98 == _T_5[9:0] ? image_1_152 : _GEN_727; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_729 = 10'h99 == _T_5[9:0] ? image_1_153 : _GEN_728; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_730 = 10'h9a == _T_5[9:0] ? image_1_154 : _GEN_729; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_731 = 10'h9b == _T_5[9:0] ? image_1_155 : _GEN_730; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_732 = 10'h9c == _T_5[9:0] ? image_1_156 : _GEN_731; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_733 = 10'h9d == _T_5[9:0] ? image_1_157 : _GEN_732; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_734 = 10'h9e == _T_5[9:0] ? image_1_158 : _GEN_733; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_735 = 10'h9f == _T_5[9:0] ? image_1_159 : _GEN_734; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_736 = 10'ha0 == _T_5[9:0] ? image_1_160 : _GEN_735; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_737 = 10'ha1 == _T_5[9:0] ? image_1_161 : _GEN_736; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_738 = 10'ha2 == _T_5[9:0] ? image_1_162 : _GEN_737; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_739 = 10'ha3 == _T_5[9:0] ? image_1_163 : _GEN_738; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_740 = 10'ha4 == _T_5[9:0] ? image_1_164 : _GEN_739; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_741 = 10'ha5 == _T_5[9:0] ? image_1_165 : _GEN_740; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_742 = 10'ha6 == _T_5[9:0] ? image_1_166 : _GEN_741; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_743 = 10'ha7 == _T_5[9:0] ? image_1_167 : _GEN_742; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_744 = 10'ha8 == _T_5[9:0] ? image_1_168 : _GEN_743; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_745 = 10'ha9 == _T_5[9:0] ? image_1_169 : _GEN_744; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_746 = 10'haa == _T_5[9:0] ? image_1_170 : _GEN_745; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_747 = 10'hab == _T_5[9:0] ? image_1_171 : _GEN_746; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_748 = 10'hac == _T_5[9:0] ? image_1_172 : _GEN_747; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_749 = 10'had == _T_5[9:0] ? image_1_173 : _GEN_748; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_750 = 10'hae == _T_5[9:0] ? image_1_174 : _GEN_749; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_751 = 10'haf == _T_5[9:0] ? image_1_175 : _GEN_750; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_752 = 10'hb0 == _T_5[9:0] ? image_1_176 : _GEN_751; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_753 = 10'hb1 == _T_5[9:0] ? image_1_177 : _GEN_752; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_754 = 10'hb2 == _T_5[9:0] ? image_1_178 : _GEN_753; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_755 = 10'hb3 == _T_5[9:0] ? image_1_179 : _GEN_754; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_756 = 10'hb4 == _T_5[9:0] ? image_1_180 : _GEN_755; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_757 = 10'hb5 == _T_5[9:0] ? image_1_181 : _GEN_756; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_758 = 10'hb6 == _T_5[9:0] ? image_1_182 : _GEN_757; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_759 = 10'hb7 == _T_5[9:0] ? image_1_183 : _GEN_758; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_760 = 10'hb8 == _T_5[9:0] ? image_1_184 : _GEN_759; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_761 = 10'hb9 == _T_5[9:0] ? image_1_185 : _GEN_760; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_762 = 10'hba == _T_5[9:0] ? image_1_186 : _GEN_761; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_763 = 10'hbb == _T_5[9:0] ? image_1_187 : _GEN_762; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_764 = 10'hbc == _T_5[9:0] ? image_1_188 : _GEN_763; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_765 = 10'hbd == _T_5[9:0] ? image_1_189 : _GEN_764; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_766 = 10'hbe == _T_5[9:0] ? image_1_190 : _GEN_765; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_767 = 10'hbf == _T_5[9:0] ? image_1_191 : _GEN_766; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_768 = 10'hc0 == _T_5[9:0] ? image_1_192 : _GEN_767; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_769 = 10'hc1 == _T_5[9:0] ? image_1_193 : _GEN_768; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_770 = 10'hc2 == _T_5[9:0] ? image_1_194 : _GEN_769; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_771 = 10'hc3 == _T_5[9:0] ? image_1_195 : _GEN_770; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_772 = 10'hc4 == _T_5[9:0] ? image_1_196 : _GEN_771; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_773 = 10'hc5 == _T_5[9:0] ? image_1_197 : _GEN_772; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_774 = 10'hc6 == _T_5[9:0] ? image_1_198 : _GEN_773; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_775 = 10'hc7 == _T_5[9:0] ? image_1_199 : _GEN_774; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_776 = 10'hc8 == _T_5[9:0] ? image_1_200 : _GEN_775; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_777 = 10'hc9 == _T_5[9:0] ? image_1_201 : _GEN_776; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_778 = 10'hca == _T_5[9:0] ? image_1_202 : _GEN_777; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_779 = 10'hcb == _T_5[9:0] ? image_1_203 : _GEN_778; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_780 = 10'hcc == _T_5[9:0] ? image_1_204 : _GEN_779; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_781 = 10'hcd == _T_5[9:0] ? image_1_205 : _GEN_780; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_782 = 10'hce == _T_5[9:0] ? image_1_206 : _GEN_781; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_783 = 10'hcf == _T_5[9:0] ? image_1_207 : _GEN_782; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_784 = 10'hd0 == _T_5[9:0] ? image_1_208 : _GEN_783; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_785 = 10'hd1 == _T_5[9:0] ? image_1_209 : _GEN_784; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_786 = 10'hd2 == _T_5[9:0] ? image_1_210 : _GEN_785; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_787 = 10'hd3 == _T_5[9:0] ? image_1_211 : _GEN_786; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_788 = 10'hd4 == _T_5[9:0] ? image_1_212 : _GEN_787; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_789 = 10'hd5 == _T_5[9:0] ? image_1_213 : _GEN_788; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_790 = 10'hd6 == _T_5[9:0] ? image_1_214 : _GEN_789; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_791 = 10'hd7 == _T_5[9:0] ? image_1_215 : _GEN_790; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_792 = 10'hd8 == _T_5[9:0] ? image_1_216 : _GEN_791; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_793 = 10'hd9 == _T_5[9:0] ? image_1_217 : _GEN_792; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_794 = 10'hda == _T_5[9:0] ? image_1_218 : _GEN_793; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_795 = 10'hdb == _T_5[9:0] ? image_1_219 : _GEN_794; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_796 = 10'hdc == _T_5[9:0] ? image_1_220 : _GEN_795; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_797 = 10'hdd == _T_5[9:0] ? image_1_221 : _GEN_796; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_798 = 10'hde == _T_5[9:0] ? image_1_222 : _GEN_797; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_799 = 10'hdf == _T_5[9:0] ? image_1_223 : _GEN_798; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_800 = 10'he0 == _T_5[9:0] ? image_1_224 : _GEN_799; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_801 = 10'he1 == _T_5[9:0] ? image_1_225 : _GEN_800; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_802 = 10'he2 == _T_5[9:0] ? image_1_226 : _GEN_801; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_803 = 10'he3 == _T_5[9:0] ? image_1_227 : _GEN_802; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_804 = 10'he4 == _T_5[9:0] ? image_1_228 : _GEN_803; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_805 = 10'he5 == _T_5[9:0] ? image_1_229 : _GEN_804; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_806 = 10'he6 == _T_5[9:0] ? image_1_230 : _GEN_805; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_807 = 10'he7 == _T_5[9:0] ? image_1_231 : _GEN_806; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_808 = 10'he8 == _T_5[9:0] ? image_1_232 : _GEN_807; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_809 = 10'he9 == _T_5[9:0] ? image_1_233 : _GEN_808; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_810 = 10'hea == _T_5[9:0] ? image_1_234 : _GEN_809; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_811 = 10'heb == _T_5[9:0] ? image_1_235 : _GEN_810; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_812 = 10'hec == _T_5[9:0] ? image_1_236 : _GEN_811; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_813 = 10'hed == _T_5[9:0] ? image_1_237 : _GEN_812; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_814 = 10'hee == _T_5[9:0] ? image_1_238 : _GEN_813; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_815 = 10'hef == _T_5[9:0] ? image_1_239 : _GEN_814; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_816 = 10'hf0 == _T_5[9:0] ? image_1_240 : _GEN_815; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_817 = 10'hf1 == _T_5[9:0] ? image_1_241 : _GEN_816; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_818 = 10'hf2 == _T_5[9:0] ? image_1_242 : _GEN_817; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_819 = 10'hf3 == _T_5[9:0] ? image_1_243 : _GEN_818; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_820 = 10'hf4 == _T_5[9:0] ? image_1_244 : _GEN_819; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_821 = 10'hf5 == _T_5[9:0] ? image_1_245 : _GEN_820; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_822 = 10'hf6 == _T_5[9:0] ? image_1_246 : _GEN_821; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_823 = 10'hf7 == _T_5[9:0] ? image_1_247 : _GEN_822; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_824 = 10'hf8 == _T_5[9:0] ? image_1_248 : _GEN_823; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_825 = 10'hf9 == _T_5[9:0] ? image_1_249 : _GEN_824; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_826 = 10'hfa == _T_5[9:0] ? image_1_250 : _GEN_825; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_827 = 10'hfb == _T_5[9:0] ? image_1_251 : _GEN_826; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_828 = 10'hfc == _T_5[9:0] ? image_1_252 : _GEN_827; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_829 = 10'hfd == _T_5[9:0] ? image_1_253 : _GEN_828; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_830 = 10'hfe == _T_5[9:0] ? image_1_254 : _GEN_829; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_831 = 10'hff == _T_5[9:0] ? image_1_255 : _GEN_830; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_832 = 10'h100 == _T_5[9:0] ? image_1_256 : _GEN_831; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_833 = 10'h101 == _T_5[9:0] ? image_1_257 : _GEN_832; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_834 = 10'h102 == _T_5[9:0] ? image_1_258 : _GEN_833; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_835 = 10'h103 == _T_5[9:0] ? image_1_259 : _GEN_834; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_836 = 10'h104 == _T_5[9:0] ? image_1_260 : _GEN_835; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_837 = 10'h105 == _T_5[9:0] ? image_1_261 : _GEN_836; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_838 = 10'h106 == _T_5[9:0] ? image_1_262 : _GEN_837; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_839 = 10'h107 == _T_5[9:0] ? image_1_263 : _GEN_838; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_840 = 10'h108 == _T_5[9:0] ? image_1_264 : _GEN_839; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_841 = 10'h109 == _T_5[9:0] ? image_1_265 : _GEN_840; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_842 = 10'h10a == _T_5[9:0] ? image_1_266 : _GEN_841; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_843 = 10'h10b == _T_5[9:0] ? image_1_267 : _GEN_842; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_844 = 10'h10c == _T_5[9:0] ? image_1_268 : _GEN_843; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_845 = 10'h10d == _T_5[9:0] ? image_1_269 : _GEN_844; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_846 = 10'h10e == _T_5[9:0] ? image_1_270 : _GEN_845; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_847 = 10'h10f == _T_5[9:0] ? image_1_271 : _GEN_846; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_848 = 10'h110 == _T_5[9:0] ? image_1_272 : _GEN_847; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_849 = 10'h111 == _T_5[9:0] ? image_1_273 : _GEN_848; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_850 = 10'h112 == _T_5[9:0] ? image_1_274 : _GEN_849; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_851 = 10'h113 == _T_5[9:0] ? image_1_275 : _GEN_850; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_852 = 10'h114 == _T_5[9:0] ? image_1_276 : _GEN_851; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_853 = 10'h115 == _T_5[9:0] ? image_1_277 : _GEN_852; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_854 = 10'h116 == _T_5[9:0] ? image_1_278 : _GEN_853; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_855 = 10'h117 == _T_5[9:0] ? image_1_279 : _GEN_854; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_856 = 10'h118 == _T_5[9:0] ? image_1_280 : _GEN_855; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_857 = 10'h119 == _T_5[9:0] ? image_1_281 : _GEN_856; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_858 = 10'h11a == _T_5[9:0] ? image_1_282 : _GEN_857; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_859 = 10'h11b == _T_5[9:0] ? image_1_283 : _GEN_858; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_860 = 10'h11c == _T_5[9:0] ? image_1_284 : _GEN_859; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_861 = 10'h11d == _T_5[9:0] ? image_1_285 : _GEN_860; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_862 = 10'h11e == _T_5[9:0] ? image_1_286 : _GEN_861; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_863 = 10'h11f == _T_5[9:0] ? image_1_287 : _GEN_862; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_864 = 10'h120 == _T_5[9:0] ? image_1_288 : _GEN_863; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_865 = 10'h121 == _T_5[9:0] ? image_1_289 : _GEN_864; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_866 = 10'h122 == _T_5[9:0] ? image_1_290 : _GEN_865; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_867 = 10'h123 == _T_5[9:0] ? image_1_291 : _GEN_866; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_868 = 10'h124 == _T_5[9:0] ? image_1_292 : _GEN_867; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_869 = 10'h125 == _T_5[9:0] ? image_1_293 : _GEN_868; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_870 = 10'h126 == _T_5[9:0] ? image_1_294 : _GEN_869; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_871 = 10'h127 == _T_5[9:0] ? image_1_295 : _GEN_870; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_872 = 10'h128 == _T_5[9:0] ? image_1_296 : _GEN_871; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_873 = 10'h129 == _T_5[9:0] ? image_1_297 : _GEN_872; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_874 = 10'h12a == _T_5[9:0] ? image_1_298 : _GEN_873; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_875 = 10'h12b == _T_5[9:0] ? image_1_299 : _GEN_874; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_876 = 10'h12c == _T_5[9:0] ? image_1_300 : _GEN_875; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_877 = 10'h12d == _T_5[9:0] ? image_1_301 : _GEN_876; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_878 = 10'h12e == _T_5[9:0] ? image_1_302 : _GEN_877; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_879 = 10'h12f == _T_5[9:0] ? image_1_303 : _GEN_878; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_880 = 10'h130 == _T_5[9:0] ? image_1_304 : _GEN_879; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_881 = 10'h131 == _T_5[9:0] ? image_1_305 : _GEN_880; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_882 = 10'h132 == _T_5[9:0] ? image_1_306 : _GEN_881; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_883 = 10'h133 == _T_5[9:0] ? image_1_307 : _GEN_882; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_884 = 10'h134 == _T_5[9:0] ? image_1_308 : _GEN_883; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_885 = 10'h135 == _T_5[9:0] ? image_1_309 : _GEN_884; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_886 = 10'h136 == _T_5[9:0] ? image_1_310 : _GEN_885; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_887 = 10'h137 == _T_5[9:0] ? image_1_311 : _GEN_886; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_888 = 10'h138 == _T_5[9:0] ? image_1_312 : _GEN_887; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_889 = 10'h139 == _T_5[9:0] ? image_1_313 : _GEN_888; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_890 = 10'h13a == _T_5[9:0] ? image_1_314 : _GEN_889; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_891 = 10'h13b == _T_5[9:0] ? image_1_315 : _GEN_890; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_892 = 10'h13c == _T_5[9:0] ? image_1_316 : _GEN_891; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_893 = 10'h13d == _T_5[9:0] ? image_1_317 : _GEN_892; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_894 = 10'h13e == _T_5[9:0] ? image_1_318 : _GEN_893; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_895 = 10'h13f == _T_5[9:0] ? image_1_319 : _GEN_894; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_896 = 10'h140 == _T_5[9:0] ? image_1_320 : _GEN_895; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_897 = 10'h141 == _T_5[9:0] ? image_1_321 : _GEN_896; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_898 = 10'h142 == _T_5[9:0] ? image_1_322 : _GEN_897; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_899 = 10'h143 == _T_5[9:0] ? image_1_323 : _GEN_898; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_900 = 10'h144 == _T_5[9:0] ? image_1_324 : _GEN_899; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_901 = 10'h145 == _T_5[9:0] ? image_1_325 : _GEN_900; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_902 = 10'h146 == _T_5[9:0] ? image_1_326 : _GEN_901; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_903 = 10'h147 == _T_5[9:0] ? image_1_327 : _GEN_902; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_904 = 10'h148 == _T_5[9:0] ? image_1_328 : _GEN_903; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_905 = 10'h149 == _T_5[9:0] ? image_1_329 : _GEN_904; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_906 = 10'h14a == _T_5[9:0] ? image_1_330 : _GEN_905; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_907 = 10'h14b == _T_5[9:0] ? image_1_331 : _GEN_906; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_908 = 10'h14c == _T_5[9:0] ? image_1_332 : _GEN_907; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_909 = 10'h14d == _T_5[9:0] ? image_1_333 : _GEN_908; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_910 = 10'h14e == _T_5[9:0] ? image_1_334 : _GEN_909; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_911 = 10'h14f == _T_5[9:0] ? image_1_335 : _GEN_910; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_912 = 10'h150 == _T_5[9:0] ? image_1_336 : _GEN_911; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_913 = 10'h151 == _T_5[9:0] ? image_1_337 : _GEN_912; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_914 = 10'h152 == _T_5[9:0] ? image_1_338 : _GEN_913; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_915 = 10'h153 == _T_5[9:0] ? image_1_339 : _GEN_914; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_916 = 10'h154 == _T_5[9:0] ? image_1_340 : _GEN_915; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_917 = 10'h155 == _T_5[9:0] ? image_1_341 : _GEN_916; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_918 = 10'h156 == _T_5[9:0] ? image_1_342 : _GEN_917; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_919 = 10'h157 == _T_5[9:0] ? image_1_343 : _GEN_918; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_920 = 10'h158 == _T_5[9:0] ? image_1_344 : _GEN_919; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_921 = 10'h159 == _T_5[9:0] ? image_1_345 : _GEN_920; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_922 = 10'h15a == _T_5[9:0] ? image_1_346 : _GEN_921; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_923 = 10'h15b == _T_5[9:0] ? image_1_347 : _GEN_922; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_924 = 10'h15c == _T_5[9:0] ? image_1_348 : _GEN_923; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_925 = 10'h15d == _T_5[9:0] ? image_1_349 : _GEN_924; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_926 = 10'h15e == _T_5[9:0] ? image_1_350 : _GEN_925; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_927 = 10'h15f == _T_5[9:0] ? image_1_351 : _GEN_926; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_928 = 10'h160 == _T_5[9:0] ? image_1_352 : _GEN_927; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_929 = 10'h161 == _T_5[9:0] ? image_1_353 : _GEN_928; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_930 = 10'h162 == _T_5[9:0] ? image_1_354 : _GEN_929; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_931 = 10'h163 == _T_5[9:0] ? image_1_355 : _GEN_930; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_932 = 10'h164 == _T_5[9:0] ? image_1_356 : _GEN_931; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_933 = 10'h165 == _T_5[9:0] ? image_1_357 : _GEN_932; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_934 = 10'h166 == _T_5[9:0] ? image_1_358 : _GEN_933; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_935 = 10'h167 == _T_5[9:0] ? image_1_359 : _GEN_934; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_936 = 10'h168 == _T_5[9:0] ? image_1_360 : _GEN_935; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_937 = 10'h169 == _T_5[9:0] ? image_1_361 : _GEN_936; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_938 = 10'h16a == _T_5[9:0] ? image_1_362 : _GEN_937; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_939 = 10'h16b == _T_5[9:0] ? image_1_363 : _GEN_938; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_940 = 10'h16c == _T_5[9:0] ? image_1_364 : _GEN_939; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_941 = 10'h16d == _T_5[9:0] ? image_1_365 : _GEN_940; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_942 = 10'h16e == _T_5[9:0] ? image_1_366 : _GEN_941; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_943 = 10'h16f == _T_5[9:0] ? image_1_367 : _GEN_942; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_944 = 10'h170 == _T_5[9:0] ? image_1_368 : _GEN_943; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_945 = 10'h171 == _T_5[9:0] ? image_1_369 : _GEN_944; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_946 = 10'h172 == _T_5[9:0] ? image_1_370 : _GEN_945; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_947 = 10'h173 == _T_5[9:0] ? image_1_371 : _GEN_946; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_948 = 10'h174 == _T_5[9:0] ? image_1_372 : _GEN_947; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_949 = 10'h175 == _T_5[9:0] ? image_1_373 : _GEN_948; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_950 = 10'h176 == _T_5[9:0] ? image_1_374 : _GEN_949; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_951 = 10'h177 == _T_5[9:0] ? image_1_375 : _GEN_950; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_952 = 10'h178 == _T_5[9:0] ? image_1_376 : _GEN_951; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_953 = 10'h179 == _T_5[9:0] ? image_1_377 : _GEN_952; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_954 = 10'h17a == _T_5[9:0] ? image_1_378 : _GEN_953; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_955 = 10'h17b == _T_5[9:0] ? image_1_379 : _GEN_954; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_956 = 10'h17c == _T_5[9:0] ? image_1_380 : _GEN_955; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_957 = 10'h17d == _T_5[9:0] ? image_1_381 : _GEN_956; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_958 = 10'h17e == _T_5[9:0] ? image_1_382 : _GEN_957; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_959 = 10'h17f == _T_5[9:0] ? image_1_383 : _GEN_958; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_960 = 10'h180 == _T_5[9:0] ? image_1_384 : _GEN_959; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_961 = 10'h181 == _T_5[9:0] ? image_1_385 : _GEN_960; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_962 = 10'h182 == _T_5[9:0] ? image_1_386 : _GEN_961; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_963 = 10'h183 == _T_5[9:0] ? image_1_387 : _GEN_962; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_964 = 10'h184 == _T_5[9:0] ? image_1_388 : _GEN_963; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_965 = 10'h185 == _T_5[9:0] ? image_1_389 : _GEN_964; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_966 = 10'h186 == _T_5[9:0] ? image_1_390 : _GEN_965; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_967 = 10'h187 == _T_5[9:0] ? image_1_391 : _GEN_966; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_968 = 10'h188 == _T_5[9:0] ? image_1_392 : _GEN_967; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_969 = 10'h189 == _T_5[9:0] ? image_1_393 : _GEN_968; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_970 = 10'h18a == _T_5[9:0] ? image_1_394 : _GEN_969; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_971 = 10'h18b == _T_5[9:0] ? image_1_395 : _GEN_970; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_972 = 10'h18c == _T_5[9:0] ? image_1_396 : _GEN_971; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_973 = 10'h18d == _T_5[9:0] ? image_1_397 : _GEN_972; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_974 = 10'h18e == _T_5[9:0] ? image_1_398 : _GEN_973; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_975 = 10'h18f == _T_5[9:0] ? image_1_399 : _GEN_974; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_976 = 10'h190 == _T_5[9:0] ? image_1_400 : _GEN_975; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_977 = 10'h191 == _T_5[9:0] ? image_1_401 : _GEN_976; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_978 = 10'h192 == _T_5[9:0] ? image_1_402 : _GEN_977; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_979 = 10'h193 == _T_5[9:0] ? image_1_403 : _GEN_978; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_980 = 10'h194 == _T_5[9:0] ? image_1_404 : _GEN_979; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_981 = 10'h195 == _T_5[9:0] ? image_1_405 : _GEN_980; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_982 = 10'h196 == _T_5[9:0] ? image_1_406 : _GEN_981; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_983 = 10'h197 == _T_5[9:0] ? image_1_407 : _GEN_982; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_984 = 10'h198 == _T_5[9:0] ? image_1_408 : _GEN_983; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_985 = 10'h199 == _T_5[9:0] ? image_1_409 : _GEN_984; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_986 = 10'h19a == _T_5[9:0] ? image_1_410 : _GEN_985; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_987 = 10'h19b == _T_5[9:0] ? image_1_411 : _GEN_986; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_988 = 10'h19c == _T_5[9:0] ? image_1_412 : _GEN_987; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_989 = 10'h19d == _T_5[9:0] ? image_1_413 : _GEN_988; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_990 = 10'h19e == _T_5[9:0] ? image_1_414 : _GEN_989; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_991 = 10'h19f == _T_5[9:0] ? image_1_415 : _GEN_990; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_992 = 10'h1a0 == _T_5[9:0] ? image_1_416 : _GEN_991; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_993 = 10'h1a1 == _T_5[9:0] ? image_1_417 : _GEN_992; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_994 = 10'h1a2 == _T_5[9:0] ? image_1_418 : _GEN_993; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_995 = 10'h1a3 == _T_5[9:0] ? image_1_419 : _GEN_994; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_996 = 10'h1a4 == _T_5[9:0] ? image_1_420 : _GEN_995; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_997 = 10'h1a5 == _T_5[9:0] ? image_1_421 : _GEN_996; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_998 = 10'h1a6 == _T_5[9:0] ? image_1_422 : _GEN_997; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_999 = 10'h1a7 == _T_5[9:0] ? image_1_423 : _GEN_998; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1000 = 10'h1a8 == _T_5[9:0] ? image_1_424 : _GEN_999; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1001 = 10'h1a9 == _T_5[9:0] ? image_1_425 : _GEN_1000; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1002 = 10'h1aa == _T_5[9:0] ? image_1_426 : _GEN_1001; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1003 = 10'h1ab == _T_5[9:0] ? image_1_427 : _GEN_1002; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1004 = 10'h1ac == _T_5[9:0] ? image_1_428 : _GEN_1003; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1005 = 10'h1ad == _T_5[9:0] ? image_1_429 : _GEN_1004; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1006 = 10'h1ae == _T_5[9:0] ? image_1_430 : _GEN_1005; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1007 = 10'h1af == _T_5[9:0] ? image_1_431 : _GEN_1006; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1008 = 10'h1b0 == _T_5[9:0] ? image_1_432 : _GEN_1007; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1009 = 10'h1b1 == _T_5[9:0] ? image_1_433 : _GEN_1008; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1010 = 10'h1b2 == _T_5[9:0] ? image_1_434 : _GEN_1009; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1011 = 10'h1b3 == _T_5[9:0] ? image_1_435 : _GEN_1010; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1012 = 10'h1b4 == _T_5[9:0] ? image_1_436 : _GEN_1011; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1013 = 10'h1b5 == _T_5[9:0] ? image_1_437 : _GEN_1012; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1014 = 10'h1b6 == _T_5[9:0] ? image_1_438 : _GEN_1013; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1015 = 10'h1b7 == _T_5[9:0] ? image_1_439 : _GEN_1014; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1016 = 10'h1b8 == _T_5[9:0] ? image_1_440 : _GEN_1015; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1017 = 10'h1b9 == _T_5[9:0] ? image_1_441 : _GEN_1016; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1018 = 10'h1ba == _T_5[9:0] ? image_1_442 : _GEN_1017; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1019 = 10'h1bb == _T_5[9:0] ? image_1_443 : _GEN_1018; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1020 = 10'h1bc == _T_5[9:0] ? image_1_444 : _GEN_1019; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1021 = 10'h1bd == _T_5[9:0] ? image_1_445 : _GEN_1020; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1022 = 10'h1be == _T_5[9:0] ? image_1_446 : _GEN_1021; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1023 = 10'h1bf == _T_5[9:0] ? image_1_447 : _GEN_1022; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1024 = 10'h1c0 == _T_5[9:0] ? image_1_448 : _GEN_1023; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1025 = 10'h1c1 == _T_5[9:0] ? image_1_449 : _GEN_1024; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1026 = 10'h1c2 == _T_5[9:0] ? image_1_450 : _GEN_1025; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1027 = 10'h1c3 == _T_5[9:0] ? image_1_451 : _GEN_1026; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1028 = 10'h1c4 == _T_5[9:0] ? image_1_452 : _GEN_1027; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1029 = 10'h1c5 == _T_5[9:0] ? image_1_453 : _GEN_1028; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1030 = 10'h1c6 == _T_5[9:0] ? image_1_454 : _GEN_1029; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1031 = 10'h1c7 == _T_5[9:0] ? image_1_455 : _GEN_1030; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1032 = 10'h1c8 == _T_5[9:0] ? image_1_456 : _GEN_1031; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1033 = 10'h1c9 == _T_5[9:0] ? image_1_457 : _GEN_1032; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1034 = 10'h1ca == _T_5[9:0] ? image_1_458 : _GEN_1033; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1035 = 10'h1cb == _T_5[9:0] ? image_1_459 : _GEN_1034; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1036 = 10'h1cc == _T_5[9:0] ? image_1_460 : _GEN_1035; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1037 = 10'h1cd == _T_5[9:0] ? image_1_461 : _GEN_1036; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1038 = 10'h1ce == _T_5[9:0] ? image_1_462 : _GEN_1037; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1039 = 10'h1cf == _T_5[9:0] ? image_1_463 : _GEN_1038; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1040 = 10'h1d0 == _T_5[9:0] ? image_1_464 : _GEN_1039; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1041 = 10'h1d1 == _T_5[9:0] ? image_1_465 : _GEN_1040; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1042 = 10'h1d2 == _T_5[9:0] ? image_1_466 : _GEN_1041; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1043 = 10'h1d3 == _T_5[9:0] ? image_1_467 : _GEN_1042; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1044 = 10'h1d4 == _T_5[9:0] ? image_1_468 : _GEN_1043; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1045 = 10'h1d5 == _T_5[9:0] ? image_1_469 : _GEN_1044; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1046 = 10'h1d6 == _T_5[9:0] ? image_1_470 : _GEN_1045; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1047 = 10'h1d7 == _T_5[9:0] ? image_1_471 : _GEN_1046; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1048 = 10'h1d8 == _T_5[9:0] ? image_1_472 : _GEN_1047; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1049 = 10'h1d9 == _T_5[9:0] ? image_1_473 : _GEN_1048; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1050 = 10'h1da == _T_5[9:0] ? image_1_474 : _GEN_1049; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1051 = 10'h1db == _T_5[9:0] ? image_1_475 : _GEN_1050; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1052 = 10'h1dc == _T_5[9:0] ? image_1_476 : _GEN_1051; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1053 = 10'h1dd == _T_5[9:0] ? image_1_477 : _GEN_1052; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1054 = 10'h1de == _T_5[9:0] ? image_1_478 : _GEN_1053; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1055 = 10'h1df == _T_5[9:0] ? image_1_479 : _GEN_1054; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1056 = 10'h1e0 == _T_5[9:0] ? image_1_480 : _GEN_1055; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1057 = 10'h1e1 == _T_5[9:0] ? image_1_481 : _GEN_1056; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1058 = 10'h1e2 == _T_5[9:0] ? image_1_482 : _GEN_1057; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1059 = 10'h1e3 == _T_5[9:0] ? image_1_483 : _GEN_1058; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1060 = 10'h1e4 == _T_5[9:0] ? image_1_484 : _GEN_1059; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1061 = 10'h1e5 == _T_5[9:0] ? image_1_485 : _GEN_1060; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1062 = 10'h1e6 == _T_5[9:0] ? image_1_486 : _GEN_1061; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1063 = 10'h1e7 == _T_5[9:0] ? image_1_487 : _GEN_1062; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1064 = 10'h1e8 == _T_5[9:0] ? image_1_488 : _GEN_1063; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1065 = 10'h1e9 == _T_5[9:0] ? image_1_489 : _GEN_1064; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1066 = 10'h1ea == _T_5[9:0] ? image_1_490 : _GEN_1065; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1067 = 10'h1eb == _T_5[9:0] ? image_1_491 : _GEN_1066; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1068 = 10'h1ec == _T_5[9:0] ? image_1_492 : _GEN_1067; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1069 = 10'h1ed == _T_5[9:0] ? image_1_493 : _GEN_1068; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1070 = 10'h1ee == _T_5[9:0] ? image_1_494 : _GEN_1069; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1071 = 10'h1ef == _T_5[9:0] ? image_1_495 : _GEN_1070; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1072 = 10'h1f0 == _T_5[9:0] ? image_1_496 : _GEN_1071; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1073 = 10'h1f1 == _T_5[9:0] ? image_1_497 : _GEN_1072; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1074 = 10'h1f2 == _T_5[9:0] ? image_1_498 : _GEN_1073; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1075 = 10'h1f3 == _T_5[9:0] ? image_1_499 : _GEN_1074; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1076 = 10'h1f4 == _T_5[9:0] ? image_1_500 : _GEN_1075; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1077 = 10'h1f5 == _T_5[9:0] ? image_1_501 : _GEN_1076; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1078 = 10'h1f6 == _T_5[9:0] ? image_1_502 : _GEN_1077; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1079 = 10'h1f7 == _T_5[9:0] ? image_1_503 : _GEN_1078; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1080 = 10'h1f8 == _T_5[9:0] ? image_1_504 : _GEN_1079; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1081 = 10'h1f9 == _T_5[9:0] ? image_1_505 : _GEN_1080; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1082 = 10'h1fa == _T_5[9:0] ? image_1_506 : _GEN_1081; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1083 = 10'h1fb == _T_5[9:0] ? image_1_507 : _GEN_1082; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1084 = 10'h1fc == _T_5[9:0] ? image_1_508 : _GEN_1083; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1085 = 10'h1fd == _T_5[9:0] ? image_1_509 : _GEN_1084; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1086 = 10'h1fe == _T_5[9:0] ? image_1_510 : _GEN_1085; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1087 = 10'h1ff == _T_5[9:0] ? image_1_511 : _GEN_1086; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1088 = 10'h200 == _T_5[9:0] ? image_1_512 : _GEN_1087; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1089 = 10'h201 == _T_5[9:0] ? image_1_513 : _GEN_1088; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1090 = 10'h202 == _T_5[9:0] ? image_1_514 : _GEN_1089; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1091 = 10'h203 == _T_5[9:0] ? image_1_515 : _GEN_1090; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1092 = 10'h204 == _T_5[9:0] ? image_1_516 : _GEN_1091; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1093 = 10'h205 == _T_5[9:0] ? image_1_517 : _GEN_1092; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1094 = 10'h206 == _T_5[9:0] ? image_1_518 : _GEN_1093; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1095 = 10'h207 == _T_5[9:0] ? image_1_519 : _GEN_1094; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1096 = 10'h208 == _T_5[9:0] ? image_1_520 : _GEN_1095; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1097 = 10'h209 == _T_5[9:0] ? image_1_521 : _GEN_1096; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1098 = 10'h20a == _T_5[9:0] ? image_1_522 : _GEN_1097; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1099 = 10'h20b == _T_5[9:0] ? image_1_523 : _GEN_1098; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1100 = 10'h20c == _T_5[9:0] ? image_1_524 : _GEN_1099; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1101 = 10'h20d == _T_5[9:0] ? image_1_525 : _GEN_1100; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1102 = 10'h20e == _T_5[9:0] ? image_1_526 : _GEN_1101; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1103 = 10'h20f == _T_5[9:0] ? image_1_527 : _GEN_1102; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1104 = 10'h210 == _T_5[9:0] ? image_1_528 : _GEN_1103; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1105 = 10'h211 == _T_5[9:0] ? image_1_529 : _GEN_1104; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1106 = 10'h212 == _T_5[9:0] ? image_1_530 : _GEN_1105; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1107 = 10'h213 == _T_5[9:0] ? image_1_531 : _GEN_1106; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1108 = 10'h214 == _T_5[9:0] ? image_1_532 : _GEN_1107; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1109 = 10'h215 == _T_5[9:0] ? image_1_533 : _GEN_1108; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1110 = 10'h216 == _T_5[9:0] ? image_1_534 : _GEN_1109; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1111 = 10'h217 == _T_5[9:0] ? image_1_535 : _GEN_1110; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1112 = 10'h218 == _T_5[9:0] ? image_1_536 : _GEN_1111; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1113 = 10'h219 == _T_5[9:0] ? image_1_537 : _GEN_1112; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1114 = 10'h21a == _T_5[9:0] ? image_1_538 : _GEN_1113; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1115 = 10'h21b == _T_5[9:0] ? image_1_539 : _GEN_1114; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1116 = 10'h21c == _T_5[9:0] ? image_1_540 : _GEN_1115; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1117 = 10'h21d == _T_5[9:0] ? image_1_541 : _GEN_1116; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1118 = 10'h21e == _T_5[9:0] ? image_1_542 : _GEN_1117; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1119 = 10'h21f == _T_5[9:0] ? image_1_543 : _GEN_1118; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1120 = 10'h220 == _T_5[9:0] ? image_1_544 : _GEN_1119; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1121 = 10'h221 == _T_5[9:0] ? image_1_545 : _GEN_1120; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1122 = 10'h222 == _T_5[9:0] ? image_1_546 : _GEN_1121; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1123 = 10'h223 == _T_5[9:0] ? image_1_547 : _GEN_1122; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1124 = 10'h224 == _T_5[9:0] ? image_1_548 : _GEN_1123; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1125 = 10'h225 == _T_5[9:0] ? image_1_549 : _GEN_1124; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1126 = 10'h226 == _T_5[9:0] ? image_1_550 : _GEN_1125; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1127 = 10'h227 == _T_5[9:0] ? image_1_551 : _GEN_1126; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1128 = 10'h228 == _T_5[9:0] ? image_1_552 : _GEN_1127; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1129 = 10'h229 == _T_5[9:0] ? image_1_553 : _GEN_1128; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1130 = 10'h22a == _T_5[9:0] ? image_1_554 : _GEN_1129; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1131 = 10'h22b == _T_5[9:0] ? image_1_555 : _GEN_1130; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1132 = 10'h22c == _T_5[9:0] ? image_1_556 : _GEN_1131; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1133 = 10'h22d == _T_5[9:0] ? image_1_557 : _GEN_1132; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1134 = 10'h22e == _T_5[9:0] ? image_1_558 : _GEN_1133; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1135 = 10'h22f == _T_5[9:0] ? image_1_559 : _GEN_1134; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1136 = 10'h230 == _T_5[9:0] ? image_1_560 : _GEN_1135; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1137 = 10'h231 == _T_5[9:0] ? image_1_561 : _GEN_1136; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1138 = 10'h232 == _T_5[9:0] ? image_1_562 : _GEN_1137; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1139 = 10'h233 == _T_5[9:0] ? image_1_563 : _GEN_1138; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1140 = 10'h234 == _T_5[9:0] ? image_1_564 : _GEN_1139; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1141 = 10'h235 == _T_5[9:0] ? image_1_565 : _GEN_1140; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1142 = 10'h236 == _T_5[9:0] ? image_1_566 : _GEN_1141; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1143 = 10'h237 == _T_5[9:0] ? image_1_567 : _GEN_1142; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1144 = 10'h238 == _T_5[9:0] ? image_1_568 : _GEN_1143; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1145 = 10'h239 == _T_5[9:0] ? image_1_569 : _GEN_1144; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1146 = 10'h23a == _T_5[9:0] ? image_1_570 : _GEN_1145; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1147 = 10'h23b == _T_5[9:0] ? image_1_571 : _GEN_1146; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1148 = 10'h23c == _T_5[9:0] ? image_1_572 : _GEN_1147; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1149 = 10'h23d == _T_5[9:0] ? image_1_573 : _GEN_1148; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1150 = 10'h23e == _T_5[9:0] ? image_1_574 : _GEN_1149; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1153 = 10'h1 == _T_5[9:0] ? image_2_1 : image_2_0; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1154 = 10'h2 == _T_5[9:0] ? image_2_2 : _GEN_1153; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1155 = 10'h3 == _T_5[9:0] ? image_2_3 : _GEN_1154; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1156 = 10'h4 == _T_5[9:0] ? image_2_4 : _GEN_1155; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1157 = 10'h5 == _T_5[9:0] ? image_2_5 : _GEN_1156; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1158 = 10'h6 == _T_5[9:0] ? image_2_6 : _GEN_1157; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1159 = 10'h7 == _T_5[9:0] ? image_2_7 : _GEN_1158; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1160 = 10'h8 == _T_5[9:0] ? image_2_8 : _GEN_1159; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1161 = 10'h9 == _T_5[9:0] ? image_2_9 : _GEN_1160; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1162 = 10'ha == _T_5[9:0] ? image_2_10 : _GEN_1161; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1163 = 10'hb == _T_5[9:0] ? image_2_11 : _GEN_1162; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1164 = 10'hc == _T_5[9:0] ? image_2_12 : _GEN_1163; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1165 = 10'hd == _T_5[9:0] ? image_2_13 : _GEN_1164; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1166 = 10'he == _T_5[9:0] ? image_2_14 : _GEN_1165; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1167 = 10'hf == _T_5[9:0] ? image_2_15 : _GEN_1166; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1168 = 10'h10 == _T_5[9:0] ? image_2_16 : _GEN_1167; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1169 = 10'h11 == _T_5[9:0] ? image_2_17 : _GEN_1168; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1170 = 10'h12 == _T_5[9:0] ? image_2_18 : _GEN_1169; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1171 = 10'h13 == _T_5[9:0] ? image_2_19 : _GEN_1170; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1172 = 10'h14 == _T_5[9:0] ? image_2_20 : _GEN_1171; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1173 = 10'h15 == _T_5[9:0] ? image_2_21 : _GEN_1172; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1174 = 10'h16 == _T_5[9:0] ? image_2_22 : _GEN_1173; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1175 = 10'h17 == _T_5[9:0] ? image_2_23 : _GEN_1174; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1176 = 10'h18 == _T_5[9:0] ? image_2_24 : _GEN_1175; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1177 = 10'h19 == _T_5[9:0] ? image_2_25 : _GEN_1176; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1178 = 10'h1a == _T_5[9:0] ? image_2_26 : _GEN_1177; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1179 = 10'h1b == _T_5[9:0] ? image_2_27 : _GEN_1178; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1180 = 10'h1c == _T_5[9:0] ? image_2_28 : _GEN_1179; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1181 = 10'h1d == _T_5[9:0] ? image_2_29 : _GEN_1180; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1182 = 10'h1e == _T_5[9:0] ? image_2_30 : _GEN_1181; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1183 = 10'h1f == _T_5[9:0] ? image_2_31 : _GEN_1182; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1184 = 10'h20 == _T_5[9:0] ? image_2_32 : _GEN_1183; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1185 = 10'h21 == _T_5[9:0] ? image_2_33 : _GEN_1184; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1186 = 10'h22 == _T_5[9:0] ? image_2_34 : _GEN_1185; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1187 = 10'h23 == _T_5[9:0] ? image_2_35 : _GEN_1186; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1188 = 10'h24 == _T_5[9:0] ? image_2_36 : _GEN_1187; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1189 = 10'h25 == _T_5[9:0] ? image_2_37 : _GEN_1188; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1190 = 10'h26 == _T_5[9:0] ? image_2_38 : _GEN_1189; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1191 = 10'h27 == _T_5[9:0] ? image_2_39 : _GEN_1190; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1192 = 10'h28 == _T_5[9:0] ? image_2_40 : _GEN_1191; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1193 = 10'h29 == _T_5[9:0] ? image_2_41 : _GEN_1192; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1194 = 10'h2a == _T_5[9:0] ? image_2_42 : _GEN_1193; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1195 = 10'h2b == _T_5[9:0] ? image_2_43 : _GEN_1194; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1196 = 10'h2c == _T_5[9:0] ? image_2_44 : _GEN_1195; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1197 = 10'h2d == _T_5[9:0] ? image_2_45 : _GEN_1196; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1198 = 10'h2e == _T_5[9:0] ? image_2_46 : _GEN_1197; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1199 = 10'h2f == _T_5[9:0] ? image_2_47 : _GEN_1198; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1200 = 10'h30 == _T_5[9:0] ? image_2_48 : _GEN_1199; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1201 = 10'h31 == _T_5[9:0] ? image_2_49 : _GEN_1200; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1202 = 10'h32 == _T_5[9:0] ? image_2_50 : _GEN_1201; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1203 = 10'h33 == _T_5[9:0] ? image_2_51 : _GEN_1202; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1204 = 10'h34 == _T_5[9:0] ? image_2_52 : _GEN_1203; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1205 = 10'h35 == _T_5[9:0] ? image_2_53 : _GEN_1204; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1206 = 10'h36 == _T_5[9:0] ? image_2_54 : _GEN_1205; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1207 = 10'h37 == _T_5[9:0] ? image_2_55 : _GEN_1206; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1208 = 10'h38 == _T_5[9:0] ? image_2_56 : _GEN_1207; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1209 = 10'h39 == _T_5[9:0] ? image_2_57 : _GEN_1208; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1210 = 10'h3a == _T_5[9:0] ? image_2_58 : _GEN_1209; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1211 = 10'h3b == _T_5[9:0] ? image_2_59 : _GEN_1210; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1212 = 10'h3c == _T_5[9:0] ? image_2_60 : _GEN_1211; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1213 = 10'h3d == _T_5[9:0] ? image_2_61 : _GEN_1212; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1214 = 10'h3e == _T_5[9:0] ? image_2_62 : _GEN_1213; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1215 = 10'h3f == _T_5[9:0] ? image_2_63 : _GEN_1214; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1216 = 10'h40 == _T_5[9:0] ? image_2_64 : _GEN_1215; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1217 = 10'h41 == _T_5[9:0] ? image_2_65 : _GEN_1216; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1218 = 10'h42 == _T_5[9:0] ? image_2_66 : _GEN_1217; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1219 = 10'h43 == _T_5[9:0] ? image_2_67 : _GEN_1218; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1220 = 10'h44 == _T_5[9:0] ? image_2_68 : _GEN_1219; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1221 = 10'h45 == _T_5[9:0] ? image_2_69 : _GEN_1220; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1222 = 10'h46 == _T_5[9:0] ? image_2_70 : _GEN_1221; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1223 = 10'h47 == _T_5[9:0] ? image_2_71 : _GEN_1222; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1224 = 10'h48 == _T_5[9:0] ? image_2_72 : _GEN_1223; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1225 = 10'h49 == _T_5[9:0] ? image_2_73 : _GEN_1224; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1226 = 10'h4a == _T_5[9:0] ? image_2_74 : _GEN_1225; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1227 = 10'h4b == _T_5[9:0] ? image_2_75 : _GEN_1226; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1228 = 10'h4c == _T_5[9:0] ? image_2_76 : _GEN_1227; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1229 = 10'h4d == _T_5[9:0] ? image_2_77 : _GEN_1228; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1230 = 10'h4e == _T_5[9:0] ? image_2_78 : _GEN_1229; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1231 = 10'h4f == _T_5[9:0] ? image_2_79 : _GEN_1230; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1232 = 10'h50 == _T_5[9:0] ? image_2_80 : _GEN_1231; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1233 = 10'h51 == _T_5[9:0] ? image_2_81 : _GEN_1232; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1234 = 10'h52 == _T_5[9:0] ? image_2_82 : _GEN_1233; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1235 = 10'h53 == _T_5[9:0] ? image_2_83 : _GEN_1234; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1236 = 10'h54 == _T_5[9:0] ? image_2_84 : _GEN_1235; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1237 = 10'h55 == _T_5[9:0] ? image_2_85 : _GEN_1236; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1238 = 10'h56 == _T_5[9:0] ? image_2_86 : _GEN_1237; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1239 = 10'h57 == _T_5[9:0] ? image_2_87 : _GEN_1238; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1240 = 10'h58 == _T_5[9:0] ? image_2_88 : _GEN_1239; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1241 = 10'h59 == _T_5[9:0] ? image_2_89 : _GEN_1240; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1242 = 10'h5a == _T_5[9:0] ? image_2_90 : _GEN_1241; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1243 = 10'h5b == _T_5[9:0] ? image_2_91 : _GEN_1242; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1244 = 10'h5c == _T_5[9:0] ? image_2_92 : _GEN_1243; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1245 = 10'h5d == _T_5[9:0] ? image_2_93 : _GEN_1244; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1246 = 10'h5e == _T_5[9:0] ? image_2_94 : _GEN_1245; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1247 = 10'h5f == _T_5[9:0] ? image_2_95 : _GEN_1246; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1248 = 10'h60 == _T_5[9:0] ? image_2_96 : _GEN_1247; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1249 = 10'h61 == _T_5[9:0] ? image_2_97 : _GEN_1248; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1250 = 10'h62 == _T_5[9:0] ? image_2_98 : _GEN_1249; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1251 = 10'h63 == _T_5[9:0] ? image_2_99 : _GEN_1250; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1252 = 10'h64 == _T_5[9:0] ? image_2_100 : _GEN_1251; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1253 = 10'h65 == _T_5[9:0] ? image_2_101 : _GEN_1252; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1254 = 10'h66 == _T_5[9:0] ? image_2_102 : _GEN_1253; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1255 = 10'h67 == _T_5[9:0] ? image_2_103 : _GEN_1254; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1256 = 10'h68 == _T_5[9:0] ? image_2_104 : _GEN_1255; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1257 = 10'h69 == _T_5[9:0] ? image_2_105 : _GEN_1256; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1258 = 10'h6a == _T_5[9:0] ? image_2_106 : _GEN_1257; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1259 = 10'h6b == _T_5[9:0] ? image_2_107 : _GEN_1258; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1260 = 10'h6c == _T_5[9:0] ? image_2_108 : _GEN_1259; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1261 = 10'h6d == _T_5[9:0] ? image_2_109 : _GEN_1260; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1262 = 10'h6e == _T_5[9:0] ? image_2_110 : _GEN_1261; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1263 = 10'h6f == _T_5[9:0] ? image_2_111 : _GEN_1262; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1264 = 10'h70 == _T_5[9:0] ? image_2_112 : _GEN_1263; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1265 = 10'h71 == _T_5[9:0] ? image_2_113 : _GEN_1264; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1266 = 10'h72 == _T_5[9:0] ? image_2_114 : _GEN_1265; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1267 = 10'h73 == _T_5[9:0] ? image_2_115 : _GEN_1266; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1268 = 10'h74 == _T_5[9:0] ? image_2_116 : _GEN_1267; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1269 = 10'h75 == _T_5[9:0] ? image_2_117 : _GEN_1268; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1270 = 10'h76 == _T_5[9:0] ? image_2_118 : _GEN_1269; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1271 = 10'h77 == _T_5[9:0] ? image_2_119 : _GEN_1270; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1272 = 10'h78 == _T_5[9:0] ? image_2_120 : _GEN_1271; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1273 = 10'h79 == _T_5[9:0] ? image_2_121 : _GEN_1272; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1274 = 10'h7a == _T_5[9:0] ? image_2_122 : _GEN_1273; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1275 = 10'h7b == _T_5[9:0] ? image_2_123 : _GEN_1274; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1276 = 10'h7c == _T_5[9:0] ? image_2_124 : _GEN_1275; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1277 = 10'h7d == _T_5[9:0] ? image_2_125 : _GEN_1276; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1278 = 10'h7e == _T_5[9:0] ? image_2_126 : _GEN_1277; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1279 = 10'h7f == _T_5[9:0] ? image_2_127 : _GEN_1278; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1280 = 10'h80 == _T_5[9:0] ? image_2_128 : _GEN_1279; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1281 = 10'h81 == _T_5[9:0] ? image_2_129 : _GEN_1280; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1282 = 10'h82 == _T_5[9:0] ? image_2_130 : _GEN_1281; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1283 = 10'h83 == _T_5[9:0] ? image_2_131 : _GEN_1282; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1284 = 10'h84 == _T_5[9:0] ? image_2_132 : _GEN_1283; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1285 = 10'h85 == _T_5[9:0] ? image_2_133 : _GEN_1284; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1286 = 10'h86 == _T_5[9:0] ? image_2_134 : _GEN_1285; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1287 = 10'h87 == _T_5[9:0] ? image_2_135 : _GEN_1286; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1288 = 10'h88 == _T_5[9:0] ? image_2_136 : _GEN_1287; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1289 = 10'h89 == _T_5[9:0] ? image_2_137 : _GEN_1288; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1290 = 10'h8a == _T_5[9:0] ? image_2_138 : _GEN_1289; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1291 = 10'h8b == _T_5[9:0] ? image_2_139 : _GEN_1290; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1292 = 10'h8c == _T_5[9:0] ? image_2_140 : _GEN_1291; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1293 = 10'h8d == _T_5[9:0] ? image_2_141 : _GEN_1292; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1294 = 10'h8e == _T_5[9:0] ? image_2_142 : _GEN_1293; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1295 = 10'h8f == _T_5[9:0] ? image_2_143 : _GEN_1294; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1296 = 10'h90 == _T_5[9:0] ? image_2_144 : _GEN_1295; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1297 = 10'h91 == _T_5[9:0] ? image_2_145 : _GEN_1296; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1298 = 10'h92 == _T_5[9:0] ? image_2_146 : _GEN_1297; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1299 = 10'h93 == _T_5[9:0] ? image_2_147 : _GEN_1298; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1300 = 10'h94 == _T_5[9:0] ? image_2_148 : _GEN_1299; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1301 = 10'h95 == _T_5[9:0] ? image_2_149 : _GEN_1300; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1302 = 10'h96 == _T_5[9:0] ? image_2_150 : _GEN_1301; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1303 = 10'h97 == _T_5[9:0] ? image_2_151 : _GEN_1302; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1304 = 10'h98 == _T_5[9:0] ? image_2_152 : _GEN_1303; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1305 = 10'h99 == _T_5[9:0] ? image_2_153 : _GEN_1304; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1306 = 10'h9a == _T_5[9:0] ? image_2_154 : _GEN_1305; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1307 = 10'h9b == _T_5[9:0] ? image_2_155 : _GEN_1306; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1308 = 10'h9c == _T_5[9:0] ? image_2_156 : _GEN_1307; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1309 = 10'h9d == _T_5[9:0] ? image_2_157 : _GEN_1308; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1310 = 10'h9e == _T_5[9:0] ? image_2_158 : _GEN_1309; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1311 = 10'h9f == _T_5[9:0] ? image_2_159 : _GEN_1310; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1312 = 10'ha0 == _T_5[9:0] ? image_2_160 : _GEN_1311; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1313 = 10'ha1 == _T_5[9:0] ? image_2_161 : _GEN_1312; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1314 = 10'ha2 == _T_5[9:0] ? image_2_162 : _GEN_1313; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1315 = 10'ha3 == _T_5[9:0] ? image_2_163 : _GEN_1314; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1316 = 10'ha4 == _T_5[9:0] ? image_2_164 : _GEN_1315; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1317 = 10'ha5 == _T_5[9:0] ? image_2_165 : _GEN_1316; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1318 = 10'ha6 == _T_5[9:0] ? image_2_166 : _GEN_1317; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1319 = 10'ha7 == _T_5[9:0] ? image_2_167 : _GEN_1318; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1320 = 10'ha8 == _T_5[9:0] ? image_2_168 : _GEN_1319; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1321 = 10'ha9 == _T_5[9:0] ? image_2_169 : _GEN_1320; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1322 = 10'haa == _T_5[9:0] ? image_2_170 : _GEN_1321; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1323 = 10'hab == _T_5[9:0] ? image_2_171 : _GEN_1322; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1324 = 10'hac == _T_5[9:0] ? image_2_172 : _GEN_1323; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1325 = 10'had == _T_5[9:0] ? image_2_173 : _GEN_1324; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1326 = 10'hae == _T_5[9:0] ? image_2_174 : _GEN_1325; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1327 = 10'haf == _T_5[9:0] ? image_2_175 : _GEN_1326; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1328 = 10'hb0 == _T_5[9:0] ? image_2_176 : _GEN_1327; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1329 = 10'hb1 == _T_5[9:0] ? image_2_177 : _GEN_1328; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1330 = 10'hb2 == _T_5[9:0] ? image_2_178 : _GEN_1329; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1331 = 10'hb3 == _T_5[9:0] ? image_2_179 : _GEN_1330; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1332 = 10'hb4 == _T_5[9:0] ? image_2_180 : _GEN_1331; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1333 = 10'hb5 == _T_5[9:0] ? image_2_181 : _GEN_1332; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1334 = 10'hb6 == _T_5[9:0] ? image_2_182 : _GEN_1333; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1335 = 10'hb7 == _T_5[9:0] ? image_2_183 : _GEN_1334; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1336 = 10'hb8 == _T_5[9:0] ? image_2_184 : _GEN_1335; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1337 = 10'hb9 == _T_5[9:0] ? image_2_185 : _GEN_1336; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1338 = 10'hba == _T_5[9:0] ? image_2_186 : _GEN_1337; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1339 = 10'hbb == _T_5[9:0] ? image_2_187 : _GEN_1338; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1340 = 10'hbc == _T_5[9:0] ? image_2_188 : _GEN_1339; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1341 = 10'hbd == _T_5[9:0] ? image_2_189 : _GEN_1340; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1342 = 10'hbe == _T_5[9:0] ? image_2_190 : _GEN_1341; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1343 = 10'hbf == _T_5[9:0] ? image_2_191 : _GEN_1342; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1344 = 10'hc0 == _T_5[9:0] ? image_2_192 : _GEN_1343; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1345 = 10'hc1 == _T_5[9:0] ? image_2_193 : _GEN_1344; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1346 = 10'hc2 == _T_5[9:0] ? image_2_194 : _GEN_1345; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1347 = 10'hc3 == _T_5[9:0] ? image_2_195 : _GEN_1346; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1348 = 10'hc4 == _T_5[9:0] ? image_2_196 : _GEN_1347; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1349 = 10'hc5 == _T_5[9:0] ? image_2_197 : _GEN_1348; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1350 = 10'hc6 == _T_5[9:0] ? image_2_198 : _GEN_1349; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1351 = 10'hc7 == _T_5[9:0] ? image_2_199 : _GEN_1350; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1352 = 10'hc8 == _T_5[9:0] ? image_2_200 : _GEN_1351; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1353 = 10'hc9 == _T_5[9:0] ? image_2_201 : _GEN_1352; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1354 = 10'hca == _T_5[9:0] ? image_2_202 : _GEN_1353; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1355 = 10'hcb == _T_5[9:0] ? image_2_203 : _GEN_1354; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1356 = 10'hcc == _T_5[9:0] ? image_2_204 : _GEN_1355; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1357 = 10'hcd == _T_5[9:0] ? image_2_205 : _GEN_1356; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1358 = 10'hce == _T_5[9:0] ? image_2_206 : _GEN_1357; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1359 = 10'hcf == _T_5[9:0] ? image_2_207 : _GEN_1358; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1360 = 10'hd0 == _T_5[9:0] ? image_2_208 : _GEN_1359; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1361 = 10'hd1 == _T_5[9:0] ? image_2_209 : _GEN_1360; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1362 = 10'hd2 == _T_5[9:0] ? image_2_210 : _GEN_1361; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1363 = 10'hd3 == _T_5[9:0] ? image_2_211 : _GEN_1362; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1364 = 10'hd4 == _T_5[9:0] ? image_2_212 : _GEN_1363; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1365 = 10'hd5 == _T_5[9:0] ? image_2_213 : _GEN_1364; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1366 = 10'hd6 == _T_5[9:0] ? image_2_214 : _GEN_1365; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1367 = 10'hd7 == _T_5[9:0] ? image_2_215 : _GEN_1366; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1368 = 10'hd8 == _T_5[9:0] ? image_2_216 : _GEN_1367; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1369 = 10'hd9 == _T_5[9:0] ? image_2_217 : _GEN_1368; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1370 = 10'hda == _T_5[9:0] ? image_2_218 : _GEN_1369; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1371 = 10'hdb == _T_5[9:0] ? image_2_219 : _GEN_1370; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1372 = 10'hdc == _T_5[9:0] ? image_2_220 : _GEN_1371; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1373 = 10'hdd == _T_5[9:0] ? image_2_221 : _GEN_1372; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1374 = 10'hde == _T_5[9:0] ? image_2_222 : _GEN_1373; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1375 = 10'hdf == _T_5[9:0] ? image_2_223 : _GEN_1374; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1376 = 10'he0 == _T_5[9:0] ? image_2_224 : _GEN_1375; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1377 = 10'he1 == _T_5[9:0] ? image_2_225 : _GEN_1376; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1378 = 10'he2 == _T_5[9:0] ? image_2_226 : _GEN_1377; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1379 = 10'he3 == _T_5[9:0] ? image_2_227 : _GEN_1378; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1380 = 10'he4 == _T_5[9:0] ? image_2_228 : _GEN_1379; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1381 = 10'he5 == _T_5[9:0] ? image_2_229 : _GEN_1380; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1382 = 10'he6 == _T_5[9:0] ? image_2_230 : _GEN_1381; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1383 = 10'he7 == _T_5[9:0] ? image_2_231 : _GEN_1382; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1384 = 10'he8 == _T_5[9:0] ? image_2_232 : _GEN_1383; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1385 = 10'he9 == _T_5[9:0] ? image_2_233 : _GEN_1384; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1386 = 10'hea == _T_5[9:0] ? image_2_234 : _GEN_1385; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1387 = 10'heb == _T_5[9:0] ? image_2_235 : _GEN_1386; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1388 = 10'hec == _T_5[9:0] ? image_2_236 : _GEN_1387; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1389 = 10'hed == _T_5[9:0] ? image_2_237 : _GEN_1388; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1390 = 10'hee == _T_5[9:0] ? image_2_238 : _GEN_1389; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1391 = 10'hef == _T_5[9:0] ? image_2_239 : _GEN_1390; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1392 = 10'hf0 == _T_5[9:0] ? image_2_240 : _GEN_1391; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1393 = 10'hf1 == _T_5[9:0] ? image_2_241 : _GEN_1392; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1394 = 10'hf2 == _T_5[9:0] ? image_2_242 : _GEN_1393; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1395 = 10'hf3 == _T_5[9:0] ? image_2_243 : _GEN_1394; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1396 = 10'hf4 == _T_5[9:0] ? image_2_244 : _GEN_1395; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1397 = 10'hf5 == _T_5[9:0] ? image_2_245 : _GEN_1396; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1398 = 10'hf6 == _T_5[9:0] ? image_2_246 : _GEN_1397; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1399 = 10'hf7 == _T_5[9:0] ? image_2_247 : _GEN_1398; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1400 = 10'hf8 == _T_5[9:0] ? image_2_248 : _GEN_1399; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1401 = 10'hf9 == _T_5[9:0] ? image_2_249 : _GEN_1400; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1402 = 10'hfa == _T_5[9:0] ? image_2_250 : _GEN_1401; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1403 = 10'hfb == _T_5[9:0] ? image_2_251 : _GEN_1402; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1404 = 10'hfc == _T_5[9:0] ? image_2_252 : _GEN_1403; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1405 = 10'hfd == _T_5[9:0] ? image_2_253 : _GEN_1404; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1406 = 10'hfe == _T_5[9:0] ? image_2_254 : _GEN_1405; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1407 = 10'hff == _T_5[9:0] ? image_2_255 : _GEN_1406; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1408 = 10'h100 == _T_5[9:0] ? image_2_256 : _GEN_1407; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1409 = 10'h101 == _T_5[9:0] ? image_2_257 : _GEN_1408; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1410 = 10'h102 == _T_5[9:0] ? image_2_258 : _GEN_1409; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1411 = 10'h103 == _T_5[9:0] ? image_2_259 : _GEN_1410; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1412 = 10'h104 == _T_5[9:0] ? image_2_260 : _GEN_1411; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1413 = 10'h105 == _T_5[9:0] ? image_2_261 : _GEN_1412; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1414 = 10'h106 == _T_5[9:0] ? image_2_262 : _GEN_1413; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1415 = 10'h107 == _T_5[9:0] ? image_2_263 : _GEN_1414; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1416 = 10'h108 == _T_5[9:0] ? image_2_264 : _GEN_1415; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1417 = 10'h109 == _T_5[9:0] ? image_2_265 : _GEN_1416; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1418 = 10'h10a == _T_5[9:0] ? image_2_266 : _GEN_1417; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1419 = 10'h10b == _T_5[9:0] ? image_2_267 : _GEN_1418; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1420 = 10'h10c == _T_5[9:0] ? image_2_268 : _GEN_1419; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1421 = 10'h10d == _T_5[9:0] ? image_2_269 : _GEN_1420; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1422 = 10'h10e == _T_5[9:0] ? image_2_270 : _GEN_1421; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1423 = 10'h10f == _T_5[9:0] ? image_2_271 : _GEN_1422; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1424 = 10'h110 == _T_5[9:0] ? image_2_272 : _GEN_1423; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1425 = 10'h111 == _T_5[9:0] ? image_2_273 : _GEN_1424; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1426 = 10'h112 == _T_5[9:0] ? image_2_274 : _GEN_1425; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1427 = 10'h113 == _T_5[9:0] ? image_2_275 : _GEN_1426; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1428 = 10'h114 == _T_5[9:0] ? image_2_276 : _GEN_1427; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1429 = 10'h115 == _T_5[9:0] ? image_2_277 : _GEN_1428; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1430 = 10'h116 == _T_5[9:0] ? image_2_278 : _GEN_1429; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1431 = 10'h117 == _T_5[9:0] ? image_2_279 : _GEN_1430; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1432 = 10'h118 == _T_5[9:0] ? image_2_280 : _GEN_1431; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1433 = 10'h119 == _T_5[9:0] ? image_2_281 : _GEN_1432; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1434 = 10'h11a == _T_5[9:0] ? image_2_282 : _GEN_1433; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1435 = 10'h11b == _T_5[9:0] ? image_2_283 : _GEN_1434; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1436 = 10'h11c == _T_5[9:0] ? image_2_284 : _GEN_1435; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1437 = 10'h11d == _T_5[9:0] ? image_2_285 : _GEN_1436; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1438 = 10'h11e == _T_5[9:0] ? image_2_286 : _GEN_1437; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1439 = 10'h11f == _T_5[9:0] ? image_2_287 : _GEN_1438; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1440 = 10'h120 == _T_5[9:0] ? image_2_288 : _GEN_1439; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1441 = 10'h121 == _T_5[9:0] ? image_2_289 : _GEN_1440; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1442 = 10'h122 == _T_5[9:0] ? image_2_290 : _GEN_1441; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1443 = 10'h123 == _T_5[9:0] ? image_2_291 : _GEN_1442; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1444 = 10'h124 == _T_5[9:0] ? image_2_292 : _GEN_1443; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1445 = 10'h125 == _T_5[9:0] ? image_2_293 : _GEN_1444; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1446 = 10'h126 == _T_5[9:0] ? image_2_294 : _GEN_1445; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1447 = 10'h127 == _T_5[9:0] ? image_2_295 : _GEN_1446; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1448 = 10'h128 == _T_5[9:0] ? image_2_296 : _GEN_1447; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1449 = 10'h129 == _T_5[9:0] ? image_2_297 : _GEN_1448; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1450 = 10'h12a == _T_5[9:0] ? image_2_298 : _GEN_1449; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1451 = 10'h12b == _T_5[9:0] ? image_2_299 : _GEN_1450; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1452 = 10'h12c == _T_5[9:0] ? image_2_300 : _GEN_1451; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1453 = 10'h12d == _T_5[9:0] ? image_2_301 : _GEN_1452; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1454 = 10'h12e == _T_5[9:0] ? image_2_302 : _GEN_1453; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1455 = 10'h12f == _T_5[9:0] ? image_2_303 : _GEN_1454; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1456 = 10'h130 == _T_5[9:0] ? image_2_304 : _GEN_1455; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1457 = 10'h131 == _T_5[9:0] ? image_2_305 : _GEN_1456; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1458 = 10'h132 == _T_5[9:0] ? image_2_306 : _GEN_1457; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1459 = 10'h133 == _T_5[9:0] ? image_2_307 : _GEN_1458; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1460 = 10'h134 == _T_5[9:0] ? image_2_308 : _GEN_1459; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1461 = 10'h135 == _T_5[9:0] ? image_2_309 : _GEN_1460; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1462 = 10'h136 == _T_5[9:0] ? image_2_310 : _GEN_1461; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1463 = 10'h137 == _T_5[9:0] ? image_2_311 : _GEN_1462; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1464 = 10'h138 == _T_5[9:0] ? image_2_312 : _GEN_1463; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1465 = 10'h139 == _T_5[9:0] ? image_2_313 : _GEN_1464; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1466 = 10'h13a == _T_5[9:0] ? image_2_314 : _GEN_1465; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1467 = 10'h13b == _T_5[9:0] ? image_2_315 : _GEN_1466; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1468 = 10'h13c == _T_5[9:0] ? image_2_316 : _GEN_1467; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1469 = 10'h13d == _T_5[9:0] ? image_2_317 : _GEN_1468; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1470 = 10'h13e == _T_5[9:0] ? image_2_318 : _GEN_1469; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1471 = 10'h13f == _T_5[9:0] ? image_2_319 : _GEN_1470; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1472 = 10'h140 == _T_5[9:0] ? image_2_320 : _GEN_1471; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1473 = 10'h141 == _T_5[9:0] ? image_2_321 : _GEN_1472; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1474 = 10'h142 == _T_5[9:0] ? image_2_322 : _GEN_1473; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1475 = 10'h143 == _T_5[9:0] ? image_2_323 : _GEN_1474; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1476 = 10'h144 == _T_5[9:0] ? image_2_324 : _GEN_1475; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1477 = 10'h145 == _T_5[9:0] ? image_2_325 : _GEN_1476; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1478 = 10'h146 == _T_5[9:0] ? image_2_326 : _GEN_1477; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1479 = 10'h147 == _T_5[9:0] ? image_2_327 : _GEN_1478; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1480 = 10'h148 == _T_5[9:0] ? image_2_328 : _GEN_1479; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1481 = 10'h149 == _T_5[9:0] ? image_2_329 : _GEN_1480; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1482 = 10'h14a == _T_5[9:0] ? image_2_330 : _GEN_1481; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1483 = 10'h14b == _T_5[9:0] ? image_2_331 : _GEN_1482; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1484 = 10'h14c == _T_5[9:0] ? image_2_332 : _GEN_1483; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1485 = 10'h14d == _T_5[9:0] ? image_2_333 : _GEN_1484; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1486 = 10'h14e == _T_5[9:0] ? image_2_334 : _GEN_1485; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1487 = 10'h14f == _T_5[9:0] ? image_2_335 : _GEN_1486; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1488 = 10'h150 == _T_5[9:0] ? image_2_336 : _GEN_1487; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1489 = 10'h151 == _T_5[9:0] ? image_2_337 : _GEN_1488; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1490 = 10'h152 == _T_5[9:0] ? image_2_338 : _GEN_1489; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1491 = 10'h153 == _T_5[9:0] ? image_2_339 : _GEN_1490; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1492 = 10'h154 == _T_5[9:0] ? image_2_340 : _GEN_1491; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1493 = 10'h155 == _T_5[9:0] ? image_2_341 : _GEN_1492; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1494 = 10'h156 == _T_5[9:0] ? image_2_342 : _GEN_1493; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1495 = 10'h157 == _T_5[9:0] ? image_2_343 : _GEN_1494; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1496 = 10'h158 == _T_5[9:0] ? image_2_344 : _GEN_1495; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1497 = 10'h159 == _T_5[9:0] ? image_2_345 : _GEN_1496; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1498 = 10'h15a == _T_5[9:0] ? image_2_346 : _GEN_1497; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1499 = 10'h15b == _T_5[9:0] ? image_2_347 : _GEN_1498; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1500 = 10'h15c == _T_5[9:0] ? image_2_348 : _GEN_1499; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1501 = 10'h15d == _T_5[9:0] ? image_2_349 : _GEN_1500; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1502 = 10'h15e == _T_5[9:0] ? image_2_350 : _GEN_1501; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1503 = 10'h15f == _T_5[9:0] ? image_2_351 : _GEN_1502; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1504 = 10'h160 == _T_5[9:0] ? image_2_352 : _GEN_1503; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1505 = 10'h161 == _T_5[9:0] ? image_2_353 : _GEN_1504; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1506 = 10'h162 == _T_5[9:0] ? image_2_354 : _GEN_1505; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1507 = 10'h163 == _T_5[9:0] ? image_2_355 : _GEN_1506; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1508 = 10'h164 == _T_5[9:0] ? image_2_356 : _GEN_1507; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1509 = 10'h165 == _T_5[9:0] ? image_2_357 : _GEN_1508; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1510 = 10'h166 == _T_5[9:0] ? image_2_358 : _GEN_1509; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1511 = 10'h167 == _T_5[9:0] ? image_2_359 : _GEN_1510; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1512 = 10'h168 == _T_5[9:0] ? image_2_360 : _GEN_1511; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1513 = 10'h169 == _T_5[9:0] ? image_2_361 : _GEN_1512; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1514 = 10'h16a == _T_5[9:0] ? image_2_362 : _GEN_1513; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1515 = 10'h16b == _T_5[9:0] ? image_2_363 : _GEN_1514; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1516 = 10'h16c == _T_5[9:0] ? image_2_364 : _GEN_1515; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1517 = 10'h16d == _T_5[9:0] ? image_2_365 : _GEN_1516; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1518 = 10'h16e == _T_5[9:0] ? image_2_366 : _GEN_1517; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1519 = 10'h16f == _T_5[9:0] ? image_2_367 : _GEN_1518; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1520 = 10'h170 == _T_5[9:0] ? image_2_368 : _GEN_1519; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1521 = 10'h171 == _T_5[9:0] ? image_2_369 : _GEN_1520; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1522 = 10'h172 == _T_5[9:0] ? image_2_370 : _GEN_1521; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1523 = 10'h173 == _T_5[9:0] ? image_2_371 : _GEN_1522; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1524 = 10'h174 == _T_5[9:0] ? image_2_372 : _GEN_1523; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1525 = 10'h175 == _T_5[9:0] ? image_2_373 : _GEN_1524; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1526 = 10'h176 == _T_5[9:0] ? image_2_374 : _GEN_1525; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1527 = 10'h177 == _T_5[9:0] ? image_2_375 : _GEN_1526; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1528 = 10'h178 == _T_5[9:0] ? image_2_376 : _GEN_1527; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1529 = 10'h179 == _T_5[9:0] ? image_2_377 : _GEN_1528; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1530 = 10'h17a == _T_5[9:0] ? image_2_378 : _GEN_1529; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1531 = 10'h17b == _T_5[9:0] ? image_2_379 : _GEN_1530; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1532 = 10'h17c == _T_5[9:0] ? image_2_380 : _GEN_1531; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1533 = 10'h17d == _T_5[9:0] ? image_2_381 : _GEN_1532; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1534 = 10'h17e == _T_5[9:0] ? image_2_382 : _GEN_1533; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1535 = 10'h17f == _T_5[9:0] ? image_2_383 : _GEN_1534; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1536 = 10'h180 == _T_5[9:0] ? image_2_384 : _GEN_1535; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1537 = 10'h181 == _T_5[9:0] ? image_2_385 : _GEN_1536; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1538 = 10'h182 == _T_5[9:0] ? image_2_386 : _GEN_1537; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1539 = 10'h183 == _T_5[9:0] ? image_2_387 : _GEN_1538; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1540 = 10'h184 == _T_5[9:0] ? image_2_388 : _GEN_1539; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1541 = 10'h185 == _T_5[9:0] ? image_2_389 : _GEN_1540; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1542 = 10'h186 == _T_5[9:0] ? image_2_390 : _GEN_1541; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1543 = 10'h187 == _T_5[9:0] ? image_2_391 : _GEN_1542; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1544 = 10'h188 == _T_5[9:0] ? image_2_392 : _GEN_1543; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1545 = 10'h189 == _T_5[9:0] ? image_2_393 : _GEN_1544; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1546 = 10'h18a == _T_5[9:0] ? image_2_394 : _GEN_1545; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1547 = 10'h18b == _T_5[9:0] ? image_2_395 : _GEN_1546; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1548 = 10'h18c == _T_5[9:0] ? image_2_396 : _GEN_1547; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1549 = 10'h18d == _T_5[9:0] ? image_2_397 : _GEN_1548; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1550 = 10'h18e == _T_5[9:0] ? image_2_398 : _GEN_1549; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1551 = 10'h18f == _T_5[9:0] ? image_2_399 : _GEN_1550; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1552 = 10'h190 == _T_5[9:0] ? image_2_400 : _GEN_1551; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1553 = 10'h191 == _T_5[9:0] ? image_2_401 : _GEN_1552; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1554 = 10'h192 == _T_5[9:0] ? image_2_402 : _GEN_1553; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1555 = 10'h193 == _T_5[9:0] ? image_2_403 : _GEN_1554; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1556 = 10'h194 == _T_5[9:0] ? image_2_404 : _GEN_1555; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1557 = 10'h195 == _T_5[9:0] ? image_2_405 : _GEN_1556; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1558 = 10'h196 == _T_5[9:0] ? image_2_406 : _GEN_1557; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1559 = 10'h197 == _T_5[9:0] ? image_2_407 : _GEN_1558; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1560 = 10'h198 == _T_5[9:0] ? image_2_408 : _GEN_1559; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1561 = 10'h199 == _T_5[9:0] ? image_2_409 : _GEN_1560; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1562 = 10'h19a == _T_5[9:0] ? image_2_410 : _GEN_1561; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1563 = 10'h19b == _T_5[9:0] ? image_2_411 : _GEN_1562; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1564 = 10'h19c == _T_5[9:0] ? image_2_412 : _GEN_1563; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1565 = 10'h19d == _T_5[9:0] ? image_2_413 : _GEN_1564; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1566 = 10'h19e == _T_5[9:0] ? image_2_414 : _GEN_1565; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1567 = 10'h19f == _T_5[9:0] ? image_2_415 : _GEN_1566; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1568 = 10'h1a0 == _T_5[9:0] ? image_2_416 : _GEN_1567; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1569 = 10'h1a1 == _T_5[9:0] ? image_2_417 : _GEN_1568; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1570 = 10'h1a2 == _T_5[9:0] ? image_2_418 : _GEN_1569; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1571 = 10'h1a3 == _T_5[9:0] ? image_2_419 : _GEN_1570; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1572 = 10'h1a4 == _T_5[9:0] ? image_2_420 : _GEN_1571; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1573 = 10'h1a5 == _T_5[9:0] ? image_2_421 : _GEN_1572; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1574 = 10'h1a6 == _T_5[9:0] ? image_2_422 : _GEN_1573; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1575 = 10'h1a7 == _T_5[9:0] ? image_2_423 : _GEN_1574; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1576 = 10'h1a8 == _T_5[9:0] ? image_2_424 : _GEN_1575; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1577 = 10'h1a9 == _T_5[9:0] ? image_2_425 : _GEN_1576; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1578 = 10'h1aa == _T_5[9:0] ? image_2_426 : _GEN_1577; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1579 = 10'h1ab == _T_5[9:0] ? image_2_427 : _GEN_1578; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1580 = 10'h1ac == _T_5[9:0] ? image_2_428 : _GEN_1579; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1581 = 10'h1ad == _T_5[9:0] ? image_2_429 : _GEN_1580; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1582 = 10'h1ae == _T_5[9:0] ? image_2_430 : _GEN_1581; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1583 = 10'h1af == _T_5[9:0] ? image_2_431 : _GEN_1582; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1584 = 10'h1b0 == _T_5[9:0] ? image_2_432 : _GEN_1583; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1585 = 10'h1b1 == _T_5[9:0] ? image_2_433 : _GEN_1584; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1586 = 10'h1b2 == _T_5[9:0] ? image_2_434 : _GEN_1585; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1587 = 10'h1b3 == _T_5[9:0] ? image_2_435 : _GEN_1586; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1588 = 10'h1b4 == _T_5[9:0] ? image_2_436 : _GEN_1587; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1589 = 10'h1b5 == _T_5[9:0] ? image_2_437 : _GEN_1588; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1590 = 10'h1b6 == _T_5[9:0] ? image_2_438 : _GEN_1589; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1591 = 10'h1b7 == _T_5[9:0] ? image_2_439 : _GEN_1590; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1592 = 10'h1b8 == _T_5[9:0] ? image_2_440 : _GEN_1591; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1593 = 10'h1b9 == _T_5[9:0] ? image_2_441 : _GEN_1592; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1594 = 10'h1ba == _T_5[9:0] ? image_2_442 : _GEN_1593; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1595 = 10'h1bb == _T_5[9:0] ? image_2_443 : _GEN_1594; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1596 = 10'h1bc == _T_5[9:0] ? image_2_444 : _GEN_1595; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1597 = 10'h1bd == _T_5[9:0] ? image_2_445 : _GEN_1596; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1598 = 10'h1be == _T_5[9:0] ? image_2_446 : _GEN_1597; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1599 = 10'h1bf == _T_5[9:0] ? image_2_447 : _GEN_1598; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1600 = 10'h1c0 == _T_5[9:0] ? image_2_448 : _GEN_1599; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1601 = 10'h1c1 == _T_5[9:0] ? image_2_449 : _GEN_1600; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1602 = 10'h1c2 == _T_5[9:0] ? image_2_450 : _GEN_1601; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1603 = 10'h1c3 == _T_5[9:0] ? image_2_451 : _GEN_1602; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1604 = 10'h1c4 == _T_5[9:0] ? image_2_452 : _GEN_1603; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1605 = 10'h1c5 == _T_5[9:0] ? image_2_453 : _GEN_1604; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1606 = 10'h1c6 == _T_5[9:0] ? image_2_454 : _GEN_1605; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1607 = 10'h1c7 == _T_5[9:0] ? image_2_455 : _GEN_1606; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1608 = 10'h1c8 == _T_5[9:0] ? image_2_456 : _GEN_1607; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1609 = 10'h1c9 == _T_5[9:0] ? image_2_457 : _GEN_1608; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1610 = 10'h1ca == _T_5[9:0] ? image_2_458 : _GEN_1609; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1611 = 10'h1cb == _T_5[9:0] ? image_2_459 : _GEN_1610; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1612 = 10'h1cc == _T_5[9:0] ? image_2_460 : _GEN_1611; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1613 = 10'h1cd == _T_5[9:0] ? image_2_461 : _GEN_1612; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1614 = 10'h1ce == _T_5[9:0] ? image_2_462 : _GEN_1613; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1615 = 10'h1cf == _T_5[9:0] ? image_2_463 : _GEN_1614; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1616 = 10'h1d0 == _T_5[9:0] ? image_2_464 : _GEN_1615; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1617 = 10'h1d1 == _T_5[9:0] ? image_2_465 : _GEN_1616; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1618 = 10'h1d2 == _T_5[9:0] ? image_2_466 : _GEN_1617; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1619 = 10'h1d3 == _T_5[9:0] ? image_2_467 : _GEN_1618; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1620 = 10'h1d4 == _T_5[9:0] ? image_2_468 : _GEN_1619; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1621 = 10'h1d5 == _T_5[9:0] ? image_2_469 : _GEN_1620; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1622 = 10'h1d6 == _T_5[9:0] ? image_2_470 : _GEN_1621; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1623 = 10'h1d7 == _T_5[9:0] ? image_2_471 : _GEN_1622; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1624 = 10'h1d8 == _T_5[9:0] ? image_2_472 : _GEN_1623; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1625 = 10'h1d9 == _T_5[9:0] ? image_2_473 : _GEN_1624; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1626 = 10'h1da == _T_5[9:0] ? image_2_474 : _GEN_1625; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1627 = 10'h1db == _T_5[9:0] ? image_2_475 : _GEN_1626; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1628 = 10'h1dc == _T_5[9:0] ? image_2_476 : _GEN_1627; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1629 = 10'h1dd == _T_5[9:0] ? image_2_477 : _GEN_1628; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1630 = 10'h1de == _T_5[9:0] ? image_2_478 : _GEN_1629; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1631 = 10'h1df == _T_5[9:0] ? image_2_479 : _GEN_1630; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1632 = 10'h1e0 == _T_5[9:0] ? image_2_480 : _GEN_1631; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1633 = 10'h1e1 == _T_5[9:0] ? image_2_481 : _GEN_1632; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1634 = 10'h1e2 == _T_5[9:0] ? image_2_482 : _GEN_1633; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1635 = 10'h1e3 == _T_5[9:0] ? image_2_483 : _GEN_1634; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1636 = 10'h1e4 == _T_5[9:0] ? image_2_484 : _GEN_1635; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1637 = 10'h1e5 == _T_5[9:0] ? image_2_485 : _GEN_1636; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1638 = 10'h1e6 == _T_5[9:0] ? image_2_486 : _GEN_1637; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1639 = 10'h1e7 == _T_5[9:0] ? image_2_487 : _GEN_1638; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1640 = 10'h1e8 == _T_5[9:0] ? image_2_488 : _GEN_1639; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1641 = 10'h1e9 == _T_5[9:0] ? image_2_489 : _GEN_1640; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1642 = 10'h1ea == _T_5[9:0] ? image_2_490 : _GEN_1641; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1643 = 10'h1eb == _T_5[9:0] ? image_2_491 : _GEN_1642; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1644 = 10'h1ec == _T_5[9:0] ? image_2_492 : _GEN_1643; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1645 = 10'h1ed == _T_5[9:0] ? image_2_493 : _GEN_1644; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1646 = 10'h1ee == _T_5[9:0] ? image_2_494 : _GEN_1645; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1647 = 10'h1ef == _T_5[9:0] ? image_2_495 : _GEN_1646; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1648 = 10'h1f0 == _T_5[9:0] ? image_2_496 : _GEN_1647; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1649 = 10'h1f1 == _T_5[9:0] ? image_2_497 : _GEN_1648; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1650 = 10'h1f2 == _T_5[9:0] ? image_2_498 : _GEN_1649; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1651 = 10'h1f3 == _T_5[9:0] ? image_2_499 : _GEN_1650; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1652 = 10'h1f4 == _T_5[9:0] ? image_2_500 : _GEN_1651; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1653 = 10'h1f5 == _T_5[9:0] ? image_2_501 : _GEN_1652; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1654 = 10'h1f6 == _T_5[9:0] ? image_2_502 : _GEN_1653; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1655 = 10'h1f7 == _T_5[9:0] ? image_2_503 : _GEN_1654; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1656 = 10'h1f8 == _T_5[9:0] ? image_2_504 : _GEN_1655; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1657 = 10'h1f9 == _T_5[9:0] ? image_2_505 : _GEN_1656; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1658 = 10'h1fa == _T_5[9:0] ? image_2_506 : _GEN_1657; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1659 = 10'h1fb == _T_5[9:0] ? image_2_507 : _GEN_1658; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1660 = 10'h1fc == _T_5[9:0] ? image_2_508 : _GEN_1659; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1661 = 10'h1fd == _T_5[9:0] ? image_2_509 : _GEN_1660; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1662 = 10'h1fe == _T_5[9:0] ? image_2_510 : _GEN_1661; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1663 = 10'h1ff == _T_5[9:0] ? image_2_511 : _GEN_1662; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1664 = 10'h200 == _T_5[9:0] ? image_2_512 : _GEN_1663; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1665 = 10'h201 == _T_5[9:0] ? image_2_513 : _GEN_1664; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1666 = 10'h202 == _T_5[9:0] ? image_2_514 : _GEN_1665; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1667 = 10'h203 == _T_5[9:0] ? image_2_515 : _GEN_1666; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1668 = 10'h204 == _T_5[9:0] ? image_2_516 : _GEN_1667; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1669 = 10'h205 == _T_5[9:0] ? image_2_517 : _GEN_1668; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1670 = 10'h206 == _T_5[9:0] ? image_2_518 : _GEN_1669; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1671 = 10'h207 == _T_5[9:0] ? image_2_519 : _GEN_1670; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1672 = 10'h208 == _T_5[9:0] ? image_2_520 : _GEN_1671; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1673 = 10'h209 == _T_5[9:0] ? image_2_521 : _GEN_1672; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1674 = 10'h20a == _T_5[9:0] ? image_2_522 : _GEN_1673; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1675 = 10'h20b == _T_5[9:0] ? image_2_523 : _GEN_1674; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1676 = 10'h20c == _T_5[9:0] ? image_2_524 : _GEN_1675; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1677 = 10'h20d == _T_5[9:0] ? image_2_525 : _GEN_1676; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1678 = 10'h20e == _T_5[9:0] ? image_2_526 : _GEN_1677; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1679 = 10'h20f == _T_5[9:0] ? image_2_527 : _GEN_1678; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1680 = 10'h210 == _T_5[9:0] ? image_2_528 : _GEN_1679; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1681 = 10'h211 == _T_5[9:0] ? image_2_529 : _GEN_1680; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1682 = 10'h212 == _T_5[9:0] ? image_2_530 : _GEN_1681; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1683 = 10'h213 == _T_5[9:0] ? image_2_531 : _GEN_1682; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1684 = 10'h214 == _T_5[9:0] ? image_2_532 : _GEN_1683; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1685 = 10'h215 == _T_5[9:0] ? image_2_533 : _GEN_1684; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1686 = 10'h216 == _T_5[9:0] ? image_2_534 : _GEN_1685; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1687 = 10'h217 == _T_5[9:0] ? image_2_535 : _GEN_1686; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1688 = 10'h218 == _T_5[9:0] ? image_2_536 : _GEN_1687; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1689 = 10'h219 == _T_5[9:0] ? image_2_537 : _GEN_1688; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1690 = 10'h21a == _T_5[9:0] ? image_2_538 : _GEN_1689; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1691 = 10'h21b == _T_5[9:0] ? image_2_539 : _GEN_1690; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1692 = 10'h21c == _T_5[9:0] ? image_2_540 : _GEN_1691; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1693 = 10'h21d == _T_5[9:0] ? image_2_541 : _GEN_1692; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1694 = 10'h21e == _T_5[9:0] ? image_2_542 : _GEN_1693; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1695 = 10'h21f == _T_5[9:0] ? image_2_543 : _GEN_1694; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1696 = 10'h220 == _T_5[9:0] ? image_2_544 : _GEN_1695; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1697 = 10'h221 == _T_5[9:0] ? image_2_545 : _GEN_1696; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1698 = 10'h222 == _T_5[9:0] ? image_2_546 : _GEN_1697; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1699 = 10'h223 == _T_5[9:0] ? image_2_547 : _GEN_1698; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1700 = 10'h224 == _T_5[9:0] ? image_2_548 : _GEN_1699; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1701 = 10'h225 == _T_5[9:0] ? image_2_549 : _GEN_1700; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1702 = 10'h226 == _T_5[9:0] ? image_2_550 : _GEN_1701; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1703 = 10'h227 == _T_5[9:0] ? image_2_551 : _GEN_1702; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1704 = 10'h228 == _T_5[9:0] ? image_2_552 : _GEN_1703; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1705 = 10'h229 == _T_5[9:0] ? image_2_553 : _GEN_1704; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1706 = 10'h22a == _T_5[9:0] ? image_2_554 : _GEN_1705; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1707 = 10'h22b == _T_5[9:0] ? image_2_555 : _GEN_1706; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1708 = 10'h22c == _T_5[9:0] ? image_2_556 : _GEN_1707; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1709 = 10'h22d == _T_5[9:0] ? image_2_557 : _GEN_1708; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1710 = 10'h22e == _T_5[9:0] ? image_2_558 : _GEN_1709; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1711 = 10'h22f == _T_5[9:0] ? image_2_559 : _GEN_1710; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1712 = 10'h230 == _T_5[9:0] ? image_2_560 : _GEN_1711; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1713 = 10'h231 == _T_5[9:0] ? image_2_561 : _GEN_1712; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1714 = 10'h232 == _T_5[9:0] ? image_2_562 : _GEN_1713; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1715 = 10'h233 == _T_5[9:0] ? image_2_563 : _GEN_1714; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1716 = 10'h234 == _T_5[9:0] ? image_2_564 : _GEN_1715; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1717 = 10'h235 == _T_5[9:0] ? image_2_565 : _GEN_1716; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1718 = 10'h236 == _T_5[9:0] ? image_2_566 : _GEN_1717; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1719 = 10'h237 == _T_5[9:0] ? image_2_567 : _GEN_1718; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1720 = 10'h238 == _T_5[9:0] ? image_2_568 : _GEN_1719; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1721 = 10'h239 == _T_5[9:0] ? image_2_569 : _GEN_1720; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1722 = 10'h23a == _T_5[9:0] ? image_2_570 : _GEN_1721; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1723 = 10'h23b == _T_5[9:0] ? image_2_571 : _GEN_1722; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1724 = 10'h23c == _T_5[9:0] ? image_2_572 : _GEN_1723; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1725 = 10'h23d == _T_5[9:0] ? image_2_573 : _GEN_1724; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1726 = 10'h23e == _T_5[9:0] ? image_2_574 : _GEN_1725; // @[VideoBuffer.scala 27:30]
  wire [32:0] _T_15 = {{1'd0}, pixelIndex}; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_19 = pixelIndex + 32'h1; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_22 = pixelIndex + 32'h2; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_25 = pixelIndex + 32'h3; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_28 = pixelIndex + 32'h4; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_31 = pixelIndex + 32'h5; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_34 = pixelIndex + 32'h6; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_37 = pixelIndex + 32'h7; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_88 = pixelIndex + 32'h8; // @[VideoBuffer.scala 36:34]
  wire [10:0] _T_89 = 6'h20 * 6'h12; // @[VideoBuffer.scala 37:42]
  wire [31:0] _GEN_17285 = {{21'd0}, _T_89}; // @[VideoBuffer.scala 37:25]
  wire  _T_90 = pixelIndex == _GEN_17285; // @[VideoBuffer.scala 37:25]
  assign io_pixelVal_out_0 = 10'h23f == _T_5[9:0] ? image_0_575 : _GEN_574; // @[VideoBuffer.scala 27:30]
  assign io_pixelVal_out_1 = 10'h23f == _T_5[9:0] ? image_1_575 : _GEN_1150; // @[VideoBuffer.scala 27:30]
  assign io_pixelVal_out_2 = 10'h23f == _T_5[9:0] ? image_2_575 : _GEN_1726; // @[VideoBuffer.scala 27:30]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  image_0_0 = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  image_0_1 = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  image_0_2 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  image_0_3 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  image_0_4 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  image_0_5 = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  image_0_6 = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  image_0_7 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  image_0_8 = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  image_0_9 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  image_0_10 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  image_0_11 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  image_0_12 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  image_0_13 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  image_0_14 = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  image_0_15 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  image_0_16 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  image_0_17 = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  image_0_18 = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  image_0_19 = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  image_0_20 = _RAND_20[3:0];
  _RAND_21 = {1{`RANDOM}};
  image_0_21 = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  image_0_22 = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  image_0_23 = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  image_0_24 = _RAND_24[3:0];
  _RAND_25 = {1{`RANDOM}};
  image_0_25 = _RAND_25[3:0];
  _RAND_26 = {1{`RANDOM}};
  image_0_26 = _RAND_26[3:0];
  _RAND_27 = {1{`RANDOM}};
  image_0_27 = _RAND_27[3:0];
  _RAND_28 = {1{`RANDOM}};
  image_0_28 = _RAND_28[3:0];
  _RAND_29 = {1{`RANDOM}};
  image_0_29 = _RAND_29[3:0];
  _RAND_30 = {1{`RANDOM}};
  image_0_30 = _RAND_30[3:0];
  _RAND_31 = {1{`RANDOM}};
  image_0_31 = _RAND_31[3:0];
  _RAND_32 = {1{`RANDOM}};
  image_0_32 = _RAND_32[3:0];
  _RAND_33 = {1{`RANDOM}};
  image_0_33 = _RAND_33[3:0];
  _RAND_34 = {1{`RANDOM}};
  image_0_34 = _RAND_34[3:0];
  _RAND_35 = {1{`RANDOM}};
  image_0_35 = _RAND_35[3:0];
  _RAND_36 = {1{`RANDOM}};
  image_0_36 = _RAND_36[3:0];
  _RAND_37 = {1{`RANDOM}};
  image_0_37 = _RAND_37[3:0];
  _RAND_38 = {1{`RANDOM}};
  image_0_38 = _RAND_38[3:0];
  _RAND_39 = {1{`RANDOM}};
  image_0_39 = _RAND_39[3:0];
  _RAND_40 = {1{`RANDOM}};
  image_0_40 = _RAND_40[3:0];
  _RAND_41 = {1{`RANDOM}};
  image_0_41 = _RAND_41[3:0];
  _RAND_42 = {1{`RANDOM}};
  image_0_42 = _RAND_42[3:0];
  _RAND_43 = {1{`RANDOM}};
  image_0_43 = _RAND_43[3:0];
  _RAND_44 = {1{`RANDOM}};
  image_0_44 = _RAND_44[3:0];
  _RAND_45 = {1{`RANDOM}};
  image_0_45 = _RAND_45[3:0];
  _RAND_46 = {1{`RANDOM}};
  image_0_46 = _RAND_46[3:0];
  _RAND_47 = {1{`RANDOM}};
  image_0_47 = _RAND_47[3:0];
  _RAND_48 = {1{`RANDOM}};
  image_0_48 = _RAND_48[3:0];
  _RAND_49 = {1{`RANDOM}};
  image_0_49 = _RAND_49[3:0];
  _RAND_50 = {1{`RANDOM}};
  image_0_50 = _RAND_50[3:0];
  _RAND_51 = {1{`RANDOM}};
  image_0_51 = _RAND_51[3:0];
  _RAND_52 = {1{`RANDOM}};
  image_0_52 = _RAND_52[3:0];
  _RAND_53 = {1{`RANDOM}};
  image_0_53 = _RAND_53[3:0];
  _RAND_54 = {1{`RANDOM}};
  image_0_54 = _RAND_54[3:0];
  _RAND_55 = {1{`RANDOM}};
  image_0_55 = _RAND_55[3:0];
  _RAND_56 = {1{`RANDOM}};
  image_0_56 = _RAND_56[3:0];
  _RAND_57 = {1{`RANDOM}};
  image_0_57 = _RAND_57[3:0];
  _RAND_58 = {1{`RANDOM}};
  image_0_58 = _RAND_58[3:0];
  _RAND_59 = {1{`RANDOM}};
  image_0_59 = _RAND_59[3:0];
  _RAND_60 = {1{`RANDOM}};
  image_0_60 = _RAND_60[3:0];
  _RAND_61 = {1{`RANDOM}};
  image_0_61 = _RAND_61[3:0];
  _RAND_62 = {1{`RANDOM}};
  image_0_62 = _RAND_62[3:0];
  _RAND_63 = {1{`RANDOM}};
  image_0_63 = _RAND_63[3:0];
  _RAND_64 = {1{`RANDOM}};
  image_0_64 = _RAND_64[3:0];
  _RAND_65 = {1{`RANDOM}};
  image_0_65 = _RAND_65[3:0];
  _RAND_66 = {1{`RANDOM}};
  image_0_66 = _RAND_66[3:0];
  _RAND_67 = {1{`RANDOM}};
  image_0_67 = _RAND_67[3:0];
  _RAND_68 = {1{`RANDOM}};
  image_0_68 = _RAND_68[3:0];
  _RAND_69 = {1{`RANDOM}};
  image_0_69 = _RAND_69[3:0];
  _RAND_70 = {1{`RANDOM}};
  image_0_70 = _RAND_70[3:0];
  _RAND_71 = {1{`RANDOM}};
  image_0_71 = _RAND_71[3:0];
  _RAND_72 = {1{`RANDOM}};
  image_0_72 = _RAND_72[3:0];
  _RAND_73 = {1{`RANDOM}};
  image_0_73 = _RAND_73[3:0];
  _RAND_74 = {1{`RANDOM}};
  image_0_74 = _RAND_74[3:0];
  _RAND_75 = {1{`RANDOM}};
  image_0_75 = _RAND_75[3:0];
  _RAND_76 = {1{`RANDOM}};
  image_0_76 = _RAND_76[3:0];
  _RAND_77 = {1{`RANDOM}};
  image_0_77 = _RAND_77[3:0];
  _RAND_78 = {1{`RANDOM}};
  image_0_78 = _RAND_78[3:0];
  _RAND_79 = {1{`RANDOM}};
  image_0_79 = _RAND_79[3:0];
  _RAND_80 = {1{`RANDOM}};
  image_0_80 = _RAND_80[3:0];
  _RAND_81 = {1{`RANDOM}};
  image_0_81 = _RAND_81[3:0];
  _RAND_82 = {1{`RANDOM}};
  image_0_82 = _RAND_82[3:0];
  _RAND_83 = {1{`RANDOM}};
  image_0_83 = _RAND_83[3:0];
  _RAND_84 = {1{`RANDOM}};
  image_0_84 = _RAND_84[3:0];
  _RAND_85 = {1{`RANDOM}};
  image_0_85 = _RAND_85[3:0];
  _RAND_86 = {1{`RANDOM}};
  image_0_86 = _RAND_86[3:0];
  _RAND_87 = {1{`RANDOM}};
  image_0_87 = _RAND_87[3:0];
  _RAND_88 = {1{`RANDOM}};
  image_0_88 = _RAND_88[3:0];
  _RAND_89 = {1{`RANDOM}};
  image_0_89 = _RAND_89[3:0];
  _RAND_90 = {1{`RANDOM}};
  image_0_90 = _RAND_90[3:0];
  _RAND_91 = {1{`RANDOM}};
  image_0_91 = _RAND_91[3:0];
  _RAND_92 = {1{`RANDOM}};
  image_0_92 = _RAND_92[3:0];
  _RAND_93 = {1{`RANDOM}};
  image_0_93 = _RAND_93[3:0];
  _RAND_94 = {1{`RANDOM}};
  image_0_94 = _RAND_94[3:0];
  _RAND_95 = {1{`RANDOM}};
  image_0_95 = _RAND_95[3:0];
  _RAND_96 = {1{`RANDOM}};
  image_0_96 = _RAND_96[3:0];
  _RAND_97 = {1{`RANDOM}};
  image_0_97 = _RAND_97[3:0];
  _RAND_98 = {1{`RANDOM}};
  image_0_98 = _RAND_98[3:0];
  _RAND_99 = {1{`RANDOM}};
  image_0_99 = _RAND_99[3:0];
  _RAND_100 = {1{`RANDOM}};
  image_0_100 = _RAND_100[3:0];
  _RAND_101 = {1{`RANDOM}};
  image_0_101 = _RAND_101[3:0];
  _RAND_102 = {1{`RANDOM}};
  image_0_102 = _RAND_102[3:0];
  _RAND_103 = {1{`RANDOM}};
  image_0_103 = _RAND_103[3:0];
  _RAND_104 = {1{`RANDOM}};
  image_0_104 = _RAND_104[3:0];
  _RAND_105 = {1{`RANDOM}};
  image_0_105 = _RAND_105[3:0];
  _RAND_106 = {1{`RANDOM}};
  image_0_106 = _RAND_106[3:0];
  _RAND_107 = {1{`RANDOM}};
  image_0_107 = _RAND_107[3:0];
  _RAND_108 = {1{`RANDOM}};
  image_0_108 = _RAND_108[3:0];
  _RAND_109 = {1{`RANDOM}};
  image_0_109 = _RAND_109[3:0];
  _RAND_110 = {1{`RANDOM}};
  image_0_110 = _RAND_110[3:0];
  _RAND_111 = {1{`RANDOM}};
  image_0_111 = _RAND_111[3:0];
  _RAND_112 = {1{`RANDOM}};
  image_0_112 = _RAND_112[3:0];
  _RAND_113 = {1{`RANDOM}};
  image_0_113 = _RAND_113[3:0];
  _RAND_114 = {1{`RANDOM}};
  image_0_114 = _RAND_114[3:0];
  _RAND_115 = {1{`RANDOM}};
  image_0_115 = _RAND_115[3:0];
  _RAND_116 = {1{`RANDOM}};
  image_0_116 = _RAND_116[3:0];
  _RAND_117 = {1{`RANDOM}};
  image_0_117 = _RAND_117[3:0];
  _RAND_118 = {1{`RANDOM}};
  image_0_118 = _RAND_118[3:0];
  _RAND_119 = {1{`RANDOM}};
  image_0_119 = _RAND_119[3:0];
  _RAND_120 = {1{`RANDOM}};
  image_0_120 = _RAND_120[3:0];
  _RAND_121 = {1{`RANDOM}};
  image_0_121 = _RAND_121[3:0];
  _RAND_122 = {1{`RANDOM}};
  image_0_122 = _RAND_122[3:0];
  _RAND_123 = {1{`RANDOM}};
  image_0_123 = _RAND_123[3:0];
  _RAND_124 = {1{`RANDOM}};
  image_0_124 = _RAND_124[3:0];
  _RAND_125 = {1{`RANDOM}};
  image_0_125 = _RAND_125[3:0];
  _RAND_126 = {1{`RANDOM}};
  image_0_126 = _RAND_126[3:0];
  _RAND_127 = {1{`RANDOM}};
  image_0_127 = _RAND_127[3:0];
  _RAND_128 = {1{`RANDOM}};
  image_0_128 = _RAND_128[3:0];
  _RAND_129 = {1{`RANDOM}};
  image_0_129 = _RAND_129[3:0];
  _RAND_130 = {1{`RANDOM}};
  image_0_130 = _RAND_130[3:0];
  _RAND_131 = {1{`RANDOM}};
  image_0_131 = _RAND_131[3:0];
  _RAND_132 = {1{`RANDOM}};
  image_0_132 = _RAND_132[3:0];
  _RAND_133 = {1{`RANDOM}};
  image_0_133 = _RAND_133[3:0];
  _RAND_134 = {1{`RANDOM}};
  image_0_134 = _RAND_134[3:0];
  _RAND_135 = {1{`RANDOM}};
  image_0_135 = _RAND_135[3:0];
  _RAND_136 = {1{`RANDOM}};
  image_0_136 = _RAND_136[3:0];
  _RAND_137 = {1{`RANDOM}};
  image_0_137 = _RAND_137[3:0];
  _RAND_138 = {1{`RANDOM}};
  image_0_138 = _RAND_138[3:0];
  _RAND_139 = {1{`RANDOM}};
  image_0_139 = _RAND_139[3:0];
  _RAND_140 = {1{`RANDOM}};
  image_0_140 = _RAND_140[3:0];
  _RAND_141 = {1{`RANDOM}};
  image_0_141 = _RAND_141[3:0];
  _RAND_142 = {1{`RANDOM}};
  image_0_142 = _RAND_142[3:0];
  _RAND_143 = {1{`RANDOM}};
  image_0_143 = _RAND_143[3:0];
  _RAND_144 = {1{`RANDOM}};
  image_0_144 = _RAND_144[3:0];
  _RAND_145 = {1{`RANDOM}};
  image_0_145 = _RAND_145[3:0];
  _RAND_146 = {1{`RANDOM}};
  image_0_146 = _RAND_146[3:0];
  _RAND_147 = {1{`RANDOM}};
  image_0_147 = _RAND_147[3:0];
  _RAND_148 = {1{`RANDOM}};
  image_0_148 = _RAND_148[3:0];
  _RAND_149 = {1{`RANDOM}};
  image_0_149 = _RAND_149[3:0];
  _RAND_150 = {1{`RANDOM}};
  image_0_150 = _RAND_150[3:0];
  _RAND_151 = {1{`RANDOM}};
  image_0_151 = _RAND_151[3:0];
  _RAND_152 = {1{`RANDOM}};
  image_0_152 = _RAND_152[3:0];
  _RAND_153 = {1{`RANDOM}};
  image_0_153 = _RAND_153[3:0];
  _RAND_154 = {1{`RANDOM}};
  image_0_154 = _RAND_154[3:0];
  _RAND_155 = {1{`RANDOM}};
  image_0_155 = _RAND_155[3:0];
  _RAND_156 = {1{`RANDOM}};
  image_0_156 = _RAND_156[3:0];
  _RAND_157 = {1{`RANDOM}};
  image_0_157 = _RAND_157[3:0];
  _RAND_158 = {1{`RANDOM}};
  image_0_158 = _RAND_158[3:0];
  _RAND_159 = {1{`RANDOM}};
  image_0_159 = _RAND_159[3:0];
  _RAND_160 = {1{`RANDOM}};
  image_0_160 = _RAND_160[3:0];
  _RAND_161 = {1{`RANDOM}};
  image_0_161 = _RAND_161[3:0];
  _RAND_162 = {1{`RANDOM}};
  image_0_162 = _RAND_162[3:0];
  _RAND_163 = {1{`RANDOM}};
  image_0_163 = _RAND_163[3:0];
  _RAND_164 = {1{`RANDOM}};
  image_0_164 = _RAND_164[3:0];
  _RAND_165 = {1{`RANDOM}};
  image_0_165 = _RAND_165[3:0];
  _RAND_166 = {1{`RANDOM}};
  image_0_166 = _RAND_166[3:0];
  _RAND_167 = {1{`RANDOM}};
  image_0_167 = _RAND_167[3:0];
  _RAND_168 = {1{`RANDOM}};
  image_0_168 = _RAND_168[3:0];
  _RAND_169 = {1{`RANDOM}};
  image_0_169 = _RAND_169[3:0];
  _RAND_170 = {1{`RANDOM}};
  image_0_170 = _RAND_170[3:0];
  _RAND_171 = {1{`RANDOM}};
  image_0_171 = _RAND_171[3:0];
  _RAND_172 = {1{`RANDOM}};
  image_0_172 = _RAND_172[3:0];
  _RAND_173 = {1{`RANDOM}};
  image_0_173 = _RAND_173[3:0];
  _RAND_174 = {1{`RANDOM}};
  image_0_174 = _RAND_174[3:0];
  _RAND_175 = {1{`RANDOM}};
  image_0_175 = _RAND_175[3:0];
  _RAND_176 = {1{`RANDOM}};
  image_0_176 = _RAND_176[3:0];
  _RAND_177 = {1{`RANDOM}};
  image_0_177 = _RAND_177[3:0];
  _RAND_178 = {1{`RANDOM}};
  image_0_178 = _RAND_178[3:0];
  _RAND_179 = {1{`RANDOM}};
  image_0_179 = _RAND_179[3:0];
  _RAND_180 = {1{`RANDOM}};
  image_0_180 = _RAND_180[3:0];
  _RAND_181 = {1{`RANDOM}};
  image_0_181 = _RAND_181[3:0];
  _RAND_182 = {1{`RANDOM}};
  image_0_182 = _RAND_182[3:0];
  _RAND_183 = {1{`RANDOM}};
  image_0_183 = _RAND_183[3:0];
  _RAND_184 = {1{`RANDOM}};
  image_0_184 = _RAND_184[3:0];
  _RAND_185 = {1{`RANDOM}};
  image_0_185 = _RAND_185[3:0];
  _RAND_186 = {1{`RANDOM}};
  image_0_186 = _RAND_186[3:0];
  _RAND_187 = {1{`RANDOM}};
  image_0_187 = _RAND_187[3:0];
  _RAND_188 = {1{`RANDOM}};
  image_0_188 = _RAND_188[3:0];
  _RAND_189 = {1{`RANDOM}};
  image_0_189 = _RAND_189[3:0];
  _RAND_190 = {1{`RANDOM}};
  image_0_190 = _RAND_190[3:0];
  _RAND_191 = {1{`RANDOM}};
  image_0_191 = _RAND_191[3:0];
  _RAND_192 = {1{`RANDOM}};
  image_0_192 = _RAND_192[3:0];
  _RAND_193 = {1{`RANDOM}};
  image_0_193 = _RAND_193[3:0];
  _RAND_194 = {1{`RANDOM}};
  image_0_194 = _RAND_194[3:0];
  _RAND_195 = {1{`RANDOM}};
  image_0_195 = _RAND_195[3:0];
  _RAND_196 = {1{`RANDOM}};
  image_0_196 = _RAND_196[3:0];
  _RAND_197 = {1{`RANDOM}};
  image_0_197 = _RAND_197[3:0];
  _RAND_198 = {1{`RANDOM}};
  image_0_198 = _RAND_198[3:0];
  _RAND_199 = {1{`RANDOM}};
  image_0_199 = _RAND_199[3:0];
  _RAND_200 = {1{`RANDOM}};
  image_0_200 = _RAND_200[3:0];
  _RAND_201 = {1{`RANDOM}};
  image_0_201 = _RAND_201[3:0];
  _RAND_202 = {1{`RANDOM}};
  image_0_202 = _RAND_202[3:0];
  _RAND_203 = {1{`RANDOM}};
  image_0_203 = _RAND_203[3:0];
  _RAND_204 = {1{`RANDOM}};
  image_0_204 = _RAND_204[3:0];
  _RAND_205 = {1{`RANDOM}};
  image_0_205 = _RAND_205[3:0];
  _RAND_206 = {1{`RANDOM}};
  image_0_206 = _RAND_206[3:0];
  _RAND_207 = {1{`RANDOM}};
  image_0_207 = _RAND_207[3:0];
  _RAND_208 = {1{`RANDOM}};
  image_0_208 = _RAND_208[3:0];
  _RAND_209 = {1{`RANDOM}};
  image_0_209 = _RAND_209[3:0];
  _RAND_210 = {1{`RANDOM}};
  image_0_210 = _RAND_210[3:0];
  _RAND_211 = {1{`RANDOM}};
  image_0_211 = _RAND_211[3:0];
  _RAND_212 = {1{`RANDOM}};
  image_0_212 = _RAND_212[3:0];
  _RAND_213 = {1{`RANDOM}};
  image_0_213 = _RAND_213[3:0];
  _RAND_214 = {1{`RANDOM}};
  image_0_214 = _RAND_214[3:0];
  _RAND_215 = {1{`RANDOM}};
  image_0_215 = _RAND_215[3:0];
  _RAND_216 = {1{`RANDOM}};
  image_0_216 = _RAND_216[3:0];
  _RAND_217 = {1{`RANDOM}};
  image_0_217 = _RAND_217[3:0];
  _RAND_218 = {1{`RANDOM}};
  image_0_218 = _RAND_218[3:0];
  _RAND_219 = {1{`RANDOM}};
  image_0_219 = _RAND_219[3:0];
  _RAND_220 = {1{`RANDOM}};
  image_0_220 = _RAND_220[3:0];
  _RAND_221 = {1{`RANDOM}};
  image_0_221 = _RAND_221[3:0];
  _RAND_222 = {1{`RANDOM}};
  image_0_222 = _RAND_222[3:0];
  _RAND_223 = {1{`RANDOM}};
  image_0_223 = _RAND_223[3:0];
  _RAND_224 = {1{`RANDOM}};
  image_0_224 = _RAND_224[3:0];
  _RAND_225 = {1{`RANDOM}};
  image_0_225 = _RAND_225[3:0];
  _RAND_226 = {1{`RANDOM}};
  image_0_226 = _RAND_226[3:0];
  _RAND_227 = {1{`RANDOM}};
  image_0_227 = _RAND_227[3:0];
  _RAND_228 = {1{`RANDOM}};
  image_0_228 = _RAND_228[3:0];
  _RAND_229 = {1{`RANDOM}};
  image_0_229 = _RAND_229[3:0];
  _RAND_230 = {1{`RANDOM}};
  image_0_230 = _RAND_230[3:0];
  _RAND_231 = {1{`RANDOM}};
  image_0_231 = _RAND_231[3:0];
  _RAND_232 = {1{`RANDOM}};
  image_0_232 = _RAND_232[3:0];
  _RAND_233 = {1{`RANDOM}};
  image_0_233 = _RAND_233[3:0];
  _RAND_234 = {1{`RANDOM}};
  image_0_234 = _RAND_234[3:0];
  _RAND_235 = {1{`RANDOM}};
  image_0_235 = _RAND_235[3:0];
  _RAND_236 = {1{`RANDOM}};
  image_0_236 = _RAND_236[3:0];
  _RAND_237 = {1{`RANDOM}};
  image_0_237 = _RAND_237[3:0];
  _RAND_238 = {1{`RANDOM}};
  image_0_238 = _RAND_238[3:0];
  _RAND_239 = {1{`RANDOM}};
  image_0_239 = _RAND_239[3:0];
  _RAND_240 = {1{`RANDOM}};
  image_0_240 = _RAND_240[3:0];
  _RAND_241 = {1{`RANDOM}};
  image_0_241 = _RAND_241[3:0];
  _RAND_242 = {1{`RANDOM}};
  image_0_242 = _RAND_242[3:0];
  _RAND_243 = {1{`RANDOM}};
  image_0_243 = _RAND_243[3:0];
  _RAND_244 = {1{`RANDOM}};
  image_0_244 = _RAND_244[3:0];
  _RAND_245 = {1{`RANDOM}};
  image_0_245 = _RAND_245[3:0];
  _RAND_246 = {1{`RANDOM}};
  image_0_246 = _RAND_246[3:0];
  _RAND_247 = {1{`RANDOM}};
  image_0_247 = _RAND_247[3:0];
  _RAND_248 = {1{`RANDOM}};
  image_0_248 = _RAND_248[3:0];
  _RAND_249 = {1{`RANDOM}};
  image_0_249 = _RAND_249[3:0];
  _RAND_250 = {1{`RANDOM}};
  image_0_250 = _RAND_250[3:0];
  _RAND_251 = {1{`RANDOM}};
  image_0_251 = _RAND_251[3:0];
  _RAND_252 = {1{`RANDOM}};
  image_0_252 = _RAND_252[3:0];
  _RAND_253 = {1{`RANDOM}};
  image_0_253 = _RAND_253[3:0];
  _RAND_254 = {1{`RANDOM}};
  image_0_254 = _RAND_254[3:0];
  _RAND_255 = {1{`RANDOM}};
  image_0_255 = _RAND_255[3:0];
  _RAND_256 = {1{`RANDOM}};
  image_0_256 = _RAND_256[3:0];
  _RAND_257 = {1{`RANDOM}};
  image_0_257 = _RAND_257[3:0];
  _RAND_258 = {1{`RANDOM}};
  image_0_258 = _RAND_258[3:0];
  _RAND_259 = {1{`RANDOM}};
  image_0_259 = _RAND_259[3:0];
  _RAND_260 = {1{`RANDOM}};
  image_0_260 = _RAND_260[3:0];
  _RAND_261 = {1{`RANDOM}};
  image_0_261 = _RAND_261[3:0];
  _RAND_262 = {1{`RANDOM}};
  image_0_262 = _RAND_262[3:0];
  _RAND_263 = {1{`RANDOM}};
  image_0_263 = _RAND_263[3:0];
  _RAND_264 = {1{`RANDOM}};
  image_0_264 = _RAND_264[3:0];
  _RAND_265 = {1{`RANDOM}};
  image_0_265 = _RAND_265[3:0];
  _RAND_266 = {1{`RANDOM}};
  image_0_266 = _RAND_266[3:0];
  _RAND_267 = {1{`RANDOM}};
  image_0_267 = _RAND_267[3:0];
  _RAND_268 = {1{`RANDOM}};
  image_0_268 = _RAND_268[3:0];
  _RAND_269 = {1{`RANDOM}};
  image_0_269 = _RAND_269[3:0];
  _RAND_270 = {1{`RANDOM}};
  image_0_270 = _RAND_270[3:0];
  _RAND_271 = {1{`RANDOM}};
  image_0_271 = _RAND_271[3:0];
  _RAND_272 = {1{`RANDOM}};
  image_0_272 = _RAND_272[3:0];
  _RAND_273 = {1{`RANDOM}};
  image_0_273 = _RAND_273[3:0];
  _RAND_274 = {1{`RANDOM}};
  image_0_274 = _RAND_274[3:0];
  _RAND_275 = {1{`RANDOM}};
  image_0_275 = _RAND_275[3:0];
  _RAND_276 = {1{`RANDOM}};
  image_0_276 = _RAND_276[3:0];
  _RAND_277 = {1{`RANDOM}};
  image_0_277 = _RAND_277[3:0];
  _RAND_278 = {1{`RANDOM}};
  image_0_278 = _RAND_278[3:0];
  _RAND_279 = {1{`RANDOM}};
  image_0_279 = _RAND_279[3:0];
  _RAND_280 = {1{`RANDOM}};
  image_0_280 = _RAND_280[3:0];
  _RAND_281 = {1{`RANDOM}};
  image_0_281 = _RAND_281[3:0];
  _RAND_282 = {1{`RANDOM}};
  image_0_282 = _RAND_282[3:0];
  _RAND_283 = {1{`RANDOM}};
  image_0_283 = _RAND_283[3:0];
  _RAND_284 = {1{`RANDOM}};
  image_0_284 = _RAND_284[3:0];
  _RAND_285 = {1{`RANDOM}};
  image_0_285 = _RAND_285[3:0];
  _RAND_286 = {1{`RANDOM}};
  image_0_286 = _RAND_286[3:0];
  _RAND_287 = {1{`RANDOM}};
  image_0_287 = _RAND_287[3:0];
  _RAND_288 = {1{`RANDOM}};
  image_0_288 = _RAND_288[3:0];
  _RAND_289 = {1{`RANDOM}};
  image_0_289 = _RAND_289[3:0];
  _RAND_290 = {1{`RANDOM}};
  image_0_290 = _RAND_290[3:0];
  _RAND_291 = {1{`RANDOM}};
  image_0_291 = _RAND_291[3:0];
  _RAND_292 = {1{`RANDOM}};
  image_0_292 = _RAND_292[3:0];
  _RAND_293 = {1{`RANDOM}};
  image_0_293 = _RAND_293[3:0];
  _RAND_294 = {1{`RANDOM}};
  image_0_294 = _RAND_294[3:0];
  _RAND_295 = {1{`RANDOM}};
  image_0_295 = _RAND_295[3:0];
  _RAND_296 = {1{`RANDOM}};
  image_0_296 = _RAND_296[3:0];
  _RAND_297 = {1{`RANDOM}};
  image_0_297 = _RAND_297[3:0];
  _RAND_298 = {1{`RANDOM}};
  image_0_298 = _RAND_298[3:0];
  _RAND_299 = {1{`RANDOM}};
  image_0_299 = _RAND_299[3:0];
  _RAND_300 = {1{`RANDOM}};
  image_0_300 = _RAND_300[3:0];
  _RAND_301 = {1{`RANDOM}};
  image_0_301 = _RAND_301[3:0];
  _RAND_302 = {1{`RANDOM}};
  image_0_302 = _RAND_302[3:0];
  _RAND_303 = {1{`RANDOM}};
  image_0_303 = _RAND_303[3:0];
  _RAND_304 = {1{`RANDOM}};
  image_0_304 = _RAND_304[3:0];
  _RAND_305 = {1{`RANDOM}};
  image_0_305 = _RAND_305[3:0];
  _RAND_306 = {1{`RANDOM}};
  image_0_306 = _RAND_306[3:0];
  _RAND_307 = {1{`RANDOM}};
  image_0_307 = _RAND_307[3:0];
  _RAND_308 = {1{`RANDOM}};
  image_0_308 = _RAND_308[3:0];
  _RAND_309 = {1{`RANDOM}};
  image_0_309 = _RAND_309[3:0];
  _RAND_310 = {1{`RANDOM}};
  image_0_310 = _RAND_310[3:0];
  _RAND_311 = {1{`RANDOM}};
  image_0_311 = _RAND_311[3:0];
  _RAND_312 = {1{`RANDOM}};
  image_0_312 = _RAND_312[3:0];
  _RAND_313 = {1{`RANDOM}};
  image_0_313 = _RAND_313[3:0];
  _RAND_314 = {1{`RANDOM}};
  image_0_314 = _RAND_314[3:0];
  _RAND_315 = {1{`RANDOM}};
  image_0_315 = _RAND_315[3:0];
  _RAND_316 = {1{`RANDOM}};
  image_0_316 = _RAND_316[3:0];
  _RAND_317 = {1{`RANDOM}};
  image_0_317 = _RAND_317[3:0];
  _RAND_318 = {1{`RANDOM}};
  image_0_318 = _RAND_318[3:0];
  _RAND_319 = {1{`RANDOM}};
  image_0_319 = _RAND_319[3:0];
  _RAND_320 = {1{`RANDOM}};
  image_0_320 = _RAND_320[3:0];
  _RAND_321 = {1{`RANDOM}};
  image_0_321 = _RAND_321[3:0];
  _RAND_322 = {1{`RANDOM}};
  image_0_322 = _RAND_322[3:0];
  _RAND_323 = {1{`RANDOM}};
  image_0_323 = _RAND_323[3:0];
  _RAND_324 = {1{`RANDOM}};
  image_0_324 = _RAND_324[3:0];
  _RAND_325 = {1{`RANDOM}};
  image_0_325 = _RAND_325[3:0];
  _RAND_326 = {1{`RANDOM}};
  image_0_326 = _RAND_326[3:0];
  _RAND_327 = {1{`RANDOM}};
  image_0_327 = _RAND_327[3:0];
  _RAND_328 = {1{`RANDOM}};
  image_0_328 = _RAND_328[3:0];
  _RAND_329 = {1{`RANDOM}};
  image_0_329 = _RAND_329[3:0];
  _RAND_330 = {1{`RANDOM}};
  image_0_330 = _RAND_330[3:0];
  _RAND_331 = {1{`RANDOM}};
  image_0_331 = _RAND_331[3:0];
  _RAND_332 = {1{`RANDOM}};
  image_0_332 = _RAND_332[3:0];
  _RAND_333 = {1{`RANDOM}};
  image_0_333 = _RAND_333[3:0];
  _RAND_334 = {1{`RANDOM}};
  image_0_334 = _RAND_334[3:0];
  _RAND_335 = {1{`RANDOM}};
  image_0_335 = _RAND_335[3:0];
  _RAND_336 = {1{`RANDOM}};
  image_0_336 = _RAND_336[3:0];
  _RAND_337 = {1{`RANDOM}};
  image_0_337 = _RAND_337[3:0];
  _RAND_338 = {1{`RANDOM}};
  image_0_338 = _RAND_338[3:0];
  _RAND_339 = {1{`RANDOM}};
  image_0_339 = _RAND_339[3:0];
  _RAND_340 = {1{`RANDOM}};
  image_0_340 = _RAND_340[3:0];
  _RAND_341 = {1{`RANDOM}};
  image_0_341 = _RAND_341[3:0];
  _RAND_342 = {1{`RANDOM}};
  image_0_342 = _RAND_342[3:0];
  _RAND_343 = {1{`RANDOM}};
  image_0_343 = _RAND_343[3:0];
  _RAND_344 = {1{`RANDOM}};
  image_0_344 = _RAND_344[3:0];
  _RAND_345 = {1{`RANDOM}};
  image_0_345 = _RAND_345[3:0];
  _RAND_346 = {1{`RANDOM}};
  image_0_346 = _RAND_346[3:0];
  _RAND_347 = {1{`RANDOM}};
  image_0_347 = _RAND_347[3:0];
  _RAND_348 = {1{`RANDOM}};
  image_0_348 = _RAND_348[3:0];
  _RAND_349 = {1{`RANDOM}};
  image_0_349 = _RAND_349[3:0];
  _RAND_350 = {1{`RANDOM}};
  image_0_350 = _RAND_350[3:0];
  _RAND_351 = {1{`RANDOM}};
  image_0_351 = _RAND_351[3:0];
  _RAND_352 = {1{`RANDOM}};
  image_0_352 = _RAND_352[3:0];
  _RAND_353 = {1{`RANDOM}};
  image_0_353 = _RAND_353[3:0];
  _RAND_354 = {1{`RANDOM}};
  image_0_354 = _RAND_354[3:0];
  _RAND_355 = {1{`RANDOM}};
  image_0_355 = _RAND_355[3:0];
  _RAND_356 = {1{`RANDOM}};
  image_0_356 = _RAND_356[3:0];
  _RAND_357 = {1{`RANDOM}};
  image_0_357 = _RAND_357[3:0];
  _RAND_358 = {1{`RANDOM}};
  image_0_358 = _RAND_358[3:0];
  _RAND_359 = {1{`RANDOM}};
  image_0_359 = _RAND_359[3:0];
  _RAND_360 = {1{`RANDOM}};
  image_0_360 = _RAND_360[3:0];
  _RAND_361 = {1{`RANDOM}};
  image_0_361 = _RAND_361[3:0];
  _RAND_362 = {1{`RANDOM}};
  image_0_362 = _RAND_362[3:0];
  _RAND_363 = {1{`RANDOM}};
  image_0_363 = _RAND_363[3:0];
  _RAND_364 = {1{`RANDOM}};
  image_0_364 = _RAND_364[3:0];
  _RAND_365 = {1{`RANDOM}};
  image_0_365 = _RAND_365[3:0];
  _RAND_366 = {1{`RANDOM}};
  image_0_366 = _RAND_366[3:0];
  _RAND_367 = {1{`RANDOM}};
  image_0_367 = _RAND_367[3:0];
  _RAND_368 = {1{`RANDOM}};
  image_0_368 = _RAND_368[3:0];
  _RAND_369 = {1{`RANDOM}};
  image_0_369 = _RAND_369[3:0];
  _RAND_370 = {1{`RANDOM}};
  image_0_370 = _RAND_370[3:0];
  _RAND_371 = {1{`RANDOM}};
  image_0_371 = _RAND_371[3:0];
  _RAND_372 = {1{`RANDOM}};
  image_0_372 = _RAND_372[3:0];
  _RAND_373 = {1{`RANDOM}};
  image_0_373 = _RAND_373[3:0];
  _RAND_374 = {1{`RANDOM}};
  image_0_374 = _RAND_374[3:0];
  _RAND_375 = {1{`RANDOM}};
  image_0_375 = _RAND_375[3:0];
  _RAND_376 = {1{`RANDOM}};
  image_0_376 = _RAND_376[3:0];
  _RAND_377 = {1{`RANDOM}};
  image_0_377 = _RAND_377[3:0];
  _RAND_378 = {1{`RANDOM}};
  image_0_378 = _RAND_378[3:0];
  _RAND_379 = {1{`RANDOM}};
  image_0_379 = _RAND_379[3:0];
  _RAND_380 = {1{`RANDOM}};
  image_0_380 = _RAND_380[3:0];
  _RAND_381 = {1{`RANDOM}};
  image_0_381 = _RAND_381[3:0];
  _RAND_382 = {1{`RANDOM}};
  image_0_382 = _RAND_382[3:0];
  _RAND_383 = {1{`RANDOM}};
  image_0_383 = _RAND_383[3:0];
  _RAND_384 = {1{`RANDOM}};
  image_0_384 = _RAND_384[3:0];
  _RAND_385 = {1{`RANDOM}};
  image_0_385 = _RAND_385[3:0];
  _RAND_386 = {1{`RANDOM}};
  image_0_386 = _RAND_386[3:0];
  _RAND_387 = {1{`RANDOM}};
  image_0_387 = _RAND_387[3:0];
  _RAND_388 = {1{`RANDOM}};
  image_0_388 = _RAND_388[3:0];
  _RAND_389 = {1{`RANDOM}};
  image_0_389 = _RAND_389[3:0];
  _RAND_390 = {1{`RANDOM}};
  image_0_390 = _RAND_390[3:0];
  _RAND_391 = {1{`RANDOM}};
  image_0_391 = _RAND_391[3:0];
  _RAND_392 = {1{`RANDOM}};
  image_0_392 = _RAND_392[3:0];
  _RAND_393 = {1{`RANDOM}};
  image_0_393 = _RAND_393[3:0];
  _RAND_394 = {1{`RANDOM}};
  image_0_394 = _RAND_394[3:0];
  _RAND_395 = {1{`RANDOM}};
  image_0_395 = _RAND_395[3:0];
  _RAND_396 = {1{`RANDOM}};
  image_0_396 = _RAND_396[3:0];
  _RAND_397 = {1{`RANDOM}};
  image_0_397 = _RAND_397[3:0];
  _RAND_398 = {1{`RANDOM}};
  image_0_398 = _RAND_398[3:0];
  _RAND_399 = {1{`RANDOM}};
  image_0_399 = _RAND_399[3:0];
  _RAND_400 = {1{`RANDOM}};
  image_0_400 = _RAND_400[3:0];
  _RAND_401 = {1{`RANDOM}};
  image_0_401 = _RAND_401[3:0];
  _RAND_402 = {1{`RANDOM}};
  image_0_402 = _RAND_402[3:0];
  _RAND_403 = {1{`RANDOM}};
  image_0_403 = _RAND_403[3:0];
  _RAND_404 = {1{`RANDOM}};
  image_0_404 = _RAND_404[3:0];
  _RAND_405 = {1{`RANDOM}};
  image_0_405 = _RAND_405[3:0];
  _RAND_406 = {1{`RANDOM}};
  image_0_406 = _RAND_406[3:0];
  _RAND_407 = {1{`RANDOM}};
  image_0_407 = _RAND_407[3:0];
  _RAND_408 = {1{`RANDOM}};
  image_0_408 = _RAND_408[3:0];
  _RAND_409 = {1{`RANDOM}};
  image_0_409 = _RAND_409[3:0];
  _RAND_410 = {1{`RANDOM}};
  image_0_410 = _RAND_410[3:0];
  _RAND_411 = {1{`RANDOM}};
  image_0_411 = _RAND_411[3:0];
  _RAND_412 = {1{`RANDOM}};
  image_0_412 = _RAND_412[3:0];
  _RAND_413 = {1{`RANDOM}};
  image_0_413 = _RAND_413[3:0];
  _RAND_414 = {1{`RANDOM}};
  image_0_414 = _RAND_414[3:0];
  _RAND_415 = {1{`RANDOM}};
  image_0_415 = _RAND_415[3:0];
  _RAND_416 = {1{`RANDOM}};
  image_0_416 = _RAND_416[3:0];
  _RAND_417 = {1{`RANDOM}};
  image_0_417 = _RAND_417[3:0];
  _RAND_418 = {1{`RANDOM}};
  image_0_418 = _RAND_418[3:0];
  _RAND_419 = {1{`RANDOM}};
  image_0_419 = _RAND_419[3:0];
  _RAND_420 = {1{`RANDOM}};
  image_0_420 = _RAND_420[3:0];
  _RAND_421 = {1{`RANDOM}};
  image_0_421 = _RAND_421[3:0];
  _RAND_422 = {1{`RANDOM}};
  image_0_422 = _RAND_422[3:0];
  _RAND_423 = {1{`RANDOM}};
  image_0_423 = _RAND_423[3:0];
  _RAND_424 = {1{`RANDOM}};
  image_0_424 = _RAND_424[3:0];
  _RAND_425 = {1{`RANDOM}};
  image_0_425 = _RAND_425[3:0];
  _RAND_426 = {1{`RANDOM}};
  image_0_426 = _RAND_426[3:0];
  _RAND_427 = {1{`RANDOM}};
  image_0_427 = _RAND_427[3:0];
  _RAND_428 = {1{`RANDOM}};
  image_0_428 = _RAND_428[3:0];
  _RAND_429 = {1{`RANDOM}};
  image_0_429 = _RAND_429[3:0];
  _RAND_430 = {1{`RANDOM}};
  image_0_430 = _RAND_430[3:0];
  _RAND_431 = {1{`RANDOM}};
  image_0_431 = _RAND_431[3:0];
  _RAND_432 = {1{`RANDOM}};
  image_0_432 = _RAND_432[3:0];
  _RAND_433 = {1{`RANDOM}};
  image_0_433 = _RAND_433[3:0];
  _RAND_434 = {1{`RANDOM}};
  image_0_434 = _RAND_434[3:0];
  _RAND_435 = {1{`RANDOM}};
  image_0_435 = _RAND_435[3:0];
  _RAND_436 = {1{`RANDOM}};
  image_0_436 = _RAND_436[3:0];
  _RAND_437 = {1{`RANDOM}};
  image_0_437 = _RAND_437[3:0];
  _RAND_438 = {1{`RANDOM}};
  image_0_438 = _RAND_438[3:0];
  _RAND_439 = {1{`RANDOM}};
  image_0_439 = _RAND_439[3:0];
  _RAND_440 = {1{`RANDOM}};
  image_0_440 = _RAND_440[3:0];
  _RAND_441 = {1{`RANDOM}};
  image_0_441 = _RAND_441[3:0];
  _RAND_442 = {1{`RANDOM}};
  image_0_442 = _RAND_442[3:0];
  _RAND_443 = {1{`RANDOM}};
  image_0_443 = _RAND_443[3:0];
  _RAND_444 = {1{`RANDOM}};
  image_0_444 = _RAND_444[3:0];
  _RAND_445 = {1{`RANDOM}};
  image_0_445 = _RAND_445[3:0];
  _RAND_446 = {1{`RANDOM}};
  image_0_446 = _RAND_446[3:0];
  _RAND_447 = {1{`RANDOM}};
  image_0_447 = _RAND_447[3:0];
  _RAND_448 = {1{`RANDOM}};
  image_0_448 = _RAND_448[3:0];
  _RAND_449 = {1{`RANDOM}};
  image_0_449 = _RAND_449[3:0];
  _RAND_450 = {1{`RANDOM}};
  image_0_450 = _RAND_450[3:0];
  _RAND_451 = {1{`RANDOM}};
  image_0_451 = _RAND_451[3:0];
  _RAND_452 = {1{`RANDOM}};
  image_0_452 = _RAND_452[3:0];
  _RAND_453 = {1{`RANDOM}};
  image_0_453 = _RAND_453[3:0];
  _RAND_454 = {1{`RANDOM}};
  image_0_454 = _RAND_454[3:0];
  _RAND_455 = {1{`RANDOM}};
  image_0_455 = _RAND_455[3:0];
  _RAND_456 = {1{`RANDOM}};
  image_0_456 = _RAND_456[3:0];
  _RAND_457 = {1{`RANDOM}};
  image_0_457 = _RAND_457[3:0];
  _RAND_458 = {1{`RANDOM}};
  image_0_458 = _RAND_458[3:0];
  _RAND_459 = {1{`RANDOM}};
  image_0_459 = _RAND_459[3:0];
  _RAND_460 = {1{`RANDOM}};
  image_0_460 = _RAND_460[3:0];
  _RAND_461 = {1{`RANDOM}};
  image_0_461 = _RAND_461[3:0];
  _RAND_462 = {1{`RANDOM}};
  image_0_462 = _RAND_462[3:0];
  _RAND_463 = {1{`RANDOM}};
  image_0_463 = _RAND_463[3:0];
  _RAND_464 = {1{`RANDOM}};
  image_0_464 = _RAND_464[3:0];
  _RAND_465 = {1{`RANDOM}};
  image_0_465 = _RAND_465[3:0];
  _RAND_466 = {1{`RANDOM}};
  image_0_466 = _RAND_466[3:0];
  _RAND_467 = {1{`RANDOM}};
  image_0_467 = _RAND_467[3:0];
  _RAND_468 = {1{`RANDOM}};
  image_0_468 = _RAND_468[3:0];
  _RAND_469 = {1{`RANDOM}};
  image_0_469 = _RAND_469[3:0];
  _RAND_470 = {1{`RANDOM}};
  image_0_470 = _RAND_470[3:0];
  _RAND_471 = {1{`RANDOM}};
  image_0_471 = _RAND_471[3:0];
  _RAND_472 = {1{`RANDOM}};
  image_0_472 = _RAND_472[3:0];
  _RAND_473 = {1{`RANDOM}};
  image_0_473 = _RAND_473[3:0];
  _RAND_474 = {1{`RANDOM}};
  image_0_474 = _RAND_474[3:0];
  _RAND_475 = {1{`RANDOM}};
  image_0_475 = _RAND_475[3:0];
  _RAND_476 = {1{`RANDOM}};
  image_0_476 = _RAND_476[3:0];
  _RAND_477 = {1{`RANDOM}};
  image_0_477 = _RAND_477[3:0];
  _RAND_478 = {1{`RANDOM}};
  image_0_478 = _RAND_478[3:0];
  _RAND_479 = {1{`RANDOM}};
  image_0_479 = _RAND_479[3:0];
  _RAND_480 = {1{`RANDOM}};
  image_0_480 = _RAND_480[3:0];
  _RAND_481 = {1{`RANDOM}};
  image_0_481 = _RAND_481[3:0];
  _RAND_482 = {1{`RANDOM}};
  image_0_482 = _RAND_482[3:0];
  _RAND_483 = {1{`RANDOM}};
  image_0_483 = _RAND_483[3:0];
  _RAND_484 = {1{`RANDOM}};
  image_0_484 = _RAND_484[3:0];
  _RAND_485 = {1{`RANDOM}};
  image_0_485 = _RAND_485[3:0];
  _RAND_486 = {1{`RANDOM}};
  image_0_486 = _RAND_486[3:0];
  _RAND_487 = {1{`RANDOM}};
  image_0_487 = _RAND_487[3:0];
  _RAND_488 = {1{`RANDOM}};
  image_0_488 = _RAND_488[3:0];
  _RAND_489 = {1{`RANDOM}};
  image_0_489 = _RAND_489[3:0];
  _RAND_490 = {1{`RANDOM}};
  image_0_490 = _RAND_490[3:0];
  _RAND_491 = {1{`RANDOM}};
  image_0_491 = _RAND_491[3:0];
  _RAND_492 = {1{`RANDOM}};
  image_0_492 = _RAND_492[3:0];
  _RAND_493 = {1{`RANDOM}};
  image_0_493 = _RAND_493[3:0];
  _RAND_494 = {1{`RANDOM}};
  image_0_494 = _RAND_494[3:0];
  _RAND_495 = {1{`RANDOM}};
  image_0_495 = _RAND_495[3:0];
  _RAND_496 = {1{`RANDOM}};
  image_0_496 = _RAND_496[3:0];
  _RAND_497 = {1{`RANDOM}};
  image_0_497 = _RAND_497[3:0];
  _RAND_498 = {1{`RANDOM}};
  image_0_498 = _RAND_498[3:0];
  _RAND_499 = {1{`RANDOM}};
  image_0_499 = _RAND_499[3:0];
  _RAND_500 = {1{`RANDOM}};
  image_0_500 = _RAND_500[3:0];
  _RAND_501 = {1{`RANDOM}};
  image_0_501 = _RAND_501[3:0];
  _RAND_502 = {1{`RANDOM}};
  image_0_502 = _RAND_502[3:0];
  _RAND_503 = {1{`RANDOM}};
  image_0_503 = _RAND_503[3:0];
  _RAND_504 = {1{`RANDOM}};
  image_0_504 = _RAND_504[3:0];
  _RAND_505 = {1{`RANDOM}};
  image_0_505 = _RAND_505[3:0];
  _RAND_506 = {1{`RANDOM}};
  image_0_506 = _RAND_506[3:0];
  _RAND_507 = {1{`RANDOM}};
  image_0_507 = _RAND_507[3:0];
  _RAND_508 = {1{`RANDOM}};
  image_0_508 = _RAND_508[3:0];
  _RAND_509 = {1{`RANDOM}};
  image_0_509 = _RAND_509[3:0];
  _RAND_510 = {1{`RANDOM}};
  image_0_510 = _RAND_510[3:0];
  _RAND_511 = {1{`RANDOM}};
  image_0_511 = _RAND_511[3:0];
  _RAND_512 = {1{`RANDOM}};
  image_0_512 = _RAND_512[3:0];
  _RAND_513 = {1{`RANDOM}};
  image_0_513 = _RAND_513[3:0];
  _RAND_514 = {1{`RANDOM}};
  image_0_514 = _RAND_514[3:0];
  _RAND_515 = {1{`RANDOM}};
  image_0_515 = _RAND_515[3:0];
  _RAND_516 = {1{`RANDOM}};
  image_0_516 = _RAND_516[3:0];
  _RAND_517 = {1{`RANDOM}};
  image_0_517 = _RAND_517[3:0];
  _RAND_518 = {1{`RANDOM}};
  image_0_518 = _RAND_518[3:0];
  _RAND_519 = {1{`RANDOM}};
  image_0_519 = _RAND_519[3:0];
  _RAND_520 = {1{`RANDOM}};
  image_0_520 = _RAND_520[3:0];
  _RAND_521 = {1{`RANDOM}};
  image_0_521 = _RAND_521[3:0];
  _RAND_522 = {1{`RANDOM}};
  image_0_522 = _RAND_522[3:0];
  _RAND_523 = {1{`RANDOM}};
  image_0_523 = _RAND_523[3:0];
  _RAND_524 = {1{`RANDOM}};
  image_0_524 = _RAND_524[3:0];
  _RAND_525 = {1{`RANDOM}};
  image_0_525 = _RAND_525[3:0];
  _RAND_526 = {1{`RANDOM}};
  image_0_526 = _RAND_526[3:0];
  _RAND_527 = {1{`RANDOM}};
  image_0_527 = _RAND_527[3:0];
  _RAND_528 = {1{`RANDOM}};
  image_0_528 = _RAND_528[3:0];
  _RAND_529 = {1{`RANDOM}};
  image_0_529 = _RAND_529[3:0];
  _RAND_530 = {1{`RANDOM}};
  image_0_530 = _RAND_530[3:0];
  _RAND_531 = {1{`RANDOM}};
  image_0_531 = _RAND_531[3:0];
  _RAND_532 = {1{`RANDOM}};
  image_0_532 = _RAND_532[3:0];
  _RAND_533 = {1{`RANDOM}};
  image_0_533 = _RAND_533[3:0];
  _RAND_534 = {1{`RANDOM}};
  image_0_534 = _RAND_534[3:0];
  _RAND_535 = {1{`RANDOM}};
  image_0_535 = _RAND_535[3:0];
  _RAND_536 = {1{`RANDOM}};
  image_0_536 = _RAND_536[3:0];
  _RAND_537 = {1{`RANDOM}};
  image_0_537 = _RAND_537[3:0];
  _RAND_538 = {1{`RANDOM}};
  image_0_538 = _RAND_538[3:0];
  _RAND_539 = {1{`RANDOM}};
  image_0_539 = _RAND_539[3:0];
  _RAND_540 = {1{`RANDOM}};
  image_0_540 = _RAND_540[3:0];
  _RAND_541 = {1{`RANDOM}};
  image_0_541 = _RAND_541[3:0];
  _RAND_542 = {1{`RANDOM}};
  image_0_542 = _RAND_542[3:0];
  _RAND_543 = {1{`RANDOM}};
  image_0_543 = _RAND_543[3:0];
  _RAND_544 = {1{`RANDOM}};
  image_0_544 = _RAND_544[3:0];
  _RAND_545 = {1{`RANDOM}};
  image_0_545 = _RAND_545[3:0];
  _RAND_546 = {1{`RANDOM}};
  image_0_546 = _RAND_546[3:0];
  _RAND_547 = {1{`RANDOM}};
  image_0_547 = _RAND_547[3:0];
  _RAND_548 = {1{`RANDOM}};
  image_0_548 = _RAND_548[3:0];
  _RAND_549 = {1{`RANDOM}};
  image_0_549 = _RAND_549[3:0];
  _RAND_550 = {1{`RANDOM}};
  image_0_550 = _RAND_550[3:0];
  _RAND_551 = {1{`RANDOM}};
  image_0_551 = _RAND_551[3:0];
  _RAND_552 = {1{`RANDOM}};
  image_0_552 = _RAND_552[3:0];
  _RAND_553 = {1{`RANDOM}};
  image_0_553 = _RAND_553[3:0];
  _RAND_554 = {1{`RANDOM}};
  image_0_554 = _RAND_554[3:0];
  _RAND_555 = {1{`RANDOM}};
  image_0_555 = _RAND_555[3:0];
  _RAND_556 = {1{`RANDOM}};
  image_0_556 = _RAND_556[3:0];
  _RAND_557 = {1{`RANDOM}};
  image_0_557 = _RAND_557[3:0];
  _RAND_558 = {1{`RANDOM}};
  image_0_558 = _RAND_558[3:0];
  _RAND_559 = {1{`RANDOM}};
  image_0_559 = _RAND_559[3:0];
  _RAND_560 = {1{`RANDOM}};
  image_0_560 = _RAND_560[3:0];
  _RAND_561 = {1{`RANDOM}};
  image_0_561 = _RAND_561[3:0];
  _RAND_562 = {1{`RANDOM}};
  image_0_562 = _RAND_562[3:0];
  _RAND_563 = {1{`RANDOM}};
  image_0_563 = _RAND_563[3:0];
  _RAND_564 = {1{`RANDOM}};
  image_0_564 = _RAND_564[3:0];
  _RAND_565 = {1{`RANDOM}};
  image_0_565 = _RAND_565[3:0];
  _RAND_566 = {1{`RANDOM}};
  image_0_566 = _RAND_566[3:0];
  _RAND_567 = {1{`RANDOM}};
  image_0_567 = _RAND_567[3:0];
  _RAND_568 = {1{`RANDOM}};
  image_0_568 = _RAND_568[3:0];
  _RAND_569 = {1{`RANDOM}};
  image_0_569 = _RAND_569[3:0];
  _RAND_570 = {1{`RANDOM}};
  image_0_570 = _RAND_570[3:0];
  _RAND_571 = {1{`RANDOM}};
  image_0_571 = _RAND_571[3:0];
  _RAND_572 = {1{`RANDOM}};
  image_0_572 = _RAND_572[3:0];
  _RAND_573 = {1{`RANDOM}};
  image_0_573 = _RAND_573[3:0];
  _RAND_574 = {1{`RANDOM}};
  image_0_574 = _RAND_574[3:0];
  _RAND_575 = {1{`RANDOM}};
  image_0_575 = _RAND_575[3:0];
  _RAND_576 = {1{`RANDOM}};
  image_1_0 = _RAND_576[3:0];
  _RAND_577 = {1{`RANDOM}};
  image_1_1 = _RAND_577[3:0];
  _RAND_578 = {1{`RANDOM}};
  image_1_2 = _RAND_578[3:0];
  _RAND_579 = {1{`RANDOM}};
  image_1_3 = _RAND_579[3:0];
  _RAND_580 = {1{`RANDOM}};
  image_1_4 = _RAND_580[3:0];
  _RAND_581 = {1{`RANDOM}};
  image_1_5 = _RAND_581[3:0];
  _RAND_582 = {1{`RANDOM}};
  image_1_6 = _RAND_582[3:0];
  _RAND_583 = {1{`RANDOM}};
  image_1_7 = _RAND_583[3:0];
  _RAND_584 = {1{`RANDOM}};
  image_1_8 = _RAND_584[3:0];
  _RAND_585 = {1{`RANDOM}};
  image_1_9 = _RAND_585[3:0];
  _RAND_586 = {1{`RANDOM}};
  image_1_10 = _RAND_586[3:0];
  _RAND_587 = {1{`RANDOM}};
  image_1_11 = _RAND_587[3:0];
  _RAND_588 = {1{`RANDOM}};
  image_1_12 = _RAND_588[3:0];
  _RAND_589 = {1{`RANDOM}};
  image_1_13 = _RAND_589[3:0];
  _RAND_590 = {1{`RANDOM}};
  image_1_14 = _RAND_590[3:0];
  _RAND_591 = {1{`RANDOM}};
  image_1_15 = _RAND_591[3:0];
  _RAND_592 = {1{`RANDOM}};
  image_1_16 = _RAND_592[3:0];
  _RAND_593 = {1{`RANDOM}};
  image_1_17 = _RAND_593[3:0];
  _RAND_594 = {1{`RANDOM}};
  image_1_18 = _RAND_594[3:0];
  _RAND_595 = {1{`RANDOM}};
  image_1_19 = _RAND_595[3:0];
  _RAND_596 = {1{`RANDOM}};
  image_1_20 = _RAND_596[3:0];
  _RAND_597 = {1{`RANDOM}};
  image_1_21 = _RAND_597[3:0];
  _RAND_598 = {1{`RANDOM}};
  image_1_22 = _RAND_598[3:0];
  _RAND_599 = {1{`RANDOM}};
  image_1_23 = _RAND_599[3:0];
  _RAND_600 = {1{`RANDOM}};
  image_1_24 = _RAND_600[3:0];
  _RAND_601 = {1{`RANDOM}};
  image_1_25 = _RAND_601[3:0];
  _RAND_602 = {1{`RANDOM}};
  image_1_26 = _RAND_602[3:0];
  _RAND_603 = {1{`RANDOM}};
  image_1_27 = _RAND_603[3:0];
  _RAND_604 = {1{`RANDOM}};
  image_1_28 = _RAND_604[3:0];
  _RAND_605 = {1{`RANDOM}};
  image_1_29 = _RAND_605[3:0];
  _RAND_606 = {1{`RANDOM}};
  image_1_30 = _RAND_606[3:0];
  _RAND_607 = {1{`RANDOM}};
  image_1_31 = _RAND_607[3:0];
  _RAND_608 = {1{`RANDOM}};
  image_1_32 = _RAND_608[3:0];
  _RAND_609 = {1{`RANDOM}};
  image_1_33 = _RAND_609[3:0];
  _RAND_610 = {1{`RANDOM}};
  image_1_34 = _RAND_610[3:0];
  _RAND_611 = {1{`RANDOM}};
  image_1_35 = _RAND_611[3:0];
  _RAND_612 = {1{`RANDOM}};
  image_1_36 = _RAND_612[3:0];
  _RAND_613 = {1{`RANDOM}};
  image_1_37 = _RAND_613[3:0];
  _RAND_614 = {1{`RANDOM}};
  image_1_38 = _RAND_614[3:0];
  _RAND_615 = {1{`RANDOM}};
  image_1_39 = _RAND_615[3:0];
  _RAND_616 = {1{`RANDOM}};
  image_1_40 = _RAND_616[3:0];
  _RAND_617 = {1{`RANDOM}};
  image_1_41 = _RAND_617[3:0];
  _RAND_618 = {1{`RANDOM}};
  image_1_42 = _RAND_618[3:0];
  _RAND_619 = {1{`RANDOM}};
  image_1_43 = _RAND_619[3:0];
  _RAND_620 = {1{`RANDOM}};
  image_1_44 = _RAND_620[3:0];
  _RAND_621 = {1{`RANDOM}};
  image_1_45 = _RAND_621[3:0];
  _RAND_622 = {1{`RANDOM}};
  image_1_46 = _RAND_622[3:0];
  _RAND_623 = {1{`RANDOM}};
  image_1_47 = _RAND_623[3:0];
  _RAND_624 = {1{`RANDOM}};
  image_1_48 = _RAND_624[3:0];
  _RAND_625 = {1{`RANDOM}};
  image_1_49 = _RAND_625[3:0];
  _RAND_626 = {1{`RANDOM}};
  image_1_50 = _RAND_626[3:0];
  _RAND_627 = {1{`RANDOM}};
  image_1_51 = _RAND_627[3:0];
  _RAND_628 = {1{`RANDOM}};
  image_1_52 = _RAND_628[3:0];
  _RAND_629 = {1{`RANDOM}};
  image_1_53 = _RAND_629[3:0];
  _RAND_630 = {1{`RANDOM}};
  image_1_54 = _RAND_630[3:0];
  _RAND_631 = {1{`RANDOM}};
  image_1_55 = _RAND_631[3:0];
  _RAND_632 = {1{`RANDOM}};
  image_1_56 = _RAND_632[3:0];
  _RAND_633 = {1{`RANDOM}};
  image_1_57 = _RAND_633[3:0];
  _RAND_634 = {1{`RANDOM}};
  image_1_58 = _RAND_634[3:0];
  _RAND_635 = {1{`RANDOM}};
  image_1_59 = _RAND_635[3:0];
  _RAND_636 = {1{`RANDOM}};
  image_1_60 = _RAND_636[3:0];
  _RAND_637 = {1{`RANDOM}};
  image_1_61 = _RAND_637[3:0];
  _RAND_638 = {1{`RANDOM}};
  image_1_62 = _RAND_638[3:0];
  _RAND_639 = {1{`RANDOM}};
  image_1_63 = _RAND_639[3:0];
  _RAND_640 = {1{`RANDOM}};
  image_1_64 = _RAND_640[3:0];
  _RAND_641 = {1{`RANDOM}};
  image_1_65 = _RAND_641[3:0];
  _RAND_642 = {1{`RANDOM}};
  image_1_66 = _RAND_642[3:0];
  _RAND_643 = {1{`RANDOM}};
  image_1_67 = _RAND_643[3:0];
  _RAND_644 = {1{`RANDOM}};
  image_1_68 = _RAND_644[3:0];
  _RAND_645 = {1{`RANDOM}};
  image_1_69 = _RAND_645[3:0];
  _RAND_646 = {1{`RANDOM}};
  image_1_70 = _RAND_646[3:0];
  _RAND_647 = {1{`RANDOM}};
  image_1_71 = _RAND_647[3:0];
  _RAND_648 = {1{`RANDOM}};
  image_1_72 = _RAND_648[3:0];
  _RAND_649 = {1{`RANDOM}};
  image_1_73 = _RAND_649[3:0];
  _RAND_650 = {1{`RANDOM}};
  image_1_74 = _RAND_650[3:0];
  _RAND_651 = {1{`RANDOM}};
  image_1_75 = _RAND_651[3:0];
  _RAND_652 = {1{`RANDOM}};
  image_1_76 = _RAND_652[3:0];
  _RAND_653 = {1{`RANDOM}};
  image_1_77 = _RAND_653[3:0];
  _RAND_654 = {1{`RANDOM}};
  image_1_78 = _RAND_654[3:0];
  _RAND_655 = {1{`RANDOM}};
  image_1_79 = _RAND_655[3:0];
  _RAND_656 = {1{`RANDOM}};
  image_1_80 = _RAND_656[3:0];
  _RAND_657 = {1{`RANDOM}};
  image_1_81 = _RAND_657[3:0];
  _RAND_658 = {1{`RANDOM}};
  image_1_82 = _RAND_658[3:0];
  _RAND_659 = {1{`RANDOM}};
  image_1_83 = _RAND_659[3:0];
  _RAND_660 = {1{`RANDOM}};
  image_1_84 = _RAND_660[3:0];
  _RAND_661 = {1{`RANDOM}};
  image_1_85 = _RAND_661[3:0];
  _RAND_662 = {1{`RANDOM}};
  image_1_86 = _RAND_662[3:0];
  _RAND_663 = {1{`RANDOM}};
  image_1_87 = _RAND_663[3:0];
  _RAND_664 = {1{`RANDOM}};
  image_1_88 = _RAND_664[3:0];
  _RAND_665 = {1{`RANDOM}};
  image_1_89 = _RAND_665[3:0];
  _RAND_666 = {1{`RANDOM}};
  image_1_90 = _RAND_666[3:0];
  _RAND_667 = {1{`RANDOM}};
  image_1_91 = _RAND_667[3:0];
  _RAND_668 = {1{`RANDOM}};
  image_1_92 = _RAND_668[3:0];
  _RAND_669 = {1{`RANDOM}};
  image_1_93 = _RAND_669[3:0];
  _RAND_670 = {1{`RANDOM}};
  image_1_94 = _RAND_670[3:0];
  _RAND_671 = {1{`RANDOM}};
  image_1_95 = _RAND_671[3:0];
  _RAND_672 = {1{`RANDOM}};
  image_1_96 = _RAND_672[3:0];
  _RAND_673 = {1{`RANDOM}};
  image_1_97 = _RAND_673[3:0];
  _RAND_674 = {1{`RANDOM}};
  image_1_98 = _RAND_674[3:0];
  _RAND_675 = {1{`RANDOM}};
  image_1_99 = _RAND_675[3:0];
  _RAND_676 = {1{`RANDOM}};
  image_1_100 = _RAND_676[3:0];
  _RAND_677 = {1{`RANDOM}};
  image_1_101 = _RAND_677[3:0];
  _RAND_678 = {1{`RANDOM}};
  image_1_102 = _RAND_678[3:0];
  _RAND_679 = {1{`RANDOM}};
  image_1_103 = _RAND_679[3:0];
  _RAND_680 = {1{`RANDOM}};
  image_1_104 = _RAND_680[3:0];
  _RAND_681 = {1{`RANDOM}};
  image_1_105 = _RAND_681[3:0];
  _RAND_682 = {1{`RANDOM}};
  image_1_106 = _RAND_682[3:0];
  _RAND_683 = {1{`RANDOM}};
  image_1_107 = _RAND_683[3:0];
  _RAND_684 = {1{`RANDOM}};
  image_1_108 = _RAND_684[3:0];
  _RAND_685 = {1{`RANDOM}};
  image_1_109 = _RAND_685[3:0];
  _RAND_686 = {1{`RANDOM}};
  image_1_110 = _RAND_686[3:0];
  _RAND_687 = {1{`RANDOM}};
  image_1_111 = _RAND_687[3:0];
  _RAND_688 = {1{`RANDOM}};
  image_1_112 = _RAND_688[3:0];
  _RAND_689 = {1{`RANDOM}};
  image_1_113 = _RAND_689[3:0];
  _RAND_690 = {1{`RANDOM}};
  image_1_114 = _RAND_690[3:0];
  _RAND_691 = {1{`RANDOM}};
  image_1_115 = _RAND_691[3:0];
  _RAND_692 = {1{`RANDOM}};
  image_1_116 = _RAND_692[3:0];
  _RAND_693 = {1{`RANDOM}};
  image_1_117 = _RAND_693[3:0];
  _RAND_694 = {1{`RANDOM}};
  image_1_118 = _RAND_694[3:0];
  _RAND_695 = {1{`RANDOM}};
  image_1_119 = _RAND_695[3:0];
  _RAND_696 = {1{`RANDOM}};
  image_1_120 = _RAND_696[3:0];
  _RAND_697 = {1{`RANDOM}};
  image_1_121 = _RAND_697[3:0];
  _RAND_698 = {1{`RANDOM}};
  image_1_122 = _RAND_698[3:0];
  _RAND_699 = {1{`RANDOM}};
  image_1_123 = _RAND_699[3:0];
  _RAND_700 = {1{`RANDOM}};
  image_1_124 = _RAND_700[3:0];
  _RAND_701 = {1{`RANDOM}};
  image_1_125 = _RAND_701[3:0];
  _RAND_702 = {1{`RANDOM}};
  image_1_126 = _RAND_702[3:0];
  _RAND_703 = {1{`RANDOM}};
  image_1_127 = _RAND_703[3:0];
  _RAND_704 = {1{`RANDOM}};
  image_1_128 = _RAND_704[3:0];
  _RAND_705 = {1{`RANDOM}};
  image_1_129 = _RAND_705[3:0];
  _RAND_706 = {1{`RANDOM}};
  image_1_130 = _RAND_706[3:0];
  _RAND_707 = {1{`RANDOM}};
  image_1_131 = _RAND_707[3:0];
  _RAND_708 = {1{`RANDOM}};
  image_1_132 = _RAND_708[3:0];
  _RAND_709 = {1{`RANDOM}};
  image_1_133 = _RAND_709[3:0];
  _RAND_710 = {1{`RANDOM}};
  image_1_134 = _RAND_710[3:0];
  _RAND_711 = {1{`RANDOM}};
  image_1_135 = _RAND_711[3:0];
  _RAND_712 = {1{`RANDOM}};
  image_1_136 = _RAND_712[3:0];
  _RAND_713 = {1{`RANDOM}};
  image_1_137 = _RAND_713[3:0];
  _RAND_714 = {1{`RANDOM}};
  image_1_138 = _RAND_714[3:0];
  _RAND_715 = {1{`RANDOM}};
  image_1_139 = _RAND_715[3:0];
  _RAND_716 = {1{`RANDOM}};
  image_1_140 = _RAND_716[3:0];
  _RAND_717 = {1{`RANDOM}};
  image_1_141 = _RAND_717[3:0];
  _RAND_718 = {1{`RANDOM}};
  image_1_142 = _RAND_718[3:0];
  _RAND_719 = {1{`RANDOM}};
  image_1_143 = _RAND_719[3:0];
  _RAND_720 = {1{`RANDOM}};
  image_1_144 = _RAND_720[3:0];
  _RAND_721 = {1{`RANDOM}};
  image_1_145 = _RAND_721[3:0];
  _RAND_722 = {1{`RANDOM}};
  image_1_146 = _RAND_722[3:0];
  _RAND_723 = {1{`RANDOM}};
  image_1_147 = _RAND_723[3:0];
  _RAND_724 = {1{`RANDOM}};
  image_1_148 = _RAND_724[3:0];
  _RAND_725 = {1{`RANDOM}};
  image_1_149 = _RAND_725[3:0];
  _RAND_726 = {1{`RANDOM}};
  image_1_150 = _RAND_726[3:0];
  _RAND_727 = {1{`RANDOM}};
  image_1_151 = _RAND_727[3:0];
  _RAND_728 = {1{`RANDOM}};
  image_1_152 = _RAND_728[3:0];
  _RAND_729 = {1{`RANDOM}};
  image_1_153 = _RAND_729[3:0];
  _RAND_730 = {1{`RANDOM}};
  image_1_154 = _RAND_730[3:0];
  _RAND_731 = {1{`RANDOM}};
  image_1_155 = _RAND_731[3:0];
  _RAND_732 = {1{`RANDOM}};
  image_1_156 = _RAND_732[3:0];
  _RAND_733 = {1{`RANDOM}};
  image_1_157 = _RAND_733[3:0];
  _RAND_734 = {1{`RANDOM}};
  image_1_158 = _RAND_734[3:0];
  _RAND_735 = {1{`RANDOM}};
  image_1_159 = _RAND_735[3:0];
  _RAND_736 = {1{`RANDOM}};
  image_1_160 = _RAND_736[3:0];
  _RAND_737 = {1{`RANDOM}};
  image_1_161 = _RAND_737[3:0];
  _RAND_738 = {1{`RANDOM}};
  image_1_162 = _RAND_738[3:0];
  _RAND_739 = {1{`RANDOM}};
  image_1_163 = _RAND_739[3:0];
  _RAND_740 = {1{`RANDOM}};
  image_1_164 = _RAND_740[3:0];
  _RAND_741 = {1{`RANDOM}};
  image_1_165 = _RAND_741[3:0];
  _RAND_742 = {1{`RANDOM}};
  image_1_166 = _RAND_742[3:0];
  _RAND_743 = {1{`RANDOM}};
  image_1_167 = _RAND_743[3:0];
  _RAND_744 = {1{`RANDOM}};
  image_1_168 = _RAND_744[3:0];
  _RAND_745 = {1{`RANDOM}};
  image_1_169 = _RAND_745[3:0];
  _RAND_746 = {1{`RANDOM}};
  image_1_170 = _RAND_746[3:0];
  _RAND_747 = {1{`RANDOM}};
  image_1_171 = _RAND_747[3:0];
  _RAND_748 = {1{`RANDOM}};
  image_1_172 = _RAND_748[3:0];
  _RAND_749 = {1{`RANDOM}};
  image_1_173 = _RAND_749[3:0];
  _RAND_750 = {1{`RANDOM}};
  image_1_174 = _RAND_750[3:0];
  _RAND_751 = {1{`RANDOM}};
  image_1_175 = _RAND_751[3:0];
  _RAND_752 = {1{`RANDOM}};
  image_1_176 = _RAND_752[3:0];
  _RAND_753 = {1{`RANDOM}};
  image_1_177 = _RAND_753[3:0];
  _RAND_754 = {1{`RANDOM}};
  image_1_178 = _RAND_754[3:0];
  _RAND_755 = {1{`RANDOM}};
  image_1_179 = _RAND_755[3:0];
  _RAND_756 = {1{`RANDOM}};
  image_1_180 = _RAND_756[3:0];
  _RAND_757 = {1{`RANDOM}};
  image_1_181 = _RAND_757[3:0];
  _RAND_758 = {1{`RANDOM}};
  image_1_182 = _RAND_758[3:0];
  _RAND_759 = {1{`RANDOM}};
  image_1_183 = _RAND_759[3:0];
  _RAND_760 = {1{`RANDOM}};
  image_1_184 = _RAND_760[3:0];
  _RAND_761 = {1{`RANDOM}};
  image_1_185 = _RAND_761[3:0];
  _RAND_762 = {1{`RANDOM}};
  image_1_186 = _RAND_762[3:0];
  _RAND_763 = {1{`RANDOM}};
  image_1_187 = _RAND_763[3:0];
  _RAND_764 = {1{`RANDOM}};
  image_1_188 = _RAND_764[3:0];
  _RAND_765 = {1{`RANDOM}};
  image_1_189 = _RAND_765[3:0];
  _RAND_766 = {1{`RANDOM}};
  image_1_190 = _RAND_766[3:0];
  _RAND_767 = {1{`RANDOM}};
  image_1_191 = _RAND_767[3:0];
  _RAND_768 = {1{`RANDOM}};
  image_1_192 = _RAND_768[3:0];
  _RAND_769 = {1{`RANDOM}};
  image_1_193 = _RAND_769[3:0];
  _RAND_770 = {1{`RANDOM}};
  image_1_194 = _RAND_770[3:0];
  _RAND_771 = {1{`RANDOM}};
  image_1_195 = _RAND_771[3:0];
  _RAND_772 = {1{`RANDOM}};
  image_1_196 = _RAND_772[3:0];
  _RAND_773 = {1{`RANDOM}};
  image_1_197 = _RAND_773[3:0];
  _RAND_774 = {1{`RANDOM}};
  image_1_198 = _RAND_774[3:0];
  _RAND_775 = {1{`RANDOM}};
  image_1_199 = _RAND_775[3:0];
  _RAND_776 = {1{`RANDOM}};
  image_1_200 = _RAND_776[3:0];
  _RAND_777 = {1{`RANDOM}};
  image_1_201 = _RAND_777[3:0];
  _RAND_778 = {1{`RANDOM}};
  image_1_202 = _RAND_778[3:0];
  _RAND_779 = {1{`RANDOM}};
  image_1_203 = _RAND_779[3:0];
  _RAND_780 = {1{`RANDOM}};
  image_1_204 = _RAND_780[3:0];
  _RAND_781 = {1{`RANDOM}};
  image_1_205 = _RAND_781[3:0];
  _RAND_782 = {1{`RANDOM}};
  image_1_206 = _RAND_782[3:0];
  _RAND_783 = {1{`RANDOM}};
  image_1_207 = _RAND_783[3:0];
  _RAND_784 = {1{`RANDOM}};
  image_1_208 = _RAND_784[3:0];
  _RAND_785 = {1{`RANDOM}};
  image_1_209 = _RAND_785[3:0];
  _RAND_786 = {1{`RANDOM}};
  image_1_210 = _RAND_786[3:0];
  _RAND_787 = {1{`RANDOM}};
  image_1_211 = _RAND_787[3:0];
  _RAND_788 = {1{`RANDOM}};
  image_1_212 = _RAND_788[3:0];
  _RAND_789 = {1{`RANDOM}};
  image_1_213 = _RAND_789[3:0];
  _RAND_790 = {1{`RANDOM}};
  image_1_214 = _RAND_790[3:0];
  _RAND_791 = {1{`RANDOM}};
  image_1_215 = _RAND_791[3:0];
  _RAND_792 = {1{`RANDOM}};
  image_1_216 = _RAND_792[3:0];
  _RAND_793 = {1{`RANDOM}};
  image_1_217 = _RAND_793[3:0];
  _RAND_794 = {1{`RANDOM}};
  image_1_218 = _RAND_794[3:0];
  _RAND_795 = {1{`RANDOM}};
  image_1_219 = _RAND_795[3:0];
  _RAND_796 = {1{`RANDOM}};
  image_1_220 = _RAND_796[3:0];
  _RAND_797 = {1{`RANDOM}};
  image_1_221 = _RAND_797[3:0];
  _RAND_798 = {1{`RANDOM}};
  image_1_222 = _RAND_798[3:0];
  _RAND_799 = {1{`RANDOM}};
  image_1_223 = _RAND_799[3:0];
  _RAND_800 = {1{`RANDOM}};
  image_1_224 = _RAND_800[3:0];
  _RAND_801 = {1{`RANDOM}};
  image_1_225 = _RAND_801[3:0];
  _RAND_802 = {1{`RANDOM}};
  image_1_226 = _RAND_802[3:0];
  _RAND_803 = {1{`RANDOM}};
  image_1_227 = _RAND_803[3:0];
  _RAND_804 = {1{`RANDOM}};
  image_1_228 = _RAND_804[3:0];
  _RAND_805 = {1{`RANDOM}};
  image_1_229 = _RAND_805[3:0];
  _RAND_806 = {1{`RANDOM}};
  image_1_230 = _RAND_806[3:0];
  _RAND_807 = {1{`RANDOM}};
  image_1_231 = _RAND_807[3:0];
  _RAND_808 = {1{`RANDOM}};
  image_1_232 = _RAND_808[3:0];
  _RAND_809 = {1{`RANDOM}};
  image_1_233 = _RAND_809[3:0];
  _RAND_810 = {1{`RANDOM}};
  image_1_234 = _RAND_810[3:0];
  _RAND_811 = {1{`RANDOM}};
  image_1_235 = _RAND_811[3:0];
  _RAND_812 = {1{`RANDOM}};
  image_1_236 = _RAND_812[3:0];
  _RAND_813 = {1{`RANDOM}};
  image_1_237 = _RAND_813[3:0];
  _RAND_814 = {1{`RANDOM}};
  image_1_238 = _RAND_814[3:0];
  _RAND_815 = {1{`RANDOM}};
  image_1_239 = _RAND_815[3:0];
  _RAND_816 = {1{`RANDOM}};
  image_1_240 = _RAND_816[3:0];
  _RAND_817 = {1{`RANDOM}};
  image_1_241 = _RAND_817[3:0];
  _RAND_818 = {1{`RANDOM}};
  image_1_242 = _RAND_818[3:0];
  _RAND_819 = {1{`RANDOM}};
  image_1_243 = _RAND_819[3:0];
  _RAND_820 = {1{`RANDOM}};
  image_1_244 = _RAND_820[3:0];
  _RAND_821 = {1{`RANDOM}};
  image_1_245 = _RAND_821[3:0];
  _RAND_822 = {1{`RANDOM}};
  image_1_246 = _RAND_822[3:0];
  _RAND_823 = {1{`RANDOM}};
  image_1_247 = _RAND_823[3:0];
  _RAND_824 = {1{`RANDOM}};
  image_1_248 = _RAND_824[3:0];
  _RAND_825 = {1{`RANDOM}};
  image_1_249 = _RAND_825[3:0];
  _RAND_826 = {1{`RANDOM}};
  image_1_250 = _RAND_826[3:0];
  _RAND_827 = {1{`RANDOM}};
  image_1_251 = _RAND_827[3:0];
  _RAND_828 = {1{`RANDOM}};
  image_1_252 = _RAND_828[3:0];
  _RAND_829 = {1{`RANDOM}};
  image_1_253 = _RAND_829[3:0];
  _RAND_830 = {1{`RANDOM}};
  image_1_254 = _RAND_830[3:0];
  _RAND_831 = {1{`RANDOM}};
  image_1_255 = _RAND_831[3:0];
  _RAND_832 = {1{`RANDOM}};
  image_1_256 = _RAND_832[3:0];
  _RAND_833 = {1{`RANDOM}};
  image_1_257 = _RAND_833[3:0];
  _RAND_834 = {1{`RANDOM}};
  image_1_258 = _RAND_834[3:0];
  _RAND_835 = {1{`RANDOM}};
  image_1_259 = _RAND_835[3:0];
  _RAND_836 = {1{`RANDOM}};
  image_1_260 = _RAND_836[3:0];
  _RAND_837 = {1{`RANDOM}};
  image_1_261 = _RAND_837[3:0];
  _RAND_838 = {1{`RANDOM}};
  image_1_262 = _RAND_838[3:0];
  _RAND_839 = {1{`RANDOM}};
  image_1_263 = _RAND_839[3:0];
  _RAND_840 = {1{`RANDOM}};
  image_1_264 = _RAND_840[3:0];
  _RAND_841 = {1{`RANDOM}};
  image_1_265 = _RAND_841[3:0];
  _RAND_842 = {1{`RANDOM}};
  image_1_266 = _RAND_842[3:0];
  _RAND_843 = {1{`RANDOM}};
  image_1_267 = _RAND_843[3:0];
  _RAND_844 = {1{`RANDOM}};
  image_1_268 = _RAND_844[3:0];
  _RAND_845 = {1{`RANDOM}};
  image_1_269 = _RAND_845[3:0];
  _RAND_846 = {1{`RANDOM}};
  image_1_270 = _RAND_846[3:0];
  _RAND_847 = {1{`RANDOM}};
  image_1_271 = _RAND_847[3:0];
  _RAND_848 = {1{`RANDOM}};
  image_1_272 = _RAND_848[3:0];
  _RAND_849 = {1{`RANDOM}};
  image_1_273 = _RAND_849[3:0];
  _RAND_850 = {1{`RANDOM}};
  image_1_274 = _RAND_850[3:0];
  _RAND_851 = {1{`RANDOM}};
  image_1_275 = _RAND_851[3:0];
  _RAND_852 = {1{`RANDOM}};
  image_1_276 = _RAND_852[3:0];
  _RAND_853 = {1{`RANDOM}};
  image_1_277 = _RAND_853[3:0];
  _RAND_854 = {1{`RANDOM}};
  image_1_278 = _RAND_854[3:0];
  _RAND_855 = {1{`RANDOM}};
  image_1_279 = _RAND_855[3:0];
  _RAND_856 = {1{`RANDOM}};
  image_1_280 = _RAND_856[3:0];
  _RAND_857 = {1{`RANDOM}};
  image_1_281 = _RAND_857[3:0];
  _RAND_858 = {1{`RANDOM}};
  image_1_282 = _RAND_858[3:0];
  _RAND_859 = {1{`RANDOM}};
  image_1_283 = _RAND_859[3:0];
  _RAND_860 = {1{`RANDOM}};
  image_1_284 = _RAND_860[3:0];
  _RAND_861 = {1{`RANDOM}};
  image_1_285 = _RAND_861[3:0];
  _RAND_862 = {1{`RANDOM}};
  image_1_286 = _RAND_862[3:0];
  _RAND_863 = {1{`RANDOM}};
  image_1_287 = _RAND_863[3:0];
  _RAND_864 = {1{`RANDOM}};
  image_1_288 = _RAND_864[3:0];
  _RAND_865 = {1{`RANDOM}};
  image_1_289 = _RAND_865[3:0];
  _RAND_866 = {1{`RANDOM}};
  image_1_290 = _RAND_866[3:0];
  _RAND_867 = {1{`RANDOM}};
  image_1_291 = _RAND_867[3:0];
  _RAND_868 = {1{`RANDOM}};
  image_1_292 = _RAND_868[3:0];
  _RAND_869 = {1{`RANDOM}};
  image_1_293 = _RAND_869[3:0];
  _RAND_870 = {1{`RANDOM}};
  image_1_294 = _RAND_870[3:0];
  _RAND_871 = {1{`RANDOM}};
  image_1_295 = _RAND_871[3:0];
  _RAND_872 = {1{`RANDOM}};
  image_1_296 = _RAND_872[3:0];
  _RAND_873 = {1{`RANDOM}};
  image_1_297 = _RAND_873[3:0];
  _RAND_874 = {1{`RANDOM}};
  image_1_298 = _RAND_874[3:0];
  _RAND_875 = {1{`RANDOM}};
  image_1_299 = _RAND_875[3:0];
  _RAND_876 = {1{`RANDOM}};
  image_1_300 = _RAND_876[3:0];
  _RAND_877 = {1{`RANDOM}};
  image_1_301 = _RAND_877[3:0];
  _RAND_878 = {1{`RANDOM}};
  image_1_302 = _RAND_878[3:0];
  _RAND_879 = {1{`RANDOM}};
  image_1_303 = _RAND_879[3:0];
  _RAND_880 = {1{`RANDOM}};
  image_1_304 = _RAND_880[3:0];
  _RAND_881 = {1{`RANDOM}};
  image_1_305 = _RAND_881[3:0];
  _RAND_882 = {1{`RANDOM}};
  image_1_306 = _RAND_882[3:0];
  _RAND_883 = {1{`RANDOM}};
  image_1_307 = _RAND_883[3:0];
  _RAND_884 = {1{`RANDOM}};
  image_1_308 = _RAND_884[3:0];
  _RAND_885 = {1{`RANDOM}};
  image_1_309 = _RAND_885[3:0];
  _RAND_886 = {1{`RANDOM}};
  image_1_310 = _RAND_886[3:0];
  _RAND_887 = {1{`RANDOM}};
  image_1_311 = _RAND_887[3:0];
  _RAND_888 = {1{`RANDOM}};
  image_1_312 = _RAND_888[3:0];
  _RAND_889 = {1{`RANDOM}};
  image_1_313 = _RAND_889[3:0];
  _RAND_890 = {1{`RANDOM}};
  image_1_314 = _RAND_890[3:0];
  _RAND_891 = {1{`RANDOM}};
  image_1_315 = _RAND_891[3:0];
  _RAND_892 = {1{`RANDOM}};
  image_1_316 = _RAND_892[3:0];
  _RAND_893 = {1{`RANDOM}};
  image_1_317 = _RAND_893[3:0];
  _RAND_894 = {1{`RANDOM}};
  image_1_318 = _RAND_894[3:0];
  _RAND_895 = {1{`RANDOM}};
  image_1_319 = _RAND_895[3:0];
  _RAND_896 = {1{`RANDOM}};
  image_1_320 = _RAND_896[3:0];
  _RAND_897 = {1{`RANDOM}};
  image_1_321 = _RAND_897[3:0];
  _RAND_898 = {1{`RANDOM}};
  image_1_322 = _RAND_898[3:0];
  _RAND_899 = {1{`RANDOM}};
  image_1_323 = _RAND_899[3:0];
  _RAND_900 = {1{`RANDOM}};
  image_1_324 = _RAND_900[3:0];
  _RAND_901 = {1{`RANDOM}};
  image_1_325 = _RAND_901[3:0];
  _RAND_902 = {1{`RANDOM}};
  image_1_326 = _RAND_902[3:0];
  _RAND_903 = {1{`RANDOM}};
  image_1_327 = _RAND_903[3:0];
  _RAND_904 = {1{`RANDOM}};
  image_1_328 = _RAND_904[3:0];
  _RAND_905 = {1{`RANDOM}};
  image_1_329 = _RAND_905[3:0];
  _RAND_906 = {1{`RANDOM}};
  image_1_330 = _RAND_906[3:0];
  _RAND_907 = {1{`RANDOM}};
  image_1_331 = _RAND_907[3:0];
  _RAND_908 = {1{`RANDOM}};
  image_1_332 = _RAND_908[3:0];
  _RAND_909 = {1{`RANDOM}};
  image_1_333 = _RAND_909[3:0];
  _RAND_910 = {1{`RANDOM}};
  image_1_334 = _RAND_910[3:0];
  _RAND_911 = {1{`RANDOM}};
  image_1_335 = _RAND_911[3:0];
  _RAND_912 = {1{`RANDOM}};
  image_1_336 = _RAND_912[3:0];
  _RAND_913 = {1{`RANDOM}};
  image_1_337 = _RAND_913[3:0];
  _RAND_914 = {1{`RANDOM}};
  image_1_338 = _RAND_914[3:0];
  _RAND_915 = {1{`RANDOM}};
  image_1_339 = _RAND_915[3:0];
  _RAND_916 = {1{`RANDOM}};
  image_1_340 = _RAND_916[3:0];
  _RAND_917 = {1{`RANDOM}};
  image_1_341 = _RAND_917[3:0];
  _RAND_918 = {1{`RANDOM}};
  image_1_342 = _RAND_918[3:0];
  _RAND_919 = {1{`RANDOM}};
  image_1_343 = _RAND_919[3:0];
  _RAND_920 = {1{`RANDOM}};
  image_1_344 = _RAND_920[3:0];
  _RAND_921 = {1{`RANDOM}};
  image_1_345 = _RAND_921[3:0];
  _RAND_922 = {1{`RANDOM}};
  image_1_346 = _RAND_922[3:0];
  _RAND_923 = {1{`RANDOM}};
  image_1_347 = _RAND_923[3:0];
  _RAND_924 = {1{`RANDOM}};
  image_1_348 = _RAND_924[3:0];
  _RAND_925 = {1{`RANDOM}};
  image_1_349 = _RAND_925[3:0];
  _RAND_926 = {1{`RANDOM}};
  image_1_350 = _RAND_926[3:0];
  _RAND_927 = {1{`RANDOM}};
  image_1_351 = _RAND_927[3:0];
  _RAND_928 = {1{`RANDOM}};
  image_1_352 = _RAND_928[3:0];
  _RAND_929 = {1{`RANDOM}};
  image_1_353 = _RAND_929[3:0];
  _RAND_930 = {1{`RANDOM}};
  image_1_354 = _RAND_930[3:0];
  _RAND_931 = {1{`RANDOM}};
  image_1_355 = _RAND_931[3:0];
  _RAND_932 = {1{`RANDOM}};
  image_1_356 = _RAND_932[3:0];
  _RAND_933 = {1{`RANDOM}};
  image_1_357 = _RAND_933[3:0];
  _RAND_934 = {1{`RANDOM}};
  image_1_358 = _RAND_934[3:0];
  _RAND_935 = {1{`RANDOM}};
  image_1_359 = _RAND_935[3:0];
  _RAND_936 = {1{`RANDOM}};
  image_1_360 = _RAND_936[3:0];
  _RAND_937 = {1{`RANDOM}};
  image_1_361 = _RAND_937[3:0];
  _RAND_938 = {1{`RANDOM}};
  image_1_362 = _RAND_938[3:0];
  _RAND_939 = {1{`RANDOM}};
  image_1_363 = _RAND_939[3:0];
  _RAND_940 = {1{`RANDOM}};
  image_1_364 = _RAND_940[3:0];
  _RAND_941 = {1{`RANDOM}};
  image_1_365 = _RAND_941[3:0];
  _RAND_942 = {1{`RANDOM}};
  image_1_366 = _RAND_942[3:0];
  _RAND_943 = {1{`RANDOM}};
  image_1_367 = _RAND_943[3:0];
  _RAND_944 = {1{`RANDOM}};
  image_1_368 = _RAND_944[3:0];
  _RAND_945 = {1{`RANDOM}};
  image_1_369 = _RAND_945[3:0];
  _RAND_946 = {1{`RANDOM}};
  image_1_370 = _RAND_946[3:0];
  _RAND_947 = {1{`RANDOM}};
  image_1_371 = _RAND_947[3:0];
  _RAND_948 = {1{`RANDOM}};
  image_1_372 = _RAND_948[3:0];
  _RAND_949 = {1{`RANDOM}};
  image_1_373 = _RAND_949[3:0];
  _RAND_950 = {1{`RANDOM}};
  image_1_374 = _RAND_950[3:0];
  _RAND_951 = {1{`RANDOM}};
  image_1_375 = _RAND_951[3:0];
  _RAND_952 = {1{`RANDOM}};
  image_1_376 = _RAND_952[3:0];
  _RAND_953 = {1{`RANDOM}};
  image_1_377 = _RAND_953[3:0];
  _RAND_954 = {1{`RANDOM}};
  image_1_378 = _RAND_954[3:0];
  _RAND_955 = {1{`RANDOM}};
  image_1_379 = _RAND_955[3:0];
  _RAND_956 = {1{`RANDOM}};
  image_1_380 = _RAND_956[3:0];
  _RAND_957 = {1{`RANDOM}};
  image_1_381 = _RAND_957[3:0];
  _RAND_958 = {1{`RANDOM}};
  image_1_382 = _RAND_958[3:0];
  _RAND_959 = {1{`RANDOM}};
  image_1_383 = _RAND_959[3:0];
  _RAND_960 = {1{`RANDOM}};
  image_1_384 = _RAND_960[3:0];
  _RAND_961 = {1{`RANDOM}};
  image_1_385 = _RAND_961[3:0];
  _RAND_962 = {1{`RANDOM}};
  image_1_386 = _RAND_962[3:0];
  _RAND_963 = {1{`RANDOM}};
  image_1_387 = _RAND_963[3:0];
  _RAND_964 = {1{`RANDOM}};
  image_1_388 = _RAND_964[3:0];
  _RAND_965 = {1{`RANDOM}};
  image_1_389 = _RAND_965[3:0];
  _RAND_966 = {1{`RANDOM}};
  image_1_390 = _RAND_966[3:0];
  _RAND_967 = {1{`RANDOM}};
  image_1_391 = _RAND_967[3:0];
  _RAND_968 = {1{`RANDOM}};
  image_1_392 = _RAND_968[3:0];
  _RAND_969 = {1{`RANDOM}};
  image_1_393 = _RAND_969[3:0];
  _RAND_970 = {1{`RANDOM}};
  image_1_394 = _RAND_970[3:0];
  _RAND_971 = {1{`RANDOM}};
  image_1_395 = _RAND_971[3:0];
  _RAND_972 = {1{`RANDOM}};
  image_1_396 = _RAND_972[3:0];
  _RAND_973 = {1{`RANDOM}};
  image_1_397 = _RAND_973[3:0];
  _RAND_974 = {1{`RANDOM}};
  image_1_398 = _RAND_974[3:0];
  _RAND_975 = {1{`RANDOM}};
  image_1_399 = _RAND_975[3:0];
  _RAND_976 = {1{`RANDOM}};
  image_1_400 = _RAND_976[3:0];
  _RAND_977 = {1{`RANDOM}};
  image_1_401 = _RAND_977[3:0];
  _RAND_978 = {1{`RANDOM}};
  image_1_402 = _RAND_978[3:0];
  _RAND_979 = {1{`RANDOM}};
  image_1_403 = _RAND_979[3:0];
  _RAND_980 = {1{`RANDOM}};
  image_1_404 = _RAND_980[3:0];
  _RAND_981 = {1{`RANDOM}};
  image_1_405 = _RAND_981[3:0];
  _RAND_982 = {1{`RANDOM}};
  image_1_406 = _RAND_982[3:0];
  _RAND_983 = {1{`RANDOM}};
  image_1_407 = _RAND_983[3:0];
  _RAND_984 = {1{`RANDOM}};
  image_1_408 = _RAND_984[3:0];
  _RAND_985 = {1{`RANDOM}};
  image_1_409 = _RAND_985[3:0];
  _RAND_986 = {1{`RANDOM}};
  image_1_410 = _RAND_986[3:0];
  _RAND_987 = {1{`RANDOM}};
  image_1_411 = _RAND_987[3:0];
  _RAND_988 = {1{`RANDOM}};
  image_1_412 = _RAND_988[3:0];
  _RAND_989 = {1{`RANDOM}};
  image_1_413 = _RAND_989[3:0];
  _RAND_990 = {1{`RANDOM}};
  image_1_414 = _RAND_990[3:0];
  _RAND_991 = {1{`RANDOM}};
  image_1_415 = _RAND_991[3:0];
  _RAND_992 = {1{`RANDOM}};
  image_1_416 = _RAND_992[3:0];
  _RAND_993 = {1{`RANDOM}};
  image_1_417 = _RAND_993[3:0];
  _RAND_994 = {1{`RANDOM}};
  image_1_418 = _RAND_994[3:0];
  _RAND_995 = {1{`RANDOM}};
  image_1_419 = _RAND_995[3:0];
  _RAND_996 = {1{`RANDOM}};
  image_1_420 = _RAND_996[3:0];
  _RAND_997 = {1{`RANDOM}};
  image_1_421 = _RAND_997[3:0];
  _RAND_998 = {1{`RANDOM}};
  image_1_422 = _RAND_998[3:0];
  _RAND_999 = {1{`RANDOM}};
  image_1_423 = _RAND_999[3:0];
  _RAND_1000 = {1{`RANDOM}};
  image_1_424 = _RAND_1000[3:0];
  _RAND_1001 = {1{`RANDOM}};
  image_1_425 = _RAND_1001[3:0];
  _RAND_1002 = {1{`RANDOM}};
  image_1_426 = _RAND_1002[3:0];
  _RAND_1003 = {1{`RANDOM}};
  image_1_427 = _RAND_1003[3:0];
  _RAND_1004 = {1{`RANDOM}};
  image_1_428 = _RAND_1004[3:0];
  _RAND_1005 = {1{`RANDOM}};
  image_1_429 = _RAND_1005[3:0];
  _RAND_1006 = {1{`RANDOM}};
  image_1_430 = _RAND_1006[3:0];
  _RAND_1007 = {1{`RANDOM}};
  image_1_431 = _RAND_1007[3:0];
  _RAND_1008 = {1{`RANDOM}};
  image_1_432 = _RAND_1008[3:0];
  _RAND_1009 = {1{`RANDOM}};
  image_1_433 = _RAND_1009[3:0];
  _RAND_1010 = {1{`RANDOM}};
  image_1_434 = _RAND_1010[3:0];
  _RAND_1011 = {1{`RANDOM}};
  image_1_435 = _RAND_1011[3:0];
  _RAND_1012 = {1{`RANDOM}};
  image_1_436 = _RAND_1012[3:0];
  _RAND_1013 = {1{`RANDOM}};
  image_1_437 = _RAND_1013[3:0];
  _RAND_1014 = {1{`RANDOM}};
  image_1_438 = _RAND_1014[3:0];
  _RAND_1015 = {1{`RANDOM}};
  image_1_439 = _RAND_1015[3:0];
  _RAND_1016 = {1{`RANDOM}};
  image_1_440 = _RAND_1016[3:0];
  _RAND_1017 = {1{`RANDOM}};
  image_1_441 = _RAND_1017[3:0];
  _RAND_1018 = {1{`RANDOM}};
  image_1_442 = _RAND_1018[3:0];
  _RAND_1019 = {1{`RANDOM}};
  image_1_443 = _RAND_1019[3:0];
  _RAND_1020 = {1{`RANDOM}};
  image_1_444 = _RAND_1020[3:0];
  _RAND_1021 = {1{`RANDOM}};
  image_1_445 = _RAND_1021[3:0];
  _RAND_1022 = {1{`RANDOM}};
  image_1_446 = _RAND_1022[3:0];
  _RAND_1023 = {1{`RANDOM}};
  image_1_447 = _RAND_1023[3:0];
  _RAND_1024 = {1{`RANDOM}};
  image_1_448 = _RAND_1024[3:0];
  _RAND_1025 = {1{`RANDOM}};
  image_1_449 = _RAND_1025[3:0];
  _RAND_1026 = {1{`RANDOM}};
  image_1_450 = _RAND_1026[3:0];
  _RAND_1027 = {1{`RANDOM}};
  image_1_451 = _RAND_1027[3:0];
  _RAND_1028 = {1{`RANDOM}};
  image_1_452 = _RAND_1028[3:0];
  _RAND_1029 = {1{`RANDOM}};
  image_1_453 = _RAND_1029[3:0];
  _RAND_1030 = {1{`RANDOM}};
  image_1_454 = _RAND_1030[3:0];
  _RAND_1031 = {1{`RANDOM}};
  image_1_455 = _RAND_1031[3:0];
  _RAND_1032 = {1{`RANDOM}};
  image_1_456 = _RAND_1032[3:0];
  _RAND_1033 = {1{`RANDOM}};
  image_1_457 = _RAND_1033[3:0];
  _RAND_1034 = {1{`RANDOM}};
  image_1_458 = _RAND_1034[3:0];
  _RAND_1035 = {1{`RANDOM}};
  image_1_459 = _RAND_1035[3:0];
  _RAND_1036 = {1{`RANDOM}};
  image_1_460 = _RAND_1036[3:0];
  _RAND_1037 = {1{`RANDOM}};
  image_1_461 = _RAND_1037[3:0];
  _RAND_1038 = {1{`RANDOM}};
  image_1_462 = _RAND_1038[3:0];
  _RAND_1039 = {1{`RANDOM}};
  image_1_463 = _RAND_1039[3:0];
  _RAND_1040 = {1{`RANDOM}};
  image_1_464 = _RAND_1040[3:0];
  _RAND_1041 = {1{`RANDOM}};
  image_1_465 = _RAND_1041[3:0];
  _RAND_1042 = {1{`RANDOM}};
  image_1_466 = _RAND_1042[3:0];
  _RAND_1043 = {1{`RANDOM}};
  image_1_467 = _RAND_1043[3:0];
  _RAND_1044 = {1{`RANDOM}};
  image_1_468 = _RAND_1044[3:0];
  _RAND_1045 = {1{`RANDOM}};
  image_1_469 = _RAND_1045[3:0];
  _RAND_1046 = {1{`RANDOM}};
  image_1_470 = _RAND_1046[3:0];
  _RAND_1047 = {1{`RANDOM}};
  image_1_471 = _RAND_1047[3:0];
  _RAND_1048 = {1{`RANDOM}};
  image_1_472 = _RAND_1048[3:0];
  _RAND_1049 = {1{`RANDOM}};
  image_1_473 = _RAND_1049[3:0];
  _RAND_1050 = {1{`RANDOM}};
  image_1_474 = _RAND_1050[3:0];
  _RAND_1051 = {1{`RANDOM}};
  image_1_475 = _RAND_1051[3:0];
  _RAND_1052 = {1{`RANDOM}};
  image_1_476 = _RAND_1052[3:0];
  _RAND_1053 = {1{`RANDOM}};
  image_1_477 = _RAND_1053[3:0];
  _RAND_1054 = {1{`RANDOM}};
  image_1_478 = _RAND_1054[3:0];
  _RAND_1055 = {1{`RANDOM}};
  image_1_479 = _RAND_1055[3:0];
  _RAND_1056 = {1{`RANDOM}};
  image_1_480 = _RAND_1056[3:0];
  _RAND_1057 = {1{`RANDOM}};
  image_1_481 = _RAND_1057[3:0];
  _RAND_1058 = {1{`RANDOM}};
  image_1_482 = _RAND_1058[3:0];
  _RAND_1059 = {1{`RANDOM}};
  image_1_483 = _RAND_1059[3:0];
  _RAND_1060 = {1{`RANDOM}};
  image_1_484 = _RAND_1060[3:0];
  _RAND_1061 = {1{`RANDOM}};
  image_1_485 = _RAND_1061[3:0];
  _RAND_1062 = {1{`RANDOM}};
  image_1_486 = _RAND_1062[3:0];
  _RAND_1063 = {1{`RANDOM}};
  image_1_487 = _RAND_1063[3:0];
  _RAND_1064 = {1{`RANDOM}};
  image_1_488 = _RAND_1064[3:0];
  _RAND_1065 = {1{`RANDOM}};
  image_1_489 = _RAND_1065[3:0];
  _RAND_1066 = {1{`RANDOM}};
  image_1_490 = _RAND_1066[3:0];
  _RAND_1067 = {1{`RANDOM}};
  image_1_491 = _RAND_1067[3:0];
  _RAND_1068 = {1{`RANDOM}};
  image_1_492 = _RAND_1068[3:0];
  _RAND_1069 = {1{`RANDOM}};
  image_1_493 = _RAND_1069[3:0];
  _RAND_1070 = {1{`RANDOM}};
  image_1_494 = _RAND_1070[3:0];
  _RAND_1071 = {1{`RANDOM}};
  image_1_495 = _RAND_1071[3:0];
  _RAND_1072 = {1{`RANDOM}};
  image_1_496 = _RAND_1072[3:0];
  _RAND_1073 = {1{`RANDOM}};
  image_1_497 = _RAND_1073[3:0];
  _RAND_1074 = {1{`RANDOM}};
  image_1_498 = _RAND_1074[3:0];
  _RAND_1075 = {1{`RANDOM}};
  image_1_499 = _RAND_1075[3:0];
  _RAND_1076 = {1{`RANDOM}};
  image_1_500 = _RAND_1076[3:0];
  _RAND_1077 = {1{`RANDOM}};
  image_1_501 = _RAND_1077[3:0];
  _RAND_1078 = {1{`RANDOM}};
  image_1_502 = _RAND_1078[3:0];
  _RAND_1079 = {1{`RANDOM}};
  image_1_503 = _RAND_1079[3:0];
  _RAND_1080 = {1{`RANDOM}};
  image_1_504 = _RAND_1080[3:0];
  _RAND_1081 = {1{`RANDOM}};
  image_1_505 = _RAND_1081[3:0];
  _RAND_1082 = {1{`RANDOM}};
  image_1_506 = _RAND_1082[3:0];
  _RAND_1083 = {1{`RANDOM}};
  image_1_507 = _RAND_1083[3:0];
  _RAND_1084 = {1{`RANDOM}};
  image_1_508 = _RAND_1084[3:0];
  _RAND_1085 = {1{`RANDOM}};
  image_1_509 = _RAND_1085[3:0];
  _RAND_1086 = {1{`RANDOM}};
  image_1_510 = _RAND_1086[3:0];
  _RAND_1087 = {1{`RANDOM}};
  image_1_511 = _RAND_1087[3:0];
  _RAND_1088 = {1{`RANDOM}};
  image_1_512 = _RAND_1088[3:0];
  _RAND_1089 = {1{`RANDOM}};
  image_1_513 = _RAND_1089[3:0];
  _RAND_1090 = {1{`RANDOM}};
  image_1_514 = _RAND_1090[3:0];
  _RAND_1091 = {1{`RANDOM}};
  image_1_515 = _RAND_1091[3:0];
  _RAND_1092 = {1{`RANDOM}};
  image_1_516 = _RAND_1092[3:0];
  _RAND_1093 = {1{`RANDOM}};
  image_1_517 = _RAND_1093[3:0];
  _RAND_1094 = {1{`RANDOM}};
  image_1_518 = _RAND_1094[3:0];
  _RAND_1095 = {1{`RANDOM}};
  image_1_519 = _RAND_1095[3:0];
  _RAND_1096 = {1{`RANDOM}};
  image_1_520 = _RAND_1096[3:0];
  _RAND_1097 = {1{`RANDOM}};
  image_1_521 = _RAND_1097[3:0];
  _RAND_1098 = {1{`RANDOM}};
  image_1_522 = _RAND_1098[3:0];
  _RAND_1099 = {1{`RANDOM}};
  image_1_523 = _RAND_1099[3:0];
  _RAND_1100 = {1{`RANDOM}};
  image_1_524 = _RAND_1100[3:0];
  _RAND_1101 = {1{`RANDOM}};
  image_1_525 = _RAND_1101[3:0];
  _RAND_1102 = {1{`RANDOM}};
  image_1_526 = _RAND_1102[3:0];
  _RAND_1103 = {1{`RANDOM}};
  image_1_527 = _RAND_1103[3:0];
  _RAND_1104 = {1{`RANDOM}};
  image_1_528 = _RAND_1104[3:0];
  _RAND_1105 = {1{`RANDOM}};
  image_1_529 = _RAND_1105[3:0];
  _RAND_1106 = {1{`RANDOM}};
  image_1_530 = _RAND_1106[3:0];
  _RAND_1107 = {1{`RANDOM}};
  image_1_531 = _RAND_1107[3:0];
  _RAND_1108 = {1{`RANDOM}};
  image_1_532 = _RAND_1108[3:0];
  _RAND_1109 = {1{`RANDOM}};
  image_1_533 = _RAND_1109[3:0];
  _RAND_1110 = {1{`RANDOM}};
  image_1_534 = _RAND_1110[3:0];
  _RAND_1111 = {1{`RANDOM}};
  image_1_535 = _RAND_1111[3:0];
  _RAND_1112 = {1{`RANDOM}};
  image_1_536 = _RAND_1112[3:0];
  _RAND_1113 = {1{`RANDOM}};
  image_1_537 = _RAND_1113[3:0];
  _RAND_1114 = {1{`RANDOM}};
  image_1_538 = _RAND_1114[3:0];
  _RAND_1115 = {1{`RANDOM}};
  image_1_539 = _RAND_1115[3:0];
  _RAND_1116 = {1{`RANDOM}};
  image_1_540 = _RAND_1116[3:0];
  _RAND_1117 = {1{`RANDOM}};
  image_1_541 = _RAND_1117[3:0];
  _RAND_1118 = {1{`RANDOM}};
  image_1_542 = _RAND_1118[3:0];
  _RAND_1119 = {1{`RANDOM}};
  image_1_543 = _RAND_1119[3:0];
  _RAND_1120 = {1{`RANDOM}};
  image_1_544 = _RAND_1120[3:0];
  _RAND_1121 = {1{`RANDOM}};
  image_1_545 = _RAND_1121[3:0];
  _RAND_1122 = {1{`RANDOM}};
  image_1_546 = _RAND_1122[3:0];
  _RAND_1123 = {1{`RANDOM}};
  image_1_547 = _RAND_1123[3:0];
  _RAND_1124 = {1{`RANDOM}};
  image_1_548 = _RAND_1124[3:0];
  _RAND_1125 = {1{`RANDOM}};
  image_1_549 = _RAND_1125[3:0];
  _RAND_1126 = {1{`RANDOM}};
  image_1_550 = _RAND_1126[3:0];
  _RAND_1127 = {1{`RANDOM}};
  image_1_551 = _RAND_1127[3:0];
  _RAND_1128 = {1{`RANDOM}};
  image_1_552 = _RAND_1128[3:0];
  _RAND_1129 = {1{`RANDOM}};
  image_1_553 = _RAND_1129[3:0];
  _RAND_1130 = {1{`RANDOM}};
  image_1_554 = _RAND_1130[3:0];
  _RAND_1131 = {1{`RANDOM}};
  image_1_555 = _RAND_1131[3:0];
  _RAND_1132 = {1{`RANDOM}};
  image_1_556 = _RAND_1132[3:0];
  _RAND_1133 = {1{`RANDOM}};
  image_1_557 = _RAND_1133[3:0];
  _RAND_1134 = {1{`RANDOM}};
  image_1_558 = _RAND_1134[3:0];
  _RAND_1135 = {1{`RANDOM}};
  image_1_559 = _RAND_1135[3:0];
  _RAND_1136 = {1{`RANDOM}};
  image_1_560 = _RAND_1136[3:0];
  _RAND_1137 = {1{`RANDOM}};
  image_1_561 = _RAND_1137[3:0];
  _RAND_1138 = {1{`RANDOM}};
  image_1_562 = _RAND_1138[3:0];
  _RAND_1139 = {1{`RANDOM}};
  image_1_563 = _RAND_1139[3:0];
  _RAND_1140 = {1{`RANDOM}};
  image_1_564 = _RAND_1140[3:0];
  _RAND_1141 = {1{`RANDOM}};
  image_1_565 = _RAND_1141[3:0];
  _RAND_1142 = {1{`RANDOM}};
  image_1_566 = _RAND_1142[3:0];
  _RAND_1143 = {1{`RANDOM}};
  image_1_567 = _RAND_1143[3:0];
  _RAND_1144 = {1{`RANDOM}};
  image_1_568 = _RAND_1144[3:0];
  _RAND_1145 = {1{`RANDOM}};
  image_1_569 = _RAND_1145[3:0];
  _RAND_1146 = {1{`RANDOM}};
  image_1_570 = _RAND_1146[3:0];
  _RAND_1147 = {1{`RANDOM}};
  image_1_571 = _RAND_1147[3:0];
  _RAND_1148 = {1{`RANDOM}};
  image_1_572 = _RAND_1148[3:0];
  _RAND_1149 = {1{`RANDOM}};
  image_1_573 = _RAND_1149[3:0];
  _RAND_1150 = {1{`RANDOM}};
  image_1_574 = _RAND_1150[3:0];
  _RAND_1151 = {1{`RANDOM}};
  image_1_575 = _RAND_1151[3:0];
  _RAND_1152 = {1{`RANDOM}};
  image_2_0 = _RAND_1152[3:0];
  _RAND_1153 = {1{`RANDOM}};
  image_2_1 = _RAND_1153[3:0];
  _RAND_1154 = {1{`RANDOM}};
  image_2_2 = _RAND_1154[3:0];
  _RAND_1155 = {1{`RANDOM}};
  image_2_3 = _RAND_1155[3:0];
  _RAND_1156 = {1{`RANDOM}};
  image_2_4 = _RAND_1156[3:0];
  _RAND_1157 = {1{`RANDOM}};
  image_2_5 = _RAND_1157[3:0];
  _RAND_1158 = {1{`RANDOM}};
  image_2_6 = _RAND_1158[3:0];
  _RAND_1159 = {1{`RANDOM}};
  image_2_7 = _RAND_1159[3:0];
  _RAND_1160 = {1{`RANDOM}};
  image_2_8 = _RAND_1160[3:0];
  _RAND_1161 = {1{`RANDOM}};
  image_2_9 = _RAND_1161[3:0];
  _RAND_1162 = {1{`RANDOM}};
  image_2_10 = _RAND_1162[3:0];
  _RAND_1163 = {1{`RANDOM}};
  image_2_11 = _RAND_1163[3:0];
  _RAND_1164 = {1{`RANDOM}};
  image_2_12 = _RAND_1164[3:0];
  _RAND_1165 = {1{`RANDOM}};
  image_2_13 = _RAND_1165[3:0];
  _RAND_1166 = {1{`RANDOM}};
  image_2_14 = _RAND_1166[3:0];
  _RAND_1167 = {1{`RANDOM}};
  image_2_15 = _RAND_1167[3:0];
  _RAND_1168 = {1{`RANDOM}};
  image_2_16 = _RAND_1168[3:0];
  _RAND_1169 = {1{`RANDOM}};
  image_2_17 = _RAND_1169[3:0];
  _RAND_1170 = {1{`RANDOM}};
  image_2_18 = _RAND_1170[3:0];
  _RAND_1171 = {1{`RANDOM}};
  image_2_19 = _RAND_1171[3:0];
  _RAND_1172 = {1{`RANDOM}};
  image_2_20 = _RAND_1172[3:0];
  _RAND_1173 = {1{`RANDOM}};
  image_2_21 = _RAND_1173[3:0];
  _RAND_1174 = {1{`RANDOM}};
  image_2_22 = _RAND_1174[3:0];
  _RAND_1175 = {1{`RANDOM}};
  image_2_23 = _RAND_1175[3:0];
  _RAND_1176 = {1{`RANDOM}};
  image_2_24 = _RAND_1176[3:0];
  _RAND_1177 = {1{`RANDOM}};
  image_2_25 = _RAND_1177[3:0];
  _RAND_1178 = {1{`RANDOM}};
  image_2_26 = _RAND_1178[3:0];
  _RAND_1179 = {1{`RANDOM}};
  image_2_27 = _RAND_1179[3:0];
  _RAND_1180 = {1{`RANDOM}};
  image_2_28 = _RAND_1180[3:0];
  _RAND_1181 = {1{`RANDOM}};
  image_2_29 = _RAND_1181[3:0];
  _RAND_1182 = {1{`RANDOM}};
  image_2_30 = _RAND_1182[3:0];
  _RAND_1183 = {1{`RANDOM}};
  image_2_31 = _RAND_1183[3:0];
  _RAND_1184 = {1{`RANDOM}};
  image_2_32 = _RAND_1184[3:0];
  _RAND_1185 = {1{`RANDOM}};
  image_2_33 = _RAND_1185[3:0];
  _RAND_1186 = {1{`RANDOM}};
  image_2_34 = _RAND_1186[3:0];
  _RAND_1187 = {1{`RANDOM}};
  image_2_35 = _RAND_1187[3:0];
  _RAND_1188 = {1{`RANDOM}};
  image_2_36 = _RAND_1188[3:0];
  _RAND_1189 = {1{`RANDOM}};
  image_2_37 = _RAND_1189[3:0];
  _RAND_1190 = {1{`RANDOM}};
  image_2_38 = _RAND_1190[3:0];
  _RAND_1191 = {1{`RANDOM}};
  image_2_39 = _RAND_1191[3:0];
  _RAND_1192 = {1{`RANDOM}};
  image_2_40 = _RAND_1192[3:0];
  _RAND_1193 = {1{`RANDOM}};
  image_2_41 = _RAND_1193[3:0];
  _RAND_1194 = {1{`RANDOM}};
  image_2_42 = _RAND_1194[3:0];
  _RAND_1195 = {1{`RANDOM}};
  image_2_43 = _RAND_1195[3:0];
  _RAND_1196 = {1{`RANDOM}};
  image_2_44 = _RAND_1196[3:0];
  _RAND_1197 = {1{`RANDOM}};
  image_2_45 = _RAND_1197[3:0];
  _RAND_1198 = {1{`RANDOM}};
  image_2_46 = _RAND_1198[3:0];
  _RAND_1199 = {1{`RANDOM}};
  image_2_47 = _RAND_1199[3:0];
  _RAND_1200 = {1{`RANDOM}};
  image_2_48 = _RAND_1200[3:0];
  _RAND_1201 = {1{`RANDOM}};
  image_2_49 = _RAND_1201[3:0];
  _RAND_1202 = {1{`RANDOM}};
  image_2_50 = _RAND_1202[3:0];
  _RAND_1203 = {1{`RANDOM}};
  image_2_51 = _RAND_1203[3:0];
  _RAND_1204 = {1{`RANDOM}};
  image_2_52 = _RAND_1204[3:0];
  _RAND_1205 = {1{`RANDOM}};
  image_2_53 = _RAND_1205[3:0];
  _RAND_1206 = {1{`RANDOM}};
  image_2_54 = _RAND_1206[3:0];
  _RAND_1207 = {1{`RANDOM}};
  image_2_55 = _RAND_1207[3:0];
  _RAND_1208 = {1{`RANDOM}};
  image_2_56 = _RAND_1208[3:0];
  _RAND_1209 = {1{`RANDOM}};
  image_2_57 = _RAND_1209[3:0];
  _RAND_1210 = {1{`RANDOM}};
  image_2_58 = _RAND_1210[3:0];
  _RAND_1211 = {1{`RANDOM}};
  image_2_59 = _RAND_1211[3:0];
  _RAND_1212 = {1{`RANDOM}};
  image_2_60 = _RAND_1212[3:0];
  _RAND_1213 = {1{`RANDOM}};
  image_2_61 = _RAND_1213[3:0];
  _RAND_1214 = {1{`RANDOM}};
  image_2_62 = _RAND_1214[3:0];
  _RAND_1215 = {1{`RANDOM}};
  image_2_63 = _RAND_1215[3:0];
  _RAND_1216 = {1{`RANDOM}};
  image_2_64 = _RAND_1216[3:0];
  _RAND_1217 = {1{`RANDOM}};
  image_2_65 = _RAND_1217[3:0];
  _RAND_1218 = {1{`RANDOM}};
  image_2_66 = _RAND_1218[3:0];
  _RAND_1219 = {1{`RANDOM}};
  image_2_67 = _RAND_1219[3:0];
  _RAND_1220 = {1{`RANDOM}};
  image_2_68 = _RAND_1220[3:0];
  _RAND_1221 = {1{`RANDOM}};
  image_2_69 = _RAND_1221[3:0];
  _RAND_1222 = {1{`RANDOM}};
  image_2_70 = _RAND_1222[3:0];
  _RAND_1223 = {1{`RANDOM}};
  image_2_71 = _RAND_1223[3:0];
  _RAND_1224 = {1{`RANDOM}};
  image_2_72 = _RAND_1224[3:0];
  _RAND_1225 = {1{`RANDOM}};
  image_2_73 = _RAND_1225[3:0];
  _RAND_1226 = {1{`RANDOM}};
  image_2_74 = _RAND_1226[3:0];
  _RAND_1227 = {1{`RANDOM}};
  image_2_75 = _RAND_1227[3:0];
  _RAND_1228 = {1{`RANDOM}};
  image_2_76 = _RAND_1228[3:0];
  _RAND_1229 = {1{`RANDOM}};
  image_2_77 = _RAND_1229[3:0];
  _RAND_1230 = {1{`RANDOM}};
  image_2_78 = _RAND_1230[3:0];
  _RAND_1231 = {1{`RANDOM}};
  image_2_79 = _RAND_1231[3:0];
  _RAND_1232 = {1{`RANDOM}};
  image_2_80 = _RAND_1232[3:0];
  _RAND_1233 = {1{`RANDOM}};
  image_2_81 = _RAND_1233[3:0];
  _RAND_1234 = {1{`RANDOM}};
  image_2_82 = _RAND_1234[3:0];
  _RAND_1235 = {1{`RANDOM}};
  image_2_83 = _RAND_1235[3:0];
  _RAND_1236 = {1{`RANDOM}};
  image_2_84 = _RAND_1236[3:0];
  _RAND_1237 = {1{`RANDOM}};
  image_2_85 = _RAND_1237[3:0];
  _RAND_1238 = {1{`RANDOM}};
  image_2_86 = _RAND_1238[3:0];
  _RAND_1239 = {1{`RANDOM}};
  image_2_87 = _RAND_1239[3:0];
  _RAND_1240 = {1{`RANDOM}};
  image_2_88 = _RAND_1240[3:0];
  _RAND_1241 = {1{`RANDOM}};
  image_2_89 = _RAND_1241[3:0];
  _RAND_1242 = {1{`RANDOM}};
  image_2_90 = _RAND_1242[3:0];
  _RAND_1243 = {1{`RANDOM}};
  image_2_91 = _RAND_1243[3:0];
  _RAND_1244 = {1{`RANDOM}};
  image_2_92 = _RAND_1244[3:0];
  _RAND_1245 = {1{`RANDOM}};
  image_2_93 = _RAND_1245[3:0];
  _RAND_1246 = {1{`RANDOM}};
  image_2_94 = _RAND_1246[3:0];
  _RAND_1247 = {1{`RANDOM}};
  image_2_95 = _RAND_1247[3:0];
  _RAND_1248 = {1{`RANDOM}};
  image_2_96 = _RAND_1248[3:0];
  _RAND_1249 = {1{`RANDOM}};
  image_2_97 = _RAND_1249[3:0];
  _RAND_1250 = {1{`RANDOM}};
  image_2_98 = _RAND_1250[3:0];
  _RAND_1251 = {1{`RANDOM}};
  image_2_99 = _RAND_1251[3:0];
  _RAND_1252 = {1{`RANDOM}};
  image_2_100 = _RAND_1252[3:0];
  _RAND_1253 = {1{`RANDOM}};
  image_2_101 = _RAND_1253[3:0];
  _RAND_1254 = {1{`RANDOM}};
  image_2_102 = _RAND_1254[3:0];
  _RAND_1255 = {1{`RANDOM}};
  image_2_103 = _RAND_1255[3:0];
  _RAND_1256 = {1{`RANDOM}};
  image_2_104 = _RAND_1256[3:0];
  _RAND_1257 = {1{`RANDOM}};
  image_2_105 = _RAND_1257[3:0];
  _RAND_1258 = {1{`RANDOM}};
  image_2_106 = _RAND_1258[3:0];
  _RAND_1259 = {1{`RANDOM}};
  image_2_107 = _RAND_1259[3:0];
  _RAND_1260 = {1{`RANDOM}};
  image_2_108 = _RAND_1260[3:0];
  _RAND_1261 = {1{`RANDOM}};
  image_2_109 = _RAND_1261[3:0];
  _RAND_1262 = {1{`RANDOM}};
  image_2_110 = _RAND_1262[3:0];
  _RAND_1263 = {1{`RANDOM}};
  image_2_111 = _RAND_1263[3:0];
  _RAND_1264 = {1{`RANDOM}};
  image_2_112 = _RAND_1264[3:0];
  _RAND_1265 = {1{`RANDOM}};
  image_2_113 = _RAND_1265[3:0];
  _RAND_1266 = {1{`RANDOM}};
  image_2_114 = _RAND_1266[3:0];
  _RAND_1267 = {1{`RANDOM}};
  image_2_115 = _RAND_1267[3:0];
  _RAND_1268 = {1{`RANDOM}};
  image_2_116 = _RAND_1268[3:0];
  _RAND_1269 = {1{`RANDOM}};
  image_2_117 = _RAND_1269[3:0];
  _RAND_1270 = {1{`RANDOM}};
  image_2_118 = _RAND_1270[3:0];
  _RAND_1271 = {1{`RANDOM}};
  image_2_119 = _RAND_1271[3:0];
  _RAND_1272 = {1{`RANDOM}};
  image_2_120 = _RAND_1272[3:0];
  _RAND_1273 = {1{`RANDOM}};
  image_2_121 = _RAND_1273[3:0];
  _RAND_1274 = {1{`RANDOM}};
  image_2_122 = _RAND_1274[3:0];
  _RAND_1275 = {1{`RANDOM}};
  image_2_123 = _RAND_1275[3:0];
  _RAND_1276 = {1{`RANDOM}};
  image_2_124 = _RAND_1276[3:0];
  _RAND_1277 = {1{`RANDOM}};
  image_2_125 = _RAND_1277[3:0];
  _RAND_1278 = {1{`RANDOM}};
  image_2_126 = _RAND_1278[3:0];
  _RAND_1279 = {1{`RANDOM}};
  image_2_127 = _RAND_1279[3:0];
  _RAND_1280 = {1{`RANDOM}};
  image_2_128 = _RAND_1280[3:0];
  _RAND_1281 = {1{`RANDOM}};
  image_2_129 = _RAND_1281[3:0];
  _RAND_1282 = {1{`RANDOM}};
  image_2_130 = _RAND_1282[3:0];
  _RAND_1283 = {1{`RANDOM}};
  image_2_131 = _RAND_1283[3:0];
  _RAND_1284 = {1{`RANDOM}};
  image_2_132 = _RAND_1284[3:0];
  _RAND_1285 = {1{`RANDOM}};
  image_2_133 = _RAND_1285[3:0];
  _RAND_1286 = {1{`RANDOM}};
  image_2_134 = _RAND_1286[3:0];
  _RAND_1287 = {1{`RANDOM}};
  image_2_135 = _RAND_1287[3:0];
  _RAND_1288 = {1{`RANDOM}};
  image_2_136 = _RAND_1288[3:0];
  _RAND_1289 = {1{`RANDOM}};
  image_2_137 = _RAND_1289[3:0];
  _RAND_1290 = {1{`RANDOM}};
  image_2_138 = _RAND_1290[3:0];
  _RAND_1291 = {1{`RANDOM}};
  image_2_139 = _RAND_1291[3:0];
  _RAND_1292 = {1{`RANDOM}};
  image_2_140 = _RAND_1292[3:0];
  _RAND_1293 = {1{`RANDOM}};
  image_2_141 = _RAND_1293[3:0];
  _RAND_1294 = {1{`RANDOM}};
  image_2_142 = _RAND_1294[3:0];
  _RAND_1295 = {1{`RANDOM}};
  image_2_143 = _RAND_1295[3:0];
  _RAND_1296 = {1{`RANDOM}};
  image_2_144 = _RAND_1296[3:0];
  _RAND_1297 = {1{`RANDOM}};
  image_2_145 = _RAND_1297[3:0];
  _RAND_1298 = {1{`RANDOM}};
  image_2_146 = _RAND_1298[3:0];
  _RAND_1299 = {1{`RANDOM}};
  image_2_147 = _RAND_1299[3:0];
  _RAND_1300 = {1{`RANDOM}};
  image_2_148 = _RAND_1300[3:0];
  _RAND_1301 = {1{`RANDOM}};
  image_2_149 = _RAND_1301[3:0];
  _RAND_1302 = {1{`RANDOM}};
  image_2_150 = _RAND_1302[3:0];
  _RAND_1303 = {1{`RANDOM}};
  image_2_151 = _RAND_1303[3:0];
  _RAND_1304 = {1{`RANDOM}};
  image_2_152 = _RAND_1304[3:0];
  _RAND_1305 = {1{`RANDOM}};
  image_2_153 = _RAND_1305[3:0];
  _RAND_1306 = {1{`RANDOM}};
  image_2_154 = _RAND_1306[3:0];
  _RAND_1307 = {1{`RANDOM}};
  image_2_155 = _RAND_1307[3:0];
  _RAND_1308 = {1{`RANDOM}};
  image_2_156 = _RAND_1308[3:0];
  _RAND_1309 = {1{`RANDOM}};
  image_2_157 = _RAND_1309[3:0];
  _RAND_1310 = {1{`RANDOM}};
  image_2_158 = _RAND_1310[3:0];
  _RAND_1311 = {1{`RANDOM}};
  image_2_159 = _RAND_1311[3:0];
  _RAND_1312 = {1{`RANDOM}};
  image_2_160 = _RAND_1312[3:0];
  _RAND_1313 = {1{`RANDOM}};
  image_2_161 = _RAND_1313[3:0];
  _RAND_1314 = {1{`RANDOM}};
  image_2_162 = _RAND_1314[3:0];
  _RAND_1315 = {1{`RANDOM}};
  image_2_163 = _RAND_1315[3:0];
  _RAND_1316 = {1{`RANDOM}};
  image_2_164 = _RAND_1316[3:0];
  _RAND_1317 = {1{`RANDOM}};
  image_2_165 = _RAND_1317[3:0];
  _RAND_1318 = {1{`RANDOM}};
  image_2_166 = _RAND_1318[3:0];
  _RAND_1319 = {1{`RANDOM}};
  image_2_167 = _RAND_1319[3:0];
  _RAND_1320 = {1{`RANDOM}};
  image_2_168 = _RAND_1320[3:0];
  _RAND_1321 = {1{`RANDOM}};
  image_2_169 = _RAND_1321[3:0];
  _RAND_1322 = {1{`RANDOM}};
  image_2_170 = _RAND_1322[3:0];
  _RAND_1323 = {1{`RANDOM}};
  image_2_171 = _RAND_1323[3:0];
  _RAND_1324 = {1{`RANDOM}};
  image_2_172 = _RAND_1324[3:0];
  _RAND_1325 = {1{`RANDOM}};
  image_2_173 = _RAND_1325[3:0];
  _RAND_1326 = {1{`RANDOM}};
  image_2_174 = _RAND_1326[3:0];
  _RAND_1327 = {1{`RANDOM}};
  image_2_175 = _RAND_1327[3:0];
  _RAND_1328 = {1{`RANDOM}};
  image_2_176 = _RAND_1328[3:0];
  _RAND_1329 = {1{`RANDOM}};
  image_2_177 = _RAND_1329[3:0];
  _RAND_1330 = {1{`RANDOM}};
  image_2_178 = _RAND_1330[3:0];
  _RAND_1331 = {1{`RANDOM}};
  image_2_179 = _RAND_1331[3:0];
  _RAND_1332 = {1{`RANDOM}};
  image_2_180 = _RAND_1332[3:0];
  _RAND_1333 = {1{`RANDOM}};
  image_2_181 = _RAND_1333[3:0];
  _RAND_1334 = {1{`RANDOM}};
  image_2_182 = _RAND_1334[3:0];
  _RAND_1335 = {1{`RANDOM}};
  image_2_183 = _RAND_1335[3:0];
  _RAND_1336 = {1{`RANDOM}};
  image_2_184 = _RAND_1336[3:0];
  _RAND_1337 = {1{`RANDOM}};
  image_2_185 = _RAND_1337[3:0];
  _RAND_1338 = {1{`RANDOM}};
  image_2_186 = _RAND_1338[3:0];
  _RAND_1339 = {1{`RANDOM}};
  image_2_187 = _RAND_1339[3:0];
  _RAND_1340 = {1{`RANDOM}};
  image_2_188 = _RAND_1340[3:0];
  _RAND_1341 = {1{`RANDOM}};
  image_2_189 = _RAND_1341[3:0];
  _RAND_1342 = {1{`RANDOM}};
  image_2_190 = _RAND_1342[3:0];
  _RAND_1343 = {1{`RANDOM}};
  image_2_191 = _RAND_1343[3:0];
  _RAND_1344 = {1{`RANDOM}};
  image_2_192 = _RAND_1344[3:0];
  _RAND_1345 = {1{`RANDOM}};
  image_2_193 = _RAND_1345[3:0];
  _RAND_1346 = {1{`RANDOM}};
  image_2_194 = _RAND_1346[3:0];
  _RAND_1347 = {1{`RANDOM}};
  image_2_195 = _RAND_1347[3:0];
  _RAND_1348 = {1{`RANDOM}};
  image_2_196 = _RAND_1348[3:0];
  _RAND_1349 = {1{`RANDOM}};
  image_2_197 = _RAND_1349[3:0];
  _RAND_1350 = {1{`RANDOM}};
  image_2_198 = _RAND_1350[3:0];
  _RAND_1351 = {1{`RANDOM}};
  image_2_199 = _RAND_1351[3:0];
  _RAND_1352 = {1{`RANDOM}};
  image_2_200 = _RAND_1352[3:0];
  _RAND_1353 = {1{`RANDOM}};
  image_2_201 = _RAND_1353[3:0];
  _RAND_1354 = {1{`RANDOM}};
  image_2_202 = _RAND_1354[3:0];
  _RAND_1355 = {1{`RANDOM}};
  image_2_203 = _RAND_1355[3:0];
  _RAND_1356 = {1{`RANDOM}};
  image_2_204 = _RAND_1356[3:0];
  _RAND_1357 = {1{`RANDOM}};
  image_2_205 = _RAND_1357[3:0];
  _RAND_1358 = {1{`RANDOM}};
  image_2_206 = _RAND_1358[3:0];
  _RAND_1359 = {1{`RANDOM}};
  image_2_207 = _RAND_1359[3:0];
  _RAND_1360 = {1{`RANDOM}};
  image_2_208 = _RAND_1360[3:0];
  _RAND_1361 = {1{`RANDOM}};
  image_2_209 = _RAND_1361[3:0];
  _RAND_1362 = {1{`RANDOM}};
  image_2_210 = _RAND_1362[3:0];
  _RAND_1363 = {1{`RANDOM}};
  image_2_211 = _RAND_1363[3:0];
  _RAND_1364 = {1{`RANDOM}};
  image_2_212 = _RAND_1364[3:0];
  _RAND_1365 = {1{`RANDOM}};
  image_2_213 = _RAND_1365[3:0];
  _RAND_1366 = {1{`RANDOM}};
  image_2_214 = _RAND_1366[3:0];
  _RAND_1367 = {1{`RANDOM}};
  image_2_215 = _RAND_1367[3:0];
  _RAND_1368 = {1{`RANDOM}};
  image_2_216 = _RAND_1368[3:0];
  _RAND_1369 = {1{`RANDOM}};
  image_2_217 = _RAND_1369[3:0];
  _RAND_1370 = {1{`RANDOM}};
  image_2_218 = _RAND_1370[3:0];
  _RAND_1371 = {1{`RANDOM}};
  image_2_219 = _RAND_1371[3:0];
  _RAND_1372 = {1{`RANDOM}};
  image_2_220 = _RAND_1372[3:0];
  _RAND_1373 = {1{`RANDOM}};
  image_2_221 = _RAND_1373[3:0];
  _RAND_1374 = {1{`RANDOM}};
  image_2_222 = _RAND_1374[3:0];
  _RAND_1375 = {1{`RANDOM}};
  image_2_223 = _RAND_1375[3:0];
  _RAND_1376 = {1{`RANDOM}};
  image_2_224 = _RAND_1376[3:0];
  _RAND_1377 = {1{`RANDOM}};
  image_2_225 = _RAND_1377[3:0];
  _RAND_1378 = {1{`RANDOM}};
  image_2_226 = _RAND_1378[3:0];
  _RAND_1379 = {1{`RANDOM}};
  image_2_227 = _RAND_1379[3:0];
  _RAND_1380 = {1{`RANDOM}};
  image_2_228 = _RAND_1380[3:0];
  _RAND_1381 = {1{`RANDOM}};
  image_2_229 = _RAND_1381[3:0];
  _RAND_1382 = {1{`RANDOM}};
  image_2_230 = _RAND_1382[3:0];
  _RAND_1383 = {1{`RANDOM}};
  image_2_231 = _RAND_1383[3:0];
  _RAND_1384 = {1{`RANDOM}};
  image_2_232 = _RAND_1384[3:0];
  _RAND_1385 = {1{`RANDOM}};
  image_2_233 = _RAND_1385[3:0];
  _RAND_1386 = {1{`RANDOM}};
  image_2_234 = _RAND_1386[3:0];
  _RAND_1387 = {1{`RANDOM}};
  image_2_235 = _RAND_1387[3:0];
  _RAND_1388 = {1{`RANDOM}};
  image_2_236 = _RAND_1388[3:0];
  _RAND_1389 = {1{`RANDOM}};
  image_2_237 = _RAND_1389[3:0];
  _RAND_1390 = {1{`RANDOM}};
  image_2_238 = _RAND_1390[3:0];
  _RAND_1391 = {1{`RANDOM}};
  image_2_239 = _RAND_1391[3:0];
  _RAND_1392 = {1{`RANDOM}};
  image_2_240 = _RAND_1392[3:0];
  _RAND_1393 = {1{`RANDOM}};
  image_2_241 = _RAND_1393[3:0];
  _RAND_1394 = {1{`RANDOM}};
  image_2_242 = _RAND_1394[3:0];
  _RAND_1395 = {1{`RANDOM}};
  image_2_243 = _RAND_1395[3:0];
  _RAND_1396 = {1{`RANDOM}};
  image_2_244 = _RAND_1396[3:0];
  _RAND_1397 = {1{`RANDOM}};
  image_2_245 = _RAND_1397[3:0];
  _RAND_1398 = {1{`RANDOM}};
  image_2_246 = _RAND_1398[3:0];
  _RAND_1399 = {1{`RANDOM}};
  image_2_247 = _RAND_1399[3:0];
  _RAND_1400 = {1{`RANDOM}};
  image_2_248 = _RAND_1400[3:0];
  _RAND_1401 = {1{`RANDOM}};
  image_2_249 = _RAND_1401[3:0];
  _RAND_1402 = {1{`RANDOM}};
  image_2_250 = _RAND_1402[3:0];
  _RAND_1403 = {1{`RANDOM}};
  image_2_251 = _RAND_1403[3:0];
  _RAND_1404 = {1{`RANDOM}};
  image_2_252 = _RAND_1404[3:0];
  _RAND_1405 = {1{`RANDOM}};
  image_2_253 = _RAND_1405[3:0];
  _RAND_1406 = {1{`RANDOM}};
  image_2_254 = _RAND_1406[3:0];
  _RAND_1407 = {1{`RANDOM}};
  image_2_255 = _RAND_1407[3:0];
  _RAND_1408 = {1{`RANDOM}};
  image_2_256 = _RAND_1408[3:0];
  _RAND_1409 = {1{`RANDOM}};
  image_2_257 = _RAND_1409[3:0];
  _RAND_1410 = {1{`RANDOM}};
  image_2_258 = _RAND_1410[3:0];
  _RAND_1411 = {1{`RANDOM}};
  image_2_259 = _RAND_1411[3:0];
  _RAND_1412 = {1{`RANDOM}};
  image_2_260 = _RAND_1412[3:0];
  _RAND_1413 = {1{`RANDOM}};
  image_2_261 = _RAND_1413[3:0];
  _RAND_1414 = {1{`RANDOM}};
  image_2_262 = _RAND_1414[3:0];
  _RAND_1415 = {1{`RANDOM}};
  image_2_263 = _RAND_1415[3:0];
  _RAND_1416 = {1{`RANDOM}};
  image_2_264 = _RAND_1416[3:0];
  _RAND_1417 = {1{`RANDOM}};
  image_2_265 = _RAND_1417[3:0];
  _RAND_1418 = {1{`RANDOM}};
  image_2_266 = _RAND_1418[3:0];
  _RAND_1419 = {1{`RANDOM}};
  image_2_267 = _RAND_1419[3:0];
  _RAND_1420 = {1{`RANDOM}};
  image_2_268 = _RAND_1420[3:0];
  _RAND_1421 = {1{`RANDOM}};
  image_2_269 = _RAND_1421[3:0];
  _RAND_1422 = {1{`RANDOM}};
  image_2_270 = _RAND_1422[3:0];
  _RAND_1423 = {1{`RANDOM}};
  image_2_271 = _RAND_1423[3:0];
  _RAND_1424 = {1{`RANDOM}};
  image_2_272 = _RAND_1424[3:0];
  _RAND_1425 = {1{`RANDOM}};
  image_2_273 = _RAND_1425[3:0];
  _RAND_1426 = {1{`RANDOM}};
  image_2_274 = _RAND_1426[3:0];
  _RAND_1427 = {1{`RANDOM}};
  image_2_275 = _RAND_1427[3:0];
  _RAND_1428 = {1{`RANDOM}};
  image_2_276 = _RAND_1428[3:0];
  _RAND_1429 = {1{`RANDOM}};
  image_2_277 = _RAND_1429[3:0];
  _RAND_1430 = {1{`RANDOM}};
  image_2_278 = _RAND_1430[3:0];
  _RAND_1431 = {1{`RANDOM}};
  image_2_279 = _RAND_1431[3:0];
  _RAND_1432 = {1{`RANDOM}};
  image_2_280 = _RAND_1432[3:0];
  _RAND_1433 = {1{`RANDOM}};
  image_2_281 = _RAND_1433[3:0];
  _RAND_1434 = {1{`RANDOM}};
  image_2_282 = _RAND_1434[3:0];
  _RAND_1435 = {1{`RANDOM}};
  image_2_283 = _RAND_1435[3:0];
  _RAND_1436 = {1{`RANDOM}};
  image_2_284 = _RAND_1436[3:0];
  _RAND_1437 = {1{`RANDOM}};
  image_2_285 = _RAND_1437[3:0];
  _RAND_1438 = {1{`RANDOM}};
  image_2_286 = _RAND_1438[3:0];
  _RAND_1439 = {1{`RANDOM}};
  image_2_287 = _RAND_1439[3:0];
  _RAND_1440 = {1{`RANDOM}};
  image_2_288 = _RAND_1440[3:0];
  _RAND_1441 = {1{`RANDOM}};
  image_2_289 = _RAND_1441[3:0];
  _RAND_1442 = {1{`RANDOM}};
  image_2_290 = _RAND_1442[3:0];
  _RAND_1443 = {1{`RANDOM}};
  image_2_291 = _RAND_1443[3:0];
  _RAND_1444 = {1{`RANDOM}};
  image_2_292 = _RAND_1444[3:0];
  _RAND_1445 = {1{`RANDOM}};
  image_2_293 = _RAND_1445[3:0];
  _RAND_1446 = {1{`RANDOM}};
  image_2_294 = _RAND_1446[3:0];
  _RAND_1447 = {1{`RANDOM}};
  image_2_295 = _RAND_1447[3:0];
  _RAND_1448 = {1{`RANDOM}};
  image_2_296 = _RAND_1448[3:0];
  _RAND_1449 = {1{`RANDOM}};
  image_2_297 = _RAND_1449[3:0];
  _RAND_1450 = {1{`RANDOM}};
  image_2_298 = _RAND_1450[3:0];
  _RAND_1451 = {1{`RANDOM}};
  image_2_299 = _RAND_1451[3:0];
  _RAND_1452 = {1{`RANDOM}};
  image_2_300 = _RAND_1452[3:0];
  _RAND_1453 = {1{`RANDOM}};
  image_2_301 = _RAND_1453[3:0];
  _RAND_1454 = {1{`RANDOM}};
  image_2_302 = _RAND_1454[3:0];
  _RAND_1455 = {1{`RANDOM}};
  image_2_303 = _RAND_1455[3:0];
  _RAND_1456 = {1{`RANDOM}};
  image_2_304 = _RAND_1456[3:0];
  _RAND_1457 = {1{`RANDOM}};
  image_2_305 = _RAND_1457[3:0];
  _RAND_1458 = {1{`RANDOM}};
  image_2_306 = _RAND_1458[3:0];
  _RAND_1459 = {1{`RANDOM}};
  image_2_307 = _RAND_1459[3:0];
  _RAND_1460 = {1{`RANDOM}};
  image_2_308 = _RAND_1460[3:0];
  _RAND_1461 = {1{`RANDOM}};
  image_2_309 = _RAND_1461[3:0];
  _RAND_1462 = {1{`RANDOM}};
  image_2_310 = _RAND_1462[3:0];
  _RAND_1463 = {1{`RANDOM}};
  image_2_311 = _RAND_1463[3:0];
  _RAND_1464 = {1{`RANDOM}};
  image_2_312 = _RAND_1464[3:0];
  _RAND_1465 = {1{`RANDOM}};
  image_2_313 = _RAND_1465[3:0];
  _RAND_1466 = {1{`RANDOM}};
  image_2_314 = _RAND_1466[3:0];
  _RAND_1467 = {1{`RANDOM}};
  image_2_315 = _RAND_1467[3:0];
  _RAND_1468 = {1{`RANDOM}};
  image_2_316 = _RAND_1468[3:0];
  _RAND_1469 = {1{`RANDOM}};
  image_2_317 = _RAND_1469[3:0];
  _RAND_1470 = {1{`RANDOM}};
  image_2_318 = _RAND_1470[3:0];
  _RAND_1471 = {1{`RANDOM}};
  image_2_319 = _RAND_1471[3:0];
  _RAND_1472 = {1{`RANDOM}};
  image_2_320 = _RAND_1472[3:0];
  _RAND_1473 = {1{`RANDOM}};
  image_2_321 = _RAND_1473[3:0];
  _RAND_1474 = {1{`RANDOM}};
  image_2_322 = _RAND_1474[3:0];
  _RAND_1475 = {1{`RANDOM}};
  image_2_323 = _RAND_1475[3:0];
  _RAND_1476 = {1{`RANDOM}};
  image_2_324 = _RAND_1476[3:0];
  _RAND_1477 = {1{`RANDOM}};
  image_2_325 = _RAND_1477[3:0];
  _RAND_1478 = {1{`RANDOM}};
  image_2_326 = _RAND_1478[3:0];
  _RAND_1479 = {1{`RANDOM}};
  image_2_327 = _RAND_1479[3:0];
  _RAND_1480 = {1{`RANDOM}};
  image_2_328 = _RAND_1480[3:0];
  _RAND_1481 = {1{`RANDOM}};
  image_2_329 = _RAND_1481[3:0];
  _RAND_1482 = {1{`RANDOM}};
  image_2_330 = _RAND_1482[3:0];
  _RAND_1483 = {1{`RANDOM}};
  image_2_331 = _RAND_1483[3:0];
  _RAND_1484 = {1{`RANDOM}};
  image_2_332 = _RAND_1484[3:0];
  _RAND_1485 = {1{`RANDOM}};
  image_2_333 = _RAND_1485[3:0];
  _RAND_1486 = {1{`RANDOM}};
  image_2_334 = _RAND_1486[3:0];
  _RAND_1487 = {1{`RANDOM}};
  image_2_335 = _RAND_1487[3:0];
  _RAND_1488 = {1{`RANDOM}};
  image_2_336 = _RAND_1488[3:0];
  _RAND_1489 = {1{`RANDOM}};
  image_2_337 = _RAND_1489[3:0];
  _RAND_1490 = {1{`RANDOM}};
  image_2_338 = _RAND_1490[3:0];
  _RAND_1491 = {1{`RANDOM}};
  image_2_339 = _RAND_1491[3:0];
  _RAND_1492 = {1{`RANDOM}};
  image_2_340 = _RAND_1492[3:0];
  _RAND_1493 = {1{`RANDOM}};
  image_2_341 = _RAND_1493[3:0];
  _RAND_1494 = {1{`RANDOM}};
  image_2_342 = _RAND_1494[3:0];
  _RAND_1495 = {1{`RANDOM}};
  image_2_343 = _RAND_1495[3:0];
  _RAND_1496 = {1{`RANDOM}};
  image_2_344 = _RAND_1496[3:0];
  _RAND_1497 = {1{`RANDOM}};
  image_2_345 = _RAND_1497[3:0];
  _RAND_1498 = {1{`RANDOM}};
  image_2_346 = _RAND_1498[3:0];
  _RAND_1499 = {1{`RANDOM}};
  image_2_347 = _RAND_1499[3:0];
  _RAND_1500 = {1{`RANDOM}};
  image_2_348 = _RAND_1500[3:0];
  _RAND_1501 = {1{`RANDOM}};
  image_2_349 = _RAND_1501[3:0];
  _RAND_1502 = {1{`RANDOM}};
  image_2_350 = _RAND_1502[3:0];
  _RAND_1503 = {1{`RANDOM}};
  image_2_351 = _RAND_1503[3:0];
  _RAND_1504 = {1{`RANDOM}};
  image_2_352 = _RAND_1504[3:0];
  _RAND_1505 = {1{`RANDOM}};
  image_2_353 = _RAND_1505[3:0];
  _RAND_1506 = {1{`RANDOM}};
  image_2_354 = _RAND_1506[3:0];
  _RAND_1507 = {1{`RANDOM}};
  image_2_355 = _RAND_1507[3:0];
  _RAND_1508 = {1{`RANDOM}};
  image_2_356 = _RAND_1508[3:0];
  _RAND_1509 = {1{`RANDOM}};
  image_2_357 = _RAND_1509[3:0];
  _RAND_1510 = {1{`RANDOM}};
  image_2_358 = _RAND_1510[3:0];
  _RAND_1511 = {1{`RANDOM}};
  image_2_359 = _RAND_1511[3:0];
  _RAND_1512 = {1{`RANDOM}};
  image_2_360 = _RAND_1512[3:0];
  _RAND_1513 = {1{`RANDOM}};
  image_2_361 = _RAND_1513[3:0];
  _RAND_1514 = {1{`RANDOM}};
  image_2_362 = _RAND_1514[3:0];
  _RAND_1515 = {1{`RANDOM}};
  image_2_363 = _RAND_1515[3:0];
  _RAND_1516 = {1{`RANDOM}};
  image_2_364 = _RAND_1516[3:0];
  _RAND_1517 = {1{`RANDOM}};
  image_2_365 = _RAND_1517[3:0];
  _RAND_1518 = {1{`RANDOM}};
  image_2_366 = _RAND_1518[3:0];
  _RAND_1519 = {1{`RANDOM}};
  image_2_367 = _RAND_1519[3:0];
  _RAND_1520 = {1{`RANDOM}};
  image_2_368 = _RAND_1520[3:0];
  _RAND_1521 = {1{`RANDOM}};
  image_2_369 = _RAND_1521[3:0];
  _RAND_1522 = {1{`RANDOM}};
  image_2_370 = _RAND_1522[3:0];
  _RAND_1523 = {1{`RANDOM}};
  image_2_371 = _RAND_1523[3:0];
  _RAND_1524 = {1{`RANDOM}};
  image_2_372 = _RAND_1524[3:0];
  _RAND_1525 = {1{`RANDOM}};
  image_2_373 = _RAND_1525[3:0];
  _RAND_1526 = {1{`RANDOM}};
  image_2_374 = _RAND_1526[3:0];
  _RAND_1527 = {1{`RANDOM}};
  image_2_375 = _RAND_1527[3:0];
  _RAND_1528 = {1{`RANDOM}};
  image_2_376 = _RAND_1528[3:0];
  _RAND_1529 = {1{`RANDOM}};
  image_2_377 = _RAND_1529[3:0];
  _RAND_1530 = {1{`RANDOM}};
  image_2_378 = _RAND_1530[3:0];
  _RAND_1531 = {1{`RANDOM}};
  image_2_379 = _RAND_1531[3:0];
  _RAND_1532 = {1{`RANDOM}};
  image_2_380 = _RAND_1532[3:0];
  _RAND_1533 = {1{`RANDOM}};
  image_2_381 = _RAND_1533[3:0];
  _RAND_1534 = {1{`RANDOM}};
  image_2_382 = _RAND_1534[3:0];
  _RAND_1535 = {1{`RANDOM}};
  image_2_383 = _RAND_1535[3:0];
  _RAND_1536 = {1{`RANDOM}};
  image_2_384 = _RAND_1536[3:0];
  _RAND_1537 = {1{`RANDOM}};
  image_2_385 = _RAND_1537[3:0];
  _RAND_1538 = {1{`RANDOM}};
  image_2_386 = _RAND_1538[3:0];
  _RAND_1539 = {1{`RANDOM}};
  image_2_387 = _RAND_1539[3:0];
  _RAND_1540 = {1{`RANDOM}};
  image_2_388 = _RAND_1540[3:0];
  _RAND_1541 = {1{`RANDOM}};
  image_2_389 = _RAND_1541[3:0];
  _RAND_1542 = {1{`RANDOM}};
  image_2_390 = _RAND_1542[3:0];
  _RAND_1543 = {1{`RANDOM}};
  image_2_391 = _RAND_1543[3:0];
  _RAND_1544 = {1{`RANDOM}};
  image_2_392 = _RAND_1544[3:0];
  _RAND_1545 = {1{`RANDOM}};
  image_2_393 = _RAND_1545[3:0];
  _RAND_1546 = {1{`RANDOM}};
  image_2_394 = _RAND_1546[3:0];
  _RAND_1547 = {1{`RANDOM}};
  image_2_395 = _RAND_1547[3:0];
  _RAND_1548 = {1{`RANDOM}};
  image_2_396 = _RAND_1548[3:0];
  _RAND_1549 = {1{`RANDOM}};
  image_2_397 = _RAND_1549[3:0];
  _RAND_1550 = {1{`RANDOM}};
  image_2_398 = _RAND_1550[3:0];
  _RAND_1551 = {1{`RANDOM}};
  image_2_399 = _RAND_1551[3:0];
  _RAND_1552 = {1{`RANDOM}};
  image_2_400 = _RAND_1552[3:0];
  _RAND_1553 = {1{`RANDOM}};
  image_2_401 = _RAND_1553[3:0];
  _RAND_1554 = {1{`RANDOM}};
  image_2_402 = _RAND_1554[3:0];
  _RAND_1555 = {1{`RANDOM}};
  image_2_403 = _RAND_1555[3:0];
  _RAND_1556 = {1{`RANDOM}};
  image_2_404 = _RAND_1556[3:0];
  _RAND_1557 = {1{`RANDOM}};
  image_2_405 = _RAND_1557[3:0];
  _RAND_1558 = {1{`RANDOM}};
  image_2_406 = _RAND_1558[3:0];
  _RAND_1559 = {1{`RANDOM}};
  image_2_407 = _RAND_1559[3:0];
  _RAND_1560 = {1{`RANDOM}};
  image_2_408 = _RAND_1560[3:0];
  _RAND_1561 = {1{`RANDOM}};
  image_2_409 = _RAND_1561[3:0];
  _RAND_1562 = {1{`RANDOM}};
  image_2_410 = _RAND_1562[3:0];
  _RAND_1563 = {1{`RANDOM}};
  image_2_411 = _RAND_1563[3:0];
  _RAND_1564 = {1{`RANDOM}};
  image_2_412 = _RAND_1564[3:0];
  _RAND_1565 = {1{`RANDOM}};
  image_2_413 = _RAND_1565[3:0];
  _RAND_1566 = {1{`RANDOM}};
  image_2_414 = _RAND_1566[3:0];
  _RAND_1567 = {1{`RANDOM}};
  image_2_415 = _RAND_1567[3:0];
  _RAND_1568 = {1{`RANDOM}};
  image_2_416 = _RAND_1568[3:0];
  _RAND_1569 = {1{`RANDOM}};
  image_2_417 = _RAND_1569[3:0];
  _RAND_1570 = {1{`RANDOM}};
  image_2_418 = _RAND_1570[3:0];
  _RAND_1571 = {1{`RANDOM}};
  image_2_419 = _RAND_1571[3:0];
  _RAND_1572 = {1{`RANDOM}};
  image_2_420 = _RAND_1572[3:0];
  _RAND_1573 = {1{`RANDOM}};
  image_2_421 = _RAND_1573[3:0];
  _RAND_1574 = {1{`RANDOM}};
  image_2_422 = _RAND_1574[3:0];
  _RAND_1575 = {1{`RANDOM}};
  image_2_423 = _RAND_1575[3:0];
  _RAND_1576 = {1{`RANDOM}};
  image_2_424 = _RAND_1576[3:0];
  _RAND_1577 = {1{`RANDOM}};
  image_2_425 = _RAND_1577[3:0];
  _RAND_1578 = {1{`RANDOM}};
  image_2_426 = _RAND_1578[3:0];
  _RAND_1579 = {1{`RANDOM}};
  image_2_427 = _RAND_1579[3:0];
  _RAND_1580 = {1{`RANDOM}};
  image_2_428 = _RAND_1580[3:0];
  _RAND_1581 = {1{`RANDOM}};
  image_2_429 = _RAND_1581[3:0];
  _RAND_1582 = {1{`RANDOM}};
  image_2_430 = _RAND_1582[3:0];
  _RAND_1583 = {1{`RANDOM}};
  image_2_431 = _RAND_1583[3:0];
  _RAND_1584 = {1{`RANDOM}};
  image_2_432 = _RAND_1584[3:0];
  _RAND_1585 = {1{`RANDOM}};
  image_2_433 = _RAND_1585[3:0];
  _RAND_1586 = {1{`RANDOM}};
  image_2_434 = _RAND_1586[3:0];
  _RAND_1587 = {1{`RANDOM}};
  image_2_435 = _RAND_1587[3:0];
  _RAND_1588 = {1{`RANDOM}};
  image_2_436 = _RAND_1588[3:0];
  _RAND_1589 = {1{`RANDOM}};
  image_2_437 = _RAND_1589[3:0];
  _RAND_1590 = {1{`RANDOM}};
  image_2_438 = _RAND_1590[3:0];
  _RAND_1591 = {1{`RANDOM}};
  image_2_439 = _RAND_1591[3:0];
  _RAND_1592 = {1{`RANDOM}};
  image_2_440 = _RAND_1592[3:0];
  _RAND_1593 = {1{`RANDOM}};
  image_2_441 = _RAND_1593[3:0];
  _RAND_1594 = {1{`RANDOM}};
  image_2_442 = _RAND_1594[3:0];
  _RAND_1595 = {1{`RANDOM}};
  image_2_443 = _RAND_1595[3:0];
  _RAND_1596 = {1{`RANDOM}};
  image_2_444 = _RAND_1596[3:0];
  _RAND_1597 = {1{`RANDOM}};
  image_2_445 = _RAND_1597[3:0];
  _RAND_1598 = {1{`RANDOM}};
  image_2_446 = _RAND_1598[3:0];
  _RAND_1599 = {1{`RANDOM}};
  image_2_447 = _RAND_1599[3:0];
  _RAND_1600 = {1{`RANDOM}};
  image_2_448 = _RAND_1600[3:0];
  _RAND_1601 = {1{`RANDOM}};
  image_2_449 = _RAND_1601[3:0];
  _RAND_1602 = {1{`RANDOM}};
  image_2_450 = _RAND_1602[3:0];
  _RAND_1603 = {1{`RANDOM}};
  image_2_451 = _RAND_1603[3:0];
  _RAND_1604 = {1{`RANDOM}};
  image_2_452 = _RAND_1604[3:0];
  _RAND_1605 = {1{`RANDOM}};
  image_2_453 = _RAND_1605[3:0];
  _RAND_1606 = {1{`RANDOM}};
  image_2_454 = _RAND_1606[3:0];
  _RAND_1607 = {1{`RANDOM}};
  image_2_455 = _RAND_1607[3:0];
  _RAND_1608 = {1{`RANDOM}};
  image_2_456 = _RAND_1608[3:0];
  _RAND_1609 = {1{`RANDOM}};
  image_2_457 = _RAND_1609[3:0];
  _RAND_1610 = {1{`RANDOM}};
  image_2_458 = _RAND_1610[3:0];
  _RAND_1611 = {1{`RANDOM}};
  image_2_459 = _RAND_1611[3:0];
  _RAND_1612 = {1{`RANDOM}};
  image_2_460 = _RAND_1612[3:0];
  _RAND_1613 = {1{`RANDOM}};
  image_2_461 = _RAND_1613[3:0];
  _RAND_1614 = {1{`RANDOM}};
  image_2_462 = _RAND_1614[3:0];
  _RAND_1615 = {1{`RANDOM}};
  image_2_463 = _RAND_1615[3:0];
  _RAND_1616 = {1{`RANDOM}};
  image_2_464 = _RAND_1616[3:0];
  _RAND_1617 = {1{`RANDOM}};
  image_2_465 = _RAND_1617[3:0];
  _RAND_1618 = {1{`RANDOM}};
  image_2_466 = _RAND_1618[3:0];
  _RAND_1619 = {1{`RANDOM}};
  image_2_467 = _RAND_1619[3:0];
  _RAND_1620 = {1{`RANDOM}};
  image_2_468 = _RAND_1620[3:0];
  _RAND_1621 = {1{`RANDOM}};
  image_2_469 = _RAND_1621[3:0];
  _RAND_1622 = {1{`RANDOM}};
  image_2_470 = _RAND_1622[3:0];
  _RAND_1623 = {1{`RANDOM}};
  image_2_471 = _RAND_1623[3:0];
  _RAND_1624 = {1{`RANDOM}};
  image_2_472 = _RAND_1624[3:0];
  _RAND_1625 = {1{`RANDOM}};
  image_2_473 = _RAND_1625[3:0];
  _RAND_1626 = {1{`RANDOM}};
  image_2_474 = _RAND_1626[3:0];
  _RAND_1627 = {1{`RANDOM}};
  image_2_475 = _RAND_1627[3:0];
  _RAND_1628 = {1{`RANDOM}};
  image_2_476 = _RAND_1628[3:0];
  _RAND_1629 = {1{`RANDOM}};
  image_2_477 = _RAND_1629[3:0];
  _RAND_1630 = {1{`RANDOM}};
  image_2_478 = _RAND_1630[3:0];
  _RAND_1631 = {1{`RANDOM}};
  image_2_479 = _RAND_1631[3:0];
  _RAND_1632 = {1{`RANDOM}};
  image_2_480 = _RAND_1632[3:0];
  _RAND_1633 = {1{`RANDOM}};
  image_2_481 = _RAND_1633[3:0];
  _RAND_1634 = {1{`RANDOM}};
  image_2_482 = _RAND_1634[3:0];
  _RAND_1635 = {1{`RANDOM}};
  image_2_483 = _RAND_1635[3:0];
  _RAND_1636 = {1{`RANDOM}};
  image_2_484 = _RAND_1636[3:0];
  _RAND_1637 = {1{`RANDOM}};
  image_2_485 = _RAND_1637[3:0];
  _RAND_1638 = {1{`RANDOM}};
  image_2_486 = _RAND_1638[3:0];
  _RAND_1639 = {1{`RANDOM}};
  image_2_487 = _RAND_1639[3:0];
  _RAND_1640 = {1{`RANDOM}};
  image_2_488 = _RAND_1640[3:0];
  _RAND_1641 = {1{`RANDOM}};
  image_2_489 = _RAND_1641[3:0];
  _RAND_1642 = {1{`RANDOM}};
  image_2_490 = _RAND_1642[3:0];
  _RAND_1643 = {1{`RANDOM}};
  image_2_491 = _RAND_1643[3:0];
  _RAND_1644 = {1{`RANDOM}};
  image_2_492 = _RAND_1644[3:0];
  _RAND_1645 = {1{`RANDOM}};
  image_2_493 = _RAND_1645[3:0];
  _RAND_1646 = {1{`RANDOM}};
  image_2_494 = _RAND_1646[3:0];
  _RAND_1647 = {1{`RANDOM}};
  image_2_495 = _RAND_1647[3:0];
  _RAND_1648 = {1{`RANDOM}};
  image_2_496 = _RAND_1648[3:0];
  _RAND_1649 = {1{`RANDOM}};
  image_2_497 = _RAND_1649[3:0];
  _RAND_1650 = {1{`RANDOM}};
  image_2_498 = _RAND_1650[3:0];
  _RAND_1651 = {1{`RANDOM}};
  image_2_499 = _RAND_1651[3:0];
  _RAND_1652 = {1{`RANDOM}};
  image_2_500 = _RAND_1652[3:0];
  _RAND_1653 = {1{`RANDOM}};
  image_2_501 = _RAND_1653[3:0];
  _RAND_1654 = {1{`RANDOM}};
  image_2_502 = _RAND_1654[3:0];
  _RAND_1655 = {1{`RANDOM}};
  image_2_503 = _RAND_1655[3:0];
  _RAND_1656 = {1{`RANDOM}};
  image_2_504 = _RAND_1656[3:0];
  _RAND_1657 = {1{`RANDOM}};
  image_2_505 = _RAND_1657[3:0];
  _RAND_1658 = {1{`RANDOM}};
  image_2_506 = _RAND_1658[3:0];
  _RAND_1659 = {1{`RANDOM}};
  image_2_507 = _RAND_1659[3:0];
  _RAND_1660 = {1{`RANDOM}};
  image_2_508 = _RAND_1660[3:0];
  _RAND_1661 = {1{`RANDOM}};
  image_2_509 = _RAND_1661[3:0];
  _RAND_1662 = {1{`RANDOM}};
  image_2_510 = _RAND_1662[3:0];
  _RAND_1663 = {1{`RANDOM}};
  image_2_511 = _RAND_1663[3:0];
  _RAND_1664 = {1{`RANDOM}};
  image_2_512 = _RAND_1664[3:0];
  _RAND_1665 = {1{`RANDOM}};
  image_2_513 = _RAND_1665[3:0];
  _RAND_1666 = {1{`RANDOM}};
  image_2_514 = _RAND_1666[3:0];
  _RAND_1667 = {1{`RANDOM}};
  image_2_515 = _RAND_1667[3:0];
  _RAND_1668 = {1{`RANDOM}};
  image_2_516 = _RAND_1668[3:0];
  _RAND_1669 = {1{`RANDOM}};
  image_2_517 = _RAND_1669[3:0];
  _RAND_1670 = {1{`RANDOM}};
  image_2_518 = _RAND_1670[3:0];
  _RAND_1671 = {1{`RANDOM}};
  image_2_519 = _RAND_1671[3:0];
  _RAND_1672 = {1{`RANDOM}};
  image_2_520 = _RAND_1672[3:0];
  _RAND_1673 = {1{`RANDOM}};
  image_2_521 = _RAND_1673[3:0];
  _RAND_1674 = {1{`RANDOM}};
  image_2_522 = _RAND_1674[3:0];
  _RAND_1675 = {1{`RANDOM}};
  image_2_523 = _RAND_1675[3:0];
  _RAND_1676 = {1{`RANDOM}};
  image_2_524 = _RAND_1676[3:0];
  _RAND_1677 = {1{`RANDOM}};
  image_2_525 = _RAND_1677[3:0];
  _RAND_1678 = {1{`RANDOM}};
  image_2_526 = _RAND_1678[3:0];
  _RAND_1679 = {1{`RANDOM}};
  image_2_527 = _RAND_1679[3:0];
  _RAND_1680 = {1{`RANDOM}};
  image_2_528 = _RAND_1680[3:0];
  _RAND_1681 = {1{`RANDOM}};
  image_2_529 = _RAND_1681[3:0];
  _RAND_1682 = {1{`RANDOM}};
  image_2_530 = _RAND_1682[3:0];
  _RAND_1683 = {1{`RANDOM}};
  image_2_531 = _RAND_1683[3:0];
  _RAND_1684 = {1{`RANDOM}};
  image_2_532 = _RAND_1684[3:0];
  _RAND_1685 = {1{`RANDOM}};
  image_2_533 = _RAND_1685[3:0];
  _RAND_1686 = {1{`RANDOM}};
  image_2_534 = _RAND_1686[3:0];
  _RAND_1687 = {1{`RANDOM}};
  image_2_535 = _RAND_1687[3:0];
  _RAND_1688 = {1{`RANDOM}};
  image_2_536 = _RAND_1688[3:0];
  _RAND_1689 = {1{`RANDOM}};
  image_2_537 = _RAND_1689[3:0];
  _RAND_1690 = {1{`RANDOM}};
  image_2_538 = _RAND_1690[3:0];
  _RAND_1691 = {1{`RANDOM}};
  image_2_539 = _RAND_1691[3:0];
  _RAND_1692 = {1{`RANDOM}};
  image_2_540 = _RAND_1692[3:0];
  _RAND_1693 = {1{`RANDOM}};
  image_2_541 = _RAND_1693[3:0];
  _RAND_1694 = {1{`RANDOM}};
  image_2_542 = _RAND_1694[3:0];
  _RAND_1695 = {1{`RANDOM}};
  image_2_543 = _RAND_1695[3:0];
  _RAND_1696 = {1{`RANDOM}};
  image_2_544 = _RAND_1696[3:0];
  _RAND_1697 = {1{`RANDOM}};
  image_2_545 = _RAND_1697[3:0];
  _RAND_1698 = {1{`RANDOM}};
  image_2_546 = _RAND_1698[3:0];
  _RAND_1699 = {1{`RANDOM}};
  image_2_547 = _RAND_1699[3:0];
  _RAND_1700 = {1{`RANDOM}};
  image_2_548 = _RAND_1700[3:0];
  _RAND_1701 = {1{`RANDOM}};
  image_2_549 = _RAND_1701[3:0];
  _RAND_1702 = {1{`RANDOM}};
  image_2_550 = _RAND_1702[3:0];
  _RAND_1703 = {1{`RANDOM}};
  image_2_551 = _RAND_1703[3:0];
  _RAND_1704 = {1{`RANDOM}};
  image_2_552 = _RAND_1704[3:0];
  _RAND_1705 = {1{`RANDOM}};
  image_2_553 = _RAND_1705[3:0];
  _RAND_1706 = {1{`RANDOM}};
  image_2_554 = _RAND_1706[3:0];
  _RAND_1707 = {1{`RANDOM}};
  image_2_555 = _RAND_1707[3:0];
  _RAND_1708 = {1{`RANDOM}};
  image_2_556 = _RAND_1708[3:0];
  _RAND_1709 = {1{`RANDOM}};
  image_2_557 = _RAND_1709[3:0];
  _RAND_1710 = {1{`RANDOM}};
  image_2_558 = _RAND_1710[3:0];
  _RAND_1711 = {1{`RANDOM}};
  image_2_559 = _RAND_1711[3:0];
  _RAND_1712 = {1{`RANDOM}};
  image_2_560 = _RAND_1712[3:0];
  _RAND_1713 = {1{`RANDOM}};
  image_2_561 = _RAND_1713[3:0];
  _RAND_1714 = {1{`RANDOM}};
  image_2_562 = _RAND_1714[3:0];
  _RAND_1715 = {1{`RANDOM}};
  image_2_563 = _RAND_1715[3:0];
  _RAND_1716 = {1{`RANDOM}};
  image_2_564 = _RAND_1716[3:0];
  _RAND_1717 = {1{`RANDOM}};
  image_2_565 = _RAND_1717[3:0];
  _RAND_1718 = {1{`RANDOM}};
  image_2_566 = _RAND_1718[3:0];
  _RAND_1719 = {1{`RANDOM}};
  image_2_567 = _RAND_1719[3:0];
  _RAND_1720 = {1{`RANDOM}};
  image_2_568 = _RAND_1720[3:0];
  _RAND_1721 = {1{`RANDOM}};
  image_2_569 = _RAND_1721[3:0];
  _RAND_1722 = {1{`RANDOM}};
  image_2_570 = _RAND_1722[3:0];
  _RAND_1723 = {1{`RANDOM}};
  image_2_571 = _RAND_1723[3:0];
  _RAND_1724 = {1{`RANDOM}};
  image_2_572 = _RAND_1724[3:0];
  _RAND_1725 = {1{`RANDOM}};
  image_2_573 = _RAND_1725[3:0];
  _RAND_1726 = {1{`RANDOM}};
  image_2_574 = _RAND_1726[3:0];
  _RAND_1727 = {1{`RANDOM}};
  image_2_575 = _RAND_1727[3:0];
  _RAND_1728 = {1{`RANDOM}};
  pixelIndex = _RAND_1728[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      image_0_0 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h0 == _T_37[9:0]) begin
        image_0_0 <= io_pixelVal_in_0_7;
      end else if (10'h0 == _T_34[9:0]) begin
        image_0_0 <= io_pixelVal_in_0_6;
      end else if (10'h0 == _T_31[9:0]) begin
        image_0_0 <= io_pixelVal_in_0_5;
      end else if (10'h0 == _T_28[9:0]) begin
        image_0_0 <= io_pixelVal_in_0_4;
      end else if (10'h0 == _T_25[9:0]) begin
        image_0_0 <= io_pixelVal_in_0_3;
      end else if (10'h0 == _T_22[9:0]) begin
        image_0_0 <= io_pixelVal_in_0_2;
      end else if (10'h0 == _T_19[9:0]) begin
        image_0_0 <= io_pixelVal_in_0_1;
      end else if (10'h0 == _T_15[9:0]) begin
        image_0_0 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_1 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1 == _T_37[9:0]) begin
        image_0_1 <= io_pixelVal_in_0_7;
      end else if (10'h1 == _T_34[9:0]) begin
        image_0_1 <= io_pixelVal_in_0_6;
      end else if (10'h1 == _T_31[9:0]) begin
        image_0_1 <= io_pixelVal_in_0_5;
      end else if (10'h1 == _T_28[9:0]) begin
        image_0_1 <= io_pixelVal_in_0_4;
      end else if (10'h1 == _T_25[9:0]) begin
        image_0_1 <= io_pixelVal_in_0_3;
      end else if (10'h1 == _T_22[9:0]) begin
        image_0_1 <= io_pixelVal_in_0_2;
      end else if (10'h1 == _T_19[9:0]) begin
        image_0_1 <= io_pixelVal_in_0_1;
      end else if (10'h1 == _T_15[9:0]) begin
        image_0_1 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_2 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h2 == _T_37[9:0]) begin
        image_0_2 <= io_pixelVal_in_0_7;
      end else if (10'h2 == _T_34[9:0]) begin
        image_0_2 <= io_pixelVal_in_0_6;
      end else if (10'h2 == _T_31[9:0]) begin
        image_0_2 <= io_pixelVal_in_0_5;
      end else if (10'h2 == _T_28[9:0]) begin
        image_0_2 <= io_pixelVal_in_0_4;
      end else if (10'h2 == _T_25[9:0]) begin
        image_0_2 <= io_pixelVal_in_0_3;
      end else if (10'h2 == _T_22[9:0]) begin
        image_0_2 <= io_pixelVal_in_0_2;
      end else if (10'h2 == _T_19[9:0]) begin
        image_0_2 <= io_pixelVal_in_0_1;
      end else if (10'h2 == _T_15[9:0]) begin
        image_0_2 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_3 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h3 == _T_37[9:0]) begin
        image_0_3 <= io_pixelVal_in_0_7;
      end else if (10'h3 == _T_34[9:0]) begin
        image_0_3 <= io_pixelVal_in_0_6;
      end else if (10'h3 == _T_31[9:0]) begin
        image_0_3 <= io_pixelVal_in_0_5;
      end else if (10'h3 == _T_28[9:0]) begin
        image_0_3 <= io_pixelVal_in_0_4;
      end else if (10'h3 == _T_25[9:0]) begin
        image_0_3 <= io_pixelVal_in_0_3;
      end else if (10'h3 == _T_22[9:0]) begin
        image_0_3 <= io_pixelVal_in_0_2;
      end else if (10'h3 == _T_19[9:0]) begin
        image_0_3 <= io_pixelVal_in_0_1;
      end else if (10'h3 == _T_15[9:0]) begin
        image_0_3 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_4 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h4 == _T_37[9:0]) begin
        image_0_4 <= io_pixelVal_in_0_7;
      end else if (10'h4 == _T_34[9:0]) begin
        image_0_4 <= io_pixelVal_in_0_6;
      end else if (10'h4 == _T_31[9:0]) begin
        image_0_4 <= io_pixelVal_in_0_5;
      end else if (10'h4 == _T_28[9:0]) begin
        image_0_4 <= io_pixelVal_in_0_4;
      end else if (10'h4 == _T_25[9:0]) begin
        image_0_4 <= io_pixelVal_in_0_3;
      end else if (10'h4 == _T_22[9:0]) begin
        image_0_4 <= io_pixelVal_in_0_2;
      end else if (10'h4 == _T_19[9:0]) begin
        image_0_4 <= io_pixelVal_in_0_1;
      end else if (10'h4 == _T_15[9:0]) begin
        image_0_4 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_5 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h5 == _T_37[9:0]) begin
        image_0_5 <= io_pixelVal_in_0_7;
      end else if (10'h5 == _T_34[9:0]) begin
        image_0_5 <= io_pixelVal_in_0_6;
      end else if (10'h5 == _T_31[9:0]) begin
        image_0_5 <= io_pixelVal_in_0_5;
      end else if (10'h5 == _T_28[9:0]) begin
        image_0_5 <= io_pixelVal_in_0_4;
      end else if (10'h5 == _T_25[9:0]) begin
        image_0_5 <= io_pixelVal_in_0_3;
      end else if (10'h5 == _T_22[9:0]) begin
        image_0_5 <= io_pixelVal_in_0_2;
      end else if (10'h5 == _T_19[9:0]) begin
        image_0_5 <= io_pixelVal_in_0_1;
      end else if (10'h5 == _T_15[9:0]) begin
        image_0_5 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_6 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h6 == _T_37[9:0]) begin
        image_0_6 <= io_pixelVal_in_0_7;
      end else if (10'h6 == _T_34[9:0]) begin
        image_0_6 <= io_pixelVal_in_0_6;
      end else if (10'h6 == _T_31[9:0]) begin
        image_0_6 <= io_pixelVal_in_0_5;
      end else if (10'h6 == _T_28[9:0]) begin
        image_0_6 <= io_pixelVal_in_0_4;
      end else if (10'h6 == _T_25[9:0]) begin
        image_0_6 <= io_pixelVal_in_0_3;
      end else if (10'h6 == _T_22[9:0]) begin
        image_0_6 <= io_pixelVal_in_0_2;
      end else if (10'h6 == _T_19[9:0]) begin
        image_0_6 <= io_pixelVal_in_0_1;
      end else if (10'h6 == _T_15[9:0]) begin
        image_0_6 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_7 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h7 == _T_37[9:0]) begin
        image_0_7 <= io_pixelVal_in_0_7;
      end else if (10'h7 == _T_34[9:0]) begin
        image_0_7 <= io_pixelVal_in_0_6;
      end else if (10'h7 == _T_31[9:0]) begin
        image_0_7 <= io_pixelVal_in_0_5;
      end else if (10'h7 == _T_28[9:0]) begin
        image_0_7 <= io_pixelVal_in_0_4;
      end else if (10'h7 == _T_25[9:0]) begin
        image_0_7 <= io_pixelVal_in_0_3;
      end else if (10'h7 == _T_22[9:0]) begin
        image_0_7 <= io_pixelVal_in_0_2;
      end else if (10'h7 == _T_19[9:0]) begin
        image_0_7 <= io_pixelVal_in_0_1;
      end else if (10'h7 == _T_15[9:0]) begin
        image_0_7 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_8 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h8 == _T_37[9:0]) begin
        image_0_8 <= io_pixelVal_in_0_7;
      end else if (10'h8 == _T_34[9:0]) begin
        image_0_8 <= io_pixelVal_in_0_6;
      end else if (10'h8 == _T_31[9:0]) begin
        image_0_8 <= io_pixelVal_in_0_5;
      end else if (10'h8 == _T_28[9:0]) begin
        image_0_8 <= io_pixelVal_in_0_4;
      end else if (10'h8 == _T_25[9:0]) begin
        image_0_8 <= io_pixelVal_in_0_3;
      end else if (10'h8 == _T_22[9:0]) begin
        image_0_8 <= io_pixelVal_in_0_2;
      end else if (10'h8 == _T_19[9:0]) begin
        image_0_8 <= io_pixelVal_in_0_1;
      end else if (10'h8 == _T_15[9:0]) begin
        image_0_8 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_9 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h9 == _T_37[9:0]) begin
        image_0_9 <= io_pixelVal_in_0_7;
      end else if (10'h9 == _T_34[9:0]) begin
        image_0_9 <= io_pixelVal_in_0_6;
      end else if (10'h9 == _T_31[9:0]) begin
        image_0_9 <= io_pixelVal_in_0_5;
      end else if (10'h9 == _T_28[9:0]) begin
        image_0_9 <= io_pixelVal_in_0_4;
      end else if (10'h9 == _T_25[9:0]) begin
        image_0_9 <= io_pixelVal_in_0_3;
      end else if (10'h9 == _T_22[9:0]) begin
        image_0_9 <= io_pixelVal_in_0_2;
      end else if (10'h9 == _T_19[9:0]) begin
        image_0_9 <= io_pixelVal_in_0_1;
      end else if (10'h9 == _T_15[9:0]) begin
        image_0_9 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_10 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'ha == _T_37[9:0]) begin
        image_0_10 <= io_pixelVal_in_0_7;
      end else if (10'ha == _T_34[9:0]) begin
        image_0_10 <= io_pixelVal_in_0_6;
      end else if (10'ha == _T_31[9:0]) begin
        image_0_10 <= io_pixelVal_in_0_5;
      end else if (10'ha == _T_28[9:0]) begin
        image_0_10 <= io_pixelVal_in_0_4;
      end else if (10'ha == _T_25[9:0]) begin
        image_0_10 <= io_pixelVal_in_0_3;
      end else if (10'ha == _T_22[9:0]) begin
        image_0_10 <= io_pixelVal_in_0_2;
      end else if (10'ha == _T_19[9:0]) begin
        image_0_10 <= io_pixelVal_in_0_1;
      end else if (10'ha == _T_15[9:0]) begin
        image_0_10 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_11 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hb == _T_37[9:0]) begin
        image_0_11 <= io_pixelVal_in_0_7;
      end else if (10'hb == _T_34[9:0]) begin
        image_0_11 <= io_pixelVal_in_0_6;
      end else if (10'hb == _T_31[9:0]) begin
        image_0_11 <= io_pixelVal_in_0_5;
      end else if (10'hb == _T_28[9:0]) begin
        image_0_11 <= io_pixelVal_in_0_4;
      end else if (10'hb == _T_25[9:0]) begin
        image_0_11 <= io_pixelVal_in_0_3;
      end else if (10'hb == _T_22[9:0]) begin
        image_0_11 <= io_pixelVal_in_0_2;
      end else if (10'hb == _T_19[9:0]) begin
        image_0_11 <= io_pixelVal_in_0_1;
      end else if (10'hb == _T_15[9:0]) begin
        image_0_11 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_12 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hc == _T_37[9:0]) begin
        image_0_12 <= io_pixelVal_in_0_7;
      end else if (10'hc == _T_34[9:0]) begin
        image_0_12 <= io_pixelVal_in_0_6;
      end else if (10'hc == _T_31[9:0]) begin
        image_0_12 <= io_pixelVal_in_0_5;
      end else if (10'hc == _T_28[9:0]) begin
        image_0_12 <= io_pixelVal_in_0_4;
      end else if (10'hc == _T_25[9:0]) begin
        image_0_12 <= io_pixelVal_in_0_3;
      end else if (10'hc == _T_22[9:0]) begin
        image_0_12 <= io_pixelVal_in_0_2;
      end else if (10'hc == _T_19[9:0]) begin
        image_0_12 <= io_pixelVal_in_0_1;
      end else if (10'hc == _T_15[9:0]) begin
        image_0_12 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_13 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hd == _T_37[9:0]) begin
        image_0_13 <= io_pixelVal_in_0_7;
      end else if (10'hd == _T_34[9:0]) begin
        image_0_13 <= io_pixelVal_in_0_6;
      end else if (10'hd == _T_31[9:0]) begin
        image_0_13 <= io_pixelVal_in_0_5;
      end else if (10'hd == _T_28[9:0]) begin
        image_0_13 <= io_pixelVal_in_0_4;
      end else if (10'hd == _T_25[9:0]) begin
        image_0_13 <= io_pixelVal_in_0_3;
      end else if (10'hd == _T_22[9:0]) begin
        image_0_13 <= io_pixelVal_in_0_2;
      end else if (10'hd == _T_19[9:0]) begin
        image_0_13 <= io_pixelVal_in_0_1;
      end else if (10'hd == _T_15[9:0]) begin
        image_0_13 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_14 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'he == _T_37[9:0]) begin
        image_0_14 <= io_pixelVal_in_0_7;
      end else if (10'he == _T_34[9:0]) begin
        image_0_14 <= io_pixelVal_in_0_6;
      end else if (10'he == _T_31[9:0]) begin
        image_0_14 <= io_pixelVal_in_0_5;
      end else if (10'he == _T_28[9:0]) begin
        image_0_14 <= io_pixelVal_in_0_4;
      end else if (10'he == _T_25[9:0]) begin
        image_0_14 <= io_pixelVal_in_0_3;
      end else if (10'he == _T_22[9:0]) begin
        image_0_14 <= io_pixelVal_in_0_2;
      end else if (10'he == _T_19[9:0]) begin
        image_0_14 <= io_pixelVal_in_0_1;
      end else if (10'he == _T_15[9:0]) begin
        image_0_14 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_15 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hf == _T_37[9:0]) begin
        image_0_15 <= io_pixelVal_in_0_7;
      end else if (10'hf == _T_34[9:0]) begin
        image_0_15 <= io_pixelVal_in_0_6;
      end else if (10'hf == _T_31[9:0]) begin
        image_0_15 <= io_pixelVal_in_0_5;
      end else if (10'hf == _T_28[9:0]) begin
        image_0_15 <= io_pixelVal_in_0_4;
      end else if (10'hf == _T_25[9:0]) begin
        image_0_15 <= io_pixelVal_in_0_3;
      end else if (10'hf == _T_22[9:0]) begin
        image_0_15 <= io_pixelVal_in_0_2;
      end else if (10'hf == _T_19[9:0]) begin
        image_0_15 <= io_pixelVal_in_0_1;
      end else if (10'hf == _T_15[9:0]) begin
        image_0_15 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_16 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h10 == _T_37[9:0]) begin
        image_0_16 <= io_pixelVal_in_0_7;
      end else if (10'h10 == _T_34[9:0]) begin
        image_0_16 <= io_pixelVal_in_0_6;
      end else if (10'h10 == _T_31[9:0]) begin
        image_0_16 <= io_pixelVal_in_0_5;
      end else if (10'h10 == _T_28[9:0]) begin
        image_0_16 <= io_pixelVal_in_0_4;
      end else if (10'h10 == _T_25[9:0]) begin
        image_0_16 <= io_pixelVal_in_0_3;
      end else if (10'h10 == _T_22[9:0]) begin
        image_0_16 <= io_pixelVal_in_0_2;
      end else if (10'h10 == _T_19[9:0]) begin
        image_0_16 <= io_pixelVal_in_0_1;
      end else if (10'h10 == _T_15[9:0]) begin
        image_0_16 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_17 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h11 == _T_37[9:0]) begin
        image_0_17 <= io_pixelVal_in_0_7;
      end else if (10'h11 == _T_34[9:0]) begin
        image_0_17 <= io_pixelVal_in_0_6;
      end else if (10'h11 == _T_31[9:0]) begin
        image_0_17 <= io_pixelVal_in_0_5;
      end else if (10'h11 == _T_28[9:0]) begin
        image_0_17 <= io_pixelVal_in_0_4;
      end else if (10'h11 == _T_25[9:0]) begin
        image_0_17 <= io_pixelVal_in_0_3;
      end else if (10'h11 == _T_22[9:0]) begin
        image_0_17 <= io_pixelVal_in_0_2;
      end else if (10'h11 == _T_19[9:0]) begin
        image_0_17 <= io_pixelVal_in_0_1;
      end else if (10'h11 == _T_15[9:0]) begin
        image_0_17 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_18 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h12 == _T_37[9:0]) begin
        image_0_18 <= io_pixelVal_in_0_7;
      end else if (10'h12 == _T_34[9:0]) begin
        image_0_18 <= io_pixelVal_in_0_6;
      end else if (10'h12 == _T_31[9:0]) begin
        image_0_18 <= io_pixelVal_in_0_5;
      end else if (10'h12 == _T_28[9:0]) begin
        image_0_18 <= io_pixelVal_in_0_4;
      end else if (10'h12 == _T_25[9:0]) begin
        image_0_18 <= io_pixelVal_in_0_3;
      end else if (10'h12 == _T_22[9:0]) begin
        image_0_18 <= io_pixelVal_in_0_2;
      end else if (10'h12 == _T_19[9:0]) begin
        image_0_18 <= io_pixelVal_in_0_1;
      end else if (10'h12 == _T_15[9:0]) begin
        image_0_18 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_19 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h13 == _T_37[9:0]) begin
        image_0_19 <= io_pixelVal_in_0_7;
      end else if (10'h13 == _T_34[9:0]) begin
        image_0_19 <= io_pixelVal_in_0_6;
      end else if (10'h13 == _T_31[9:0]) begin
        image_0_19 <= io_pixelVal_in_0_5;
      end else if (10'h13 == _T_28[9:0]) begin
        image_0_19 <= io_pixelVal_in_0_4;
      end else if (10'h13 == _T_25[9:0]) begin
        image_0_19 <= io_pixelVal_in_0_3;
      end else if (10'h13 == _T_22[9:0]) begin
        image_0_19 <= io_pixelVal_in_0_2;
      end else if (10'h13 == _T_19[9:0]) begin
        image_0_19 <= io_pixelVal_in_0_1;
      end else if (10'h13 == _T_15[9:0]) begin
        image_0_19 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_20 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h14 == _T_37[9:0]) begin
        image_0_20 <= io_pixelVal_in_0_7;
      end else if (10'h14 == _T_34[9:0]) begin
        image_0_20 <= io_pixelVal_in_0_6;
      end else if (10'h14 == _T_31[9:0]) begin
        image_0_20 <= io_pixelVal_in_0_5;
      end else if (10'h14 == _T_28[9:0]) begin
        image_0_20 <= io_pixelVal_in_0_4;
      end else if (10'h14 == _T_25[9:0]) begin
        image_0_20 <= io_pixelVal_in_0_3;
      end else if (10'h14 == _T_22[9:0]) begin
        image_0_20 <= io_pixelVal_in_0_2;
      end else if (10'h14 == _T_19[9:0]) begin
        image_0_20 <= io_pixelVal_in_0_1;
      end else if (10'h14 == _T_15[9:0]) begin
        image_0_20 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_21 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h15 == _T_37[9:0]) begin
        image_0_21 <= io_pixelVal_in_0_7;
      end else if (10'h15 == _T_34[9:0]) begin
        image_0_21 <= io_pixelVal_in_0_6;
      end else if (10'h15 == _T_31[9:0]) begin
        image_0_21 <= io_pixelVal_in_0_5;
      end else if (10'h15 == _T_28[9:0]) begin
        image_0_21 <= io_pixelVal_in_0_4;
      end else if (10'h15 == _T_25[9:0]) begin
        image_0_21 <= io_pixelVal_in_0_3;
      end else if (10'h15 == _T_22[9:0]) begin
        image_0_21 <= io_pixelVal_in_0_2;
      end else if (10'h15 == _T_19[9:0]) begin
        image_0_21 <= io_pixelVal_in_0_1;
      end else if (10'h15 == _T_15[9:0]) begin
        image_0_21 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_22 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h16 == _T_37[9:0]) begin
        image_0_22 <= io_pixelVal_in_0_7;
      end else if (10'h16 == _T_34[9:0]) begin
        image_0_22 <= io_pixelVal_in_0_6;
      end else if (10'h16 == _T_31[9:0]) begin
        image_0_22 <= io_pixelVal_in_0_5;
      end else if (10'h16 == _T_28[9:0]) begin
        image_0_22 <= io_pixelVal_in_0_4;
      end else if (10'h16 == _T_25[9:0]) begin
        image_0_22 <= io_pixelVal_in_0_3;
      end else if (10'h16 == _T_22[9:0]) begin
        image_0_22 <= io_pixelVal_in_0_2;
      end else if (10'h16 == _T_19[9:0]) begin
        image_0_22 <= io_pixelVal_in_0_1;
      end else if (10'h16 == _T_15[9:0]) begin
        image_0_22 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_23 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h17 == _T_37[9:0]) begin
        image_0_23 <= io_pixelVal_in_0_7;
      end else if (10'h17 == _T_34[9:0]) begin
        image_0_23 <= io_pixelVal_in_0_6;
      end else if (10'h17 == _T_31[9:0]) begin
        image_0_23 <= io_pixelVal_in_0_5;
      end else if (10'h17 == _T_28[9:0]) begin
        image_0_23 <= io_pixelVal_in_0_4;
      end else if (10'h17 == _T_25[9:0]) begin
        image_0_23 <= io_pixelVal_in_0_3;
      end else if (10'h17 == _T_22[9:0]) begin
        image_0_23 <= io_pixelVal_in_0_2;
      end else if (10'h17 == _T_19[9:0]) begin
        image_0_23 <= io_pixelVal_in_0_1;
      end else if (10'h17 == _T_15[9:0]) begin
        image_0_23 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_24 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h18 == _T_37[9:0]) begin
        image_0_24 <= io_pixelVal_in_0_7;
      end else if (10'h18 == _T_34[9:0]) begin
        image_0_24 <= io_pixelVal_in_0_6;
      end else if (10'h18 == _T_31[9:0]) begin
        image_0_24 <= io_pixelVal_in_0_5;
      end else if (10'h18 == _T_28[9:0]) begin
        image_0_24 <= io_pixelVal_in_0_4;
      end else if (10'h18 == _T_25[9:0]) begin
        image_0_24 <= io_pixelVal_in_0_3;
      end else if (10'h18 == _T_22[9:0]) begin
        image_0_24 <= io_pixelVal_in_0_2;
      end else if (10'h18 == _T_19[9:0]) begin
        image_0_24 <= io_pixelVal_in_0_1;
      end else if (10'h18 == _T_15[9:0]) begin
        image_0_24 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_25 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h19 == _T_37[9:0]) begin
        image_0_25 <= io_pixelVal_in_0_7;
      end else if (10'h19 == _T_34[9:0]) begin
        image_0_25 <= io_pixelVal_in_0_6;
      end else if (10'h19 == _T_31[9:0]) begin
        image_0_25 <= io_pixelVal_in_0_5;
      end else if (10'h19 == _T_28[9:0]) begin
        image_0_25 <= io_pixelVal_in_0_4;
      end else if (10'h19 == _T_25[9:0]) begin
        image_0_25 <= io_pixelVal_in_0_3;
      end else if (10'h19 == _T_22[9:0]) begin
        image_0_25 <= io_pixelVal_in_0_2;
      end else if (10'h19 == _T_19[9:0]) begin
        image_0_25 <= io_pixelVal_in_0_1;
      end else if (10'h19 == _T_15[9:0]) begin
        image_0_25 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_26 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1a == _T_37[9:0]) begin
        image_0_26 <= io_pixelVal_in_0_7;
      end else if (10'h1a == _T_34[9:0]) begin
        image_0_26 <= io_pixelVal_in_0_6;
      end else if (10'h1a == _T_31[9:0]) begin
        image_0_26 <= io_pixelVal_in_0_5;
      end else if (10'h1a == _T_28[9:0]) begin
        image_0_26 <= io_pixelVal_in_0_4;
      end else if (10'h1a == _T_25[9:0]) begin
        image_0_26 <= io_pixelVal_in_0_3;
      end else if (10'h1a == _T_22[9:0]) begin
        image_0_26 <= io_pixelVal_in_0_2;
      end else if (10'h1a == _T_19[9:0]) begin
        image_0_26 <= io_pixelVal_in_0_1;
      end else if (10'h1a == _T_15[9:0]) begin
        image_0_26 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_27 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1b == _T_37[9:0]) begin
        image_0_27 <= io_pixelVal_in_0_7;
      end else if (10'h1b == _T_34[9:0]) begin
        image_0_27 <= io_pixelVal_in_0_6;
      end else if (10'h1b == _T_31[9:0]) begin
        image_0_27 <= io_pixelVal_in_0_5;
      end else if (10'h1b == _T_28[9:0]) begin
        image_0_27 <= io_pixelVal_in_0_4;
      end else if (10'h1b == _T_25[9:0]) begin
        image_0_27 <= io_pixelVal_in_0_3;
      end else if (10'h1b == _T_22[9:0]) begin
        image_0_27 <= io_pixelVal_in_0_2;
      end else if (10'h1b == _T_19[9:0]) begin
        image_0_27 <= io_pixelVal_in_0_1;
      end else if (10'h1b == _T_15[9:0]) begin
        image_0_27 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_28 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1c == _T_37[9:0]) begin
        image_0_28 <= io_pixelVal_in_0_7;
      end else if (10'h1c == _T_34[9:0]) begin
        image_0_28 <= io_pixelVal_in_0_6;
      end else if (10'h1c == _T_31[9:0]) begin
        image_0_28 <= io_pixelVal_in_0_5;
      end else if (10'h1c == _T_28[9:0]) begin
        image_0_28 <= io_pixelVal_in_0_4;
      end else if (10'h1c == _T_25[9:0]) begin
        image_0_28 <= io_pixelVal_in_0_3;
      end else if (10'h1c == _T_22[9:0]) begin
        image_0_28 <= io_pixelVal_in_0_2;
      end else if (10'h1c == _T_19[9:0]) begin
        image_0_28 <= io_pixelVal_in_0_1;
      end else if (10'h1c == _T_15[9:0]) begin
        image_0_28 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_29 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1d == _T_37[9:0]) begin
        image_0_29 <= io_pixelVal_in_0_7;
      end else if (10'h1d == _T_34[9:0]) begin
        image_0_29 <= io_pixelVal_in_0_6;
      end else if (10'h1d == _T_31[9:0]) begin
        image_0_29 <= io_pixelVal_in_0_5;
      end else if (10'h1d == _T_28[9:0]) begin
        image_0_29 <= io_pixelVal_in_0_4;
      end else if (10'h1d == _T_25[9:0]) begin
        image_0_29 <= io_pixelVal_in_0_3;
      end else if (10'h1d == _T_22[9:0]) begin
        image_0_29 <= io_pixelVal_in_0_2;
      end else if (10'h1d == _T_19[9:0]) begin
        image_0_29 <= io_pixelVal_in_0_1;
      end else if (10'h1d == _T_15[9:0]) begin
        image_0_29 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_30 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1e == _T_37[9:0]) begin
        image_0_30 <= io_pixelVal_in_0_7;
      end else if (10'h1e == _T_34[9:0]) begin
        image_0_30 <= io_pixelVal_in_0_6;
      end else if (10'h1e == _T_31[9:0]) begin
        image_0_30 <= io_pixelVal_in_0_5;
      end else if (10'h1e == _T_28[9:0]) begin
        image_0_30 <= io_pixelVal_in_0_4;
      end else if (10'h1e == _T_25[9:0]) begin
        image_0_30 <= io_pixelVal_in_0_3;
      end else if (10'h1e == _T_22[9:0]) begin
        image_0_30 <= io_pixelVal_in_0_2;
      end else if (10'h1e == _T_19[9:0]) begin
        image_0_30 <= io_pixelVal_in_0_1;
      end else if (10'h1e == _T_15[9:0]) begin
        image_0_30 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_31 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1f == _T_37[9:0]) begin
        image_0_31 <= io_pixelVal_in_0_7;
      end else if (10'h1f == _T_34[9:0]) begin
        image_0_31 <= io_pixelVal_in_0_6;
      end else if (10'h1f == _T_31[9:0]) begin
        image_0_31 <= io_pixelVal_in_0_5;
      end else if (10'h1f == _T_28[9:0]) begin
        image_0_31 <= io_pixelVal_in_0_4;
      end else if (10'h1f == _T_25[9:0]) begin
        image_0_31 <= io_pixelVal_in_0_3;
      end else if (10'h1f == _T_22[9:0]) begin
        image_0_31 <= io_pixelVal_in_0_2;
      end else if (10'h1f == _T_19[9:0]) begin
        image_0_31 <= io_pixelVal_in_0_1;
      end else if (10'h1f == _T_15[9:0]) begin
        image_0_31 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_32 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h20 == _T_37[9:0]) begin
        image_0_32 <= io_pixelVal_in_0_7;
      end else if (10'h20 == _T_34[9:0]) begin
        image_0_32 <= io_pixelVal_in_0_6;
      end else if (10'h20 == _T_31[9:0]) begin
        image_0_32 <= io_pixelVal_in_0_5;
      end else if (10'h20 == _T_28[9:0]) begin
        image_0_32 <= io_pixelVal_in_0_4;
      end else if (10'h20 == _T_25[9:0]) begin
        image_0_32 <= io_pixelVal_in_0_3;
      end else if (10'h20 == _T_22[9:0]) begin
        image_0_32 <= io_pixelVal_in_0_2;
      end else if (10'h20 == _T_19[9:0]) begin
        image_0_32 <= io_pixelVal_in_0_1;
      end else if (10'h20 == _T_15[9:0]) begin
        image_0_32 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_33 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h21 == _T_37[9:0]) begin
        image_0_33 <= io_pixelVal_in_0_7;
      end else if (10'h21 == _T_34[9:0]) begin
        image_0_33 <= io_pixelVal_in_0_6;
      end else if (10'h21 == _T_31[9:0]) begin
        image_0_33 <= io_pixelVal_in_0_5;
      end else if (10'h21 == _T_28[9:0]) begin
        image_0_33 <= io_pixelVal_in_0_4;
      end else if (10'h21 == _T_25[9:0]) begin
        image_0_33 <= io_pixelVal_in_0_3;
      end else if (10'h21 == _T_22[9:0]) begin
        image_0_33 <= io_pixelVal_in_0_2;
      end else if (10'h21 == _T_19[9:0]) begin
        image_0_33 <= io_pixelVal_in_0_1;
      end else if (10'h21 == _T_15[9:0]) begin
        image_0_33 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_34 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h22 == _T_37[9:0]) begin
        image_0_34 <= io_pixelVal_in_0_7;
      end else if (10'h22 == _T_34[9:0]) begin
        image_0_34 <= io_pixelVal_in_0_6;
      end else if (10'h22 == _T_31[9:0]) begin
        image_0_34 <= io_pixelVal_in_0_5;
      end else if (10'h22 == _T_28[9:0]) begin
        image_0_34 <= io_pixelVal_in_0_4;
      end else if (10'h22 == _T_25[9:0]) begin
        image_0_34 <= io_pixelVal_in_0_3;
      end else if (10'h22 == _T_22[9:0]) begin
        image_0_34 <= io_pixelVal_in_0_2;
      end else if (10'h22 == _T_19[9:0]) begin
        image_0_34 <= io_pixelVal_in_0_1;
      end else if (10'h22 == _T_15[9:0]) begin
        image_0_34 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_35 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h23 == _T_37[9:0]) begin
        image_0_35 <= io_pixelVal_in_0_7;
      end else if (10'h23 == _T_34[9:0]) begin
        image_0_35 <= io_pixelVal_in_0_6;
      end else if (10'h23 == _T_31[9:0]) begin
        image_0_35 <= io_pixelVal_in_0_5;
      end else if (10'h23 == _T_28[9:0]) begin
        image_0_35 <= io_pixelVal_in_0_4;
      end else if (10'h23 == _T_25[9:0]) begin
        image_0_35 <= io_pixelVal_in_0_3;
      end else if (10'h23 == _T_22[9:0]) begin
        image_0_35 <= io_pixelVal_in_0_2;
      end else if (10'h23 == _T_19[9:0]) begin
        image_0_35 <= io_pixelVal_in_0_1;
      end else if (10'h23 == _T_15[9:0]) begin
        image_0_35 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_36 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h24 == _T_37[9:0]) begin
        image_0_36 <= io_pixelVal_in_0_7;
      end else if (10'h24 == _T_34[9:0]) begin
        image_0_36 <= io_pixelVal_in_0_6;
      end else if (10'h24 == _T_31[9:0]) begin
        image_0_36 <= io_pixelVal_in_0_5;
      end else if (10'h24 == _T_28[9:0]) begin
        image_0_36 <= io_pixelVal_in_0_4;
      end else if (10'h24 == _T_25[9:0]) begin
        image_0_36 <= io_pixelVal_in_0_3;
      end else if (10'h24 == _T_22[9:0]) begin
        image_0_36 <= io_pixelVal_in_0_2;
      end else if (10'h24 == _T_19[9:0]) begin
        image_0_36 <= io_pixelVal_in_0_1;
      end else if (10'h24 == _T_15[9:0]) begin
        image_0_36 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_37 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h25 == _T_37[9:0]) begin
        image_0_37 <= io_pixelVal_in_0_7;
      end else if (10'h25 == _T_34[9:0]) begin
        image_0_37 <= io_pixelVal_in_0_6;
      end else if (10'h25 == _T_31[9:0]) begin
        image_0_37 <= io_pixelVal_in_0_5;
      end else if (10'h25 == _T_28[9:0]) begin
        image_0_37 <= io_pixelVal_in_0_4;
      end else if (10'h25 == _T_25[9:0]) begin
        image_0_37 <= io_pixelVal_in_0_3;
      end else if (10'h25 == _T_22[9:0]) begin
        image_0_37 <= io_pixelVal_in_0_2;
      end else if (10'h25 == _T_19[9:0]) begin
        image_0_37 <= io_pixelVal_in_0_1;
      end else if (10'h25 == _T_15[9:0]) begin
        image_0_37 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_38 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h26 == _T_37[9:0]) begin
        image_0_38 <= io_pixelVal_in_0_7;
      end else if (10'h26 == _T_34[9:0]) begin
        image_0_38 <= io_pixelVal_in_0_6;
      end else if (10'h26 == _T_31[9:0]) begin
        image_0_38 <= io_pixelVal_in_0_5;
      end else if (10'h26 == _T_28[9:0]) begin
        image_0_38 <= io_pixelVal_in_0_4;
      end else if (10'h26 == _T_25[9:0]) begin
        image_0_38 <= io_pixelVal_in_0_3;
      end else if (10'h26 == _T_22[9:0]) begin
        image_0_38 <= io_pixelVal_in_0_2;
      end else if (10'h26 == _T_19[9:0]) begin
        image_0_38 <= io_pixelVal_in_0_1;
      end else if (10'h26 == _T_15[9:0]) begin
        image_0_38 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_39 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h27 == _T_37[9:0]) begin
        image_0_39 <= io_pixelVal_in_0_7;
      end else if (10'h27 == _T_34[9:0]) begin
        image_0_39 <= io_pixelVal_in_0_6;
      end else if (10'h27 == _T_31[9:0]) begin
        image_0_39 <= io_pixelVal_in_0_5;
      end else if (10'h27 == _T_28[9:0]) begin
        image_0_39 <= io_pixelVal_in_0_4;
      end else if (10'h27 == _T_25[9:0]) begin
        image_0_39 <= io_pixelVal_in_0_3;
      end else if (10'h27 == _T_22[9:0]) begin
        image_0_39 <= io_pixelVal_in_0_2;
      end else if (10'h27 == _T_19[9:0]) begin
        image_0_39 <= io_pixelVal_in_0_1;
      end else if (10'h27 == _T_15[9:0]) begin
        image_0_39 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_40 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h28 == _T_37[9:0]) begin
        image_0_40 <= io_pixelVal_in_0_7;
      end else if (10'h28 == _T_34[9:0]) begin
        image_0_40 <= io_pixelVal_in_0_6;
      end else if (10'h28 == _T_31[9:0]) begin
        image_0_40 <= io_pixelVal_in_0_5;
      end else if (10'h28 == _T_28[9:0]) begin
        image_0_40 <= io_pixelVal_in_0_4;
      end else if (10'h28 == _T_25[9:0]) begin
        image_0_40 <= io_pixelVal_in_0_3;
      end else if (10'h28 == _T_22[9:0]) begin
        image_0_40 <= io_pixelVal_in_0_2;
      end else if (10'h28 == _T_19[9:0]) begin
        image_0_40 <= io_pixelVal_in_0_1;
      end else if (10'h28 == _T_15[9:0]) begin
        image_0_40 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_41 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h29 == _T_37[9:0]) begin
        image_0_41 <= io_pixelVal_in_0_7;
      end else if (10'h29 == _T_34[9:0]) begin
        image_0_41 <= io_pixelVal_in_0_6;
      end else if (10'h29 == _T_31[9:0]) begin
        image_0_41 <= io_pixelVal_in_0_5;
      end else if (10'h29 == _T_28[9:0]) begin
        image_0_41 <= io_pixelVal_in_0_4;
      end else if (10'h29 == _T_25[9:0]) begin
        image_0_41 <= io_pixelVal_in_0_3;
      end else if (10'h29 == _T_22[9:0]) begin
        image_0_41 <= io_pixelVal_in_0_2;
      end else if (10'h29 == _T_19[9:0]) begin
        image_0_41 <= io_pixelVal_in_0_1;
      end else if (10'h29 == _T_15[9:0]) begin
        image_0_41 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_42 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h2a == _T_37[9:0]) begin
        image_0_42 <= io_pixelVal_in_0_7;
      end else if (10'h2a == _T_34[9:0]) begin
        image_0_42 <= io_pixelVal_in_0_6;
      end else if (10'h2a == _T_31[9:0]) begin
        image_0_42 <= io_pixelVal_in_0_5;
      end else if (10'h2a == _T_28[9:0]) begin
        image_0_42 <= io_pixelVal_in_0_4;
      end else if (10'h2a == _T_25[9:0]) begin
        image_0_42 <= io_pixelVal_in_0_3;
      end else if (10'h2a == _T_22[9:0]) begin
        image_0_42 <= io_pixelVal_in_0_2;
      end else if (10'h2a == _T_19[9:0]) begin
        image_0_42 <= io_pixelVal_in_0_1;
      end else if (10'h2a == _T_15[9:0]) begin
        image_0_42 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_43 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h2b == _T_37[9:0]) begin
        image_0_43 <= io_pixelVal_in_0_7;
      end else if (10'h2b == _T_34[9:0]) begin
        image_0_43 <= io_pixelVal_in_0_6;
      end else if (10'h2b == _T_31[9:0]) begin
        image_0_43 <= io_pixelVal_in_0_5;
      end else if (10'h2b == _T_28[9:0]) begin
        image_0_43 <= io_pixelVal_in_0_4;
      end else if (10'h2b == _T_25[9:0]) begin
        image_0_43 <= io_pixelVal_in_0_3;
      end else if (10'h2b == _T_22[9:0]) begin
        image_0_43 <= io_pixelVal_in_0_2;
      end else if (10'h2b == _T_19[9:0]) begin
        image_0_43 <= io_pixelVal_in_0_1;
      end else if (10'h2b == _T_15[9:0]) begin
        image_0_43 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_44 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h2c == _T_37[9:0]) begin
        image_0_44 <= io_pixelVal_in_0_7;
      end else if (10'h2c == _T_34[9:0]) begin
        image_0_44 <= io_pixelVal_in_0_6;
      end else if (10'h2c == _T_31[9:0]) begin
        image_0_44 <= io_pixelVal_in_0_5;
      end else if (10'h2c == _T_28[9:0]) begin
        image_0_44 <= io_pixelVal_in_0_4;
      end else if (10'h2c == _T_25[9:0]) begin
        image_0_44 <= io_pixelVal_in_0_3;
      end else if (10'h2c == _T_22[9:0]) begin
        image_0_44 <= io_pixelVal_in_0_2;
      end else if (10'h2c == _T_19[9:0]) begin
        image_0_44 <= io_pixelVal_in_0_1;
      end else if (10'h2c == _T_15[9:0]) begin
        image_0_44 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_45 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h2d == _T_37[9:0]) begin
        image_0_45 <= io_pixelVal_in_0_7;
      end else if (10'h2d == _T_34[9:0]) begin
        image_0_45 <= io_pixelVal_in_0_6;
      end else if (10'h2d == _T_31[9:0]) begin
        image_0_45 <= io_pixelVal_in_0_5;
      end else if (10'h2d == _T_28[9:0]) begin
        image_0_45 <= io_pixelVal_in_0_4;
      end else if (10'h2d == _T_25[9:0]) begin
        image_0_45 <= io_pixelVal_in_0_3;
      end else if (10'h2d == _T_22[9:0]) begin
        image_0_45 <= io_pixelVal_in_0_2;
      end else if (10'h2d == _T_19[9:0]) begin
        image_0_45 <= io_pixelVal_in_0_1;
      end else if (10'h2d == _T_15[9:0]) begin
        image_0_45 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_46 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h2e == _T_37[9:0]) begin
        image_0_46 <= io_pixelVal_in_0_7;
      end else if (10'h2e == _T_34[9:0]) begin
        image_0_46 <= io_pixelVal_in_0_6;
      end else if (10'h2e == _T_31[9:0]) begin
        image_0_46 <= io_pixelVal_in_0_5;
      end else if (10'h2e == _T_28[9:0]) begin
        image_0_46 <= io_pixelVal_in_0_4;
      end else if (10'h2e == _T_25[9:0]) begin
        image_0_46 <= io_pixelVal_in_0_3;
      end else if (10'h2e == _T_22[9:0]) begin
        image_0_46 <= io_pixelVal_in_0_2;
      end else if (10'h2e == _T_19[9:0]) begin
        image_0_46 <= io_pixelVal_in_0_1;
      end else if (10'h2e == _T_15[9:0]) begin
        image_0_46 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_47 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h2f == _T_37[9:0]) begin
        image_0_47 <= io_pixelVal_in_0_7;
      end else if (10'h2f == _T_34[9:0]) begin
        image_0_47 <= io_pixelVal_in_0_6;
      end else if (10'h2f == _T_31[9:0]) begin
        image_0_47 <= io_pixelVal_in_0_5;
      end else if (10'h2f == _T_28[9:0]) begin
        image_0_47 <= io_pixelVal_in_0_4;
      end else if (10'h2f == _T_25[9:0]) begin
        image_0_47 <= io_pixelVal_in_0_3;
      end else if (10'h2f == _T_22[9:0]) begin
        image_0_47 <= io_pixelVal_in_0_2;
      end else if (10'h2f == _T_19[9:0]) begin
        image_0_47 <= io_pixelVal_in_0_1;
      end else if (10'h2f == _T_15[9:0]) begin
        image_0_47 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_48 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h30 == _T_37[9:0]) begin
        image_0_48 <= io_pixelVal_in_0_7;
      end else if (10'h30 == _T_34[9:0]) begin
        image_0_48 <= io_pixelVal_in_0_6;
      end else if (10'h30 == _T_31[9:0]) begin
        image_0_48 <= io_pixelVal_in_0_5;
      end else if (10'h30 == _T_28[9:0]) begin
        image_0_48 <= io_pixelVal_in_0_4;
      end else if (10'h30 == _T_25[9:0]) begin
        image_0_48 <= io_pixelVal_in_0_3;
      end else if (10'h30 == _T_22[9:0]) begin
        image_0_48 <= io_pixelVal_in_0_2;
      end else if (10'h30 == _T_19[9:0]) begin
        image_0_48 <= io_pixelVal_in_0_1;
      end else if (10'h30 == _T_15[9:0]) begin
        image_0_48 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_49 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h31 == _T_37[9:0]) begin
        image_0_49 <= io_pixelVal_in_0_7;
      end else if (10'h31 == _T_34[9:0]) begin
        image_0_49 <= io_pixelVal_in_0_6;
      end else if (10'h31 == _T_31[9:0]) begin
        image_0_49 <= io_pixelVal_in_0_5;
      end else if (10'h31 == _T_28[9:0]) begin
        image_0_49 <= io_pixelVal_in_0_4;
      end else if (10'h31 == _T_25[9:0]) begin
        image_0_49 <= io_pixelVal_in_0_3;
      end else if (10'h31 == _T_22[9:0]) begin
        image_0_49 <= io_pixelVal_in_0_2;
      end else if (10'h31 == _T_19[9:0]) begin
        image_0_49 <= io_pixelVal_in_0_1;
      end else if (10'h31 == _T_15[9:0]) begin
        image_0_49 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_50 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h32 == _T_37[9:0]) begin
        image_0_50 <= io_pixelVal_in_0_7;
      end else if (10'h32 == _T_34[9:0]) begin
        image_0_50 <= io_pixelVal_in_0_6;
      end else if (10'h32 == _T_31[9:0]) begin
        image_0_50 <= io_pixelVal_in_0_5;
      end else if (10'h32 == _T_28[9:0]) begin
        image_0_50 <= io_pixelVal_in_0_4;
      end else if (10'h32 == _T_25[9:0]) begin
        image_0_50 <= io_pixelVal_in_0_3;
      end else if (10'h32 == _T_22[9:0]) begin
        image_0_50 <= io_pixelVal_in_0_2;
      end else if (10'h32 == _T_19[9:0]) begin
        image_0_50 <= io_pixelVal_in_0_1;
      end else if (10'h32 == _T_15[9:0]) begin
        image_0_50 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_51 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h33 == _T_37[9:0]) begin
        image_0_51 <= io_pixelVal_in_0_7;
      end else if (10'h33 == _T_34[9:0]) begin
        image_0_51 <= io_pixelVal_in_0_6;
      end else if (10'h33 == _T_31[9:0]) begin
        image_0_51 <= io_pixelVal_in_0_5;
      end else if (10'h33 == _T_28[9:0]) begin
        image_0_51 <= io_pixelVal_in_0_4;
      end else if (10'h33 == _T_25[9:0]) begin
        image_0_51 <= io_pixelVal_in_0_3;
      end else if (10'h33 == _T_22[9:0]) begin
        image_0_51 <= io_pixelVal_in_0_2;
      end else if (10'h33 == _T_19[9:0]) begin
        image_0_51 <= io_pixelVal_in_0_1;
      end else if (10'h33 == _T_15[9:0]) begin
        image_0_51 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_52 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h34 == _T_37[9:0]) begin
        image_0_52 <= io_pixelVal_in_0_7;
      end else if (10'h34 == _T_34[9:0]) begin
        image_0_52 <= io_pixelVal_in_0_6;
      end else if (10'h34 == _T_31[9:0]) begin
        image_0_52 <= io_pixelVal_in_0_5;
      end else if (10'h34 == _T_28[9:0]) begin
        image_0_52 <= io_pixelVal_in_0_4;
      end else if (10'h34 == _T_25[9:0]) begin
        image_0_52 <= io_pixelVal_in_0_3;
      end else if (10'h34 == _T_22[9:0]) begin
        image_0_52 <= io_pixelVal_in_0_2;
      end else if (10'h34 == _T_19[9:0]) begin
        image_0_52 <= io_pixelVal_in_0_1;
      end else if (10'h34 == _T_15[9:0]) begin
        image_0_52 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_53 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h35 == _T_37[9:0]) begin
        image_0_53 <= io_pixelVal_in_0_7;
      end else if (10'h35 == _T_34[9:0]) begin
        image_0_53 <= io_pixelVal_in_0_6;
      end else if (10'h35 == _T_31[9:0]) begin
        image_0_53 <= io_pixelVal_in_0_5;
      end else if (10'h35 == _T_28[9:0]) begin
        image_0_53 <= io_pixelVal_in_0_4;
      end else if (10'h35 == _T_25[9:0]) begin
        image_0_53 <= io_pixelVal_in_0_3;
      end else if (10'h35 == _T_22[9:0]) begin
        image_0_53 <= io_pixelVal_in_0_2;
      end else if (10'h35 == _T_19[9:0]) begin
        image_0_53 <= io_pixelVal_in_0_1;
      end else if (10'h35 == _T_15[9:0]) begin
        image_0_53 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_54 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h36 == _T_37[9:0]) begin
        image_0_54 <= io_pixelVal_in_0_7;
      end else if (10'h36 == _T_34[9:0]) begin
        image_0_54 <= io_pixelVal_in_0_6;
      end else if (10'h36 == _T_31[9:0]) begin
        image_0_54 <= io_pixelVal_in_0_5;
      end else if (10'h36 == _T_28[9:0]) begin
        image_0_54 <= io_pixelVal_in_0_4;
      end else if (10'h36 == _T_25[9:0]) begin
        image_0_54 <= io_pixelVal_in_0_3;
      end else if (10'h36 == _T_22[9:0]) begin
        image_0_54 <= io_pixelVal_in_0_2;
      end else if (10'h36 == _T_19[9:0]) begin
        image_0_54 <= io_pixelVal_in_0_1;
      end else if (10'h36 == _T_15[9:0]) begin
        image_0_54 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_55 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h37 == _T_37[9:0]) begin
        image_0_55 <= io_pixelVal_in_0_7;
      end else if (10'h37 == _T_34[9:0]) begin
        image_0_55 <= io_pixelVal_in_0_6;
      end else if (10'h37 == _T_31[9:0]) begin
        image_0_55 <= io_pixelVal_in_0_5;
      end else if (10'h37 == _T_28[9:0]) begin
        image_0_55 <= io_pixelVal_in_0_4;
      end else if (10'h37 == _T_25[9:0]) begin
        image_0_55 <= io_pixelVal_in_0_3;
      end else if (10'h37 == _T_22[9:0]) begin
        image_0_55 <= io_pixelVal_in_0_2;
      end else if (10'h37 == _T_19[9:0]) begin
        image_0_55 <= io_pixelVal_in_0_1;
      end else if (10'h37 == _T_15[9:0]) begin
        image_0_55 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_56 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h38 == _T_37[9:0]) begin
        image_0_56 <= io_pixelVal_in_0_7;
      end else if (10'h38 == _T_34[9:0]) begin
        image_0_56 <= io_pixelVal_in_0_6;
      end else if (10'h38 == _T_31[9:0]) begin
        image_0_56 <= io_pixelVal_in_0_5;
      end else if (10'h38 == _T_28[9:0]) begin
        image_0_56 <= io_pixelVal_in_0_4;
      end else if (10'h38 == _T_25[9:0]) begin
        image_0_56 <= io_pixelVal_in_0_3;
      end else if (10'h38 == _T_22[9:0]) begin
        image_0_56 <= io_pixelVal_in_0_2;
      end else if (10'h38 == _T_19[9:0]) begin
        image_0_56 <= io_pixelVal_in_0_1;
      end else if (10'h38 == _T_15[9:0]) begin
        image_0_56 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_57 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h39 == _T_37[9:0]) begin
        image_0_57 <= io_pixelVal_in_0_7;
      end else if (10'h39 == _T_34[9:0]) begin
        image_0_57 <= io_pixelVal_in_0_6;
      end else if (10'h39 == _T_31[9:0]) begin
        image_0_57 <= io_pixelVal_in_0_5;
      end else if (10'h39 == _T_28[9:0]) begin
        image_0_57 <= io_pixelVal_in_0_4;
      end else if (10'h39 == _T_25[9:0]) begin
        image_0_57 <= io_pixelVal_in_0_3;
      end else if (10'h39 == _T_22[9:0]) begin
        image_0_57 <= io_pixelVal_in_0_2;
      end else if (10'h39 == _T_19[9:0]) begin
        image_0_57 <= io_pixelVal_in_0_1;
      end else if (10'h39 == _T_15[9:0]) begin
        image_0_57 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_58 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h3a == _T_37[9:0]) begin
        image_0_58 <= io_pixelVal_in_0_7;
      end else if (10'h3a == _T_34[9:0]) begin
        image_0_58 <= io_pixelVal_in_0_6;
      end else if (10'h3a == _T_31[9:0]) begin
        image_0_58 <= io_pixelVal_in_0_5;
      end else if (10'h3a == _T_28[9:0]) begin
        image_0_58 <= io_pixelVal_in_0_4;
      end else if (10'h3a == _T_25[9:0]) begin
        image_0_58 <= io_pixelVal_in_0_3;
      end else if (10'h3a == _T_22[9:0]) begin
        image_0_58 <= io_pixelVal_in_0_2;
      end else if (10'h3a == _T_19[9:0]) begin
        image_0_58 <= io_pixelVal_in_0_1;
      end else if (10'h3a == _T_15[9:0]) begin
        image_0_58 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_59 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h3b == _T_37[9:0]) begin
        image_0_59 <= io_pixelVal_in_0_7;
      end else if (10'h3b == _T_34[9:0]) begin
        image_0_59 <= io_pixelVal_in_0_6;
      end else if (10'h3b == _T_31[9:0]) begin
        image_0_59 <= io_pixelVal_in_0_5;
      end else if (10'h3b == _T_28[9:0]) begin
        image_0_59 <= io_pixelVal_in_0_4;
      end else if (10'h3b == _T_25[9:0]) begin
        image_0_59 <= io_pixelVal_in_0_3;
      end else if (10'h3b == _T_22[9:0]) begin
        image_0_59 <= io_pixelVal_in_0_2;
      end else if (10'h3b == _T_19[9:0]) begin
        image_0_59 <= io_pixelVal_in_0_1;
      end else if (10'h3b == _T_15[9:0]) begin
        image_0_59 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_60 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h3c == _T_37[9:0]) begin
        image_0_60 <= io_pixelVal_in_0_7;
      end else if (10'h3c == _T_34[9:0]) begin
        image_0_60 <= io_pixelVal_in_0_6;
      end else if (10'h3c == _T_31[9:0]) begin
        image_0_60 <= io_pixelVal_in_0_5;
      end else if (10'h3c == _T_28[9:0]) begin
        image_0_60 <= io_pixelVal_in_0_4;
      end else if (10'h3c == _T_25[9:0]) begin
        image_0_60 <= io_pixelVal_in_0_3;
      end else if (10'h3c == _T_22[9:0]) begin
        image_0_60 <= io_pixelVal_in_0_2;
      end else if (10'h3c == _T_19[9:0]) begin
        image_0_60 <= io_pixelVal_in_0_1;
      end else if (10'h3c == _T_15[9:0]) begin
        image_0_60 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_61 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h3d == _T_37[9:0]) begin
        image_0_61 <= io_pixelVal_in_0_7;
      end else if (10'h3d == _T_34[9:0]) begin
        image_0_61 <= io_pixelVal_in_0_6;
      end else if (10'h3d == _T_31[9:0]) begin
        image_0_61 <= io_pixelVal_in_0_5;
      end else if (10'h3d == _T_28[9:0]) begin
        image_0_61 <= io_pixelVal_in_0_4;
      end else if (10'h3d == _T_25[9:0]) begin
        image_0_61 <= io_pixelVal_in_0_3;
      end else if (10'h3d == _T_22[9:0]) begin
        image_0_61 <= io_pixelVal_in_0_2;
      end else if (10'h3d == _T_19[9:0]) begin
        image_0_61 <= io_pixelVal_in_0_1;
      end else if (10'h3d == _T_15[9:0]) begin
        image_0_61 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_62 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h3e == _T_37[9:0]) begin
        image_0_62 <= io_pixelVal_in_0_7;
      end else if (10'h3e == _T_34[9:0]) begin
        image_0_62 <= io_pixelVal_in_0_6;
      end else if (10'h3e == _T_31[9:0]) begin
        image_0_62 <= io_pixelVal_in_0_5;
      end else if (10'h3e == _T_28[9:0]) begin
        image_0_62 <= io_pixelVal_in_0_4;
      end else if (10'h3e == _T_25[9:0]) begin
        image_0_62 <= io_pixelVal_in_0_3;
      end else if (10'h3e == _T_22[9:0]) begin
        image_0_62 <= io_pixelVal_in_0_2;
      end else if (10'h3e == _T_19[9:0]) begin
        image_0_62 <= io_pixelVal_in_0_1;
      end else if (10'h3e == _T_15[9:0]) begin
        image_0_62 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_63 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h3f == _T_37[9:0]) begin
        image_0_63 <= io_pixelVal_in_0_7;
      end else if (10'h3f == _T_34[9:0]) begin
        image_0_63 <= io_pixelVal_in_0_6;
      end else if (10'h3f == _T_31[9:0]) begin
        image_0_63 <= io_pixelVal_in_0_5;
      end else if (10'h3f == _T_28[9:0]) begin
        image_0_63 <= io_pixelVal_in_0_4;
      end else if (10'h3f == _T_25[9:0]) begin
        image_0_63 <= io_pixelVal_in_0_3;
      end else if (10'h3f == _T_22[9:0]) begin
        image_0_63 <= io_pixelVal_in_0_2;
      end else if (10'h3f == _T_19[9:0]) begin
        image_0_63 <= io_pixelVal_in_0_1;
      end else if (10'h3f == _T_15[9:0]) begin
        image_0_63 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_64 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h40 == _T_37[9:0]) begin
        image_0_64 <= io_pixelVal_in_0_7;
      end else if (10'h40 == _T_34[9:0]) begin
        image_0_64 <= io_pixelVal_in_0_6;
      end else if (10'h40 == _T_31[9:0]) begin
        image_0_64 <= io_pixelVal_in_0_5;
      end else if (10'h40 == _T_28[9:0]) begin
        image_0_64 <= io_pixelVal_in_0_4;
      end else if (10'h40 == _T_25[9:0]) begin
        image_0_64 <= io_pixelVal_in_0_3;
      end else if (10'h40 == _T_22[9:0]) begin
        image_0_64 <= io_pixelVal_in_0_2;
      end else if (10'h40 == _T_19[9:0]) begin
        image_0_64 <= io_pixelVal_in_0_1;
      end else if (10'h40 == _T_15[9:0]) begin
        image_0_64 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_65 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h41 == _T_37[9:0]) begin
        image_0_65 <= io_pixelVal_in_0_7;
      end else if (10'h41 == _T_34[9:0]) begin
        image_0_65 <= io_pixelVal_in_0_6;
      end else if (10'h41 == _T_31[9:0]) begin
        image_0_65 <= io_pixelVal_in_0_5;
      end else if (10'h41 == _T_28[9:0]) begin
        image_0_65 <= io_pixelVal_in_0_4;
      end else if (10'h41 == _T_25[9:0]) begin
        image_0_65 <= io_pixelVal_in_0_3;
      end else if (10'h41 == _T_22[9:0]) begin
        image_0_65 <= io_pixelVal_in_0_2;
      end else if (10'h41 == _T_19[9:0]) begin
        image_0_65 <= io_pixelVal_in_0_1;
      end else if (10'h41 == _T_15[9:0]) begin
        image_0_65 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_66 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h42 == _T_37[9:0]) begin
        image_0_66 <= io_pixelVal_in_0_7;
      end else if (10'h42 == _T_34[9:0]) begin
        image_0_66 <= io_pixelVal_in_0_6;
      end else if (10'h42 == _T_31[9:0]) begin
        image_0_66 <= io_pixelVal_in_0_5;
      end else if (10'h42 == _T_28[9:0]) begin
        image_0_66 <= io_pixelVal_in_0_4;
      end else if (10'h42 == _T_25[9:0]) begin
        image_0_66 <= io_pixelVal_in_0_3;
      end else if (10'h42 == _T_22[9:0]) begin
        image_0_66 <= io_pixelVal_in_0_2;
      end else if (10'h42 == _T_19[9:0]) begin
        image_0_66 <= io_pixelVal_in_0_1;
      end else if (10'h42 == _T_15[9:0]) begin
        image_0_66 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_67 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h43 == _T_37[9:0]) begin
        image_0_67 <= io_pixelVal_in_0_7;
      end else if (10'h43 == _T_34[9:0]) begin
        image_0_67 <= io_pixelVal_in_0_6;
      end else if (10'h43 == _T_31[9:0]) begin
        image_0_67 <= io_pixelVal_in_0_5;
      end else if (10'h43 == _T_28[9:0]) begin
        image_0_67 <= io_pixelVal_in_0_4;
      end else if (10'h43 == _T_25[9:0]) begin
        image_0_67 <= io_pixelVal_in_0_3;
      end else if (10'h43 == _T_22[9:0]) begin
        image_0_67 <= io_pixelVal_in_0_2;
      end else if (10'h43 == _T_19[9:0]) begin
        image_0_67 <= io_pixelVal_in_0_1;
      end else if (10'h43 == _T_15[9:0]) begin
        image_0_67 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_68 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h44 == _T_37[9:0]) begin
        image_0_68 <= io_pixelVal_in_0_7;
      end else if (10'h44 == _T_34[9:0]) begin
        image_0_68 <= io_pixelVal_in_0_6;
      end else if (10'h44 == _T_31[9:0]) begin
        image_0_68 <= io_pixelVal_in_0_5;
      end else if (10'h44 == _T_28[9:0]) begin
        image_0_68 <= io_pixelVal_in_0_4;
      end else if (10'h44 == _T_25[9:0]) begin
        image_0_68 <= io_pixelVal_in_0_3;
      end else if (10'h44 == _T_22[9:0]) begin
        image_0_68 <= io_pixelVal_in_0_2;
      end else if (10'h44 == _T_19[9:0]) begin
        image_0_68 <= io_pixelVal_in_0_1;
      end else if (10'h44 == _T_15[9:0]) begin
        image_0_68 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_69 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h45 == _T_37[9:0]) begin
        image_0_69 <= io_pixelVal_in_0_7;
      end else if (10'h45 == _T_34[9:0]) begin
        image_0_69 <= io_pixelVal_in_0_6;
      end else if (10'h45 == _T_31[9:0]) begin
        image_0_69 <= io_pixelVal_in_0_5;
      end else if (10'h45 == _T_28[9:0]) begin
        image_0_69 <= io_pixelVal_in_0_4;
      end else if (10'h45 == _T_25[9:0]) begin
        image_0_69 <= io_pixelVal_in_0_3;
      end else if (10'h45 == _T_22[9:0]) begin
        image_0_69 <= io_pixelVal_in_0_2;
      end else if (10'h45 == _T_19[9:0]) begin
        image_0_69 <= io_pixelVal_in_0_1;
      end else if (10'h45 == _T_15[9:0]) begin
        image_0_69 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_70 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h46 == _T_37[9:0]) begin
        image_0_70 <= io_pixelVal_in_0_7;
      end else if (10'h46 == _T_34[9:0]) begin
        image_0_70 <= io_pixelVal_in_0_6;
      end else if (10'h46 == _T_31[9:0]) begin
        image_0_70 <= io_pixelVal_in_0_5;
      end else if (10'h46 == _T_28[9:0]) begin
        image_0_70 <= io_pixelVal_in_0_4;
      end else if (10'h46 == _T_25[9:0]) begin
        image_0_70 <= io_pixelVal_in_0_3;
      end else if (10'h46 == _T_22[9:0]) begin
        image_0_70 <= io_pixelVal_in_0_2;
      end else if (10'h46 == _T_19[9:0]) begin
        image_0_70 <= io_pixelVal_in_0_1;
      end else if (10'h46 == _T_15[9:0]) begin
        image_0_70 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_71 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h47 == _T_37[9:0]) begin
        image_0_71 <= io_pixelVal_in_0_7;
      end else if (10'h47 == _T_34[9:0]) begin
        image_0_71 <= io_pixelVal_in_0_6;
      end else if (10'h47 == _T_31[9:0]) begin
        image_0_71 <= io_pixelVal_in_0_5;
      end else if (10'h47 == _T_28[9:0]) begin
        image_0_71 <= io_pixelVal_in_0_4;
      end else if (10'h47 == _T_25[9:0]) begin
        image_0_71 <= io_pixelVal_in_0_3;
      end else if (10'h47 == _T_22[9:0]) begin
        image_0_71 <= io_pixelVal_in_0_2;
      end else if (10'h47 == _T_19[9:0]) begin
        image_0_71 <= io_pixelVal_in_0_1;
      end else if (10'h47 == _T_15[9:0]) begin
        image_0_71 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_72 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h48 == _T_37[9:0]) begin
        image_0_72 <= io_pixelVal_in_0_7;
      end else if (10'h48 == _T_34[9:0]) begin
        image_0_72 <= io_pixelVal_in_0_6;
      end else if (10'h48 == _T_31[9:0]) begin
        image_0_72 <= io_pixelVal_in_0_5;
      end else if (10'h48 == _T_28[9:0]) begin
        image_0_72 <= io_pixelVal_in_0_4;
      end else if (10'h48 == _T_25[9:0]) begin
        image_0_72 <= io_pixelVal_in_0_3;
      end else if (10'h48 == _T_22[9:0]) begin
        image_0_72 <= io_pixelVal_in_0_2;
      end else if (10'h48 == _T_19[9:0]) begin
        image_0_72 <= io_pixelVal_in_0_1;
      end else if (10'h48 == _T_15[9:0]) begin
        image_0_72 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_73 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h49 == _T_37[9:0]) begin
        image_0_73 <= io_pixelVal_in_0_7;
      end else if (10'h49 == _T_34[9:0]) begin
        image_0_73 <= io_pixelVal_in_0_6;
      end else if (10'h49 == _T_31[9:0]) begin
        image_0_73 <= io_pixelVal_in_0_5;
      end else if (10'h49 == _T_28[9:0]) begin
        image_0_73 <= io_pixelVal_in_0_4;
      end else if (10'h49 == _T_25[9:0]) begin
        image_0_73 <= io_pixelVal_in_0_3;
      end else if (10'h49 == _T_22[9:0]) begin
        image_0_73 <= io_pixelVal_in_0_2;
      end else if (10'h49 == _T_19[9:0]) begin
        image_0_73 <= io_pixelVal_in_0_1;
      end else if (10'h49 == _T_15[9:0]) begin
        image_0_73 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_74 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h4a == _T_37[9:0]) begin
        image_0_74 <= io_pixelVal_in_0_7;
      end else if (10'h4a == _T_34[9:0]) begin
        image_0_74 <= io_pixelVal_in_0_6;
      end else if (10'h4a == _T_31[9:0]) begin
        image_0_74 <= io_pixelVal_in_0_5;
      end else if (10'h4a == _T_28[9:0]) begin
        image_0_74 <= io_pixelVal_in_0_4;
      end else if (10'h4a == _T_25[9:0]) begin
        image_0_74 <= io_pixelVal_in_0_3;
      end else if (10'h4a == _T_22[9:0]) begin
        image_0_74 <= io_pixelVal_in_0_2;
      end else if (10'h4a == _T_19[9:0]) begin
        image_0_74 <= io_pixelVal_in_0_1;
      end else if (10'h4a == _T_15[9:0]) begin
        image_0_74 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_75 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h4b == _T_37[9:0]) begin
        image_0_75 <= io_pixelVal_in_0_7;
      end else if (10'h4b == _T_34[9:0]) begin
        image_0_75 <= io_pixelVal_in_0_6;
      end else if (10'h4b == _T_31[9:0]) begin
        image_0_75 <= io_pixelVal_in_0_5;
      end else if (10'h4b == _T_28[9:0]) begin
        image_0_75 <= io_pixelVal_in_0_4;
      end else if (10'h4b == _T_25[9:0]) begin
        image_0_75 <= io_pixelVal_in_0_3;
      end else if (10'h4b == _T_22[9:0]) begin
        image_0_75 <= io_pixelVal_in_0_2;
      end else if (10'h4b == _T_19[9:0]) begin
        image_0_75 <= io_pixelVal_in_0_1;
      end else if (10'h4b == _T_15[9:0]) begin
        image_0_75 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_76 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h4c == _T_37[9:0]) begin
        image_0_76 <= io_pixelVal_in_0_7;
      end else if (10'h4c == _T_34[9:0]) begin
        image_0_76 <= io_pixelVal_in_0_6;
      end else if (10'h4c == _T_31[9:0]) begin
        image_0_76 <= io_pixelVal_in_0_5;
      end else if (10'h4c == _T_28[9:0]) begin
        image_0_76 <= io_pixelVal_in_0_4;
      end else if (10'h4c == _T_25[9:0]) begin
        image_0_76 <= io_pixelVal_in_0_3;
      end else if (10'h4c == _T_22[9:0]) begin
        image_0_76 <= io_pixelVal_in_0_2;
      end else if (10'h4c == _T_19[9:0]) begin
        image_0_76 <= io_pixelVal_in_0_1;
      end else if (10'h4c == _T_15[9:0]) begin
        image_0_76 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_77 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h4d == _T_37[9:0]) begin
        image_0_77 <= io_pixelVal_in_0_7;
      end else if (10'h4d == _T_34[9:0]) begin
        image_0_77 <= io_pixelVal_in_0_6;
      end else if (10'h4d == _T_31[9:0]) begin
        image_0_77 <= io_pixelVal_in_0_5;
      end else if (10'h4d == _T_28[9:0]) begin
        image_0_77 <= io_pixelVal_in_0_4;
      end else if (10'h4d == _T_25[9:0]) begin
        image_0_77 <= io_pixelVal_in_0_3;
      end else if (10'h4d == _T_22[9:0]) begin
        image_0_77 <= io_pixelVal_in_0_2;
      end else if (10'h4d == _T_19[9:0]) begin
        image_0_77 <= io_pixelVal_in_0_1;
      end else if (10'h4d == _T_15[9:0]) begin
        image_0_77 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_78 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h4e == _T_37[9:0]) begin
        image_0_78 <= io_pixelVal_in_0_7;
      end else if (10'h4e == _T_34[9:0]) begin
        image_0_78 <= io_pixelVal_in_0_6;
      end else if (10'h4e == _T_31[9:0]) begin
        image_0_78 <= io_pixelVal_in_0_5;
      end else if (10'h4e == _T_28[9:0]) begin
        image_0_78 <= io_pixelVal_in_0_4;
      end else if (10'h4e == _T_25[9:0]) begin
        image_0_78 <= io_pixelVal_in_0_3;
      end else if (10'h4e == _T_22[9:0]) begin
        image_0_78 <= io_pixelVal_in_0_2;
      end else if (10'h4e == _T_19[9:0]) begin
        image_0_78 <= io_pixelVal_in_0_1;
      end else if (10'h4e == _T_15[9:0]) begin
        image_0_78 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_79 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h4f == _T_37[9:0]) begin
        image_0_79 <= io_pixelVal_in_0_7;
      end else if (10'h4f == _T_34[9:0]) begin
        image_0_79 <= io_pixelVal_in_0_6;
      end else if (10'h4f == _T_31[9:0]) begin
        image_0_79 <= io_pixelVal_in_0_5;
      end else if (10'h4f == _T_28[9:0]) begin
        image_0_79 <= io_pixelVal_in_0_4;
      end else if (10'h4f == _T_25[9:0]) begin
        image_0_79 <= io_pixelVal_in_0_3;
      end else if (10'h4f == _T_22[9:0]) begin
        image_0_79 <= io_pixelVal_in_0_2;
      end else if (10'h4f == _T_19[9:0]) begin
        image_0_79 <= io_pixelVal_in_0_1;
      end else if (10'h4f == _T_15[9:0]) begin
        image_0_79 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_80 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h50 == _T_37[9:0]) begin
        image_0_80 <= io_pixelVal_in_0_7;
      end else if (10'h50 == _T_34[9:0]) begin
        image_0_80 <= io_pixelVal_in_0_6;
      end else if (10'h50 == _T_31[9:0]) begin
        image_0_80 <= io_pixelVal_in_0_5;
      end else if (10'h50 == _T_28[9:0]) begin
        image_0_80 <= io_pixelVal_in_0_4;
      end else if (10'h50 == _T_25[9:0]) begin
        image_0_80 <= io_pixelVal_in_0_3;
      end else if (10'h50 == _T_22[9:0]) begin
        image_0_80 <= io_pixelVal_in_0_2;
      end else if (10'h50 == _T_19[9:0]) begin
        image_0_80 <= io_pixelVal_in_0_1;
      end else if (10'h50 == _T_15[9:0]) begin
        image_0_80 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_81 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h51 == _T_37[9:0]) begin
        image_0_81 <= io_pixelVal_in_0_7;
      end else if (10'h51 == _T_34[9:0]) begin
        image_0_81 <= io_pixelVal_in_0_6;
      end else if (10'h51 == _T_31[9:0]) begin
        image_0_81 <= io_pixelVal_in_0_5;
      end else if (10'h51 == _T_28[9:0]) begin
        image_0_81 <= io_pixelVal_in_0_4;
      end else if (10'h51 == _T_25[9:0]) begin
        image_0_81 <= io_pixelVal_in_0_3;
      end else if (10'h51 == _T_22[9:0]) begin
        image_0_81 <= io_pixelVal_in_0_2;
      end else if (10'h51 == _T_19[9:0]) begin
        image_0_81 <= io_pixelVal_in_0_1;
      end else if (10'h51 == _T_15[9:0]) begin
        image_0_81 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_82 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h52 == _T_37[9:0]) begin
        image_0_82 <= io_pixelVal_in_0_7;
      end else if (10'h52 == _T_34[9:0]) begin
        image_0_82 <= io_pixelVal_in_0_6;
      end else if (10'h52 == _T_31[9:0]) begin
        image_0_82 <= io_pixelVal_in_0_5;
      end else if (10'h52 == _T_28[9:0]) begin
        image_0_82 <= io_pixelVal_in_0_4;
      end else if (10'h52 == _T_25[9:0]) begin
        image_0_82 <= io_pixelVal_in_0_3;
      end else if (10'h52 == _T_22[9:0]) begin
        image_0_82 <= io_pixelVal_in_0_2;
      end else if (10'h52 == _T_19[9:0]) begin
        image_0_82 <= io_pixelVal_in_0_1;
      end else if (10'h52 == _T_15[9:0]) begin
        image_0_82 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_83 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h53 == _T_37[9:0]) begin
        image_0_83 <= io_pixelVal_in_0_7;
      end else if (10'h53 == _T_34[9:0]) begin
        image_0_83 <= io_pixelVal_in_0_6;
      end else if (10'h53 == _T_31[9:0]) begin
        image_0_83 <= io_pixelVal_in_0_5;
      end else if (10'h53 == _T_28[9:0]) begin
        image_0_83 <= io_pixelVal_in_0_4;
      end else if (10'h53 == _T_25[9:0]) begin
        image_0_83 <= io_pixelVal_in_0_3;
      end else if (10'h53 == _T_22[9:0]) begin
        image_0_83 <= io_pixelVal_in_0_2;
      end else if (10'h53 == _T_19[9:0]) begin
        image_0_83 <= io_pixelVal_in_0_1;
      end else if (10'h53 == _T_15[9:0]) begin
        image_0_83 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_84 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h54 == _T_37[9:0]) begin
        image_0_84 <= io_pixelVal_in_0_7;
      end else if (10'h54 == _T_34[9:0]) begin
        image_0_84 <= io_pixelVal_in_0_6;
      end else if (10'h54 == _T_31[9:0]) begin
        image_0_84 <= io_pixelVal_in_0_5;
      end else if (10'h54 == _T_28[9:0]) begin
        image_0_84 <= io_pixelVal_in_0_4;
      end else if (10'h54 == _T_25[9:0]) begin
        image_0_84 <= io_pixelVal_in_0_3;
      end else if (10'h54 == _T_22[9:0]) begin
        image_0_84 <= io_pixelVal_in_0_2;
      end else if (10'h54 == _T_19[9:0]) begin
        image_0_84 <= io_pixelVal_in_0_1;
      end else if (10'h54 == _T_15[9:0]) begin
        image_0_84 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_85 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h55 == _T_37[9:0]) begin
        image_0_85 <= io_pixelVal_in_0_7;
      end else if (10'h55 == _T_34[9:0]) begin
        image_0_85 <= io_pixelVal_in_0_6;
      end else if (10'h55 == _T_31[9:0]) begin
        image_0_85 <= io_pixelVal_in_0_5;
      end else if (10'h55 == _T_28[9:0]) begin
        image_0_85 <= io_pixelVal_in_0_4;
      end else if (10'h55 == _T_25[9:0]) begin
        image_0_85 <= io_pixelVal_in_0_3;
      end else if (10'h55 == _T_22[9:0]) begin
        image_0_85 <= io_pixelVal_in_0_2;
      end else if (10'h55 == _T_19[9:0]) begin
        image_0_85 <= io_pixelVal_in_0_1;
      end else if (10'h55 == _T_15[9:0]) begin
        image_0_85 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_86 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h56 == _T_37[9:0]) begin
        image_0_86 <= io_pixelVal_in_0_7;
      end else if (10'h56 == _T_34[9:0]) begin
        image_0_86 <= io_pixelVal_in_0_6;
      end else if (10'h56 == _T_31[9:0]) begin
        image_0_86 <= io_pixelVal_in_0_5;
      end else if (10'h56 == _T_28[9:0]) begin
        image_0_86 <= io_pixelVal_in_0_4;
      end else if (10'h56 == _T_25[9:0]) begin
        image_0_86 <= io_pixelVal_in_0_3;
      end else if (10'h56 == _T_22[9:0]) begin
        image_0_86 <= io_pixelVal_in_0_2;
      end else if (10'h56 == _T_19[9:0]) begin
        image_0_86 <= io_pixelVal_in_0_1;
      end else if (10'h56 == _T_15[9:0]) begin
        image_0_86 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_87 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h57 == _T_37[9:0]) begin
        image_0_87 <= io_pixelVal_in_0_7;
      end else if (10'h57 == _T_34[9:0]) begin
        image_0_87 <= io_pixelVal_in_0_6;
      end else if (10'h57 == _T_31[9:0]) begin
        image_0_87 <= io_pixelVal_in_0_5;
      end else if (10'h57 == _T_28[9:0]) begin
        image_0_87 <= io_pixelVal_in_0_4;
      end else if (10'h57 == _T_25[9:0]) begin
        image_0_87 <= io_pixelVal_in_0_3;
      end else if (10'h57 == _T_22[9:0]) begin
        image_0_87 <= io_pixelVal_in_0_2;
      end else if (10'h57 == _T_19[9:0]) begin
        image_0_87 <= io_pixelVal_in_0_1;
      end else if (10'h57 == _T_15[9:0]) begin
        image_0_87 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_88 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h58 == _T_37[9:0]) begin
        image_0_88 <= io_pixelVal_in_0_7;
      end else if (10'h58 == _T_34[9:0]) begin
        image_0_88 <= io_pixelVal_in_0_6;
      end else if (10'h58 == _T_31[9:0]) begin
        image_0_88 <= io_pixelVal_in_0_5;
      end else if (10'h58 == _T_28[9:0]) begin
        image_0_88 <= io_pixelVal_in_0_4;
      end else if (10'h58 == _T_25[9:0]) begin
        image_0_88 <= io_pixelVal_in_0_3;
      end else if (10'h58 == _T_22[9:0]) begin
        image_0_88 <= io_pixelVal_in_0_2;
      end else if (10'h58 == _T_19[9:0]) begin
        image_0_88 <= io_pixelVal_in_0_1;
      end else if (10'h58 == _T_15[9:0]) begin
        image_0_88 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_89 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h59 == _T_37[9:0]) begin
        image_0_89 <= io_pixelVal_in_0_7;
      end else if (10'h59 == _T_34[9:0]) begin
        image_0_89 <= io_pixelVal_in_0_6;
      end else if (10'h59 == _T_31[9:0]) begin
        image_0_89 <= io_pixelVal_in_0_5;
      end else if (10'h59 == _T_28[9:0]) begin
        image_0_89 <= io_pixelVal_in_0_4;
      end else if (10'h59 == _T_25[9:0]) begin
        image_0_89 <= io_pixelVal_in_0_3;
      end else if (10'h59 == _T_22[9:0]) begin
        image_0_89 <= io_pixelVal_in_0_2;
      end else if (10'h59 == _T_19[9:0]) begin
        image_0_89 <= io_pixelVal_in_0_1;
      end else if (10'h59 == _T_15[9:0]) begin
        image_0_89 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_90 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h5a == _T_37[9:0]) begin
        image_0_90 <= io_pixelVal_in_0_7;
      end else if (10'h5a == _T_34[9:0]) begin
        image_0_90 <= io_pixelVal_in_0_6;
      end else if (10'h5a == _T_31[9:0]) begin
        image_0_90 <= io_pixelVal_in_0_5;
      end else if (10'h5a == _T_28[9:0]) begin
        image_0_90 <= io_pixelVal_in_0_4;
      end else if (10'h5a == _T_25[9:0]) begin
        image_0_90 <= io_pixelVal_in_0_3;
      end else if (10'h5a == _T_22[9:0]) begin
        image_0_90 <= io_pixelVal_in_0_2;
      end else if (10'h5a == _T_19[9:0]) begin
        image_0_90 <= io_pixelVal_in_0_1;
      end else if (10'h5a == _T_15[9:0]) begin
        image_0_90 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_91 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h5b == _T_37[9:0]) begin
        image_0_91 <= io_pixelVal_in_0_7;
      end else if (10'h5b == _T_34[9:0]) begin
        image_0_91 <= io_pixelVal_in_0_6;
      end else if (10'h5b == _T_31[9:0]) begin
        image_0_91 <= io_pixelVal_in_0_5;
      end else if (10'h5b == _T_28[9:0]) begin
        image_0_91 <= io_pixelVal_in_0_4;
      end else if (10'h5b == _T_25[9:0]) begin
        image_0_91 <= io_pixelVal_in_0_3;
      end else if (10'h5b == _T_22[9:0]) begin
        image_0_91 <= io_pixelVal_in_0_2;
      end else if (10'h5b == _T_19[9:0]) begin
        image_0_91 <= io_pixelVal_in_0_1;
      end else if (10'h5b == _T_15[9:0]) begin
        image_0_91 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_92 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h5c == _T_37[9:0]) begin
        image_0_92 <= io_pixelVal_in_0_7;
      end else if (10'h5c == _T_34[9:0]) begin
        image_0_92 <= io_pixelVal_in_0_6;
      end else if (10'h5c == _T_31[9:0]) begin
        image_0_92 <= io_pixelVal_in_0_5;
      end else if (10'h5c == _T_28[9:0]) begin
        image_0_92 <= io_pixelVal_in_0_4;
      end else if (10'h5c == _T_25[9:0]) begin
        image_0_92 <= io_pixelVal_in_0_3;
      end else if (10'h5c == _T_22[9:0]) begin
        image_0_92 <= io_pixelVal_in_0_2;
      end else if (10'h5c == _T_19[9:0]) begin
        image_0_92 <= io_pixelVal_in_0_1;
      end else if (10'h5c == _T_15[9:0]) begin
        image_0_92 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_93 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h5d == _T_37[9:0]) begin
        image_0_93 <= io_pixelVal_in_0_7;
      end else if (10'h5d == _T_34[9:0]) begin
        image_0_93 <= io_pixelVal_in_0_6;
      end else if (10'h5d == _T_31[9:0]) begin
        image_0_93 <= io_pixelVal_in_0_5;
      end else if (10'h5d == _T_28[9:0]) begin
        image_0_93 <= io_pixelVal_in_0_4;
      end else if (10'h5d == _T_25[9:0]) begin
        image_0_93 <= io_pixelVal_in_0_3;
      end else if (10'h5d == _T_22[9:0]) begin
        image_0_93 <= io_pixelVal_in_0_2;
      end else if (10'h5d == _T_19[9:0]) begin
        image_0_93 <= io_pixelVal_in_0_1;
      end else if (10'h5d == _T_15[9:0]) begin
        image_0_93 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_94 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h5e == _T_37[9:0]) begin
        image_0_94 <= io_pixelVal_in_0_7;
      end else if (10'h5e == _T_34[9:0]) begin
        image_0_94 <= io_pixelVal_in_0_6;
      end else if (10'h5e == _T_31[9:0]) begin
        image_0_94 <= io_pixelVal_in_0_5;
      end else if (10'h5e == _T_28[9:0]) begin
        image_0_94 <= io_pixelVal_in_0_4;
      end else if (10'h5e == _T_25[9:0]) begin
        image_0_94 <= io_pixelVal_in_0_3;
      end else if (10'h5e == _T_22[9:0]) begin
        image_0_94 <= io_pixelVal_in_0_2;
      end else if (10'h5e == _T_19[9:0]) begin
        image_0_94 <= io_pixelVal_in_0_1;
      end else if (10'h5e == _T_15[9:0]) begin
        image_0_94 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_95 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h5f == _T_37[9:0]) begin
        image_0_95 <= io_pixelVal_in_0_7;
      end else if (10'h5f == _T_34[9:0]) begin
        image_0_95 <= io_pixelVal_in_0_6;
      end else if (10'h5f == _T_31[9:0]) begin
        image_0_95 <= io_pixelVal_in_0_5;
      end else if (10'h5f == _T_28[9:0]) begin
        image_0_95 <= io_pixelVal_in_0_4;
      end else if (10'h5f == _T_25[9:0]) begin
        image_0_95 <= io_pixelVal_in_0_3;
      end else if (10'h5f == _T_22[9:0]) begin
        image_0_95 <= io_pixelVal_in_0_2;
      end else if (10'h5f == _T_19[9:0]) begin
        image_0_95 <= io_pixelVal_in_0_1;
      end else if (10'h5f == _T_15[9:0]) begin
        image_0_95 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_96 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h60 == _T_37[9:0]) begin
        image_0_96 <= io_pixelVal_in_0_7;
      end else if (10'h60 == _T_34[9:0]) begin
        image_0_96 <= io_pixelVal_in_0_6;
      end else if (10'h60 == _T_31[9:0]) begin
        image_0_96 <= io_pixelVal_in_0_5;
      end else if (10'h60 == _T_28[9:0]) begin
        image_0_96 <= io_pixelVal_in_0_4;
      end else if (10'h60 == _T_25[9:0]) begin
        image_0_96 <= io_pixelVal_in_0_3;
      end else if (10'h60 == _T_22[9:0]) begin
        image_0_96 <= io_pixelVal_in_0_2;
      end else if (10'h60 == _T_19[9:0]) begin
        image_0_96 <= io_pixelVal_in_0_1;
      end else if (10'h60 == _T_15[9:0]) begin
        image_0_96 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_97 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h61 == _T_37[9:0]) begin
        image_0_97 <= io_pixelVal_in_0_7;
      end else if (10'h61 == _T_34[9:0]) begin
        image_0_97 <= io_pixelVal_in_0_6;
      end else if (10'h61 == _T_31[9:0]) begin
        image_0_97 <= io_pixelVal_in_0_5;
      end else if (10'h61 == _T_28[9:0]) begin
        image_0_97 <= io_pixelVal_in_0_4;
      end else if (10'h61 == _T_25[9:0]) begin
        image_0_97 <= io_pixelVal_in_0_3;
      end else if (10'h61 == _T_22[9:0]) begin
        image_0_97 <= io_pixelVal_in_0_2;
      end else if (10'h61 == _T_19[9:0]) begin
        image_0_97 <= io_pixelVal_in_0_1;
      end else if (10'h61 == _T_15[9:0]) begin
        image_0_97 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_98 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h62 == _T_37[9:0]) begin
        image_0_98 <= io_pixelVal_in_0_7;
      end else if (10'h62 == _T_34[9:0]) begin
        image_0_98 <= io_pixelVal_in_0_6;
      end else if (10'h62 == _T_31[9:0]) begin
        image_0_98 <= io_pixelVal_in_0_5;
      end else if (10'h62 == _T_28[9:0]) begin
        image_0_98 <= io_pixelVal_in_0_4;
      end else if (10'h62 == _T_25[9:0]) begin
        image_0_98 <= io_pixelVal_in_0_3;
      end else if (10'h62 == _T_22[9:0]) begin
        image_0_98 <= io_pixelVal_in_0_2;
      end else if (10'h62 == _T_19[9:0]) begin
        image_0_98 <= io_pixelVal_in_0_1;
      end else if (10'h62 == _T_15[9:0]) begin
        image_0_98 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_99 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h63 == _T_37[9:0]) begin
        image_0_99 <= io_pixelVal_in_0_7;
      end else if (10'h63 == _T_34[9:0]) begin
        image_0_99 <= io_pixelVal_in_0_6;
      end else if (10'h63 == _T_31[9:0]) begin
        image_0_99 <= io_pixelVal_in_0_5;
      end else if (10'h63 == _T_28[9:0]) begin
        image_0_99 <= io_pixelVal_in_0_4;
      end else if (10'h63 == _T_25[9:0]) begin
        image_0_99 <= io_pixelVal_in_0_3;
      end else if (10'h63 == _T_22[9:0]) begin
        image_0_99 <= io_pixelVal_in_0_2;
      end else if (10'h63 == _T_19[9:0]) begin
        image_0_99 <= io_pixelVal_in_0_1;
      end else if (10'h63 == _T_15[9:0]) begin
        image_0_99 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_100 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h64 == _T_37[9:0]) begin
        image_0_100 <= io_pixelVal_in_0_7;
      end else if (10'h64 == _T_34[9:0]) begin
        image_0_100 <= io_pixelVal_in_0_6;
      end else if (10'h64 == _T_31[9:0]) begin
        image_0_100 <= io_pixelVal_in_0_5;
      end else if (10'h64 == _T_28[9:0]) begin
        image_0_100 <= io_pixelVal_in_0_4;
      end else if (10'h64 == _T_25[9:0]) begin
        image_0_100 <= io_pixelVal_in_0_3;
      end else if (10'h64 == _T_22[9:0]) begin
        image_0_100 <= io_pixelVal_in_0_2;
      end else if (10'h64 == _T_19[9:0]) begin
        image_0_100 <= io_pixelVal_in_0_1;
      end else if (10'h64 == _T_15[9:0]) begin
        image_0_100 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_101 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h65 == _T_37[9:0]) begin
        image_0_101 <= io_pixelVal_in_0_7;
      end else if (10'h65 == _T_34[9:0]) begin
        image_0_101 <= io_pixelVal_in_0_6;
      end else if (10'h65 == _T_31[9:0]) begin
        image_0_101 <= io_pixelVal_in_0_5;
      end else if (10'h65 == _T_28[9:0]) begin
        image_0_101 <= io_pixelVal_in_0_4;
      end else if (10'h65 == _T_25[9:0]) begin
        image_0_101 <= io_pixelVal_in_0_3;
      end else if (10'h65 == _T_22[9:0]) begin
        image_0_101 <= io_pixelVal_in_0_2;
      end else if (10'h65 == _T_19[9:0]) begin
        image_0_101 <= io_pixelVal_in_0_1;
      end else if (10'h65 == _T_15[9:0]) begin
        image_0_101 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_102 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h66 == _T_37[9:0]) begin
        image_0_102 <= io_pixelVal_in_0_7;
      end else if (10'h66 == _T_34[9:0]) begin
        image_0_102 <= io_pixelVal_in_0_6;
      end else if (10'h66 == _T_31[9:0]) begin
        image_0_102 <= io_pixelVal_in_0_5;
      end else if (10'h66 == _T_28[9:0]) begin
        image_0_102 <= io_pixelVal_in_0_4;
      end else if (10'h66 == _T_25[9:0]) begin
        image_0_102 <= io_pixelVal_in_0_3;
      end else if (10'h66 == _T_22[9:0]) begin
        image_0_102 <= io_pixelVal_in_0_2;
      end else if (10'h66 == _T_19[9:0]) begin
        image_0_102 <= io_pixelVal_in_0_1;
      end else if (10'h66 == _T_15[9:0]) begin
        image_0_102 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_103 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h67 == _T_37[9:0]) begin
        image_0_103 <= io_pixelVal_in_0_7;
      end else if (10'h67 == _T_34[9:0]) begin
        image_0_103 <= io_pixelVal_in_0_6;
      end else if (10'h67 == _T_31[9:0]) begin
        image_0_103 <= io_pixelVal_in_0_5;
      end else if (10'h67 == _T_28[9:0]) begin
        image_0_103 <= io_pixelVal_in_0_4;
      end else if (10'h67 == _T_25[9:0]) begin
        image_0_103 <= io_pixelVal_in_0_3;
      end else if (10'h67 == _T_22[9:0]) begin
        image_0_103 <= io_pixelVal_in_0_2;
      end else if (10'h67 == _T_19[9:0]) begin
        image_0_103 <= io_pixelVal_in_0_1;
      end else if (10'h67 == _T_15[9:0]) begin
        image_0_103 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_104 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h68 == _T_37[9:0]) begin
        image_0_104 <= io_pixelVal_in_0_7;
      end else if (10'h68 == _T_34[9:0]) begin
        image_0_104 <= io_pixelVal_in_0_6;
      end else if (10'h68 == _T_31[9:0]) begin
        image_0_104 <= io_pixelVal_in_0_5;
      end else if (10'h68 == _T_28[9:0]) begin
        image_0_104 <= io_pixelVal_in_0_4;
      end else if (10'h68 == _T_25[9:0]) begin
        image_0_104 <= io_pixelVal_in_0_3;
      end else if (10'h68 == _T_22[9:0]) begin
        image_0_104 <= io_pixelVal_in_0_2;
      end else if (10'h68 == _T_19[9:0]) begin
        image_0_104 <= io_pixelVal_in_0_1;
      end else if (10'h68 == _T_15[9:0]) begin
        image_0_104 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_105 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h69 == _T_37[9:0]) begin
        image_0_105 <= io_pixelVal_in_0_7;
      end else if (10'h69 == _T_34[9:0]) begin
        image_0_105 <= io_pixelVal_in_0_6;
      end else if (10'h69 == _T_31[9:0]) begin
        image_0_105 <= io_pixelVal_in_0_5;
      end else if (10'h69 == _T_28[9:0]) begin
        image_0_105 <= io_pixelVal_in_0_4;
      end else if (10'h69 == _T_25[9:0]) begin
        image_0_105 <= io_pixelVal_in_0_3;
      end else if (10'h69 == _T_22[9:0]) begin
        image_0_105 <= io_pixelVal_in_0_2;
      end else if (10'h69 == _T_19[9:0]) begin
        image_0_105 <= io_pixelVal_in_0_1;
      end else if (10'h69 == _T_15[9:0]) begin
        image_0_105 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_106 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h6a == _T_37[9:0]) begin
        image_0_106 <= io_pixelVal_in_0_7;
      end else if (10'h6a == _T_34[9:0]) begin
        image_0_106 <= io_pixelVal_in_0_6;
      end else if (10'h6a == _T_31[9:0]) begin
        image_0_106 <= io_pixelVal_in_0_5;
      end else if (10'h6a == _T_28[9:0]) begin
        image_0_106 <= io_pixelVal_in_0_4;
      end else if (10'h6a == _T_25[9:0]) begin
        image_0_106 <= io_pixelVal_in_0_3;
      end else if (10'h6a == _T_22[9:0]) begin
        image_0_106 <= io_pixelVal_in_0_2;
      end else if (10'h6a == _T_19[9:0]) begin
        image_0_106 <= io_pixelVal_in_0_1;
      end else if (10'h6a == _T_15[9:0]) begin
        image_0_106 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_107 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h6b == _T_37[9:0]) begin
        image_0_107 <= io_pixelVal_in_0_7;
      end else if (10'h6b == _T_34[9:0]) begin
        image_0_107 <= io_pixelVal_in_0_6;
      end else if (10'h6b == _T_31[9:0]) begin
        image_0_107 <= io_pixelVal_in_0_5;
      end else if (10'h6b == _T_28[9:0]) begin
        image_0_107 <= io_pixelVal_in_0_4;
      end else if (10'h6b == _T_25[9:0]) begin
        image_0_107 <= io_pixelVal_in_0_3;
      end else if (10'h6b == _T_22[9:0]) begin
        image_0_107 <= io_pixelVal_in_0_2;
      end else if (10'h6b == _T_19[9:0]) begin
        image_0_107 <= io_pixelVal_in_0_1;
      end else if (10'h6b == _T_15[9:0]) begin
        image_0_107 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_108 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h6c == _T_37[9:0]) begin
        image_0_108 <= io_pixelVal_in_0_7;
      end else if (10'h6c == _T_34[9:0]) begin
        image_0_108 <= io_pixelVal_in_0_6;
      end else if (10'h6c == _T_31[9:0]) begin
        image_0_108 <= io_pixelVal_in_0_5;
      end else if (10'h6c == _T_28[9:0]) begin
        image_0_108 <= io_pixelVal_in_0_4;
      end else if (10'h6c == _T_25[9:0]) begin
        image_0_108 <= io_pixelVal_in_0_3;
      end else if (10'h6c == _T_22[9:0]) begin
        image_0_108 <= io_pixelVal_in_0_2;
      end else if (10'h6c == _T_19[9:0]) begin
        image_0_108 <= io_pixelVal_in_0_1;
      end else if (10'h6c == _T_15[9:0]) begin
        image_0_108 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_109 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h6d == _T_37[9:0]) begin
        image_0_109 <= io_pixelVal_in_0_7;
      end else if (10'h6d == _T_34[9:0]) begin
        image_0_109 <= io_pixelVal_in_0_6;
      end else if (10'h6d == _T_31[9:0]) begin
        image_0_109 <= io_pixelVal_in_0_5;
      end else if (10'h6d == _T_28[9:0]) begin
        image_0_109 <= io_pixelVal_in_0_4;
      end else if (10'h6d == _T_25[9:0]) begin
        image_0_109 <= io_pixelVal_in_0_3;
      end else if (10'h6d == _T_22[9:0]) begin
        image_0_109 <= io_pixelVal_in_0_2;
      end else if (10'h6d == _T_19[9:0]) begin
        image_0_109 <= io_pixelVal_in_0_1;
      end else if (10'h6d == _T_15[9:0]) begin
        image_0_109 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_110 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h6e == _T_37[9:0]) begin
        image_0_110 <= io_pixelVal_in_0_7;
      end else if (10'h6e == _T_34[9:0]) begin
        image_0_110 <= io_pixelVal_in_0_6;
      end else if (10'h6e == _T_31[9:0]) begin
        image_0_110 <= io_pixelVal_in_0_5;
      end else if (10'h6e == _T_28[9:0]) begin
        image_0_110 <= io_pixelVal_in_0_4;
      end else if (10'h6e == _T_25[9:0]) begin
        image_0_110 <= io_pixelVal_in_0_3;
      end else if (10'h6e == _T_22[9:0]) begin
        image_0_110 <= io_pixelVal_in_0_2;
      end else if (10'h6e == _T_19[9:0]) begin
        image_0_110 <= io_pixelVal_in_0_1;
      end else if (10'h6e == _T_15[9:0]) begin
        image_0_110 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_111 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h6f == _T_37[9:0]) begin
        image_0_111 <= io_pixelVal_in_0_7;
      end else if (10'h6f == _T_34[9:0]) begin
        image_0_111 <= io_pixelVal_in_0_6;
      end else if (10'h6f == _T_31[9:0]) begin
        image_0_111 <= io_pixelVal_in_0_5;
      end else if (10'h6f == _T_28[9:0]) begin
        image_0_111 <= io_pixelVal_in_0_4;
      end else if (10'h6f == _T_25[9:0]) begin
        image_0_111 <= io_pixelVal_in_0_3;
      end else if (10'h6f == _T_22[9:0]) begin
        image_0_111 <= io_pixelVal_in_0_2;
      end else if (10'h6f == _T_19[9:0]) begin
        image_0_111 <= io_pixelVal_in_0_1;
      end else if (10'h6f == _T_15[9:0]) begin
        image_0_111 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_112 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h70 == _T_37[9:0]) begin
        image_0_112 <= io_pixelVal_in_0_7;
      end else if (10'h70 == _T_34[9:0]) begin
        image_0_112 <= io_pixelVal_in_0_6;
      end else if (10'h70 == _T_31[9:0]) begin
        image_0_112 <= io_pixelVal_in_0_5;
      end else if (10'h70 == _T_28[9:0]) begin
        image_0_112 <= io_pixelVal_in_0_4;
      end else if (10'h70 == _T_25[9:0]) begin
        image_0_112 <= io_pixelVal_in_0_3;
      end else if (10'h70 == _T_22[9:0]) begin
        image_0_112 <= io_pixelVal_in_0_2;
      end else if (10'h70 == _T_19[9:0]) begin
        image_0_112 <= io_pixelVal_in_0_1;
      end else if (10'h70 == _T_15[9:0]) begin
        image_0_112 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_113 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h71 == _T_37[9:0]) begin
        image_0_113 <= io_pixelVal_in_0_7;
      end else if (10'h71 == _T_34[9:0]) begin
        image_0_113 <= io_pixelVal_in_0_6;
      end else if (10'h71 == _T_31[9:0]) begin
        image_0_113 <= io_pixelVal_in_0_5;
      end else if (10'h71 == _T_28[9:0]) begin
        image_0_113 <= io_pixelVal_in_0_4;
      end else if (10'h71 == _T_25[9:0]) begin
        image_0_113 <= io_pixelVal_in_0_3;
      end else if (10'h71 == _T_22[9:0]) begin
        image_0_113 <= io_pixelVal_in_0_2;
      end else if (10'h71 == _T_19[9:0]) begin
        image_0_113 <= io_pixelVal_in_0_1;
      end else if (10'h71 == _T_15[9:0]) begin
        image_0_113 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_114 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h72 == _T_37[9:0]) begin
        image_0_114 <= io_pixelVal_in_0_7;
      end else if (10'h72 == _T_34[9:0]) begin
        image_0_114 <= io_pixelVal_in_0_6;
      end else if (10'h72 == _T_31[9:0]) begin
        image_0_114 <= io_pixelVal_in_0_5;
      end else if (10'h72 == _T_28[9:0]) begin
        image_0_114 <= io_pixelVal_in_0_4;
      end else if (10'h72 == _T_25[9:0]) begin
        image_0_114 <= io_pixelVal_in_0_3;
      end else if (10'h72 == _T_22[9:0]) begin
        image_0_114 <= io_pixelVal_in_0_2;
      end else if (10'h72 == _T_19[9:0]) begin
        image_0_114 <= io_pixelVal_in_0_1;
      end else if (10'h72 == _T_15[9:0]) begin
        image_0_114 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_115 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h73 == _T_37[9:0]) begin
        image_0_115 <= io_pixelVal_in_0_7;
      end else if (10'h73 == _T_34[9:0]) begin
        image_0_115 <= io_pixelVal_in_0_6;
      end else if (10'h73 == _T_31[9:0]) begin
        image_0_115 <= io_pixelVal_in_0_5;
      end else if (10'h73 == _T_28[9:0]) begin
        image_0_115 <= io_pixelVal_in_0_4;
      end else if (10'h73 == _T_25[9:0]) begin
        image_0_115 <= io_pixelVal_in_0_3;
      end else if (10'h73 == _T_22[9:0]) begin
        image_0_115 <= io_pixelVal_in_0_2;
      end else if (10'h73 == _T_19[9:0]) begin
        image_0_115 <= io_pixelVal_in_0_1;
      end else if (10'h73 == _T_15[9:0]) begin
        image_0_115 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_116 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h74 == _T_37[9:0]) begin
        image_0_116 <= io_pixelVal_in_0_7;
      end else if (10'h74 == _T_34[9:0]) begin
        image_0_116 <= io_pixelVal_in_0_6;
      end else if (10'h74 == _T_31[9:0]) begin
        image_0_116 <= io_pixelVal_in_0_5;
      end else if (10'h74 == _T_28[9:0]) begin
        image_0_116 <= io_pixelVal_in_0_4;
      end else if (10'h74 == _T_25[9:0]) begin
        image_0_116 <= io_pixelVal_in_0_3;
      end else if (10'h74 == _T_22[9:0]) begin
        image_0_116 <= io_pixelVal_in_0_2;
      end else if (10'h74 == _T_19[9:0]) begin
        image_0_116 <= io_pixelVal_in_0_1;
      end else if (10'h74 == _T_15[9:0]) begin
        image_0_116 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_117 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h75 == _T_37[9:0]) begin
        image_0_117 <= io_pixelVal_in_0_7;
      end else if (10'h75 == _T_34[9:0]) begin
        image_0_117 <= io_pixelVal_in_0_6;
      end else if (10'h75 == _T_31[9:0]) begin
        image_0_117 <= io_pixelVal_in_0_5;
      end else if (10'h75 == _T_28[9:0]) begin
        image_0_117 <= io_pixelVal_in_0_4;
      end else if (10'h75 == _T_25[9:0]) begin
        image_0_117 <= io_pixelVal_in_0_3;
      end else if (10'h75 == _T_22[9:0]) begin
        image_0_117 <= io_pixelVal_in_0_2;
      end else if (10'h75 == _T_19[9:0]) begin
        image_0_117 <= io_pixelVal_in_0_1;
      end else if (10'h75 == _T_15[9:0]) begin
        image_0_117 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_118 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h76 == _T_37[9:0]) begin
        image_0_118 <= io_pixelVal_in_0_7;
      end else if (10'h76 == _T_34[9:0]) begin
        image_0_118 <= io_pixelVal_in_0_6;
      end else if (10'h76 == _T_31[9:0]) begin
        image_0_118 <= io_pixelVal_in_0_5;
      end else if (10'h76 == _T_28[9:0]) begin
        image_0_118 <= io_pixelVal_in_0_4;
      end else if (10'h76 == _T_25[9:0]) begin
        image_0_118 <= io_pixelVal_in_0_3;
      end else if (10'h76 == _T_22[9:0]) begin
        image_0_118 <= io_pixelVal_in_0_2;
      end else if (10'h76 == _T_19[9:0]) begin
        image_0_118 <= io_pixelVal_in_0_1;
      end else if (10'h76 == _T_15[9:0]) begin
        image_0_118 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_119 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h77 == _T_37[9:0]) begin
        image_0_119 <= io_pixelVal_in_0_7;
      end else if (10'h77 == _T_34[9:0]) begin
        image_0_119 <= io_pixelVal_in_0_6;
      end else if (10'h77 == _T_31[9:0]) begin
        image_0_119 <= io_pixelVal_in_0_5;
      end else if (10'h77 == _T_28[9:0]) begin
        image_0_119 <= io_pixelVal_in_0_4;
      end else if (10'h77 == _T_25[9:0]) begin
        image_0_119 <= io_pixelVal_in_0_3;
      end else if (10'h77 == _T_22[9:0]) begin
        image_0_119 <= io_pixelVal_in_0_2;
      end else if (10'h77 == _T_19[9:0]) begin
        image_0_119 <= io_pixelVal_in_0_1;
      end else if (10'h77 == _T_15[9:0]) begin
        image_0_119 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_120 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h78 == _T_37[9:0]) begin
        image_0_120 <= io_pixelVal_in_0_7;
      end else if (10'h78 == _T_34[9:0]) begin
        image_0_120 <= io_pixelVal_in_0_6;
      end else if (10'h78 == _T_31[9:0]) begin
        image_0_120 <= io_pixelVal_in_0_5;
      end else if (10'h78 == _T_28[9:0]) begin
        image_0_120 <= io_pixelVal_in_0_4;
      end else if (10'h78 == _T_25[9:0]) begin
        image_0_120 <= io_pixelVal_in_0_3;
      end else if (10'h78 == _T_22[9:0]) begin
        image_0_120 <= io_pixelVal_in_0_2;
      end else if (10'h78 == _T_19[9:0]) begin
        image_0_120 <= io_pixelVal_in_0_1;
      end else if (10'h78 == _T_15[9:0]) begin
        image_0_120 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_121 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h79 == _T_37[9:0]) begin
        image_0_121 <= io_pixelVal_in_0_7;
      end else if (10'h79 == _T_34[9:0]) begin
        image_0_121 <= io_pixelVal_in_0_6;
      end else if (10'h79 == _T_31[9:0]) begin
        image_0_121 <= io_pixelVal_in_0_5;
      end else if (10'h79 == _T_28[9:0]) begin
        image_0_121 <= io_pixelVal_in_0_4;
      end else if (10'h79 == _T_25[9:0]) begin
        image_0_121 <= io_pixelVal_in_0_3;
      end else if (10'h79 == _T_22[9:0]) begin
        image_0_121 <= io_pixelVal_in_0_2;
      end else if (10'h79 == _T_19[9:0]) begin
        image_0_121 <= io_pixelVal_in_0_1;
      end else if (10'h79 == _T_15[9:0]) begin
        image_0_121 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_122 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h7a == _T_37[9:0]) begin
        image_0_122 <= io_pixelVal_in_0_7;
      end else if (10'h7a == _T_34[9:0]) begin
        image_0_122 <= io_pixelVal_in_0_6;
      end else if (10'h7a == _T_31[9:0]) begin
        image_0_122 <= io_pixelVal_in_0_5;
      end else if (10'h7a == _T_28[9:0]) begin
        image_0_122 <= io_pixelVal_in_0_4;
      end else if (10'h7a == _T_25[9:0]) begin
        image_0_122 <= io_pixelVal_in_0_3;
      end else if (10'h7a == _T_22[9:0]) begin
        image_0_122 <= io_pixelVal_in_0_2;
      end else if (10'h7a == _T_19[9:0]) begin
        image_0_122 <= io_pixelVal_in_0_1;
      end else if (10'h7a == _T_15[9:0]) begin
        image_0_122 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_123 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h7b == _T_37[9:0]) begin
        image_0_123 <= io_pixelVal_in_0_7;
      end else if (10'h7b == _T_34[9:0]) begin
        image_0_123 <= io_pixelVal_in_0_6;
      end else if (10'h7b == _T_31[9:0]) begin
        image_0_123 <= io_pixelVal_in_0_5;
      end else if (10'h7b == _T_28[9:0]) begin
        image_0_123 <= io_pixelVal_in_0_4;
      end else if (10'h7b == _T_25[9:0]) begin
        image_0_123 <= io_pixelVal_in_0_3;
      end else if (10'h7b == _T_22[9:0]) begin
        image_0_123 <= io_pixelVal_in_0_2;
      end else if (10'h7b == _T_19[9:0]) begin
        image_0_123 <= io_pixelVal_in_0_1;
      end else if (10'h7b == _T_15[9:0]) begin
        image_0_123 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_124 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h7c == _T_37[9:0]) begin
        image_0_124 <= io_pixelVal_in_0_7;
      end else if (10'h7c == _T_34[9:0]) begin
        image_0_124 <= io_pixelVal_in_0_6;
      end else if (10'h7c == _T_31[9:0]) begin
        image_0_124 <= io_pixelVal_in_0_5;
      end else if (10'h7c == _T_28[9:0]) begin
        image_0_124 <= io_pixelVal_in_0_4;
      end else if (10'h7c == _T_25[9:0]) begin
        image_0_124 <= io_pixelVal_in_0_3;
      end else if (10'h7c == _T_22[9:0]) begin
        image_0_124 <= io_pixelVal_in_0_2;
      end else if (10'h7c == _T_19[9:0]) begin
        image_0_124 <= io_pixelVal_in_0_1;
      end else if (10'h7c == _T_15[9:0]) begin
        image_0_124 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_125 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h7d == _T_37[9:0]) begin
        image_0_125 <= io_pixelVal_in_0_7;
      end else if (10'h7d == _T_34[9:0]) begin
        image_0_125 <= io_pixelVal_in_0_6;
      end else if (10'h7d == _T_31[9:0]) begin
        image_0_125 <= io_pixelVal_in_0_5;
      end else if (10'h7d == _T_28[9:0]) begin
        image_0_125 <= io_pixelVal_in_0_4;
      end else if (10'h7d == _T_25[9:0]) begin
        image_0_125 <= io_pixelVal_in_0_3;
      end else if (10'h7d == _T_22[9:0]) begin
        image_0_125 <= io_pixelVal_in_0_2;
      end else if (10'h7d == _T_19[9:0]) begin
        image_0_125 <= io_pixelVal_in_0_1;
      end else if (10'h7d == _T_15[9:0]) begin
        image_0_125 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_126 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h7e == _T_37[9:0]) begin
        image_0_126 <= io_pixelVal_in_0_7;
      end else if (10'h7e == _T_34[9:0]) begin
        image_0_126 <= io_pixelVal_in_0_6;
      end else if (10'h7e == _T_31[9:0]) begin
        image_0_126 <= io_pixelVal_in_0_5;
      end else if (10'h7e == _T_28[9:0]) begin
        image_0_126 <= io_pixelVal_in_0_4;
      end else if (10'h7e == _T_25[9:0]) begin
        image_0_126 <= io_pixelVal_in_0_3;
      end else if (10'h7e == _T_22[9:0]) begin
        image_0_126 <= io_pixelVal_in_0_2;
      end else if (10'h7e == _T_19[9:0]) begin
        image_0_126 <= io_pixelVal_in_0_1;
      end else if (10'h7e == _T_15[9:0]) begin
        image_0_126 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_127 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h7f == _T_37[9:0]) begin
        image_0_127 <= io_pixelVal_in_0_7;
      end else if (10'h7f == _T_34[9:0]) begin
        image_0_127 <= io_pixelVal_in_0_6;
      end else if (10'h7f == _T_31[9:0]) begin
        image_0_127 <= io_pixelVal_in_0_5;
      end else if (10'h7f == _T_28[9:0]) begin
        image_0_127 <= io_pixelVal_in_0_4;
      end else if (10'h7f == _T_25[9:0]) begin
        image_0_127 <= io_pixelVal_in_0_3;
      end else if (10'h7f == _T_22[9:0]) begin
        image_0_127 <= io_pixelVal_in_0_2;
      end else if (10'h7f == _T_19[9:0]) begin
        image_0_127 <= io_pixelVal_in_0_1;
      end else if (10'h7f == _T_15[9:0]) begin
        image_0_127 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_128 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h80 == _T_37[9:0]) begin
        image_0_128 <= io_pixelVal_in_0_7;
      end else if (10'h80 == _T_34[9:0]) begin
        image_0_128 <= io_pixelVal_in_0_6;
      end else if (10'h80 == _T_31[9:0]) begin
        image_0_128 <= io_pixelVal_in_0_5;
      end else if (10'h80 == _T_28[9:0]) begin
        image_0_128 <= io_pixelVal_in_0_4;
      end else if (10'h80 == _T_25[9:0]) begin
        image_0_128 <= io_pixelVal_in_0_3;
      end else if (10'h80 == _T_22[9:0]) begin
        image_0_128 <= io_pixelVal_in_0_2;
      end else if (10'h80 == _T_19[9:0]) begin
        image_0_128 <= io_pixelVal_in_0_1;
      end else if (10'h80 == _T_15[9:0]) begin
        image_0_128 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_129 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h81 == _T_37[9:0]) begin
        image_0_129 <= io_pixelVal_in_0_7;
      end else if (10'h81 == _T_34[9:0]) begin
        image_0_129 <= io_pixelVal_in_0_6;
      end else if (10'h81 == _T_31[9:0]) begin
        image_0_129 <= io_pixelVal_in_0_5;
      end else if (10'h81 == _T_28[9:0]) begin
        image_0_129 <= io_pixelVal_in_0_4;
      end else if (10'h81 == _T_25[9:0]) begin
        image_0_129 <= io_pixelVal_in_0_3;
      end else if (10'h81 == _T_22[9:0]) begin
        image_0_129 <= io_pixelVal_in_0_2;
      end else if (10'h81 == _T_19[9:0]) begin
        image_0_129 <= io_pixelVal_in_0_1;
      end else if (10'h81 == _T_15[9:0]) begin
        image_0_129 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_130 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h82 == _T_37[9:0]) begin
        image_0_130 <= io_pixelVal_in_0_7;
      end else if (10'h82 == _T_34[9:0]) begin
        image_0_130 <= io_pixelVal_in_0_6;
      end else if (10'h82 == _T_31[9:0]) begin
        image_0_130 <= io_pixelVal_in_0_5;
      end else if (10'h82 == _T_28[9:0]) begin
        image_0_130 <= io_pixelVal_in_0_4;
      end else if (10'h82 == _T_25[9:0]) begin
        image_0_130 <= io_pixelVal_in_0_3;
      end else if (10'h82 == _T_22[9:0]) begin
        image_0_130 <= io_pixelVal_in_0_2;
      end else if (10'h82 == _T_19[9:0]) begin
        image_0_130 <= io_pixelVal_in_0_1;
      end else if (10'h82 == _T_15[9:0]) begin
        image_0_130 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_131 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h83 == _T_37[9:0]) begin
        image_0_131 <= io_pixelVal_in_0_7;
      end else if (10'h83 == _T_34[9:0]) begin
        image_0_131 <= io_pixelVal_in_0_6;
      end else if (10'h83 == _T_31[9:0]) begin
        image_0_131 <= io_pixelVal_in_0_5;
      end else if (10'h83 == _T_28[9:0]) begin
        image_0_131 <= io_pixelVal_in_0_4;
      end else if (10'h83 == _T_25[9:0]) begin
        image_0_131 <= io_pixelVal_in_0_3;
      end else if (10'h83 == _T_22[9:0]) begin
        image_0_131 <= io_pixelVal_in_0_2;
      end else if (10'h83 == _T_19[9:0]) begin
        image_0_131 <= io_pixelVal_in_0_1;
      end else if (10'h83 == _T_15[9:0]) begin
        image_0_131 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_132 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h84 == _T_37[9:0]) begin
        image_0_132 <= io_pixelVal_in_0_7;
      end else if (10'h84 == _T_34[9:0]) begin
        image_0_132 <= io_pixelVal_in_0_6;
      end else if (10'h84 == _T_31[9:0]) begin
        image_0_132 <= io_pixelVal_in_0_5;
      end else if (10'h84 == _T_28[9:0]) begin
        image_0_132 <= io_pixelVal_in_0_4;
      end else if (10'h84 == _T_25[9:0]) begin
        image_0_132 <= io_pixelVal_in_0_3;
      end else if (10'h84 == _T_22[9:0]) begin
        image_0_132 <= io_pixelVal_in_0_2;
      end else if (10'h84 == _T_19[9:0]) begin
        image_0_132 <= io_pixelVal_in_0_1;
      end else if (10'h84 == _T_15[9:0]) begin
        image_0_132 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_133 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h85 == _T_37[9:0]) begin
        image_0_133 <= io_pixelVal_in_0_7;
      end else if (10'h85 == _T_34[9:0]) begin
        image_0_133 <= io_pixelVal_in_0_6;
      end else if (10'h85 == _T_31[9:0]) begin
        image_0_133 <= io_pixelVal_in_0_5;
      end else if (10'h85 == _T_28[9:0]) begin
        image_0_133 <= io_pixelVal_in_0_4;
      end else if (10'h85 == _T_25[9:0]) begin
        image_0_133 <= io_pixelVal_in_0_3;
      end else if (10'h85 == _T_22[9:0]) begin
        image_0_133 <= io_pixelVal_in_0_2;
      end else if (10'h85 == _T_19[9:0]) begin
        image_0_133 <= io_pixelVal_in_0_1;
      end else if (10'h85 == _T_15[9:0]) begin
        image_0_133 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_134 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h86 == _T_37[9:0]) begin
        image_0_134 <= io_pixelVal_in_0_7;
      end else if (10'h86 == _T_34[9:0]) begin
        image_0_134 <= io_pixelVal_in_0_6;
      end else if (10'h86 == _T_31[9:0]) begin
        image_0_134 <= io_pixelVal_in_0_5;
      end else if (10'h86 == _T_28[9:0]) begin
        image_0_134 <= io_pixelVal_in_0_4;
      end else if (10'h86 == _T_25[9:0]) begin
        image_0_134 <= io_pixelVal_in_0_3;
      end else if (10'h86 == _T_22[9:0]) begin
        image_0_134 <= io_pixelVal_in_0_2;
      end else if (10'h86 == _T_19[9:0]) begin
        image_0_134 <= io_pixelVal_in_0_1;
      end else if (10'h86 == _T_15[9:0]) begin
        image_0_134 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_135 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h87 == _T_37[9:0]) begin
        image_0_135 <= io_pixelVal_in_0_7;
      end else if (10'h87 == _T_34[9:0]) begin
        image_0_135 <= io_pixelVal_in_0_6;
      end else if (10'h87 == _T_31[9:0]) begin
        image_0_135 <= io_pixelVal_in_0_5;
      end else if (10'h87 == _T_28[9:0]) begin
        image_0_135 <= io_pixelVal_in_0_4;
      end else if (10'h87 == _T_25[9:0]) begin
        image_0_135 <= io_pixelVal_in_0_3;
      end else if (10'h87 == _T_22[9:0]) begin
        image_0_135 <= io_pixelVal_in_0_2;
      end else if (10'h87 == _T_19[9:0]) begin
        image_0_135 <= io_pixelVal_in_0_1;
      end else if (10'h87 == _T_15[9:0]) begin
        image_0_135 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_136 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h88 == _T_37[9:0]) begin
        image_0_136 <= io_pixelVal_in_0_7;
      end else if (10'h88 == _T_34[9:0]) begin
        image_0_136 <= io_pixelVal_in_0_6;
      end else if (10'h88 == _T_31[9:0]) begin
        image_0_136 <= io_pixelVal_in_0_5;
      end else if (10'h88 == _T_28[9:0]) begin
        image_0_136 <= io_pixelVal_in_0_4;
      end else if (10'h88 == _T_25[9:0]) begin
        image_0_136 <= io_pixelVal_in_0_3;
      end else if (10'h88 == _T_22[9:0]) begin
        image_0_136 <= io_pixelVal_in_0_2;
      end else if (10'h88 == _T_19[9:0]) begin
        image_0_136 <= io_pixelVal_in_0_1;
      end else if (10'h88 == _T_15[9:0]) begin
        image_0_136 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_137 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h89 == _T_37[9:0]) begin
        image_0_137 <= io_pixelVal_in_0_7;
      end else if (10'h89 == _T_34[9:0]) begin
        image_0_137 <= io_pixelVal_in_0_6;
      end else if (10'h89 == _T_31[9:0]) begin
        image_0_137 <= io_pixelVal_in_0_5;
      end else if (10'h89 == _T_28[9:0]) begin
        image_0_137 <= io_pixelVal_in_0_4;
      end else if (10'h89 == _T_25[9:0]) begin
        image_0_137 <= io_pixelVal_in_0_3;
      end else if (10'h89 == _T_22[9:0]) begin
        image_0_137 <= io_pixelVal_in_0_2;
      end else if (10'h89 == _T_19[9:0]) begin
        image_0_137 <= io_pixelVal_in_0_1;
      end else if (10'h89 == _T_15[9:0]) begin
        image_0_137 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_138 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h8a == _T_37[9:0]) begin
        image_0_138 <= io_pixelVal_in_0_7;
      end else if (10'h8a == _T_34[9:0]) begin
        image_0_138 <= io_pixelVal_in_0_6;
      end else if (10'h8a == _T_31[9:0]) begin
        image_0_138 <= io_pixelVal_in_0_5;
      end else if (10'h8a == _T_28[9:0]) begin
        image_0_138 <= io_pixelVal_in_0_4;
      end else if (10'h8a == _T_25[9:0]) begin
        image_0_138 <= io_pixelVal_in_0_3;
      end else if (10'h8a == _T_22[9:0]) begin
        image_0_138 <= io_pixelVal_in_0_2;
      end else if (10'h8a == _T_19[9:0]) begin
        image_0_138 <= io_pixelVal_in_0_1;
      end else if (10'h8a == _T_15[9:0]) begin
        image_0_138 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_139 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h8b == _T_37[9:0]) begin
        image_0_139 <= io_pixelVal_in_0_7;
      end else if (10'h8b == _T_34[9:0]) begin
        image_0_139 <= io_pixelVal_in_0_6;
      end else if (10'h8b == _T_31[9:0]) begin
        image_0_139 <= io_pixelVal_in_0_5;
      end else if (10'h8b == _T_28[9:0]) begin
        image_0_139 <= io_pixelVal_in_0_4;
      end else if (10'h8b == _T_25[9:0]) begin
        image_0_139 <= io_pixelVal_in_0_3;
      end else if (10'h8b == _T_22[9:0]) begin
        image_0_139 <= io_pixelVal_in_0_2;
      end else if (10'h8b == _T_19[9:0]) begin
        image_0_139 <= io_pixelVal_in_0_1;
      end else if (10'h8b == _T_15[9:0]) begin
        image_0_139 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_140 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h8c == _T_37[9:0]) begin
        image_0_140 <= io_pixelVal_in_0_7;
      end else if (10'h8c == _T_34[9:0]) begin
        image_0_140 <= io_pixelVal_in_0_6;
      end else if (10'h8c == _T_31[9:0]) begin
        image_0_140 <= io_pixelVal_in_0_5;
      end else if (10'h8c == _T_28[9:0]) begin
        image_0_140 <= io_pixelVal_in_0_4;
      end else if (10'h8c == _T_25[9:0]) begin
        image_0_140 <= io_pixelVal_in_0_3;
      end else if (10'h8c == _T_22[9:0]) begin
        image_0_140 <= io_pixelVal_in_0_2;
      end else if (10'h8c == _T_19[9:0]) begin
        image_0_140 <= io_pixelVal_in_0_1;
      end else if (10'h8c == _T_15[9:0]) begin
        image_0_140 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_141 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h8d == _T_37[9:0]) begin
        image_0_141 <= io_pixelVal_in_0_7;
      end else if (10'h8d == _T_34[9:0]) begin
        image_0_141 <= io_pixelVal_in_0_6;
      end else if (10'h8d == _T_31[9:0]) begin
        image_0_141 <= io_pixelVal_in_0_5;
      end else if (10'h8d == _T_28[9:0]) begin
        image_0_141 <= io_pixelVal_in_0_4;
      end else if (10'h8d == _T_25[9:0]) begin
        image_0_141 <= io_pixelVal_in_0_3;
      end else if (10'h8d == _T_22[9:0]) begin
        image_0_141 <= io_pixelVal_in_0_2;
      end else if (10'h8d == _T_19[9:0]) begin
        image_0_141 <= io_pixelVal_in_0_1;
      end else if (10'h8d == _T_15[9:0]) begin
        image_0_141 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_142 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h8e == _T_37[9:0]) begin
        image_0_142 <= io_pixelVal_in_0_7;
      end else if (10'h8e == _T_34[9:0]) begin
        image_0_142 <= io_pixelVal_in_0_6;
      end else if (10'h8e == _T_31[9:0]) begin
        image_0_142 <= io_pixelVal_in_0_5;
      end else if (10'h8e == _T_28[9:0]) begin
        image_0_142 <= io_pixelVal_in_0_4;
      end else if (10'h8e == _T_25[9:0]) begin
        image_0_142 <= io_pixelVal_in_0_3;
      end else if (10'h8e == _T_22[9:0]) begin
        image_0_142 <= io_pixelVal_in_0_2;
      end else if (10'h8e == _T_19[9:0]) begin
        image_0_142 <= io_pixelVal_in_0_1;
      end else if (10'h8e == _T_15[9:0]) begin
        image_0_142 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_143 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h8f == _T_37[9:0]) begin
        image_0_143 <= io_pixelVal_in_0_7;
      end else if (10'h8f == _T_34[9:0]) begin
        image_0_143 <= io_pixelVal_in_0_6;
      end else if (10'h8f == _T_31[9:0]) begin
        image_0_143 <= io_pixelVal_in_0_5;
      end else if (10'h8f == _T_28[9:0]) begin
        image_0_143 <= io_pixelVal_in_0_4;
      end else if (10'h8f == _T_25[9:0]) begin
        image_0_143 <= io_pixelVal_in_0_3;
      end else if (10'h8f == _T_22[9:0]) begin
        image_0_143 <= io_pixelVal_in_0_2;
      end else if (10'h8f == _T_19[9:0]) begin
        image_0_143 <= io_pixelVal_in_0_1;
      end else if (10'h8f == _T_15[9:0]) begin
        image_0_143 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_144 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h90 == _T_37[9:0]) begin
        image_0_144 <= io_pixelVal_in_0_7;
      end else if (10'h90 == _T_34[9:0]) begin
        image_0_144 <= io_pixelVal_in_0_6;
      end else if (10'h90 == _T_31[9:0]) begin
        image_0_144 <= io_pixelVal_in_0_5;
      end else if (10'h90 == _T_28[9:0]) begin
        image_0_144 <= io_pixelVal_in_0_4;
      end else if (10'h90 == _T_25[9:0]) begin
        image_0_144 <= io_pixelVal_in_0_3;
      end else if (10'h90 == _T_22[9:0]) begin
        image_0_144 <= io_pixelVal_in_0_2;
      end else if (10'h90 == _T_19[9:0]) begin
        image_0_144 <= io_pixelVal_in_0_1;
      end else if (10'h90 == _T_15[9:0]) begin
        image_0_144 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_145 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h91 == _T_37[9:0]) begin
        image_0_145 <= io_pixelVal_in_0_7;
      end else if (10'h91 == _T_34[9:0]) begin
        image_0_145 <= io_pixelVal_in_0_6;
      end else if (10'h91 == _T_31[9:0]) begin
        image_0_145 <= io_pixelVal_in_0_5;
      end else if (10'h91 == _T_28[9:0]) begin
        image_0_145 <= io_pixelVal_in_0_4;
      end else if (10'h91 == _T_25[9:0]) begin
        image_0_145 <= io_pixelVal_in_0_3;
      end else if (10'h91 == _T_22[9:0]) begin
        image_0_145 <= io_pixelVal_in_0_2;
      end else if (10'h91 == _T_19[9:0]) begin
        image_0_145 <= io_pixelVal_in_0_1;
      end else if (10'h91 == _T_15[9:0]) begin
        image_0_145 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_146 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h92 == _T_37[9:0]) begin
        image_0_146 <= io_pixelVal_in_0_7;
      end else if (10'h92 == _T_34[9:0]) begin
        image_0_146 <= io_pixelVal_in_0_6;
      end else if (10'h92 == _T_31[9:0]) begin
        image_0_146 <= io_pixelVal_in_0_5;
      end else if (10'h92 == _T_28[9:0]) begin
        image_0_146 <= io_pixelVal_in_0_4;
      end else if (10'h92 == _T_25[9:0]) begin
        image_0_146 <= io_pixelVal_in_0_3;
      end else if (10'h92 == _T_22[9:0]) begin
        image_0_146 <= io_pixelVal_in_0_2;
      end else if (10'h92 == _T_19[9:0]) begin
        image_0_146 <= io_pixelVal_in_0_1;
      end else if (10'h92 == _T_15[9:0]) begin
        image_0_146 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_147 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h93 == _T_37[9:0]) begin
        image_0_147 <= io_pixelVal_in_0_7;
      end else if (10'h93 == _T_34[9:0]) begin
        image_0_147 <= io_pixelVal_in_0_6;
      end else if (10'h93 == _T_31[9:0]) begin
        image_0_147 <= io_pixelVal_in_0_5;
      end else if (10'h93 == _T_28[9:0]) begin
        image_0_147 <= io_pixelVal_in_0_4;
      end else if (10'h93 == _T_25[9:0]) begin
        image_0_147 <= io_pixelVal_in_0_3;
      end else if (10'h93 == _T_22[9:0]) begin
        image_0_147 <= io_pixelVal_in_0_2;
      end else if (10'h93 == _T_19[9:0]) begin
        image_0_147 <= io_pixelVal_in_0_1;
      end else if (10'h93 == _T_15[9:0]) begin
        image_0_147 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_148 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h94 == _T_37[9:0]) begin
        image_0_148 <= io_pixelVal_in_0_7;
      end else if (10'h94 == _T_34[9:0]) begin
        image_0_148 <= io_pixelVal_in_0_6;
      end else if (10'h94 == _T_31[9:0]) begin
        image_0_148 <= io_pixelVal_in_0_5;
      end else if (10'h94 == _T_28[9:0]) begin
        image_0_148 <= io_pixelVal_in_0_4;
      end else if (10'h94 == _T_25[9:0]) begin
        image_0_148 <= io_pixelVal_in_0_3;
      end else if (10'h94 == _T_22[9:0]) begin
        image_0_148 <= io_pixelVal_in_0_2;
      end else if (10'h94 == _T_19[9:0]) begin
        image_0_148 <= io_pixelVal_in_0_1;
      end else if (10'h94 == _T_15[9:0]) begin
        image_0_148 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_149 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h95 == _T_37[9:0]) begin
        image_0_149 <= io_pixelVal_in_0_7;
      end else if (10'h95 == _T_34[9:0]) begin
        image_0_149 <= io_pixelVal_in_0_6;
      end else if (10'h95 == _T_31[9:0]) begin
        image_0_149 <= io_pixelVal_in_0_5;
      end else if (10'h95 == _T_28[9:0]) begin
        image_0_149 <= io_pixelVal_in_0_4;
      end else if (10'h95 == _T_25[9:0]) begin
        image_0_149 <= io_pixelVal_in_0_3;
      end else if (10'h95 == _T_22[9:0]) begin
        image_0_149 <= io_pixelVal_in_0_2;
      end else if (10'h95 == _T_19[9:0]) begin
        image_0_149 <= io_pixelVal_in_0_1;
      end else if (10'h95 == _T_15[9:0]) begin
        image_0_149 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_150 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h96 == _T_37[9:0]) begin
        image_0_150 <= io_pixelVal_in_0_7;
      end else if (10'h96 == _T_34[9:0]) begin
        image_0_150 <= io_pixelVal_in_0_6;
      end else if (10'h96 == _T_31[9:0]) begin
        image_0_150 <= io_pixelVal_in_0_5;
      end else if (10'h96 == _T_28[9:0]) begin
        image_0_150 <= io_pixelVal_in_0_4;
      end else if (10'h96 == _T_25[9:0]) begin
        image_0_150 <= io_pixelVal_in_0_3;
      end else if (10'h96 == _T_22[9:0]) begin
        image_0_150 <= io_pixelVal_in_0_2;
      end else if (10'h96 == _T_19[9:0]) begin
        image_0_150 <= io_pixelVal_in_0_1;
      end else if (10'h96 == _T_15[9:0]) begin
        image_0_150 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_151 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h97 == _T_37[9:0]) begin
        image_0_151 <= io_pixelVal_in_0_7;
      end else if (10'h97 == _T_34[9:0]) begin
        image_0_151 <= io_pixelVal_in_0_6;
      end else if (10'h97 == _T_31[9:0]) begin
        image_0_151 <= io_pixelVal_in_0_5;
      end else if (10'h97 == _T_28[9:0]) begin
        image_0_151 <= io_pixelVal_in_0_4;
      end else if (10'h97 == _T_25[9:0]) begin
        image_0_151 <= io_pixelVal_in_0_3;
      end else if (10'h97 == _T_22[9:0]) begin
        image_0_151 <= io_pixelVal_in_0_2;
      end else if (10'h97 == _T_19[9:0]) begin
        image_0_151 <= io_pixelVal_in_0_1;
      end else if (10'h97 == _T_15[9:0]) begin
        image_0_151 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_152 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h98 == _T_37[9:0]) begin
        image_0_152 <= io_pixelVal_in_0_7;
      end else if (10'h98 == _T_34[9:0]) begin
        image_0_152 <= io_pixelVal_in_0_6;
      end else if (10'h98 == _T_31[9:0]) begin
        image_0_152 <= io_pixelVal_in_0_5;
      end else if (10'h98 == _T_28[9:0]) begin
        image_0_152 <= io_pixelVal_in_0_4;
      end else if (10'h98 == _T_25[9:0]) begin
        image_0_152 <= io_pixelVal_in_0_3;
      end else if (10'h98 == _T_22[9:0]) begin
        image_0_152 <= io_pixelVal_in_0_2;
      end else if (10'h98 == _T_19[9:0]) begin
        image_0_152 <= io_pixelVal_in_0_1;
      end else if (10'h98 == _T_15[9:0]) begin
        image_0_152 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_153 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h99 == _T_37[9:0]) begin
        image_0_153 <= io_pixelVal_in_0_7;
      end else if (10'h99 == _T_34[9:0]) begin
        image_0_153 <= io_pixelVal_in_0_6;
      end else if (10'h99 == _T_31[9:0]) begin
        image_0_153 <= io_pixelVal_in_0_5;
      end else if (10'h99 == _T_28[9:0]) begin
        image_0_153 <= io_pixelVal_in_0_4;
      end else if (10'h99 == _T_25[9:0]) begin
        image_0_153 <= io_pixelVal_in_0_3;
      end else if (10'h99 == _T_22[9:0]) begin
        image_0_153 <= io_pixelVal_in_0_2;
      end else if (10'h99 == _T_19[9:0]) begin
        image_0_153 <= io_pixelVal_in_0_1;
      end else if (10'h99 == _T_15[9:0]) begin
        image_0_153 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_154 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h9a == _T_37[9:0]) begin
        image_0_154 <= io_pixelVal_in_0_7;
      end else if (10'h9a == _T_34[9:0]) begin
        image_0_154 <= io_pixelVal_in_0_6;
      end else if (10'h9a == _T_31[9:0]) begin
        image_0_154 <= io_pixelVal_in_0_5;
      end else if (10'h9a == _T_28[9:0]) begin
        image_0_154 <= io_pixelVal_in_0_4;
      end else if (10'h9a == _T_25[9:0]) begin
        image_0_154 <= io_pixelVal_in_0_3;
      end else if (10'h9a == _T_22[9:0]) begin
        image_0_154 <= io_pixelVal_in_0_2;
      end else if (10'h9a == _T_19[9:0]) begin
        image_0_154 <= io_pixelVal_in_0_1;
      end else if (10'h9a == _T_15[9:0]) begin
        image_0_154 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_155 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h9b == _T_37[9:0]) begin
        image_0_155 <= io_pixelVal_in_0_7;
      end else if (10'h9b == _T_34[9:0]) begin
        image_0_155 <= io_pixelVal_in_0_6;
      end else if (10'h9b == _T_31[9:0]) begin
        image_0_155 <= io_pixelVal_in_0_5;
      end else if (10'h9b == _T_28[9:0]) begin
        image_0_155 <= io_pixelVal_in_0_4;
      end else if (10'h9b == _T_25[9:0]) begin
        image_0_155 <= io_pixelVal_in_0_3;
      end else if (10'h9b == _T_22[9:0]) begin
        image_0_155 <= io_pixelVal_in_0_2;
      end else if (10'h9b == _T_19[9:0]) begin
        image_0_155 <= io_pixelVal_in_0_1;
      end else if (10'h9b == _T_15[9:0]) begin
        image_0_155 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_156 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h9c == _T_37[9:0]) begin
        image_0_156 <= io_pixelVal_in_0_7;
      end else if (10'h9c == _T_34[9:0]) begin
        image_0_156 <= io_pixelVal_in_0_6;
      end else if (10'h9c == _T_31[9:0]) begin
        image_0_156 <= io_pixelVal_in_0_5;
      end else if (10'h9c == _T_28[9:0]) begin
        image_0_156 <= io_pixelVal_in_0_4;
      end else if (10'h9c == _T_25[9:0]) begin
        image_0_156 <= io_pixelVal_in_0_3;
      end else if (10'h9c == _T_22[9:0]) begin
        image_0_156 <= io_pixelVal_in_0_2;
      end else if (10'h9c == _T_19[9:0]) begin
        image_0_156 <= io_pixelVal_in_0_1;
      end else if (10'h9c == _T_15[9:0]) begin
        image_0_156 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_157 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h9d == _T_37[9:0]) begin
        image_0_157 <= io_pixelVal_in_0_7;
      end else if (10'h9d == _T_34[9:0]) begin
        image_0_157 <= io_pixelVal_in_0_6;
      end else if (10'h9d == _T_31[9:0]) begin
        image_0_157 <= io_pixelVal_in_0_5;
      end else if (10'h9d == _T_28[9:0]) begin
        image_0_157 <= io_pixelVal_in_0_4;
      end else if (10'h9d == _T_25[9:0]) begin
        image_0_157 <= io_pixelVal_in_0_3;
      end else if (10'h9d == _T_22[9:0]) begin
        image_0_157 <= io_pixelVal_in_0_2;
      end else if (10'h9d == _T_19[9:0]) begin
        image_0_157 <= io_pixelVal_in_0_1;
      end else if (10'h9d == _T_15[9:0]) begin
        image_0_157 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_158 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h9e == _T_37[9:0]) begin
        image_0_158 <= io_pixelVal_in_0_7;
      end else if (10'h9e == _T_34[9:0]) begin
        image_0_158 <= io_pixelVal_in_0_6;
      end else if (10'h9e == _T_31[9:0]) begin
        image_0_158 <= io_pixelVal_in_0_5;
      end else if (10'h9e == _T_28[9:0]) begin
        image_0_158 <= io_pixelVal_in_0_4;
      end else if (10'h9e == _T_25[9:0]) begin
        image_0_158 <= io_pixelVal_in_0_3;
      end else if (10'h9e == _T_22[9:0]) begin
        image_0_158 <= io_pixelVal_in_0_2;
      end else if (10'h9e == _T_19[9:0]) begin
        image_0_158 <= io_pixelVal_in_0_1;
      end else if (10'h9e == _T_15[9:0]) begin
        image_0_158 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_159 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h9f == _T_37[9:0]) begin
        image_0_159 <= io_pixelVal_in_0_7;
      end else if (10'h9f == _T_34[9:0]) begin
        image_0_159 <= io_pixelVal_in_0_6;
      end else if (10'h9f == _T_31[9:0]) begin
        image_0_159 <= io_pixelVal_in_0_5;
      end else if (10'h9f == _T_28[9:0]) begin
        image_0_159 <= io_pixelVal_in_0_4;
      end else if (10'h9f == _T_25[9:0]) begin
        image_0_159 <= io_pixelVal_in_0_3;
      end else if (10'h9f == _T_22[9:0]) begin
        image_0_159 <= io_pixelVal_in_0_2;
      end else if (10'h9f == _T_19[9:0]) begin
        image_0_159 <= io_pixelVal_in_0_1;
      end else if (10'h9f == _T_15[9:0]) begin
        image_0_159 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_160 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'ha0 == _T_37[9:0]) begin
        image_0_160 <= io_pixelVal_in_0_7;
      end else if (10'ha0 == _T_34[9:0]) begin
        image_0_160 <= io_pixelVal_in_0_6;
      end else if (10'ha0 == _T_31[9:0]) begin
        image_0_160 <= io_pixelVal_in_0_5;
      end else if (10'ha0 == _T_28[9:0]) begin
        image_0_160 <= io_pixelVal_in_0_4;
      end else if (10'ha0 == _T_25[9:0]) begin
        image_0_160 <= io_pixelVal_in_0_3;
      end else if (10'ha0 == _T_22[9:0]) begin
        image_0_160 <= io_pixelVal_in_0_2;
      end else if (10'ha0 == _T_19[9:0]) begin
        image_0_160 <= io_pixelVal_in_0_1;
      end else if (10'ha0 == _T_15[9:0]) begin
        image_0_160 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_161 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'ha1 == _T_37[9:0]) begin
        image_0_161 <= io_pixelVal_in_0_7;
      end else if (10'ha1 == _T_34[9:0]) begin
        image_0_161 <= io_pixelVal_in_0_6;
      end else if (10'ha1 == _T_31[9:0]) begin
        image_0_161 <= io_pixelVal_in_0_5;
      end else if (10'ha1 == _T_28[9:0]) begin
        image_0_161 <= io_pixelVal_in_0_4;
      end else if (10'ha1 == _T_25[9:0]) begin
        image_0_161 <= io_pixelVal_in_0_3;
      end else if (10'ha1 == _T_22[9:0]) begin
        image_0_161 <= io_pixelVal_in_0_2;
      end else if (10'ha1 == _T_19[9:0]) begin
        image_0_161 <= io_pixelVal_in_0_1;
      end else if (10'ha1 == _T_15[9:0]) begin
        image_0_161 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_162 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'ha2 == _T_37[9:0]) begin
        image_0_162 <= io_pixelVal_in_0_7;
      end else if (10'ha2 == _T_34[9:0]) begin
        image_0_162 <= io_pixelVal_in_0_6;
      end else if (10'ha2 == _T_31[9:0]) begin
        image_0_162 <= io_pixelVal_in_0_5;
      end else if (10'ha2 == _T_28[9:0]) begin
        image_0_162 <= io_pixelVal_in_0_4;
      end else if (10'ha2 == _T_25[9:0]) begin
        image_0_162 <= io_pixelVal_in_0_3;
      end else if (10'ha2 == _T_22[9:0]) begin
        image_0_162 <= io_pixelVal_in_0_2;
      end else if (10'ha2 == _T_19[9:0]) begin
        image_0_162 <= io_pixelVal_in_0_1;
      end else if (10'ha2 == _T_15[9:0]) begin
        image_0_162 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_163 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'ha3 == _T_37[9:0]) begin
        image_0_163 <= io_pixelVal_in_0_7;
      end else if (10'ha3 == _T_34[9:0]) begin
        image_0_163 <= io_pixelVal_in_0_6;
      end else if (10'ha3 == _T_31[9:0]) begin
        image_0_163 <= io_pixelVal_in_0_5;
      end else if (10'ha3 == _T_28[9:0]) begin
        image_0_163 <= io_pixelVal_in_0_4;
      end else if (10'ha3 == _T_25[9:0]) begin
        image_0_163 <= io_pixelVal_in_0_3;
      end else if (10'ha3 == _T_22[9:0]) begin
        image_0_163 <= io_pixelVal_in_0_2;
      end else if (10'ha3 == _T_19[9:0]) begin
        image_0_163 <= io_pixelVal_in_0_1;
      end else if (10'ha3 == _T_15[9:0]) begin
        image_0_163 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_164 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'ha4 == _T_37[9:0]) begin
        image_0_164 <= io_pixelVal_in_0_7;
      end else if (10'ha4 == _T_34[9:0]) begin
        image_0_164 <= io_pixelVal_in_0_6;
      end else if (10'ha4 == _T_31[9:0]) begin
        image_0_164 <= io_pixelVal_in_0_5;
      end else if (10'ha4 == _T_28[9:0]) begin
        image_0_164 <= io_pixelVal_in_0_4;
      end else if (10'ha4 == _T_25[9:0]) begin
        image_0_164 <= io_pixelVal_in_0_3;
      end else if (10'ha4 == _T_22[9:0]) begin
        image_0_164 <= io_pixelVal_in_0_2;
      end else if (10'ha4 == _T_19[9:0]) begin
        image_0_164 <= io_pixelVal_in_0_1;
      end else if (10'ha4 == _T_15[9:0]) begin
        image_0_164 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_165 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'ha5 == _T_37[9:0]) begin
        image_0_165 <= io_pixelVal_in_0_7;
      end else if (10'ha5 == _T_34[9:0]) begin
        image_0_165 <= io_pixelVal_in_0_6;
      end else if (10'ha5 == _T_31[9:0]) begin
        image_0_165 <= io_pixelVal_in_0_5;
      end else if (10'ha5 == _T_28[9:0]) begin
        image_0_165 <= io_pixelVal_in_0_4;
      end else if (10'ha5 == _T_25[9:0]) begin
        image_0_165 <= io_pixelVal_in_0_3;
      end else if (10'ha5 == _T_22[9:0]) begin
        image_0_165 <= io_pixelVal_in_0_2;
      end else if (10'ha5 == _T_19[9:0]) begin
        image_0_165 <= io_pixelVal_in_0_1;
      end else if (10'ha5 == _T_15[9:0]) begin
        image_0_165 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_166 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'ha6 == _T_37[9:0]) begin
        image_0_166 <= io_pixelVal_in_0_7;
      end else if (10'ha6 == _T_34[9:0]) begin
        image_0_166 <= io_pixelVal_in_0_6;
      end else if (10'ha6 == _T_31[9:0]) begin
        image_0_166 <= io_pixelVal_in_0_5;
      end else if (10'ha6 == _T_28[9:0]) begin
        image_0_166 <= io_pixelVal_in_0_4;
      end else if (10'ha6 == _T_25[9:0]) begin
        image_0_166 <= io_pixelVal_in_0_3;
      end else if (10'ha6 == _T_22[9:0]) begin
        image_0_166 <= io_pixelVal_in_0_2;
      end else if (10'ha6 == _T_19[9:0]) begin
        image_0_166 <= io_pixelVal_in_0_1;
      end else if (10'ha6 == _T_15[9:0]) begin
        image_0_166 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_167 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'ha7 == _T_37[9:0]) begin
        image_0_167 <= io_pixelVal_in_0_7;
      end else if (10'ha7 == _T_34[9:0]) begin
        image_0_167 <= io_pixelVal_in_0_6;
      end else if (10'ha7 == _T_31[9:0]) begin
        image_0_167 <= io_pixelVal_in_0_5;
      end else if (10'ha7 == _T_28[9:0]) begin
        image_0_167 <= io_pixelVal_in_0_4;
      end else if (10'ha7 == _T_25[9:0]) begin
        image_0_167 <= io_pixelVal_in_0_3;
      end else if (10'ha7 == _T_22[9:0]) begin
        image_0_167 <= io_pixelVal_in_0_2;
      end else if (10'ha7 == _T_19[9:0]) begin
        image_0_167 <= io_pixelVal_in_0_1;
      end else if (10'ha7 == _T_15[9:0]) begin
        image_0_167 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_168 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'ha8 == _T_37[9:0]) begin
        image_0_168 <= io_pixelVal_in_0_7;
      end else if (10'ha8 == _T_34[9:0]) begin
        image_0_168 <= io_pixelVal_in_0_6;
      end else if (10'ha8 == _T_31[9:0]) begin
        image_0_168 <= io_pixelVal_in_0_5;
      end else if (10'ha8 == _T_28[9:0]) begin
        image_0_168 <= io_pixelVal_in_0_4;
      end else if (10'ha8 == _T_25[9:0]) begin
        image_0_168 <= io_pixelVal_in_0_3;
      end else if (10'ha8 == _T_22[9:0]) begin
        image_0_168 <= io_pixelVal_in_0_2;
      end else if (10'ha8 == _T_19[9:0]) begin
        image_0_168 <= io_pixelVal_in_0_1;
      end else if (10'ha8 == _T_15[9:0]) begin
        image_0_168 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_169 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'ha9 == _T_37[9:0]) begin
        image_0_169 <= io_pixelVal_in_0_7;
      end else if (10'ha9 == _T_34[9:0]) begin
        image_0_169 <= io_pixelVal_in_0_6;
      end else if (10'ha9 == _T_31[9:0]) begin
        image_0_169 <= io_pixelVal_in_0_5;
      end else if (10'ha9 == _T_28[9:0]) begin
        image_0_169 <= io_pixelVal_in_0_4;
      end else if (10'ha9 == _T_25[9:0]) begin
        image_0_169 <= io_pixelVal_in_0_3;
      end else if (10'ha9 == _T_22[9:0]) begin
        image_0_169 <= io_pixelVal_in_0_2;
      end else if (10'ha9 == _T_19[9:0]) begin
        image_0_169 <= io_pixelVal_in_0_1;
      end else if (10'ha9 == _T_15[9:0]) begin
        image_0_169 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_170 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'haa == _T_37[9:0]) begin
        image_0_170 <= io_pixelVal_in_0_7;
      end else if (10'haa == _T_34[9:0]) begin
        image_0_170 <= io_pixelVal_in_0_6;
      end else if (10'haa == _T_31[9:0]) begin
        image_0_170 <= io_pixelVal_in_0_5;
      end else if (10'haa == _T_28[9:0]) begin
        image_0_170 <= io_pixelVal_in_0_4;
      end else if (10'haa == _T_25[9:0]) begin
        image_0_170 <= io_pixelVal_in_0_3;
      end else if (10'haa == _T_22[9:0]) begin
        image_0_170 <= io_pixelVal_in_0_2;
      end else if (10'haa == _T_19[9:0]) begin
        image_0_170 <= io_pixelVal_in_0_1;
      end else if (10'haa == _T_15[9:0]) begin
        image_0_170 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_171 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hab == _T_37[9:0]) begin
        image_0_171 <= io_pixelVal_in_0_7;
      end else if (10'hab == _T_34[9:0]) begin
        image_0_171 <= io_pixelVal_in_0_6;
      end else if (10'hab == _T_31[9:0]) begin
        image_0_171 <= io_pixelVal_in_0_5;
      end else if (10'hab == _T_28[9:0]) begin
        image_0_171 <= io_pixelVal_in_0_4;
      end else if (10'hab == _T_25[9:0]) begin
        image_0_171 <= io_pixelVal_in_0_3;
      end else if (10'hab == _T_22[9:0]) begin
        image_0_171 <= io_pixelVal_in_0_2;
      end else if (10'hab == _T_19[9:0]) begin
        image_0_171 <= io_pixelVal_in_0_1;
      end else if (10'hab == _T_15[9:0]) begin
        image_0_171 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_172 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hac == _T_37[9:0]) begin
        image_0_172 <= io_pixelVal_in_0_7;
      end else if (10'hac == _T_34[9:0]) begin
        image_0_172 <= io_pixelVal_in_0_6;
      end else if (10'hac == _T_31[9:0]) begin
        image_0_172 <= io_pixelVal_in_0_5;
      end else if (10'hac == _T_28[9:0]) begin
        image_0_172 <= io_pixelVal_in_0_4;
      end else if (10'hac == _T_25[9:0]) begin
        image_0_172 <= io_pixelVal_in_0_3;
      end else if (10'hac == _T_22[9:0]) begin
        image_0_172 <= io_pixelVal_in_0_2;
      end else if (10'hac == _T_19[9:0]) begin
        image_0_172 <= io_pixelVal_in_0_1;
      end else if (10'hac == _T_15[9:0]) begin
        image_0_172 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_173 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'had == _T_37[9:0]) begin
        image_0_173 <= io_pixelVal_in_0_7;
      end else if (10'had == _T_34[9:0]) begin
        image_0_173 <= io_pixelVal_in_0_6;
      end else if (10'had == _T_31[9:0]) begin
        image_0_173 <= io_pixelVal_in_0_5;
      end else if (10'had == _T_28[9:0]) begin
        image_0_173 <= io_pixelVal_in_0_4;
      end else if (10'had == _T_25[9:0]) begin
        image_0_173 <= io_pixelVal_in_0_3;
      end else if (10'had == _T_22[9:0]) begin
        image_0_173 <= io_pixelVal_in_0_2;
      end else if (10'had == _T_19[9:0]) begin
        image_0_173 <= io_pixelVal_in_0_1;
      end else if (10'had == _T_15[9:0]) begin
        image_0_173 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_174 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hae == _T_37[9:0]) begin
        image_0_174 <= io_pixelVal_in_0_7;
      end else if (10'hae == _T_34[9:0]) begin
        image_0_174 <= io_pixelVal_in_0_6;
      end else if (10'hae == _T_31[9:0]) begin
        image_0_174 <= io_pixelVal_in_0_5;
      end else if (10'hae == _T_28[9:0]) begin
        image_0_174 <= io_pixelVal_in_0_4;
      end else if (10'hae == _T_25[9:0]) begin
        image_0_174 <= io_pixelVal_in_0_3;
      end else if (10'hae == _T_22[9:0]) begin
        image_0_174 <= io_pixelVal_in_0_2;
      end else if (10'hae == _T_19[9:0]) begin
        image_0_174 <= io_pixelVal_in_0_1;
      end else if (10'hae == _T_15[9:0]) begin
        image_0_174 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_175 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'haf == _T_37[9:0]) begin
        image_0_175 <= io_pixelVal_in_0_7;
      end else if (10'haf == _T_34[9:0]) begin
        image_0_175 <= io_pixelVal_in_0_6;
      end else if (10'haf == _T_31[9:0]) begin
        image_0_175 <= io_pixelVal_in_0_5;
      end else if (10'haf == _T_28[9:0]) begin
        image_0_175 <= io_pixelVal_in_0_4;
      end else if (10'haf == _T_25[9:0]) begin
        image_0_175 <= io_pixelVal_in_0_3;
      end else if (10'haf == _T_22[9:0]) begin
        image_0_175 <= io_pixelVal_in_0_2;
      end else if (10'haf == _T_19[9:0]) begin
        image_0_175 <= io_pixelVal_in_0_1;
      end else if (10'haf == _T_15[9:0]) begin
        image_0_175 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_176 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hb0 == _T_37[9:0]) begin
        image_0_176 <= io_pixelVal_in_0_7;
      end else if (10'hb0 == _T_34[9:0]) begin
        image_0_176 <= io_pixelVal_in_0_6;
      end else if (10'hb0 == _T_31[9:0]) begin
        image_0_176 <= io_pixelVal_in_0_5;
      end else if (10'hb0 == _T_28[9:0]) begin
        image_0_176 <= io_pixelVal_in_0_4;
      end else if (10'hb0 == _T_25[9:0]) begin
        image_0_176 <= io_pixelVal_in_0_3;
      end else if (10'hb0 == _T_22[9:0]) begin
        image_0_176 <= io_pixelVal_in_0_2;
      end else if (10'hb0 == _T_19[9:0]) begin
        image_0_176 <= io_pixelVal_in_0_1;
      end else if (10'hb0 == _T_15[9:0]) begin
        image_0_176 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_177 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hb1 == _T_37[9:0]) begin
        image_0_177 <= io_pixelVal_in_0_7;
      end else if (10'hb1 == _T_34[9:0]) begin
        image_0_177 <= io_pixelVal_in_0_6;
      end else if (10'hb1 == _T_31[9:0]) begin
        image_0_177 <= io_pixelVal_in_0_5;
      end else if (10'hb1 == _T_28[9:0]) begin
        image_0_177 <= io_pixelVal_in_0_4;
      end else if (10'hb1 == _T_25[9:0]) begin
        image_0_177 <= io_pixelVal_in_0_3;
      end else if (10'hb1 == _T_22[9:0]) begin
        image_0_177 <= io_pixelVal_in_0_2;
      end else if (10'hb1 == _T_19[9:0]) begin
        image_0_177 <= io_pixelVal_in_0_1;
      end else if (10'hb1 == _T_15[9:0]) begin
        image_0_177 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_178 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hb2 == _T_37[9:0]) begin
        image_0_178 <= io_pixelVal_in_0_7;
      end else if (10'hb2 == _T_34[9:0]) begin
        image_0_178 <= io_pixelVal_in_0_6;
      end else if (10'hb2 == _T_31[9:0]) begin
        image_0_178 <= io_pixelVal_in_0_5;
      end else if (10'hb2 == _T_28[9:0]) begin
        image_0_178 <= io_pixelVal_in_0_4;
      end else if (10'hb2 == _T_25[9:0]) begin
        image_0_178 <= io_pixelVal_in_0_3;
      end else if (10'hb2 == _T_22[9:0]) begin
        image_0_178 <= io_pixelVal_in_0_2;
      end else if (10'hb2 == _T_19[9:0]) begin
        image_0_178 <= io_pixelVal_in_0_1;
      end else if (10'hb2 == _T_15[9:0]) begin
        image_0_178 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_179 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hb3 == _T_37[9:0]) begin
        image_0_179 <= io_pixelVal_in_0_7;
      end else if (10'hb3 == _T_34[9:0]) begin
        image_0_179 <= io_pixelVal_in_0_6;
      end else if (10'hb3 == _T_31[9:0]) begin
        image_0_179 <= io_pixelVal_in_0_5;
      end else if (10'hb3 == _T_28[9:0]) begin
        image_0_179 <= io_pixelVal_in_0_4;
      end else if (10'hb3 == _T_25[9:0]) begin
        image_0_179 <= io_pixelVal_in_0_3;
      end else if (10'hb3 == _T_22[9:0]) begin
        image_0_179 <= io_pixelVal_in_0_2;
      end else if (10'hb3 == _T_19[9:0]) begin
        image_0_179 <= io_pixelVal_in_0_1;
      end else if (10'hb3 == _T_15[9:0]) begin
        image_0_179 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_180 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hb4 == _T_37[9:0]) begin
        image_0_180 <= io_pixelVal_in_0_7;
      end else if (10'hb4 == _T_34[9:0]) begin
        image_0_180 <= io_pixelVal_in_0_6;
      end else if (10'hb4 == _T_31[9:0]) begin
        image_0_180 <= io_pixelVal_in_0_5;
      end else if (10'hb4 == _T_28[9:0]) begin
        image_0_180 <= io_pixelVal_in_0_4;
      end else if (10'hb4 == _T_25[9:0]) begin
        image_0_180 <= io_pixelVal_in_0_3;
      end else if (10'hb4 == _T_22[9:0]) begin
        image_0_180 <= io_pixelVal_in_0_2;
      end else if (10'hb4 == _T_19[9:0]) begin
        image_0_180 <= io_pixelVal_in_0_1;
      end else if (10'hb4 == _T_15[9:0]) begin
        image_0_180 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_181 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hb5 == _T_37[9:0]) begin
        image_0_181 <= io_pixelVal_in_0_7;
      end else if (10'hb5 == _T_34[9:0]) begin
        image_0_181 <= io_pixelVal_in_0_6;
      end else if (10'hb5 == _T_31[9:0]) begin
        image_0_181 <= io_pixelVal_in_0_5;
      end else if (10'hb5 == _T_28[9:0]) begin
        image_0_181 <= io_pixelVal_in_0_4;
      end else if (10'hb5 == _T_25[9:0]) begin
        image_0_181 <= io_pixelVal_in_0_3;
      end else if (10'hb5 == _T_22[9:0]) begin
        image_0_181 <= io_pixelVal_in_0_2;
      end else if (10'hb5 == _T_19[9:0]) begin
        image_0_181 <= io_pixelVal_in_0_1;
      end else if (10'hb5 == _T_15[9:0]) begin
        image_0_181 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_182 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hb6 == _T_37[9:0]) begin
        image_0_182 <= io_pixelVal_in_0_7;
      end else if (10'hb6 == _T_34[9:0]) begin
        image_0_182 <= io_pixelVal_in_0_6;
      end else if (10'hb6 == _T_31[9:0]) begin
        image_0_182 <= io_pixelVal_in_0_5;
      end else if (10'hb6 == _T_28[9:0]) begin
        image_0_182 <= io_pixelVal_in_0_4;
      end else if (10'hb6 == _T_25[9:0]) begin
        image_0_182 <= io_pixelVal_in_0_3;
      end else if (10'hb6 == _T_22[9:0]) begin
        image_0_182 <= io_pixelVal_in_0_2;
      end else if (10'hb6 == _T_19[9:0]) begin
        image_0_182 <= io_pixelVal_in_0_1;
      end else if (10'hb6 == _T_15[9:0]) begin
        image_0_182 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_183 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hb7 == _T_37[9:0]) begin
        image_0_183 <= io_pixelVal_in_0_7;
      end else if (10'hb7 == _T_34[9:0]) begin
        image_0_183 <= io_pixelVal_in_0_6;
      end else if (10'hb7 == _T_31[9:0]) begin
        image_0_183 <= io_pixelVal_in_0_5;
      end else if (10'hb7 == _T_28[9:0]) begin
        image_0_183 <= io_pixelVal_in_0_4;
      end else if (10'hb7 == _T_25[9:0]) begin
        image_0_183 <= io_pixelVal_in_0_3;
      end else if (10'hb7 == _T_22[9:0]) begin
        image_0_183 <= io_pixelVal_in_0_2;
      end else if (10'hb7 == _T_19[9:0]) begin
        image_0_183 <= io_pixelVal_in_0_1;
      end else if (10'hb7 == _T_15[9:0]) begin
        image_0_183 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_184 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hb8 == _T_37[9:0]) begin
        image_0_184 <= io_pixelVal_in_0_7;
      end else if (10'hb8 == _T_34[9:0]) begin
        image_0_184 <= io_pixelVal_in_0_6;
      end else if (10'hb8 == _T_31[9:0]) begin
        image_0_184 <= io_pixelVal_in_0_5;
      end else if (10'hb8 == _T_28[9:0]) begin
        image_0_184 <= io_pixelVal_in_0_4;
      end else if (10'hb8 == _T_25[9:0]) begin
        image_0_184 <= io_pixelVal_in_0_3;
      end else if (10'hb8 == _T_22[9:0]) begin
        image_0_184 <= io_pixelVal_in_0_2;
      end else if (10'hb8 == _T_19[9:0]) begin
        image_0_184 <= io_pixelVal_in_0_1;
      end else if (10'hb8 == _T_15[9:0]) begin
        image_0_184 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_185 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hb9 == _T_37[9:0]) begin
        image_0_185 <= io_pixelVal_in_0_7;
      end else if (10'hb9 == _T_34[9:0]) begin
        image_0_185 <= io_pixelVal_in_0_6;
      end else if (10'hb9 == _T_31[9:0]) begin
        image_0_185 <= io_pixelVal_in_0_5;
      end else if (10'hb9 == _T_28[9:0]) begin
        image_0_185 <= io_pixelVal_in_0_4;
      end else if (10'hb9 == _T_25[9:0]) begin
        image_0_185 <= io_pixelVal_in_0_3;
      end else if (10'hb9 == _T_22[9:0]) begin
        image_0_185 <= io_pixelVal_in_0_2;
      end else if (10'hb9 == _T_19[9:0]) begin
        image_0_185 <= io_pixelVal_in_0_1;
      end else if (10'hb9 == _T_15[9:0]) begin
        image_0_185 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_186 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hba == _T_37[9:0]) begin
        image_0_186 <= io_pixelVal_in_0_7;
      end else if (10'hba == _T_34[9:0]) begin
        image_0_186 <= io_pixelVal_in_0_6;
      end else if (10'hba == _T_31[9:0]) begin
        image_0_186 <= io_pixelVal_in_0_5;
      end else if (10'hba == _T_28[9:0]) begin
        image_0_186 <= io_pixelVal_in_0_4;
      end else if (10'hba == _T_25[9:0]) begin
        image_0_186 <= io_pixelVal_in_0_3;
      end else if (10'hba == _T_22[9:0]) begin
        image_0_186 <= io_pixelVal_in_0_2;
      end else if (10'hba == _T_19[9:0]) begin
        image_0_186 <= io_pixelVal_in_0_1;
      end else if (10'hba == _T_15[9:0]) begin
        image_0_186 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_187 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hbb == _T_37[9:0]) begin
        image_0_187 <= io_pixelVal_in_0_7;
      end else if (10'hbb == _T_34[9:0]) begin
        image_0_187 <= io_pixelVal_in_0_6;
      end else if (10'hbb == _T_31[9:0]) begin
        image_0_187 <= io_pixelVal_in_0_5;
      end else if (10'hbb == _T_28[9:0]) begin
        image_0_187 <= io_pixelVal_in_0_4;
      end else if (10'hbb == _T_25[9:0]) begin
        image_0_187 <= io_pixelVal_in_0_3;
      end else if (10'hbb == _T_22[9:0]) begin
        image_0_187 <= io_pixelVal_in_0_2;
      end else if (10'hbb == _T_19[9:0]) begin
        image_0_187 <= io_pixelVal_in_0_1;
      end else if (10'hbb == _T_15[9:0]) begin
        image_0_187 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_188 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hbc == _T_37[9:0]) begin
        image_0_188 <= io_pixelVal_in_0_7;
      end else if (10'hbc == _T_34[9:0]) begin
        image_0_188 <= io_pixelVal_in_0_6;
      end else if (10'hbc == _T_31[9:0]) begin
        image_0_188 <= io_pixelVal_in_0_5;
      end else if (10'hbc == _T_28[9:0]) begin
        image_0_188 <= io_pixelVal_in_0_4;
      end else if (10'hbc == _T_25[9:0]) begin
        image_0_188 <= io_pixelVal_in_0_3;
      end else if (10'hbc == _T_22[9:0]) begin
        image_0_188 <= io_pixelVal_in_0_2;
      end else if (10'hbc == _T_19[9:0]) begin
        image_0_188 <= io_pixelVal_in_0_1;
      end else if (10'hbc == _T_15[9:0]) begin
        image_0_188 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_189 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hbd == _T_37[9:0]) begin
        image_0_189 <= io_pixelVal_in_0_7;
      end else if (10'hbd == _T_34[9:0]) begin
        image_0_189 <= io_pixelVal_in_0_6;
      end else if (10'hbd == _T_31[9:0]) begin
        image_0_189 <= io_pixelVal_in_0_5;
      end else if (10'hbd == _T_28[9:0]) begin
        image_0_189 <= io_pixelVal_in_0_4;
      end else if (10'hbd == _T_25[9:0]) begin
        image_0_189 <= io_pixelVal_in_0_3;
      end else if (10'hbd == _T_22[9:0]) begin
        image_0_189 <= io_pixelVal_in_0_2;
      end else if (10'hbd == _T_19[9:0]) begin
        image_0_189 <= io_pixelVal_in_0_1;
      end else if (10'hbd == _T_15[9:0]) begin
        image_0_189 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_190 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hbe == _T_37[9:0]) begin
        image_0_190 <= io_pixelVal_in_0_7;
      end else if (10'hbe == _T_34[9:0]) begin
        image_0_190 <= io_pixelVal_in_0_6;
      end else if (10'hbe == _T_31[9:0]) begin
        image_0_190 <= io_pixelVal_in_0_5;
      end else if (10'hbe == _T_28[9:0]) begin
        image_0_190 <= io_pixelVal_in_0_4;
      end else if (10'hbe == _T_25[9:0]) begin
        image_0_190 <= io_pixelVal_in_0_3;
      end else if (10'hbe == _T_22[9:0]) begin
        image_0_190 <= io_pixelVal_in_0_2;
      end else if (10'hbe == _T_19[9:0]) begin
        image_0_190 <= io_pixelVal_in_0_1;
      end else if (10'hbe == _T_15[9:0]) begin
        image_0_190 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_191 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hbf == _T_37[9:0]) begin
        image_0_191 <= io_pixelVal_in_0_7;
      end else if (10'hbf == _T_34[9:0]) begin
        image_0_191 <= io_pixelVal_in_0_6;
      end else if (10'hbf == _T_31[9:0]) begin
        image_0_191 <= io_pixelVal_in_0_5;
      end else if (10'hbf == _T_28[9:0]) begin
        image_0_191 <= io_pixelVal_in_0_4;
      end else if (10'hbf == _T_25[9:0]) begin
        image_0_191 <= io_pixelVal_in_0_3;
      end else if (10'hbf == _T_22[9:0]) begin
        image_0_191 <= io_pixelVal_in_0_2;
      end else if (10'hbf == _T_19[9:0]) begin
        image_0_191 <= io_pixelVal_in_0_1;
      end else if (10'hbf == _T_15[9:0]) begin
        image_0_191 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_192 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hc0 == _T_37[9:0]) begin
        image_0_192 <= io_pixelVal_in_0_7;
      end else if (10'hc0 == _T_34[9:0]) begin
        image_0_192 <= io_pixelVal_in_0_6;
      end else if (10'hc0 == _T_31[9:0]) begin
        image_0_192 <= io_pixelVal_in_0_5;
      end else if (10'hc0 == _T_28[9:0]) begin
        image_0_192 <= io_pixelVal_in_0_4;
      end else if (10'hc0 == _T_25[9:0]) begin
        image_0_192 <= io_pixelVal_in_0_3;
      end else if (10'hc0 == _T_22[9:0]) begin
        image_0_192 <= io_pixelVal_in_0_2;
      end else if (10'hc0 == _T_19[9:0]) begin
        image_0_192 <= io_pixelVal_in_0_1;
      end else if (10'hc0 == _T_15[9:0]) begin
        image_0_192 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_193 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hc1 == _T_37[9:0]) begin
        image_0_193 <= io_pixelVal_in_0_7;
      end else if (10'hc1 == _T_34[9:0]) begin
        image_0_193 <= io_pixelVal_in_0_6;
      end else if (10'hc1 == _T_31[9:0]) begin
        image_0_193 <= io_pixelVal_in_0_5;
      end else if (10'hc1 == _T_28[9:0]) begin
        image_0_193 <= io_pixelVal_in_0_4;
      end else if (10'hc1 == _T_25[9:0]) begin
        image_0_193 <= io_pixelVal_in_0_3;
      end else if (10'hc1 == _T_22[9:0]) begin
        image_0_193 <= io_pixelVal_in_0_2;
      end else if (10'hc1 == _T_19[9:0]) begin
        image_0_193 <= io_pixelVal_in_0_1;
      end else if (10'hc1 == _T_15[9:0]) begin
        image_0_193 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_194 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hc2 == _T_37[9:0]) begin
        image_0_194 <= io_pixelVal_in_0_7;
      end else if (10'hc2 == _T_34[9:0]) begin
        image_0_194 <= io_pixelVal_in_0_6;
      end else if (10'hc2 == _T_31[9:0]) begin
        image_0_194 <= io_pixelVal_in_0_5;
      end else if (10'hc2 == _T_28[9:0]) begin
        image_0_194 <= io_pixelVal_in_0_4;
      end else if (10'hc2 == _T_25[9:0]) begin
        image_0_194 <= io_pixelVal_in_0_3;
      end else if (10'hc2 == _T_22[9:0]) begin
        image_0_194 <= io_pixelVal_in_0_2;
      end else if (10'hc2 == _T_19[9:0]) begin
        image_0_194 <= io_pixelVal_in_0_1;
      end else if (10'hc2 == _T_15[9:0]) begin
        image_0_194 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_195 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hc3 == _T_37[9:0]) begin
        image_0_195 <= io_pixelVal_in_0_7;
      end else if (10'hc3 == _T_34[9:0]) begin
        image_0_195 <= io_pixelVal_in_0_6;
      end else if (10'hc3 == _T_31[9:0]) begin
        image_0_195 <= io_pixelVal_in_0_5;
      end else if (10'hc3 == _T_28[9:0]) begin
        image_0_195 <= io_pixelVal_in_0_4;
      end else if (10'hc3 == _T_25[9:0]) begin
        image_0_195 <= io_pixelVal_in_0_3;
      end else if (10'hc3 == _T_22[9:0]) begin
        image_0_195 <= io_pixelVal_in_0_2;
      end else if (10'hc3 == _T_19[9:0]) begin
        image_0_195 <= io_pixelVal_in_0_1;
      end else if (10'hc3 == _T_15[9:0]) begin
        image_0_195 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_196 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hc4 == _T_37[9:0]) begin
        image_0_196 <= io_pixelVal_in_0_7;
      end else if (10'hc4 == _T_34[9:0]) begin
        image_0_196 <= io_pixelVal_in_0_6;
      end else if (10'hc4 == _T_31[9:0]) begin
        image_0_196 <= io_pixelVal_in_0_5;
      end else if (10'hc4 == _T_28[9:0]) begin
        image_0_196 <= io_pixelVal_in_0_4;
      end else if (10'hc4 == _T_25[9:0]) begin
        image_0_196 <= io_pixelVal_in_0_3;
      end else if (10'hc4 == _T_22[9:0]) begin
        image_0_196 <= io_pixelVal_in_0_2;
      end else if (10'hc4 == _T_19[9:0]) begin
        image_0_196 <= io_pixelVal_in_0_1;
      end else if (10'hc4 == _T_15[9:0]) begin
        image_0_196 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_197 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hc5 == _T_37[9:0]) begin
        image_0_197 <= io_pixelVal_in_0_7;
      end else if (10'hc5 == _T_34[9:0]) begin
        image_0_197 <= io_pixelVal_in_0_6;
      end else if (10'hc5 == _T_31[9:0]) begin
        image_0_197 <= io_pixelVal_in_0_5;
      end else if (10'hc5 == _T_28[9:0]) begin
        image_0_197 <= io_pixelVal_in_0_4;
      end else if (10'hc5 == _T_25[9:0]) begin
        image_0_197 <= io_pixelVal_in_0_3;
      end else if (10'hc5 == _T_22[9:0]) begin
        image_0_197 <= io_pixelVal_in_0_2;
      end else if (10'hc5 == _T_19[9:0]) begin
        image_0_197 <= io_pixelVal_in_0_1;
      end else if (10'hc5 == _T_15[9:0]) begin
        image_0_197 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_198 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hc6 == _T_37[9:0]) begin
        image_0_198 <= io_pixelVal_in_0_7;
      end else if (10'hc6 == _T_34[9:0]) begin
        image_0_198 <= io_pixelVal_in_0_6;
      end else if (10'hc6 == _T_31[9:0]) begin
        image_0_198 <= io_pixelVal_in_0_5;
      end else if (10'hc6 == _T_28[9:0]) begin
        image_0_198 <= io_pixelVal_in_0_4;
      end else if (10'hc6 == _T_25[9:0]) begin
        image_0_198 <= io_pixelVal_in_0_3;
      end else if (10'hc6 == _T_22[9:0]) begin
        image_0_198 <= io_pixelVal_in_0_2;
      end else if (10'hc6 == _T_19[9:0]) begin
        image_0_198 <= io_pixelVal_in_0_1;
      end else if (10'hc6 == _T_15[9:0]) begin
        image_0_198 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_199 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hc7 == _T_37[9:0]) begin
        image_0_199 <= io_pixelVal_in_0_7;
      end else if (10'hc7 == _T_34[9:0]) begin
        image_0_199 <= io_pixelVal_in_0_6;
      end else if (10'hc7 == _T_31[9:0]) begin
        image_0_199 <= io_pixelVal_in_0_5;
      end else if (10'hc7 == _T_28[9:0]) begin
        image_0_199 <= io_pixelVal_in_0_4;
      end else if (10'hc7 == _T_25[9:0]) begin
        image_0_199 <= io_pixelVal_in_0_3;
      end else if (10'hc7 == _T_22[9:0]) begin
        image_0_199 <= io_pixelVal_in_0_2;
      end else if (10'hc7 == _T_19[9:0]) begin
        image_0_199 <= io_pixelVal_in_0_1;
      end else if (10'hc7 == _T_15[9:0]) begin
        image_0_199 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_200 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hc8 == _T_37[9:0]) begin
        image_0_200 <= io_pixelVal_in_0_7;
      end else if (10'hc8 == _T_34[9:0]) begin
        image_0_200 <= io_pixelVal_in_0_6;
      end else if (10'hc8 == _T_31[9:0]) begin
        image_0_200 <= io_pixelVal_in_0_5;
      end else if (10'hc8 == _T_28[9:0]) begin
        image_0_200 <= io_pixelVal_in_0_4;
      end else if (10'hc8 == _T_25[9:0]) begin
        image_0_200 <= io_pixelVal_in_0_3;
      end else if (10'hc8 == _T_22[9:0]) begin
        image_0_200 <= io_pixelVal_in_0_2;
      end else if (10'hc8 == _T_19[9:0]) begin
        image_0_200 <= io_pixelVal_in_0_1;
      end else if (10'hc8 == _T_15[9:0]) begin
        image_0_200 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_201 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hc9 == _T_37[9:0]) begin
        image_0_201 <= io_pixelVal_in_0_7;
      end else if (10'hc9 == _T_34[9:0]) begin
        image_0_201 <= io_pixelVal_in_0_6;
      end else if (10'hc9 == _T_31[9:0]) begin
        image_0_201 <= io_pixelVal_in_0_5;
      end else if (10'hc9 == _T_28[9:0]) begin
        image_0_201 <= io_pixelVal_in_0_4;
      end else if (10'hc9 == _T_25[9:0]) begin
        image_0_201 <= io_pixelVal_in_0_3;
      end else if (10'hc9 == _T_22[9:0]) begin
        image_0_201 <= io_pixelVal_in_0_2;
      end else if (10'hc9 == _T_19[9:0]) begin
        image_0_201 <= io_pixelVal_in_0_1;
      end else if (10'hc9 == _T_15[9:0]) begin
        image_0_201 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_202 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hca == _T_37[9:0]) begin
        image_0_202 <= io_pixelVal_in_0_7;
      end else if (10'hca == _T_34[9:0]) begin
        image_0_202 <= io_pixelVal_in_0_6;
      end else if (10'hca == _T_31[9:0]) begin
        image_0_202 <= io_pixelVal_in_0_5;
      end else if (10'hca == _T_28[9:0]) begin
        image_0_202 <= io_pixelVal_in_0_4;
      end else if (10'hca == _T_25[9:0]) begin
        image_0_202 <= io_pixelVal_in_0_3;
      end else if (10'hca == _T_22[9:0]) begin
        image_0_202 <= io_pixelVal_in_0_2;
      end else if (10'hca == _T_19[9:0]) begin
        image_0_202 <= io_pixelVal_in_0_1;
      end else if (10'hca == _T_15[9:0]) begin
        image_0_202 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_203 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hcb == _T_37[9:0]) begin
        image_0_203 <= io_pixelVal_in_0_7;
      end else if (10'hcb == _T_34[9:0]) begin
        image_0_203 <= io_pixelVal_in_0_6;
      end else if (10'hcb == _T_31[9:0]) begin
        image_0_203 <= io_pixelVal_in_0_5;
      end else if (10'hcb == _T_28[9:0]) begin
        image_0_203 <= io_pixelVal_in_0_4;
      end else if (10'hcb == _T_25[9:0]) begin
        image_0_203 <= io_pixelVal_in_0_3;
      end else if (10'hcb == _T_22[9:0]) begin
        image_0_203 <= io_pixelVal_in_0_2;
      end else if (10'hcb == _T_19[9:0]) begin
        image_0_203 <= io_pixelVal_in_0_1;
      end else if (10'hcb == _T_15[9:0]) begin
        image_0_203 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_204 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hcc == _T_37[9:0]) begin
        image_0_204 <= io_pixelVal_in_0_7;
      end else if (10'hcc == _T_34[9:0]) begin
        image_0_204 <= io_pixelVal_in_0_6;
      end else if (10'hcc == _T_31[9:0]) begin
        image_0_204 <= io_pixelVal_in_0_5;
      end else if (10'hcc == _T_28[9:0]) begin
        image_0_204 <= io_pixelVal_in_0_4;
      end else if (10'hcc == _T_25[9:0]) begin
        image_0_204 <= io_pixelVal_in_0_3;
      end else if (10'hcc == _T_22[9:0]) begin
        image_0_204 <= io_pixelVal_in_0_2;
      end else if (10'hcc == _T_19[9:0]) begin
        image_0_204 <= io_pixelVal_in_0_1;
      end else if (10'hcc == _T_15[9:0]) begin
        image_0_204 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_205 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hcd == _T_37[9:0]) begin
        image_0_205 <= io_pixelVal_in_0_7;
      end else if (10'hcd == _T_34[9:0]) begin
        image_0_205 <= io_pixelVal_in_0_6;
      end else if (10'hcd == _T_31[9:0]) begin
        image_0_205 <= io_pixelVal_in_0_5;
      end else if (10'hcd == _T_28[9:0]) begin
        image_0_205 <= io_pixelVal_in_0_4;
      end else if (10'hcd == _T_25[9:0]) begin
        image_0_205 <= io_pixelVal_in_0_3;
      end else if (10'hcd == _T_22[9:0]) begin
        image_0_205 <= io_pixelVal_in_0_2;
      end else if (10'hcd == _T_19[9:0]) begin
        image_0_205 <= io_pixelVal_in_0_1;
      end else if (10'hcd == _T_15[9:0]) begin
        image_0_205 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_206 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hce == _T_37[9:0]) begin
        image_0_206 <= io_pixelVal_in_0_7;
      end else if (10'hce == _T_34[9:0]) begin
        image_0_206 <= io_pixelVal_in_0_6;
      end else if (10'hce == _T_31[9:0]) begin
        image_0_206 <= io_pixelVal_in_0_5;
      end else if (10'hce == _T_28[9:0]) begin
        image_0_206 <= io_pixelVal_in_0_4;
      end else if (10'hce == _T_25[9:0]) begin
        image_0_206 <= io_pixelVal_in_0_3;
      end else if (10'hce == _T_22[9:0]) begin
        image_0_206 <= io_pixelVal_in_0_2;
      end else if (10'hce == _T_19[9:0]) begin
        image_0_206 <= io_pixelVal_in_0_1;
      end else if (10'hce == _T_15[9:0]) begin
        image_0_206 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_207 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hcf == _T_37[9:0]) begin
        image_0_207 <= io_pixelVal_in_0_7;
      end else if (10'hcf == _T_34[9:0]) begin
        image_0_207 <= io_pixelVal_in_0_6;
      end else if (10'hcf == _T_31[9:0]) begin
        image_0_207 <= io_pixelVal_in_0_5;
      end else if (10'hcf == _T_28[9:0]) begin
        image_0_207 <= io_pixelVal_in_0_4;
      end else if (10'hcf == _T_25[9:0]) begin
        image_0_207 <= io_pixelVal_in_0_3;
      end else if (10'hcf == _T_22[9:0]) begin
        image_0_207 <= io_pixelVal_in_0_2;
      end else if (10'hcf == _T_19[9:0]) begin
        image_0_207 <= io_pixelVal_in_0_1;
      end else if (10'hcf == _T_15[9:0]) begin
        image_0_207 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_208 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hd0 == _T_37[9:0]) begin
        image_0_208 <= io_pixelVal_in_0_7;
      end else if (10'hd0 == _T_34[9:0]) begin
        image_0_208 <= io_pixelVal_in_0_6;
      end else if (10'hd0 == _T_31[9:0]) begin
        image_0_208 <= io_pixelVal_in_0_5;
      end else if (10'hd0 == _T_28[9:0]) begin
        image_0_208 <= io_pixelVal_in_0_4;
      end else if (10'hd0 == _T_25[9:0]) begin
        image_0_208 <= io_pixelVal_in_0_3;
      end else if (10'hd0 == _T_22[9:0]) begin
        image_0_208 <= io_pixelVal_in_0_2;
      end else if (10'hd0 == _T_19[9:0]) begin
        image_0_208 <= io_pixelVal_in_0_1;
      end else if (10'hd0 == _T_15[9:0]) begin
        image_0_208 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_209 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hd1 == _T_37[9:0]) begin
        image_0_209 <= io_pixelVal_in_0_7;
      end else if (10'hd1 == _T_34[9:0]) begin
        image_0_209 <= io_pixelVal_in_0_6;
      end else if (10'hd1 == _T_31[9:0]) begin
        image_0_209 <= io_pixelVal_in_0_5;
      end else if (10'hd1 == _T_28[9:0]) begin
        image_0_209 <= io_pixelVal_in_0_4;
      end else if (10'hd1 == _T_25[9:0]) begin
        image_0_209 <= io_pixelVal_in_0_3;
      end else if (10'hd1 == _T_22[9:0]) begin
        image_0_209 <= io_pixelVal_in_0_2;
      end else if (10'hd1 == _T_19[9:0]) begin
        image_0_209 <= io_pixelVal_in_0_1;
      end else if (10'hd1 == _T_15[9:0]) begin
        image_0_209 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_210 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hd2 == _T_37[9:0]) begin
        image_0_210 <= io_pixelVal_in_0_7;
      end else if (10'hd2 == _T_34[9:0]) begin
        image_0_210 <= io_pixelVal_in_0_6;
      end else if (10'hd2 == _T_31[9:0]) begin
        image_0_210 <= io_pixelVal_in_0_5;
      end else if (10'hd2 == _T_28[9:0]) begin
        image_0_210 <= io_pixelVal_in_0_4;
      end else if (10'hd2 == _T_25[9:0]) begin
        image_0_210 <= io_pixelVal_in_0_3;
      end else if (10'hd2 == _T_22[9:0]) begin
        image_0_210 <= io_pixelVal_in_0_2;
      end else if (10'hd2 == _T_19[9:0]) begin
        image_0_210 <= io_pixelVal_in_0_1;
      end else if (10'hd2 == _T_15[9:0]) begin
        image_0_210 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_211 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hd3 == _T_37[9:0]) begin
        image_0_211 <= io_pixelVal_in_0_7;
      end else if (10'hd3 == _T_34[9:0]) begin
        image_0_211 <= io_pixelVal_in_0_6;
      end else if (10'hd3 == _T_31[9:0]) begin
        image_0_211 <= io_pixelVal_in_0_5;
      end else if (10'hd3 == _T_28[9:0]) begin
        image_0_211 <= io_pixelVal_in_0_4;
      end else if (10'hd3 == _T_25[9:0]) begin
        image_0_211 <= io_pixelVal_in_0_3;
      end else if (10'hd3 == _T_22[9:0]) begin
        image_0_211 <= io_pixelVal_in_0_2;
      end else if (10'hd3 == _T_19[9:0]) begin
        image_0_211 <= io_pixelVal_in_0_1;
      end else if (10'hd3 == _T_15[9:0]) begin
        image_0_211 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_212 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hd4 == _T_37[9:0]) begin
        image_0_212 <= io_pixelVal_in_0_7;
      end else if (10'hd4 == _T_34[9:0]) begin
        image_0_212 <= io_pixelVal_in_0_6;
      end else if (10'hd4 == _T_31[9:0]) begin
        image_0_212 <= io_pixelVal_in_0_5;
      end else if (10'hd4 == _T_28[9:0]) begin
        image_0_212 <= io_pixelVal_in_0_4;
      end else if (10'hd4 == _T_25[9:0]) begin
        image_0_212 <= io_pixelVal_in_0_3;
      end else if (10'hd4 == _T_22[9:0]) begin
        image_0_212 <= io_pixelVal_in_0_2;
      end else if (10'hd4 == _T_19[9:0]) begin
        image_0_212 <= io_pixelVal_in_0_1;
      end else if (10'hd4 == _T_15[9:0]) begin
        image_0_212 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_213 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hd5 == _T_37[9:0]) begin
        image_0_213 <= io_pixelVal_in_0_7;
      end else if (10'hd5 == _T_34[9:0]) begin
        image_0_213 <= io_pixelVal_in_0_6;
      end else if (10'hd5 == _T_31[9:0]) begin
        image_0_213 <= io_pixelVal_in_0_5;
      end else if (10'hd5 == _T_28[9:0]) begin
        image_0_213 <= io_pixelVal_in_0_4;
      end else if (10'hd5 == _T_25[9:0]) begin
        image_0_213 <= io_pixelVal_in_0_3;
      end else if (10'hd5 == _T_22[9:0]) begin
        image_0_213 <= io_pixelVal_in_0_2;
      end else if (10'hd5 == _T_19[9:0]) begin
        image_0_213 <= io_pixelVal_in_0_1;
      end else if (10'hd5 == _T_15[9:0]) begin
        image_0_213 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_214 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hd6 == _T_37[9:0]) begin
        image_0_214 <= io_pixelVal_in_0_7;
      end else if (10'hd6 == _T_34[9:0]) begin
        image_0_214 <= io_pixelVal_in_0_6;
      end else if (10'hd6 == _T_31[9:0]) begin
        image_0_214 <= io_pixelVal_in_0_5;
      end else if (10'hd6 == _T_28[9:0]) begin
        image_0_214 <= io_pixelVal_in_0_4;
      end else if (10'hd6 == _T_25[9:0]) begin
        image_0_214 <= io_pixelVal_in_0_3;
      end else if (10'hd6 == _T_22[9:0]) begin
        image_0_214 <= io_pixelVal_in_0_2;
      end else if (10'hd6 == _T_19[9:0]) begin
        image_0_214 <= io_pixelVal_in_0_1;
      end else if (10'hd6 == _T_15[9:0]) begin
        image_0_214 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_215 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hd7 == _T_37[9:0]) begin
        image_0_215 <= io_pixelVal_in_0_7;
      end else if (10'hd7 == _T_34[9:0]) begin
        image_0_215 <= io_pixelVal_in_0_6;
      end else if (10'hd7 == _T_31[9:0]) begin
        image_0_215 <= io_pixelVal_in_0_5;
      end else if (10'hd7 == _T_28[9:0]) begin
        image_0_215 <= io_pixelVal_in_0_4;
      end else if (10'hd7 == _T_25[9:0]) begin
        image_0_215 <= io_pixelVal_in_0_3;
      end else if (10'hd7 == _T_22[9:0]) begin
        image_0_215 <= io_pixelVal_in_0_2;
      end else if (10'hd7 == _T_19[9:0]) begin
        image_0_215 <= io_pixelVal_in_0_1;
      end else if (10'hd7 == _T_15[9:0]) begin
        image_0_215 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_216 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hd8 == _T_37[9:0]) begin
        image_0_216 <= io_pixelVal_in_0_7;
      end else if (10'hd8 == _T_34[9:0]) begin
        image_0_216 <= io_pixelVal_in_0_6;
      end else if (10'hd8 == _T_31[9:0]) begin
        image_0_216 <= io_pixelVal_in_0_5;
      end else if (10'hd8 == _T_28[9:0]) begin
        image_0_216 <= io_pixelVal_in_0_4;
      end else if (10'hd8 == _T_25[9:0]) begin
        image_0_216 <= io_pixelVal_in_0_3;
      end else if (10'hd8 == _T_22[9:0]) begin
        image_0_216 <= io_pixelVal_in_0_2;
      end else if (10'hd8 == _T_19[9:0]) begin
        image_0_216 <= io_pixelVal_in_0_1;
      end else if (10'hd8 == _T_15[9:0]) begin
        image_0_216 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_217 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hd9 == _T_37[9:0]) begin
        image_0_217 <= io_pixelVal_in_0_7;
      end else if (10'hd9 == _T_34[9:0]) begin
        image_0_217 <= io_pixelVal_in_0_6;
      end else if (10'hd9 == _T_31[9:0]) begin
        image_0_217 <= io_pixelVal_in_0_5;
      end else if (10'hd9 == _T_28[9:0]) begin
        image_0_217 <= io_pixelVal_in_0_4;
      end else if (10'hd9 == _T_25[9:0]) begin
        image_0_217 <= io_pixelVal_in_0_3;
      end else if (10'hd9 == _T_22[9:0]) begin
        image_0_217 <= io_pixelVal_in_0_2;
      end else if (10'hd9 == _T_19[9:0]) begin
        image_0_217 <= io_pixelVal_in_0_1;
      end else if (10'hd9 == _T_15[9:0]) begin
        image_0_217 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_218 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hda == _T_37[9:0]) begin
        image_0_218 <= io_pixelVal_in_0_7;
      end else if (10'hda == _T_34[9:0]) begin
        image_0_218 <= io_pixelVal_in_0_6;
      end else if (10'hda == _T_31[9:0]) begin
        image_0_218 <= io_pixelVal_in_0_5;
      end else if (10'hda == _T_28[9:0]) begin
        image_0_218 <= io_pixelVal_in_0_4;
      end else if (10'hda == _T_25[9:0]) begin
        image_0_218 <= io_pixelVal_in_0_3;
      end else if (10'hda == _T_22[9:0]) begin
        image_0_218 <= io_pixelVal_in_0_2;
      end else if (10'hda == _T_19[9:0]) begin
        image_0_218 <= io_pixelVal_in_0_1;
      end else if (10'hda == _T_15[9:0]) begin
        image_0_218 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_219 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hdb == _T_37[9:0]) begin
        image_0_219 <= io_pixelVal_in_0_7;
      end else if (10'hdb == _T_34[9:0]) begin
        image_0_219 <= io_pixelVal_in_0_6;
      end else if (10'hdb == _T_31[9:0]) begin
        image_0_219 <= io_pixelVal_in_0_5;
      end else if (10'hdb == _T_28[9:0]) begin
        image_0_219 <= io_pixelVal_in_0_4;
      end else if (10'hdb == _T_25[9:0]) begin
        image_0_219 <= io_pixelVal_in_0_3;
      end else if (10'hdb == _T_22[9:0]) begin
        image_0_219 <= io_pixelVal_in_0_2;
      end else if (10'hdb == _T_19[9:0]) begin
        image_0_219 <= io_pixelVal_in_0_1;
      end else if (10'hdb == _T_15[9:0]) begin
        image_0_219 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_220 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hdc == _T_37[9:0]) begin
        image_0_220 <= io_pixelVal_in_0_7;
      end else if (10'hdc == _T_34[9:0]) begin
        image_0_220 <= io_pixelVal_in_0_6;
      end else if (10'hdc == _T_31[9:0]) begin
        image_0_220 <= io_pixelVal_in_0_5;
      end else if (10'hdc == _T_28[9:0]) begin
        image_0_220 <= io_pixelVal_in_0_4;
      end else if (10'hdc == _T_25[9:0]) begin
        image_0_220 <= io_pixelVal_in_0_3;
      end else if (10'hdc == _T_22[9:0]) begin
        image_0_220 <= io_pixelVal_in_0_2;
      end else if (10'hdc == _T_19[9:0]) begin
        image_0_220 <= io_pixelVal_in_0_1;
      end else if (10'hdc == _T_15[9:0]) begin
        image_0_220 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_221 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hdd == _T_37[9:0]) begin
        image_0_221 <= io_pixelVal_in_0_7;
      end else if (10'hdd == _T_34[9:0]) begin
        image_0_221 <= io_pixelVal_in_0_6;
      end else if (10'hdd == _T_31[9:0]) begin
        image_0_221 <= io_pixelVal_in_0_5;
      end else if (10'hdd == _T_28[9:0]) begin
        image_0_221 <= io_pixelVal_in_0_4;
      end else if (10'hdd == _T_25[9:0]) begin
        image_0_221 <= io_pixelVal_in_0_3;
      end else if (10'hdd == _T_22[9:0]) begin
        image_0_221 <= io_pixelVal_in_0_2;
      end else if (10'hdd == _T_19[9:0]) begin
        image_0_221 <= io_pixelVal_in_0_1;
      end else if (10'hdd == _T_15[9:0]) begin
        image_0_221 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_222 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hde == _T_37[9:0]) begin
        image_0_222 <= io_pixelVal_in_0_7;
      end else if (10'hde == _T_34[9:0]) begin
        image_0_222 <= io_pixelVal_in_0_6;
      end else if (10'hde == _T_31[9:0]) begin
        image_0_222 <= io_pixelVal_in_0_5;
      end else if (10'hde == _T_28[9:0]) begin
        image_0_222 <= io_pixelVal_in_0_4;
      end else if (10'hde == _T_25[9:0]) begin
        image_0_222 <= io_pixelVal_in_0_3;
      end else if (10'hde == _T_22[9:0]) begin
        image_0_222 <= io_pixelVal_in_0_2;
      end else if (10'hde == _T_19[9:0]) begin
        image_0_222 <= io_pixelVal_in_0_1;
      end else if (10'hde == _T_15[9:0]) begin
        image_0_222 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_223 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hdf == _T_37[9:0]) begin
        image_0_223 <= io_pixelVal_in_0_7;
      end else if (10'hdf == _T_34[9:0]) begin
        image_0_223 <= io_pixelVal_in_0_6;
      end else if (10'hdf == _T_31[9:0]) begin
        image_0_223 <= io_pixelVal_in_0_5;
      end else if (10'hdf == _T_28[9:0]) begin
        image_0_223 <= io_pixelVal_in_0_4;
      end else if (10'hdf == _T_25[9:0]) begin
        image_0_223 <= io_pixelVal_in_0_3;
      end else if (10'hdf == _T_22[9:0]) begin
        image_0_223 <= io_pixelVal_in_0_2;
      end else if (10'hdf == _T_19[9:0]) begin
        image_0_223 <= io_pixelVal_in_0_1;
      end else if (10'hdf == _T_15[9:0]) begin
        image_0_223 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_224 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'he0 == _T_37[9:0]) begin
        image_0_224 <= io_pixelVal_in_0_7;
      end else if (10'he0 == _T_34[9:0]) begin
        image_0_224 <= io_pixelVal_in_0_6;
      end else if (10'he0 == _T_31[9:0]) begin
        image_0_224 <= io_pixelVal_in_0_5;
      end else if (10'he0 == _T_28[9:0]) begin
        image_0_224 <= io_pixelVal_in_0_4;
      end else if (10'he0 == _T_25[9:0]) begin
        image_0_224 <= io_pixelVal_in_0_3;
      end else if (10'he0 == _T_22[9:0]) begin
        image_0_224 <= io_pixelVal_in_0_2;
      end else if (10'he0 == _T_19[9:0]) begin
        image_0_224 <= io_pixelVal_in_0_1;
      end else if (10'he0 == _T_15[9:0]) begin
        image_0_224 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_225 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'he1 == _T_37[9:0]) begin
        image_0_225 <= io_pixelVal_in_0_7;
      end else if (10'he1 == _T_34[9:0]) begin
        image_0_225 <= io_pixelVal_in_0_6;
      end else if (10'he1 == _T_31[9:0]) begin
        image_0_225 <= io_pixelVal_in_0_5;
      end else if (10'he1 == _T_28[9:0]) begin
        image_0_225 <= io_pixelVal_in_0_4;
      end else if (10'he1 == _T_25[9:0]) begin
        image_0_225 <= io_pixelVal_in_0_3;
      end else if (10'he1 == _T_22[9:0]) begin
        image_0_225 <= io_pixelVal_in_0_2;
      end else if (10'he1 == _T_19[9:0]) begin
        image_0_225 <= io_pixelVal_in_0_1;
      end else if (10'he1 == _T_15[9:0]) begin
        image_0_225 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_226 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'he2 == _T_37[9:0]) begin
        image_0_226 <= io_pixelVal_in_0_7;
      end else if (10'he2 == _T_34[9:0]) begin
        image_0_226 <= io_pixelVal_in_0_6;
      end else if (10'he2 == _T_31[9:0]) begin
        image_0_226 <= io_pixelVal_in_0_5;
      end else if (10'he2 == _T_28[9:0]) begin
        image_0_226 <= io_pixelVal_in_0_4;
      end else if (10'he2 == _T_25[9:0]) begin
        image_0_226 <= io_pixelVal_in_0_3;
      end else if (10'he2 == _T_22[9:0]) begin
        image_0_226 <= io_pixelVal_in_0_2;
      end else if (10'he2 == _T_19[9:0]) begin
        image_0_226 <= io_pixelVal_in_0_1;
      end else if (10'he2 == _T_15[9:0]) begin
        image_0_226 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_227 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'he3 == _T_37[9:0]) begin
        image_0_227 <= io_pixelVal_in_0_7;
      end else if (10'he3 == _T_34[9:0]) begin
        image_0_227 <= io_pixelVal_in_0_6;
      end else if (10'he3 == _T_31[9:0]) begin
        image_0_227 <= io_pixelVal_in_0_5;
      end else if (10'he3 == _T_28[9:0]) begin
        image_0_227 <= io_pixelVal_in_0_4;
      end else if (10'he3 == _T_25[9:0]) begin
        image_0_227 <= io_pixelVal_in_0_3;
      end else if (10'he3 == _T_22[9:0]) begin
        image_0_227 <= io_pixelVal_in_0_2;
      end else if (10'he3 == _T_19[9:0]) begin
        image_0_227 <= io_pixelVal_in_0_1;
      end else if (10'he3 == _T_15[9:0]) begin
        image_0_227 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_228 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'he4 == _T_37[9:0]) begin
        image_0_228 <= io_pixelVal_in_0_7;
      end else if (10'he4 == _T_34[9:0]) begin
        image_0_228 <= io_pixelVal_in_0_6;
      end else if (10'he4 == _T_31[9:0]) begin
        image_0_228 <= io_pixelVal_in_0_5;
      end else if (10'he4 == _T_28[9:0]) begin
        image_0_228 <= io_pixelVal_in_0_4;
      end else if (10'he4 == _T_25[9:0]) begin
        image_0_228 <= io_pixelVal_in_0_3;
      end else if (10'he4 == _T_22[9:0]) begin
        image_0_228 <= io_pixelVal_in_0_2;
      end else if (10'he4 == _T_19[9:0]) begin
        image_0_228 <= io_pixelVal_in_0_1;
      end else if (10'he4 == _T_15[9:0]) begin
        image_0_228 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_229 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'he5 == _T_37[9:0]) begin
        image_0_229 <= io_pixelVal_in_0_7;
      end else if (10'he5 == _T_34[9:0]) begin
        image_0_229 <= io_pixelVal_in_0_6;
      end else if (10'he5 == _T_31[9:0]) begin
        image_0_229 <= io_pixelVal_in_0_5;
      end else if (10'he5 == _T_28[9:0]) begin
        image_0_229 <= io_pixelVal_in_0_4;
      end else if (10'he5 == _T_25[9:0]) begin
        image_0_229 <= io_pixelVal_in_0_3;
      end else if (10'he5 == _T_22[9:0]) begin
        image_0_229 <= io_pixelVal_in_0_2;
      end else if (10'he5 == _T_19[9:0]) begin
        image_0_229 <= io_pixelVal_in_0_1;
      end else if (10'he5 == _T_15[9:0]) begin
        image_0_229 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_230 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'he6 == _T_37[9:0]) begin
        image_0_230 <= io_pixelVal_in_0_7;
      end else if (10'he6 == _T_34[9:0]) begin
        image_0_230 <= io_pixelVal_in_0_6;
      end else if (10'he6 == _T_31[9:0]) begin
        image_0_230 <= io_pixelVal_in_0_5;
      end else if (10'he6 == _T_28[9:0]) begin
        image_0_230 <= io_pixelVal_in_0_4;
      end else if (10'he6 == _T_25[9:0]) begin
        image_0_230 <= io_pixelVal_in_0_3;
      end else if (10'he6 == _T_22[9:0]) begin
        image_0_230 <= io_pixelVal_in_0_2;
      end else if (10'he6 == _T_19[9:0]) begin
        image_0_230 <= io_pixelVal_in_0_1;
      end else if (10'he6 == _T_15[9:0]) begin
        image_0_230 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_231 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'he7 == _T_37[9:0]) begin
        image_0_231 <= io_pixelVal_in_0_7;
      end else if (10'he7 == _T_34[9:0]) begin
        image_0_231 <= io_pixelVal_in_0_6;
      end else if (10'he7 == _T_31[9:0]) begin
        image_0_231 <= io_pixelVal_in_0_5;
      end else if (10'he7 == _T_28[9:0]) begin
        image_0_231 <= io_pixelVal_in_0_4;
      end else if (10'he7 == _T_25[9:0]) begin
        image_0_231 <= io_pixelVal_in_0_3;
      end else if (10'he7 == _T_22[9:0]) begin
        image_0_231 <= io_pixelVal_in_0_2;
      end else if (10'he7 == _T_19[9:0]) begin
        image_0_231 <= io_pixelVal_in_0_1;
      end else if (10'he7 == _T_15[9:0]) begin
        image_0_231 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_232 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'he8 == _T_37[9:0]) begin
        image_0_232 <= io_pixelVal_in_0_7;
      end else if (10'he8 == _T_34[9:0]) begin
        image_0_232 <= io_pixelVal_in_0_6;
      end else if (10'he8 == _T_31[9:0]) begin
        image_0_232 <= io_pixelVal_in_0_5;
      end else if (10'he8 == _T_28[9:0]) begin
        image_0_232 <= io_pixelVal_in_0_4;
      end else if (10'he8 == _T_25[9:0]) begin
        image_0_232 <= io_pixelVal_in_0_3;
      end else if (10'he8 == _T_22[9:0]) begin
        image_0_232 <= io_pixelVal_in_0_2;
      end else if (10'he8 == _T_19[9:0]) begin
        image_0_232 <= io_pixelVal_in_0_1;
      end else if (10'he8 == _T_15[9:0]) begin
        image_0_232 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_233 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'he9 == _T_37[9:0]) begin
        image_0_233 <= io_pixelVal_in_0_7;
      end else if (10'he9 == _T_34[9:0]) begin
        image_0_233 <= io_pixelVal_in_0_6;
      end else if (10'he9 == _T_31[9:0]) begin
        image_0_233 <= io_pixelVal_in_0_5;
      end else if (10'he9 == _T_28[9:0]) begin
        image_0_233 <= io_pixelVal_in_0_4;
      end else if (10'he9 == _T_25[9:0]) begin
        image_0_233 <= io_pixelVal_in_0_3;
      end else if (10'he9 == _T_22[9:0]) begin
        image_0_233 <= io_pixelVal_in_0_2;
      end else if (10'he9 == _T_19[9:0]) begin
        image_0_233 <= io_pixelVal_in_0_1;
      end else if (10'he9 == _T_15[9:0]) begin
        image_0_233 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_234 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hea == _T_37[9:0]) begin
        image_0_234 <= io_pixelVal_in_0_7;
      end else if (10'hea == _T_34[9:0]) begin
        image_0_234 <= io_pixelVal_in_0_6;
      end else if (10'hea == _T_31[9:0]) begin
        image_0_234 <= io_pixelVal_in_0_5;
      end else if (10'hea == _T_28[9:0]) begin
        image_0_234 <= io_pixelVal_in_0_4;
      end else if (10'hea == _T_25[9:0]) begin
        image_0_234 <= io_pixelVal_in_0_3;
      end else if (10'hea == _T_22[9:0]) begin
        image_0_234 <= io_pixelVal_in_0_2;
      end else if (10'hea == _T_19[9:0]) begin
        image_0_234 <= io_pixelVal_in_0_1;
      end else if (10'hea == _T_15[9:0]) begin
        image_0_234 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_235 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'heb == _T_37[9:0]) begin
        image_0_235 <= io_pixelVal_in_0_7;
      end else if (10'heb == _T_34[9:0]) begin
        image_0_235 <= io_pixelVal_in_0_6;
      end else if (10'heb == _T_31[9:0]) begin
        image_0_235 <= io_pixelVal_in_0_5;
      end else if (10'heb == _T_28[9:0]) begin
        image_0_235 <= io_pixelVal_in_0_4;
      end else if (10'heb == _T_25[9:0]) begin
        image_0_235 <= io_pixelVal_in_0_3;
      end else if (10'heb == _T_22[9:0]) begin
        image_0_235 <= io_pixelVal_in_0_2;
      end else if (10'heb == _T_19[9:0]) begin
        image_0_235 <= io_pixelVal_in_0_1;
      end else if (10'heb == _T_15[9:0]) begin
        image_0_235 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_236 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hec == _T_37[9:0]) begin
        image_0_236 <= io_pixelVal_in_0_7;
      end else if (10'hec == _T_34[9:0]) begin
        image_0_236 <= io_pixelVal_in_0_6;
      end else if (10'hec == _T_31[9:0]) begin
        image_0_236 <= io_pixelVal_in_0_5;
      end else if (10'hec == _T_28[9:0]) begin
        image_0_236 <= io_pixelVal_in_0_4;
      end else if (10'hec == _T_25[9:0]) begin
        image_0_236 <= io_pixelVal_in_0_3;
      end else if (10'hec == _T_22[9:0]) begin
        image_0_236 <= io_pixelVal_in_0_2;
      end else if (10'hec == _T_19[9:0]) begin
        image_0_236 <= io_pixelVal_in_0_1;
      end else if (10'hec == _T_15[9:0]) begin
        image_0_236 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_237 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hed == _T_37[9:0]) begin
        image_0_237 <= io_pixelVal_in_0_7;
      end else if (10'hed == _T_34[9:0]) begin
        image_0_237 <= io_pixelVal_in_0_6;
      end else if (10'hed == _T_31[9:0]) begin
        image_0_237 <= io_pixelVal_in_0_5;
      end else if (10'hed == _T_28[9:0]) begin
        image_0_237 <= io_pixelVal_in_0_4;
      end else if (10'hed == _T_25[9:0]) begin
        image_0_237 <= io_pixelVal_in_0_3;
      end else if (10'hed == _T_22[9:0]) begin
        image_0_237 <= io_pixelVal_in_0_2;
      end else if (10'hed == _T_19[9:0]) begin
        image_0_237 <= io_pixelVal_in_0_1;
      end else if (10'hed == _T_15[9:0]) begin
        image_0_237 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_238 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hee == _T_37[9:0]) begin
        image_0_238 <= io_pixelVal_in_0_7;
      end else if (10'hee == _T_34[9:0]) begin
        image_0_238 <= io_pixelVal_in_0_6;
      end else if (10'hee == _T_31[9:0]) begin
        image_0_238 <= io_pixelVal_in_0_5;
      end else if (10'hee == _T_28[9:0]) begin
        image_0_238 <= io_pixelVal_in_0_4;
      end else if (10'hee == _T_25[9:0]) begin
        image_0_238 <= io_pixelVal_in_0_3;
      end else if (10'hee == _T_22[9:0]) begin
        image_0_238 <= io_pixelVal_in_0_2;
      end else if (10'hee == _T_19[9:0]) begin
        image_0_238 <= io_pixelVal_in_0_1;
      end else if (10'hee == _T_15[9:0]) begin
        image_0_238 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_239 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hef == _T_37[9:0]) begin
        image_0_239 <= io_pixelVal_in_0_7;
      end else if (10'hef == _T_34[9:0]) begin
        image_0_239 <= io_pixelVal_in_0_6;
      end else if (10'hef == _T_31[9:0]) begin
        image_0_239 <= io_pixelVal_in_0_5;
      end else if (10'hef == _T_28[9:0]) begin
        image_0_239 <= io_pixelVal_in_0_4;
      end else if (10'hef == _T_25[9:0]) begin
        image_0_239 <= io_pixelVal_in_0_3;
      end else if (10'hef == _T_22[9:0]) begin
        image_0_239 <= io_pixelVal_in_0_2;
      end else if (10'hef == _T_19[9:0]) begin
        image_0_239 <= io_pixelVal_in_0_1;
      end else if (10'hef == _T_15[9:0]) begin
        image_0_239 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_240 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hf0 == _T_37[9:0]) begin
        image_0_240 <= io_pixelVal_in_0_7;
      end else if (10'hf0 == _T_34[9:0]) begin
        image_0_240 <= io_pixelVal_in_0_6;
      end else if (10'hf0 == _T_31[9:0]) begin
        image_0_240 <= io_pixelVal_in_0_5;
      end else if (10'hf0 == _T_28[9:0]) begin
        image_0_240 <= io_pixelVal_in_0_4;
      end else if (10'hf0 == _T_25[9:0]) begin
        image_0_240 <= io_pixelVal_in_0_3;
      end else if (10'hf0 == _T_22[9:0]) begin
        image_0_240 <= io_pixelVal_in_0_2;
      end else if (10'hf0 == _T_19[9:0]) begin
        image_0_240 <= io_pixelVal_in_0_1;
      end else if (10'hf0 == _T_15[9:0]) begin
        image_0_240 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_241 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hf1 == _T_37[9:0]) begin
        image_0_241 <= io_pixelVal_in_0_7;
      end else if (10'hf1 == _T_34[9:0]) begin
        image_0_241 <= io_pixelVal_in_0_6;
      end else if (10'hf1 == _T_31[9:0]) begin
        image_0_241 <= io_pixelVal_in_0_5;
      end else if (10'hf1 == _T_28[9:0]) begin
        image_0_241 <= io_pixelVal_in_0_4;
      end else if (10'hf1 == _T_25[9:0]) begin
        image_0_241 <= io_pixelVal_in_0_3;
      end else if (10'hf1 == _T_22[9:0]) begin
        image_0_241 <= io_pixelVal_in_0_2;
      end else if (10'hf1 == _T_19[9:0]) begin
        image_0_241 <= io_pixelVal_in_0_1;
      end else if (10'hf1 == _T_15[9:0]) begin
        image_0_241 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_242 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hf2 == _T_37[9:0]) begin
        image_0_242 <= io_pixelVal_in_0_7;
      end else if (10'hf2 == _T_34[9:0]) begin
        image_0_242 <= io_pixelVal_in_0_6;
      end else if (10'hf2 == _T_31[9:0]) begin
        image_0_242 <= io_pixelVal_in_0_5;
      end else if (10'hf2 == _T_28[9:0]) begin
        image_0_242 <= io_pixelVal_in_0_4;
      end else if (10'hf2 == _T_25[9:0]) begin
        image_0_242 <= io_pixelVal_in_0_3;
      end else if (10'hf2 == _T_22[9:0]) begin
        image_0_242 <= io_pixelVal_in_0_2;
      end else if (10'hf2 == _T_19[9:0]) begin
        image_0_242 <= io_pixelVal_in_0_1;
      end else if (10'hf2 == _T_15[9:0]) begin
        image_0_242 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_243 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hf3 == _T_37[9:0]) begin
        image_0_243 <= io_pixelVal_in_0_7;
      end else if (10'hf3 == _T_34[9:0]) begin
        image_0_243 <= io_pixelVal_in_0_6;
      end else if (10'hf3 == _T_31[9:0]) begin
        image_0_243 <= io_pixelVal_in_0_5;
      end else if (10'hf3 == _T_28[9:0]) begin
        image_0_243 <= io_pixelVal_in_0_4;
      end else if (10'hf3 == _T_25[9:0]) begin
        image_0_243 <= io_pixelVal_in_0_3;
      end else if (10'hf3 == _T_22[9:0]) begin
        image_0_243 <= io_pixelVal_in_0_2;
      end else if (10'hf3 == _T_19[9:0]) begin
        image_0_243 <= io_pixelVal_in_0_1;
      end else if (10'hf3 == _T_15[9:0]) begin
        image_0_243 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_244 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hf4 == _T_37[9:0]) begin
        image_0_244 <= io_pixelVal_in_0_7;
      end else if (10'hf4 == _T_34[9:0]) begin
        image_0_244 <= io_pixelVal_in_0_6;
      end else if (10'hf4 == _T_31[9:0]) begin
        image_0_244 <= io_pixelVal_in_0_5;
      end else if (10'hf4 == _T_28[9:0]) begin
        image_0_244 <= io_pixelVal_in_0_4;
      end else if (10'hf4 == _T_25[9:0]) begin
        image_0_244 <= io_pixelVal_in_0_3;
      end else if (10'hf4 == _T_22[9:0]) begin
        image_0_244 <= io_pixelVal_in_0_2;
      end else if (10'hf4 == _T_19[9:0]) begin
        image_0_244 <= io_pixelVal_in_0_1;
      end else if (10'hf4 == _T_15[9:0]) begin
        image_0_244 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_245 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hf5 == _T_37[9:0]) begin
        image_0_245 <= io_pixelVal_in_0_7;
      end else if (10'hf5 == _T_34[9:0]) begin
        image_0_245 <= io_pixelVal_in_0_6;
      end else if (10'hf5 == _T_31[9:0]) begin
        image_0_245 <= io_pixelVal_in_0_5;
      end else if (10'hf5 == _T_28[9:0]) begin
        image_0_245 <= io_pixelVal_in_0_4;
      end else if (10'hf5 == _T_25[9:0]) begin
        image_0_245 <= io_pixelVal_in_0_3;
      end else if (10'hf5 == _T_22[9:0]) begin
        image_0_245 <= io_pixelVal_in_0_2;
      end else if (10'hf5 == _T_19[9:0]) begin
        image_0_245 <= io_pixelVal_in_0_1;
      end else if (10'hf5 == _T_15[9:0]) begin
        image_0_245 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_246 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hf6 == _T_37[9:0]) begin
        image_0_246 <= io_pixelVal_in_0_7;
      end else if (10'hf6 == _T_34[9:0]) begin
        image_0_246 <= io_pixelVal_in_0_6;
      end else if (10'hf6 == _T_31[9:0]) begin
        image_0_246 <= io_pixelVal_in_0_5;
      end else if (10'hf6 == _T_28[9:0]) begin
        image_0_246 <= io_pixelVal_in_0_4;
      end else if (10'hf6 == _T_25[9:0]) begin
        image_0_246 <= io_pixelVal_in_0_3;
      end else if (10'hf6 == _T_22[9:0]) begin
        image_0_246 <= io_pixelVal_in_0_2;
      end else if (10'hf6 == _T_19[9:0]) begin
        image_0_246 <= io_pixelVal_in_0_1;
      end else if (10'hf6 == _T_15[9:0]) begin
        image_0_246 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_247 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hf7 == _T_37[9:0]) begin
        image_0_247 <= io_pixelVal_in_0_7;
      end else if (10'hf7 == _T_34[9:0]) begin
        image_0_247 <= io_pixelVal_in_0_6;
      end else if (10'hf7 == _T_31[9:0]) begin
        image_0_247 <= io_pixelVal_in_0_5;
      end else if (10'hf7 == _T_28[9:0]) begin
        image_0_247 <= io_pixelVal_in_0_4;
      end else if (10'hf7 == _T_25[9:0]) begin
        image_0_247 <= io_pixelVal_in_0_3;
      end else if (10'hf7 == _T_22[9:0]) begin
        image_0_247 <= io_pixelVal_in_0_2;
      end else if (10'hf7 == _T_19[9:0]) begin
        image_0_247 <= io_pixelVal_in_0_1;
      end else if (10'hf7 == _T_15[9:0]) begin
        image_0_247 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_248 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hf8 == _T_37[9:0]) begin
        image_0_248 <= io_pixelVal_in_0_7;
      end else if (10'hf8 == _T_34[9:0]) begin
        image_0_248 <= io_pixelVal_in_0_6;
      end else if (10'hf8 == _T_31[9:0]) begin
        image_0_248 <= io_pixelVal_in_0_5;
      end else if (10'hf8 == _T_28[9:0]) begin
        image_0_248 <= io_pixelVal_in_0_4;
      end else if (10'hf8 == _T_25[9:0]) begin
        image_0_248 <= io_pixelVal_in_0_3;
      end else if (10'hf8 == _T_22[9:0]) begin
        image_0_248 <= io_pixelVal_in_0_2;
      end else if (10'hf8 == _T_19[9:0]) begin
        image_0_248 <= io_pixelVal_in_0_1;
      end else if (10'hf8 == _T_15[9:0]) begin
        image_0_248 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_249 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hf9 == _T_37[9:0]) begin
        image_0_249 <= io_pixelVal_in_0_7;
      end else if (10'hf9 == _T_34[9:0]) begin
        image_0_249 <= io_pixelVal_in_0_6;
      end else if (10'hf9 == _T_31[9:0]) begin
        image_0_249 <= io_pixelVal_in_0_5;
      end else if (10'hf9 == _T_28[9:0]) begin
        image_0_249 <= io_pixelVal_in_0_4;
      end else if (10'hf9 == _T_25[9:0]) begin
        image_0_249 <= io_pixelVal_in_0_3;
      end else if (10'hf9 == _T_22[9:0]) begin
        image_0_249 <= io_pixelVal_in_0_2;
      end else if (10'hf9 == _T_19[9:0]) begin
        image_0_249 <= io_pixelVal_in_0_1;
      end else if (10'hf9 == _T_15[9:0]) begin
        image_0_249 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_250 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hfa == _T_37[9:0]) begin
        image_0_250 <= io_pixelVal_in_0_7;
      end else if (10'hfa == _T_34[9:0]) begin
        image_0_250 <= io_pixelVal_in_0_6;
      end else if (10'hfa == _T_31[9:0]) begin
        image_0_250 <= io_pixelVal_in_0_5;
      end else if (10'hfa == _T_28[9:0]) begin
        image_0_250 <= io_pixelVal_in_0_4;
      end else if (10'hfa == _T_25[9:0]) begin
        image_0_250 <= io_pixelVal_in_0_3;
      end else if (10'hfa == _T_22[9:0]) begin
        image_0_250 <= io_pixelVal_in_0_2;
      end else if (10'hfa == _T_19[9:0]) begin
        image_0_250 <= io_pixelVal_in_0_1;
      end else if (10'hfa == _T_15[9:0]) begin
        image_0_250 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_251 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hfb == _T_37[9:0]) begin
        image_0_251 <= io_pixelVal_in_0_7;
      end else if (10'hfb == _T_34[9:0]) begin
        image_0_251 <= io_pixelVal_in_0_6;
      end else if (10'hfb == _T_31[9:0]) begin
        image_0_251 <= io_pixelVal_in_0_5;
      end else if (10'hfb == _T_28[9:0]) begin
        image_0_251 <= io_pixelVal_in_0_4;
      end else if (10'hfb == _T_25[9:0]) begin
        image_0_251 <= io_pixelVal_in_0_3;
      end else if (10'hfb == _T_22[9:0]) begin
        image_0_251 <= io_pixelVal_in_0_2;
      end else if (10'hfb == _T_19[9:0]) begin
        image_0_251 <= io_pixelVal_in_0_1;
      end else if (10'hfb == _T_15[9:0]) begin
        image_0_251 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_252 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hfc == _T_37[9:0]) begin
        image_0_252 <= io_pixelVal_in_0_7;
      end else if (10'hfc == _T_34[9:0]) begin
        image_0_252 <= io_pixelVal_in_0_6;
      end else if (10'hfc == _T_31[9:0]) begin
        image_0_252 <= io_pixelVal_in_0_5;
      end else if (10'hfc == _T_28[9:0]) begin
        image_0_252 <= io_pixelVal_in_0_4;
      end else if (10'hfc == _T_25[9:0]) begin
        image_0_252 <= io_pixelVal_in_0_3;
      end else if (10'hfc == _T_22[9:0]) begin
        image_0_252 <= io_pixelVal_in_0_2;
      end else if (10'hfc == _T_19[9:0]) begin
        image_0_252 <= io_pixelVal_in_0_1;
      end else if (10'hfc == _T_15[9:0]) begin
        image_0_252 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_253 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hfd == _T_37[9:0]) begin
        image_0_253 <= io_pixelVal_in_0_7;
      end else if (10'hfd == _T_34[9:0]) begin
        image_0_253 <= io_pixelVal_in_0_6;
      end else if (10'hfd == _T_31[9:0]) begin
        image_0_253 <= io_pixelVal_in_0_5;
      end else if (10'hfd == _T_28[9:0]) begin
        image_0_253 <= io_pixelVal_in_0_4;
      end else if (10'hfd == _T_25[9:0]) begin
        image_0_253 <= io_pixelVal_in_0_3;
      end else if (10'hfd == _T_22[9:0]) begin
        image_0_253 <= io_pixelVal_in_0_2;
      end else if (10'hfd == _T_19[9:0]) begin
        image_0_253 <= io_pixelVal_in_0_1;
      end else if (10'hfd == _T_15[9:0]) begin
        image_0_253 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_254 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hfe == _T_37[9:0]) begin
        image_0_254 <= io_pixelVal_in_0_7;
      end else if (10'hfe == _T_34[9:0]) begin
        image_0_254 <= io_pixelVal_in_0_6;
      end else if (10'hfe == _T_31[9:0]) begin
        image_0_254 <= io_pixelVal_in_0_5;
      end else if (10'hfe == _T_28[9:0]) begin
        image_0_254 <= io_pixelVal_in_0_4;
      end else if (10'hfe == _T_25[9:0]) begin
        image_0_254 <= io_pixelVal_in_0_3;
      end else if (10'hfe == _T_22[9:0]) begin
        image_0_254 <= io_pixelVal_in_0_2;
      end else if (10'hfe == _T_19[9:0]) begin
        image_0_254 <= io_pixelVal_in_0_1;
      end else if (10'hfe == _T_15[9:0]) begin
        image_0_254 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_255 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hff == _T_37[9:0]) begin
        image_0_255 <= io_pixelVal_in_0_7;
      end else if (10'hff == _T_34[9:0]) begin
        image_0_255 <= io_pixelVal_in_0_6;
      end else if (10'hff == _T_31[9:0]) begin
        image_0_255 <= io_pixelVal_in_0_5;
      end else if (10'hff == _T_28[9:0]) begin
        image_0_255 <= io_pixelVal_in_0_4;
      end else if (10'hff == _T_25[9:0]) begin
        image_0_255 <= io_pixelVal_in_0_3;
      end else if (10'hff == _T_22[9:0]) begin
        image_0_255 <= io_pixelVal_in_0_2;
      end else if (10'hff == _T_19[9:0]) begin
        image_0_255 <= io_pixelVal_in_0_1;
      end else if (10'hff == _T_15[9:0]) begin
        image_0_255 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_256 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h100 == _T_37[9:0]) begin
        image_0_256 <= io_pixelVal_in_0_7;
      end else if (10'h100 == _T_34[9:0]) begin
        image_0_256 <= io_pixelVal_in_0_6;
      end else if (10'h100 == _T_31[9:0]) begin
        image_0_256 <= io_pixelVal_in_0_5;
      end else if (10'h100 == _T_28[9:0]) begin
        image_0_256 <= io_pixelVal_in_0_4;
      end else if (10'h100 == _T_25[9:0]) begin
        image_0_256 <= io_pixelVal_in_0_3;
      end else if (10'h100 == _T_22[9:0]) begin
        image_0_256 <= io_pixelVal_in_0_2;
      end else if (10'h100 == _T_19[9:0]) begin
        image_0_256 <= io_pixelVal_in_0_1;
      end else if (10'h100 == _T_15[9:0]) begin
        image_0_256 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_257 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h101 == _T_37[9:0]) begin
        image_0_257 <= io_pixelVal_in_0_7;
      end else if (10'h101 == _T_34[9:0]) begin
        image_0_257 <= io_pixelVal_in_0_6;
      end else if (10'h101 == _T_31[9:0]) begin
        image_0_257 <= io_pixelVal_in_0_5;
      end else if (10'h101 == _T_28[9:0]) begin
        image_0_257 <= io_pixelVal_in_0_4;
      end else if (10'h101 == _T_25[9:0]) begin
        image_0_257 <= io_pixelVal_in_0_3;
      end else if (10'h101 == _T_22[9:0]) begin
        image_0_257 <= io_pixelVal_in_0_2;
      end else if (10'h101 == _T_19[9:0]) begin
        image_0_257 <= io_pixelVal_in_0_1;
      end else if (10'h101 == _T_15[9:0]) begin
        image_0_257 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_258 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h102 == _T_37[9:0]) begin
        image_0_258 <= io_pixelVal_in_0_7;
      end else if (10'h102 == _T_34[9:0]) begin
        image_0_258 <= io_pixelVal_in_0_6;
      end else if (10'h102 == _T_31[9:0]) begin
        image_0_258 <= io_pixelVal_in_0_5;
      end else if (10'h102 == _T_28[9:0]) begin
        image_0_258 <= io_pixelVal_in_0_4;
      end else if (10'h102 == _T_25[9:0]) begin
        image_0_258 <= io_pixelVal_in_0_3;
      end else if (10'h102 == _T_22[9:0]) begin
        image_0_258 <= io_pixelVal_in_0_2;
      end else if (10'h102 == _T_19[9:0]) begin
        image_0_258 <= io_pixelVal_in_0_1;
      end else if (10'h102 == _T_15[9:0]) begin
        image_0_258 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_259 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h103 == _T_37[9:0]) begin
        image_0_259 <= io_pixelVal_in_0_7;
      end else if (10'h103 == _T_34[9:0]) begin
        image_0_259 <= io_pixelVal_in_0_6;
      end else if (10'h103 == _T_31[9:0]) begin
        image_0_259 <= io_pixelVal_in_0_5;
      end else if (10'h103 == _T_28[9:0]) begin
        image_0_259 <= io_pixelVal_in_0_4;
      end else if (10'h103 == _T_25[9:0]) begin
        image_0_259 <= io_pixelVal_in_0_3;
      end else if (10'h103 == _T_22[9:0]) begin
        image_0_259 <= io_pixelVal_in_0_2;
      end else if (10'h103 == _T_19[9:0]) begin
        image_0_259 <= io_pixelVal_in_0_1;
      end else if (10'h103 == _T_15[9:0]) begin
        image_0_259 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_260 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h104 == _T_37[9:0]) begin
        image_0_260 <= io_pixelVal_in_0_7;
      end else if (10'h104 == _T_34[9:0]) begin
        image_0_260 <= io_pixelVal_in_0_6;
      end else if (10'h104 == _T_31[9:0]) begin
        image_0_260 <= io_pixelVal_in_0_5;
      end else if (10'h104 == _T_28[9:0]) begin
        image_0_260 <= io_pixelVal_in_0_4;
      end else if (10'h104 == _T_25[9:0]) begin
        image_0_260 <= io_pixelVal_in_0_3;
      end else if (10'h104 == _T_22[9:0]) begin
        image_0_260 <= io_pixelVal_in_0_2;
      end else if (10'h104 == _T_19[9:0]) begin
        image_0_260 <= io_pixelVal_in_0_1;
      end else if (10'h104 == _T_15[9:0]) begin
        image_0_260 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_261 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h105 == _T_37[9:0]) begin
        image_0_261 <= io_pixelVal_in_0_7;
      end else if (10'h105 == _T_34[9:0]) begin
        image_0_261 <= io_pixelVal_in_0_6;
      end else if (10'h105 == _T_31[9:0]) begin
        image_0_261 <= io_pixelVal_in_0_5;
      end else if (10'h105 == _T_28[9:0]) begin
        image_0_261 <= io_pixelVal_in_0_4;
      end else if (10'h105 == _T_25[9:0]) begin
        image_0_261 <= io_pixelVal_in_0_3;
      end else if (10'h105 == _T_22[9:0]) begin
        image_0_261 <= io_pixelVal_in_0_2;
      end else if (10'h105 == _T_19[9:0]) begin
        image_0_261 <= io_pixelVal_in_0_1;
      end else if (10'h105 == _T_15[9:0]) begin
        image_0_261 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_262 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h106 == _T_37[9:0]) begin
        image_0_262 <= io_pixelVal_in_0_7;
      end else if (10'h106 == _T_34[9:0]) begin
        image_0_262 <= io_pixelVal_in_0_6;
      end else if (10'h106 == _T_31[9:0]) begin
        image_0_262 <= io_pixelVal_in_0_5;
      end else if (10'h106 == _T_28[9:0]) begin
        image_0_262 <= io_pixelVal_in_0_4;
      end else if (10'h106 == _T_25[9:0]) begin
        image_0_262 <= io_pixelVal_in_0_3;
      end else if (10'h106 == _T_22[9:0]) begin
        image_0_262 <= io_pixelVal_in_0_2;
      end else if (10'h106 == _T_19[9:0]) begin
        image_0_262 <= io_pixelVal_in_0_1;
      end else if (10'h106 == _T_15[9:0]) begin
        image_0_262 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_263 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h107 == _T_37[9:0]) begin
        image_0_263 <= io_pixelVal_in_0_7;
      end else if (10'h107 == _T_34[9:0]) begin
        image_0_263 <= io_pixelVal_in_0_6;
      end else if (10'h107 == _T_31[9:0]) begin
        image_0_263 <= io_pixelVal_in_0_5;
      end else if (10'h107 == _T_28[9:0]) begin
        image_0_263 <= io_pixelVal_in_0_4;
      end else if (10'h107 == _T_25[9:0]) begin
        image_0_263 <= io_pixelVal_in_0_3;
      end else if (10'h107 == _T_22[9:0]) begin
        image_0_263 <= io_pixelVal_in_0_2;
      end else if (10'h107 == _T_19[9:0]) begin
        image_0_263 <= io_pixelVal_in_0_1;
      end else if (10'h107 == _T_15[9:0]) begin
        image_0_263 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_264 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h108 == _T_37[9:0]) begin
        image_0_264 <= io_pixelVal_in_0_7;
      end else if (10'h108 == _T_34[9:0]) begin
        image_0_264 <= io_pixelVal_in_0_6;
      end else if (10'h108 == _T_31[9:0]) begin
        image_0_264 <= io_pixelVal_in_0_5;
      end else if (10'h108 == _T_28[9:0]) begin
        image_0_264 <= io_pixelVal_in_0_4;
      end else if (10'h108 == _T_25[9:0]) begin
        image_0_264 <= io_pixelVal_in_0_3;
      end else if (10'h108 == _T_22[9:0]) begin
        image_0_264 <= io_pixelVal_in_0_2;
      end else if (10'h108 == _T_19[9:0]) begin
        image_0_264 <= io_pixelVal_in_0_1;
      end else if (10'h108 == _T_15[9:0]) begin
        image_0_264 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_265 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h109 == _T_37[9:0]) begin
        image_0_265 <= io_pixelVal_in_0_7;
      end else if (10'h109 == _T_34[9:0]) begin
        image_0_265 <= io_pixelVal_in_0_6;
      end else if (10'h109 == _T_31[9:0]) begin
        image_0_265 <= io_pixelVal_in_0_5;
      end else if (10'h109 == _T_28[9:0]) begin
        image_0_265 <= io_pixelVal_in_0_4;
      end else if (10'h109 == _T_25[9:0]) begin
        image_0_265 <= io_pixelVal_in_0_3;
      end else if (10'h109 == _T_22[9:0]) begin
        image_0_265 <= io_pixelVal_in_0_2;
      end else if (10'h109 == _T_19[9:0]) begin
        image_0_265 <= io_pixelVal_in_0_1;
      end else if (10'h109 == _T_15[9:0]) begin
        image_0_265 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_266 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h10a == _T_37[9:0]) begin
        image_0_266 <= io_pixelVal_in_0_7;
      end else if (10'h10a == _T_34[9:0]) begin
        image_0_266 <= io_pixelVal_in_0_6;
      end else if (10'h10a == _T_31[9:0]) begin
        image_0_266 <= io_pixelVal_in_0_5;
      end else if (10'h10a == _T_28[9:0]) begin
        image_0_266 <= io_pixelVal_in_0_4;
      end else if (10'h10a == _T_25[9:0]) begin
        image_0_266 <= io_pixelVal_in_0_3;
      end else if (10'h10a == _T_22[9:0]) begin
        image_0_266 <= io_pixelVal_in_0_2;
      end else if (10'h10a == _T_19[9:0]) begin
        image_0_266 <= io_pixelVal_in_0_1;
      end else if (10'h10a == _T_15[9:0]) begin
        image_0_266 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_267 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h10b == _T_37[9:0]) begin
        image_0_267 <= io_pixelVal_in_0_7;
      end else if (10'h10b == _T_34[9:0]) begin
        image_0_267 <= io_pixelVal_in_0_6;
      end else if (10'h10b == _T_31[9:0]) begin
        image_0_267 <= io_pixelVal_in_0_5;
      end else if (10'h10b == _T_28[9:0]) begin
        image_0_267 <= io_pixelVal_in_0_4;
      end else if (10'h10b == _T_25[9:0]) begin
        image_0_267 <= io_pixelVal_in_0_3;
      end else if (10'h10b == _T_22[9:0]) begin
        image_0_267 <= io_pixelVal_in_0_2;
      end else if (10'h10b == _T_19[9:0]) begin
        image_0_267 <= io_pixelVal_in_0_1;
      end else if (10'h10b == _T_15[9:0]) begin
        image_0_267 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_268 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h10c == _T_37[9:0]) begin
        image_0_268 <= io_pixelVal_in_0_7;
      end else if (10'h10c == _T_34[9:0]) begin
        image_0_268 <= io_pixelVal_in_0_6;
      end else if (10'h10c == _T_31[9:0]) begin
        image_0_268 <= io_pixelVal_in_0_5;
      end else if (10'h10c == _T_28[9:0]) begin
        image_0_268 <= io_pixelVal_in_0_4;
      end else if (10'h10c == _T_25[9:0]) begin
        image_0_268 <= io_pixelVal_in_0_3;
      end else if (10'h10c == _T_22[9:0]) begin
        image_0_268 <= io_pixelVal_in_0_2;
      end else if (10'h10c == _T_19[9:0]) begin
        image_0_268 <= io_pixelVal_in_0_1;
      end else if (10'h10c == _T_15[9:0]) begin
        image_0_268 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_269 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h10d == _T_37[9:0]) begin
        image_0_269 <= io_pixelVal_in_0_7;
      end else if (10'h10d == _T_34[9:0]) begin
        image_0_269 <= io_pixelVal_in_0_6;
      end else if (10'h10d == _T_31[9:0]) begin
        image_0_269 <= io_pixelVal_in_0_5;
      end else if (10'h10d == _T_28[9:0]) begin
        image_0_269 <= io_pixelVal_in_0_4;
      end else if (10'h10d == _T_25[9:0]) begin
        image_0_269 <= io_pixelVal_in_0_3;
      end else if (10'h10d == _T_22[9:0]) begin
        image_0_269 <= io_pixelVal_in_0_2;
      end else if (10'h10d == _T_19[9:0]) begin
        image_0_269 <= io_pixelVal_in_0_1;
      end else if (10'h10d == _T_15[9:0]) begin
        image_0_269 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_270 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h10e == _T_37[9:0]) begin
        image_0_270 <= io_pixelVal_in_0_7;
      end else if (10'h10e == _T_34[9:0]) begin
        image_0_270 <= io_pixelVal_in_0_6;
      end else if (10'h10e == _T_31[9:0]) begin
        image_0_270 <= io_pixelVal_in_0_5;
      end else if (10'h10e == _T_28[9:0]) begin
        image_0_270 <= io_pixelVal_in_0_4;
      end else if (10'h10e == _T_25[9:0]) begin
        image_0_270 <= io_pixelVal_in_0_3;
      end else if (10'h10e == _T_22[9:0]) begin
        image_0_270 <= io_pixelVal_in_0_2;
      end else if (10'h10e == _T_19[9:0]) begin
        image_0_270 <= io_pixelVal_in_0_1;
      end else if (10'h10e == _T_15[9:0]) begin
        image_0_270 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_271 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h10f == _T_37[9:0]) begin
        image_0_271 <= io_pixelVal_in_0_7;
      end else if (10'h10f == _T_34[9:0]) begin
        image_0_271 <= io_pixelVal_in_0_6;
      end else if (10'h10f == _T_31[9:0]) begin
        image_0_271 <= io_pixelVal_in_0_5;
      end else if (10'h10f == _T_28[9:0]) begin
        image_0_271 <= io_pixelVal_in_0_4;
      end else if (10'h10f == _T_25[9:0]) begin
        image_0_271 <= io_pixelVal_in_0_3;
      end else if (10'h10f == _T_22[9:0]) begin
        image_0_271 <= io_pixelVal_in_0_2;
      end else if (10'h10f == _T_19[9:0]) begin
        image_0_271 <= io_pixelVal_in_0_1;
      end else if (10'h10f == _T_15[9:0]) begin
        image_0_271 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_272 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h110 == _T_37[9:0]) begin
        image_0_272 <= io_pixelVal_in_0_7;
      end else if (10'h110 == _T_34[9:0]) begin
        image_0_272 <= io_pixelVal_in_0_6;
      end else if (10'h110 == _T_31[9:0]) begin
        image_0_272 <= io_pixelVal_in_0_5;
      end else if (10'h110 == _T_28[9:0]) begin
        image_0_272 <= io_pixelVal_in_0_4;
      end else if (10'h110 == _T_25[9:0]) begin
        image_0_272 <= io_pixelVal_in_0_3;
      end else if (10'h110 == _T_22[9:0]) begin
        image_0_272 <= io_pixelVal_in_0_2;
      end else if (10'h110 == _T_19[9:0]) begin
        image_0_272 <= io_pixelVal_in_0_1;
      end else if (10'h110 == _T_15[9:0]) begin
        image_0_272 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_273 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h111 == _T_37[9:0]) begin
        image_0_273 <= io_pixelVal_in_0_7;
      end else if (10'h111 == _T_34[9:0]) begin
        image_0_273 <= io_pixelVal_in_0_6;
      end else if (10'h111 == _T_31[9:0]) begin
        image_0_273 <= io_pixelVal_in_0_5;
      end else if (10'h111 == _T_28[9:0]) begin
        image_0_273 <= io_pixelVal_in_0_4;
      end else if (10'h111 == _T_25[9:0]) begin
        image_0_273 <= io_pixelVal_in_0_3;
      end else if (10'h111 == _T_22[9:0]) begin
        image_0_273 <= io_pixelVal_in_0_2;
      end else if (10'h111 == _T_19[9:0]) begin
        image_0_273 <= io_pixelVal_in_0_1;
      end else if (10'h111 == _T_15[9:0]) begin
        image_0_273 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_274 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h112 == _T_37[9:0]) begin
        image_0_274 <= io_pixelVal_in_0_7;
      end else if (10'h112 == _T_34[9:0]) begin
        image_0_274 <= io_pixelVal_in_0_6;
      end else if (10'h112 == _T_31[9:0]) begin
        image_0_274 <= io_pixelVal_in_0_5;
      end else if (10'h112 == _T_28[9:0]) begin
        image_0_274 <= io_pixelVal_in_0_4;
      end else if (10'h112 == _T_25[9:0]) begin
        image_0_274 <= io_pixelVal_in_0_3;
      end else if (10'h112 == _T_22[9:0]) begin
        image_0_274 <= io_pixelVal_in_0_2;
      end else if (10'h112 == _T_19[9:0]) begin
        image_0_274 <= io_pixelVal_in_0_1;
      end else if (10'h112 == _T_15[9:0]) begin
        image_0_274 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_275 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h113 == _T_37[9:0]) begin
        image_0_275 <= io_pixelVal_in_0_7;
      end else if (10'h113 == _T_34[9:0]) begin
        image_0_275 <= io_pixelVal_in_0_6;
      end else if (10'h113 == _T_31[9:0]) begin
        image_0_275 <= io_pixelVal_in_0_5;
      end else if (10'h113 == _T_28[9:0]) begin
        image_0_275 <= io_pixelVal_in_0_4;
      end else if (10'h113 == _T_25[9:0]) begin
        image_0_275 <= io_pixelVal_in_0_3;
      end else if (10'h113 == _T_22[9:0]) begin
        image_0_275 <= io_pixelVal_in_0_2;
      end else if (10'h113 == _T_19[9:0]) begin
        image_0_275 <= io_pixelVal_in_0_1;
      end else if (10'h113 == _T_15[9:0]) begin
        image_0_275 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_276 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h114 == _T_37[9:0]) begin
        image_0_276 <= io_pixelVal_in_0_7;
      end else if (10'h114 == _T_34[9:0]) begin
        image_0_276 <= io_pixelVal_in_0_6;
      end else if (10'h114 == _T_31[9:0]) begin
        image_0_276 <= io_pixelVal_in_0_5;
      end else if (10'h114 == _T_28[9:0]) begin
        image_0_276 <= io_pixelVal_in_0_4;
      end else if (10'h114 == _T_25[9:0]) begin
        image_0_276 <= io_pixelVal_in_0_3;
      end else if (10'h114 == _T_22[9:0]) begin
        image_0_276 <= io_pixelVal_in_0_2;
      end else if (10'h114 == _T_19[9:0]) begin
        image_0_276 <= io_pixelVal_in_0_1;
      end else if (10'h114 == _T_15[9:0]) begin
        image_0_276 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_277 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h115 == _T_37[9:0]) begin
        image_0_277 <= io_pixelVal_in_0_7;
      end else if (10'h115 == _T_34[9:0]) begin
        image_0_277 <= io_pixelVal_in_0_6;
      end else if (10'h115 == _T_31[9:0]) begin
        image_0_277 <= io_pixelVal_in_0_5;
      end else if (10'h115 == _T_28[9:0]) begin
        image_0_277 <= io_pixelVal_in_0_4;
      end else if (10'h115 == _T_25[9:0]) begin
        image_0_277 <= io_pixelVal_in_0_3;
      end else if (10'h115 == _T_22[9:0]) begin
        image_0_277 <= io_pixelVal_in_0_2;
      end else if (10'h115 == _T_19[9:0]) begin
        image_0_277 <= io_pixelVal_in_0_1;
      end else if (10'h115 == _T_15[9:0]) begin
        image_0_277 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_278 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h116 == _T_37[9:0]) begin
        image_0_278 <= io_pixelVal_in_0_7;
      end else if (10'h116 == _T_34[9:0]) begin
        image_0_278 <= io_pixelVal_in_0_6;
      end else if (10'h116 == _T_31[9:0]) begin
        image_0_278 <= io_pixelVal_in_0_5;
      end else if (10'h116 == _T_28[9:0]) begin
        image_0_278 <= io_pixelVal_in_0_4;
      end else if (10'h116 == _T_25[9:0]) begin
        image_0_278 <= io_pixelVal_in_0_3;
      end else if (10'h116 == _T_22[9:0]) begin
        image_0_278 <= io_pixelVal_in_0_2;
      end else if (10'h116 == _T_19[9:0]) begin
        image_0_278 <= io_pixelVal_in_0_1;
      end else if (10'h116 == _T_15[9:0]) begin
        image_0_278 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_279 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h117 == _T_37[9:0]) begin
        image_0_279 <= io_pixelVal_in_0_7;
      end else if (10'h117 == _T_34[9:0]) begin
        image_0_279 <= io_pixelVal_in_0_6;
      end else if (10'h117 == _T_31[9:0]) begin
        image_0_279 <= io_pixelVal_in_0_5;
      end else if (10'h117 == _T_28[9:0]) begin
        image_0_279 <= io_pixelVal_in_0_4;
      end else if (10'h117 == _T_25[9:0]) begin
        image_0_279 <= io_pixelVal_in_0_3;
      end else if (10'h117 == _T_22[9:0]) begin
        image_0_279 <= io_pixelVal_in_0_2;
      end else if (10'h117 == _T_19[9:0]) begin
        image_0_279 <= io_pixelVal_in_0_1;
      end else if (10'h117 == _T_15[9:0]) begin
        image_0_279 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_280 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h118 == _T_37[9:0]) begin
        image_0_280 <= io_pixelVal_in_0_7;
      end else if (10'h118 == _T_34[9:0]) begin
        image_0_280 <= io_pixelVal_in_0_6;
      end else if (10'h118 == _T_31[9:0]) begin
        image_0_280 <= io_pixelVal_in_0_5;
      end else if (10'h118 == _T_28[9:0]) begin
        image_0_280 <= io_pixelVal_in_0_4;
      end else if (10'h118 == _T_25[9:0]) begin
        image_0_280 <= io_pixelVal_in_0_3;
      end else if (10'h118 == _T_22[9:0]) begin
        image_0_280 <= io_pixelVal_in_0_2;
      end else if (10'h118 == _T_19[9:0]) begin
        image_0_280 <= io_pixelVal_in_0_1;
      end else if (10'h118 == _T_15[9:0]) begin
        image_0_280 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_281 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h119 == _T_37[9:0]) begin
        image_0_281 <= io_pixelVal_in_0_7;
      end else if (10'h119 == _T_34[9:0]) begin
        image_0_281 <= io_pixelVal_in_0_6;
      end else if (10'h119 == _T_31[9:0]) begin
        image_0_281 <= io_pixelVal_in_0_5;
      end else if (10'h119 == _T_28[9:0]) begin
        image_0_281 <= io_pixelVal_in_0_4;
      end else if (10'h119 == _T_25[9:0]) begin
        image_0_281 <= io_pixelVal_in_0_3;
      end else if (10'h119 == _T_22[9:0]) begin
        image_0_281 <= io_pixelVal_in_0_2;
      end else if (10'h119 == _T_19[9:0]) begin
        image_0_281 <= io_pixelVal_in_0_1;
      end else if (10'h119 == _T_15[9:0]) begin
        image_0_281 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_282 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h11a == _T_37[9:0]) begin
        image_0_282 <= io_pixelVal_in_0_7;
      end else if (10'h11a == _T_34[9:0]) begin
        image_0_282 <= io_pixelVal_in_0_6;
      end else if (10'h11a == _T_31[9:0]) begin
        image_0_282 <= io_pixelVal_in_0_5;
      end else if (10'h11a == _T_28[9:0]) begin
        image_0_282 <= io_pixelVal_in_0_4;
      end else if (10'h11a == _T_25[9:0]) begin
        image_0_282 <= io_pixelVal_in_0_3;
      end else if (10'h11a == _T_22[9:0]) begin
        image_0_282 <= io_pixelVal_in_0_2;
      end else if (10'h11a == _T_19[9:0]) begin
        image_0_282 <= io_pixelVal_in_0_1;
      end else if (10'h11a == _T_15[9:0]) begin
        image_0_282 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_283 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h11b == _T_37[9:0]) begin
        image_0_283 <= io_pixelVal_in_0_7;
      end else if (10'h11b == _T_34[9:0]) begin
        image_0_283 <= io_pixelVal_in_0_6;
      end else if (10'h11b == _T_31[9:0]) begin
        image_0_283 <= io_pixelVal_in_0_5;
      end else if (10'h11b == _T_28[9:0]) begin
        image_0_283 <= io_pixelVal_in_0_4;
      end else if (10'h11b == _T_25[9:0]) begin
        image_0_283 <= io_pixelVal_in_0_3;
      end else if (10'h11b == _T_22[9:0]) begin
        image_0_283 <= io_pixelVal_in_0_2;
      end else if (10'h11b == _T_19[9:0]) begin
        image_0_283 <= io_pixelVal_in_0_1;
      end else if (10'h11b == _T_15[9:0]) begin
        image_0_283 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_284 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h11c == _T_37[9:0]) begin
        image_0_284 <= io_pixelVal_in_0_7;
      end else if (10'h11c == _T_34[9:0]) begin
        image_0_284 <= io_pixelVal_in_0_6;
      end else if (10'h11c == _T_31[9:0]) begin
        image_0_284 <= io_pixelVal_in_0_5;
      end else if (10'h11c == _T_28[9:0]) begin
        image_0_284 <= io_pixelVal_in_0_4;
      end else if (10'h11c == _T_25[9:0]) begin
        image_0_284 <= io_pixelVal_in_0_3;
      end else if (10'h11c == _T_22[9:0]) begin
        image_0_284 <= io_pixelVal_in_0_2;
      end else if (10'h11c == _T_19[9:0]) begin
        image_0_284 <= io_pixelVal_in_0_1;
      end else if (10'h11c == _T_15[9:0]) begin
        image_0_284 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_285 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h11d == _T_37[9:0]) begin
        image_0_285 <= io_pixelVal_in_0_7;
      end else if (10'h11d == _T_34[9:0]) begin
        image_0_285 <= io_pixelVal_in_0_6;
      end else if (10'h11d == _T_31[9:0]) begin
        image_0_285 <= io_pixelVal_in_0_5;
      end else if (10'h11d == _T_28[9:0]) begin
        image_0_285 <= io_pixelVal_in_0_4;
      end else if (10'h11d == _T_25[9:0]) begin
        image_0_285 <= io_pixelVal_in_0_3;
      end else if (10'h11d == _T_22[9:0]) begin
        image_0_285 <= io_pixelVal_in_0_2;
      end else if (10'h11d == _T_19[9:0]) begin
        image_0_285 <= io_pixelVal_in_0_1;
      end else if (10'h11d == _T_15[9:0]) begin
        image_0_285 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_286 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h11e == _T_37[9:0]) begin
        image_0_286 <= io_pixelVal_in_0_7;
      end else if (10'h11e == _T_34[9:0]) begin
        image_0_286 <= io_pixelVal_in_0_6;
      end else if (10'h11e == _T_31[9:0]) begin
        image_0_286 <= io_pixelVal_in_0_5;
      end else if (10'h11e == _T_28[9:0]) begin
        image_0_286 <= io_pixelVal_in_0_4;
      end else if (10'h11e == _T_25[9:0]) begin
        image_0_286 <= io_pixelVal_in_0_3;
      end else if (10'h11e == _T_22[9:0]) begin
        image_0_286 <= io_pixelVal_in_0_2;
      end else if (10'h11e == _T_19[9:0]) begin
        image_0_286 <= io_pixelVal_in_0_1;
      end else if (10'h11e == _T_15[9:0]) begin
        image_0_286 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_287 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h11f == _T_37[9:0]) begin
        image_0_287 <= io_pixelVal_in_0_7;
      end else if (10'h11f == _T_34[9:0]) begin
        image_0_287 <= io_pixelVal_in_0_6;
      end else if (10'h11f == _T_31[9:0]) begin
        image_0_287 <= io_pixelVal_in_0_5;
      end else if (10'h11f == _T_28[9:0]) begin
        image_0_287 <= io_pixelVal_in_0_4;
      end else if (10'h11f == _T_25[9:0]) begin
        image_0_287 <= io_pixelVal_in_0_3;
      end else if (10'h11f == _T_22[9:0]) begin
        image_0_287 <= io_pixelVal_in_0_2;
      end else if (10'h11f == _T_19[9:0]) begin
        image_0_287 <= io_pixelVal_in_0_1;
      end else if (10'h11f == _T_15[9:0]) begin
        image_0_287 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_288 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h120 == _T_37[9:0]) begin
        image_0_288 <= io_pixelVal_in_0_7;
      end else if (10'h120 == _T_34[9:0]) begin
        image_0_288 <= io_pixelVal_in_0_6;
      end else if (10'h120 == _T_31[9:0]) begin
        image_0_288 <= io_pixelVal_in_0_5;
      end else if (10'h120 == _T_28[9:0]) begin
        image_0_288 <= io_pixelVal_in_0_4;
      end else if (10'h120 == _T_25[9:0]) begin
        image_0_288 <= io_pixelVal_in_0_3;
      end else if (10'h120 == _T_22[9:0]) begin
        image_0_288 <= io_pixelVal_in_0_2;
      end else if (10'h120 == _T_19[9:0]) begin
        image_0_288 <= io_pixelVal_in_0_1;
      end else if (10'h120 == _T_15[9:0]) begin
        image_0_288 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_289 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h121 == _T_37[9:0]) begin
        image_0_289 <= io_pixelVal_in_0_7;
      end else if (10'h121 == _T_34[9:0]) begin
        image_0_289 <= io_pixelVal_in_0_6;
      end else if (10'h121 == _T_31[9:0]) begin
        image_0_289 <= io_pixelVal_in_0_5;
      end else if (10'h121 == _T_28[9:0]) begin
        image_0_289 <= io_pixelVal_in_0_4;
      end else if (10'h121 == _T_25[9:0]) begin
        image_0_289 <= io_pixelVal_in_0_3;
      end else if (10'h121 == _T_22[9:0]) begin
        image_0_289 <= io_pixelVal_in_0_2;
      end else if (10'h121 == _T_19[9:0]) begin
        image_0_289 <= io_pixelVal_in_0_1;
      end else if (10'h121 == _T_15[9:0]) begin
        image_0_289 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_290 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h122 == _T_37[9:0]) begin
        image_0_290 <= io_pixelVal_in_0_7;
      end else if (10'h122 == _T_34[9:0]) begin
        image_0_290 <= io_pixelVal_in_0_6;
      end else if (10'h122 == _T_31[9:0]) begin
        image_0_290 <= io_pixelVal_in_0_5;
      end else if (10'h122 == _T_28[9:0]) begin
        image_0_290 <= io_pixelVal_in_0_4;
      end else if (10'h122 == _T_25[9:0]) begin
        image_0_290 <= io_pixelVal_in_0_3;
      end else if (10'h122 == _T_22[9:0]) begin
        image_0_290 <= io_pixelVal_in_0_2;
      end else if (10'h122 == _T_19[9:0]) begin
        image_0_290 <= io_pixelVal_in_0_1;
      end else if (10'h122 == _T_15[9:0]) begin
        image_0_290 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_291 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h123 == _T_37[9:0]) begin
        image_0_291 <= io_pixelVal_in_0_7;
      end else if (10'h123 == _T_34[9:0]) begin
        image_0_291 <= io_pixelVal_in_0_6;
      end else if (10'h123 == _T_31[9:0]) begin
        image_0_291 <= io_pixelVal_in_0_5;
      end else if (10'h123 == _T_28[9:0]) begin
        image_0_291 <= io_pixelVal_in_0_4;
      end else if (10'h123 == _T_25[9:0]) begin
        image_0_291 <= io_pixelVal_in_0_3;
      end else if (10'h123 == _T_22[9:0]) begin
        image_0_291 <= io_pixelVal_in_0_2;
      end else if (10'h123 == _T_19[9:0]) begin
        image_0_291 <= io_pixelVal_in_0_1;
      end else if (10'h123 == _T_15[9:0]) begin
        image_0_291 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_292 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h124 == _T_37[9:0]) begin
        image_0_292 <= io_pixelVal_in_0_7;
      end else if (10'h124 == _T_34[9:0]) begin
        image_0_292 <= io_pixelVal_in_0_6;
      end else if (10'h124 == _T_31[9:0]) begin
        image_0_292 <= io_pixelVal_in_0_5;
      end else if (10'h124 == _T_28[9:0]) begin
        image_0_292 <= io_pixelVal_in_0_4;
      end else if (10'h124 == _T_25[9:0]) begin
        image_0_292 <= io_pixelVal_in_0_3;
      end else if (10'h124 == _T_22[9:0]) begin
        image_0_292 <= io_pixelVal_in_0_2;
      end else if (10'h124 == _T_19[9:0]) begin
        image_0_292 <= io_pixelVal_in_0_1;
      end else if (10'h124 == _T_15[9:0]) begin
        image_0_292 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_293 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h125 == _T_37[9:0]) begin
        image_0_293 <= io_pixelVal_in_0_7;
      end else if (10'h125 == _T_34[9:0]) begin
        image_0_293 <= io_pixelVal_in_0_6;
      end else if (10'h125 == _T_31[9:0]) begin
        image_0_293 <= io_pixelVal_in_0_5;
      end else if (10'h125 == _T_28[9:0]) begin
        image_0_293 <= io_pixelVal_in_0_4;
      end else if (10'h125 == _T_25[9:0]) begin
        image_0_293 <= io_pixelVal_in_0_3;
      end else if (10'h125 == _T_22[9:0]) begin
        image_0_293 <= io_pixelVal_in_0_2;
      end else if (10'h125 == _T_19[9:0]) begin
        image_0_293 <= io_pixelVal_in_0_1;
      end else if (10'h125 == _T_15[9:0]) begin
        image_0_293 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_294 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h126 == _T_37[9:0]) begin
        image_0_294 <= io_pixelVal_in_0_7;
      end else if (10'h126 == _T_34[9:0]) begin
        image_0_294 <= io_pixelVal_in_0_6;
      end else if (10'h126 == _T_31[9:0]) begin
        image_0_294 <= io_pixelVal_in_0_5;
      end else if (10'h126 == _T_28[9:0]) begin
        image_0_294 <= io_pixelVal_in_0_4;
      end else if (10'h126 == _T_25[9:0]) begin
        image_0_294 <= io_pixelVal_in_0_3;
      end else if (10'h126 == _T_22[9:0]) begin
        image_0_294 <= io_pixelVal_in_0_2;
      end else if (10'h126 == _T_19[9:0]) begin
        image_0_294 <= io_pixelVal_in_0_1;
      end else if (10'h126 == _T_15[9:0]) begin
        image_0_294 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_295 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h127 == _T_37[9:0]) begin
        image_0_295 <= io_pixelVal_in_0_7;
      end else if (10'h127 == _T_34[9:0]) begin
        image_0_295 <= io_pixelVal_in_0_6;
      end else if (10'h127 == _T_31[9:0]) begin
        image_0_295 <= io_pixelVal_in_0_5;
      end else if (10'h127 == _T_28[9:0]) begin
        image_0_295 <= io_pixelVal_in_0_4;
      end else if (10'h127 == _T_25[9:0]) begin
        image_0_295 <= io_pixelVal_in_0_3;
      end else if (10'h127 == _T_22[9:0]) begin
        image_0_295 <= io_pixelVal_in_0_2;
      end else if (10'h127 == _T_19[9:0]) begin
        image_0_295 <= io_pixelVal_in_0_1;
      end else if (10'h127 == _T_15[9:0]) begin
        image_0_295 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_296 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h128 == _T_37[9:0]) begin
        image_0_296 <= io_pixelVal_in_0_7;
      end else if (10'h128 == _T_34[9:0]) begin
        image_0_296 <= io_pixelVal_in_0_6;
      end else if (10'h128 == _T_31[9:0]) begin
        image_0_296 <= io_pixelVal_in_0_5;
      end else if (10'h128 == _T_28[9:0]) begin
        image_0_296 <= io_pixelVal_in_0_4;
      end else if (10'h128 == _T_25[9:0]) begin
        image_0_296 <= io_pixelVal_in_0_3;
      end else if (10'h128 == _T_22[9:0]) begin
        image_0_296 <= io_pixelVal_in_0_2;
      end else if (10'h128 == _T_19[9:0]) begin
        image_0_296 <= io_pixelVal_in_0_1;
      end else if (10'h128 == _T_15[9:0]) begin
        image_0_296 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_297 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h129 == _T_37[9:0]) begin
        image_0_297 <= io_pixelVal_in_0_7;
      end else if (10'h129 == _T_34[9:0]) begin
        image_0_297 <= io_pixelVal_in_0_6;
      end else if (10'h129 == _T_31[9:0]) begin
        image_0_297 <= io_pixelVal_in_0_5;
      end else if (10'h129 == _T_28[9:0]) begin
        image_0_297 <= io_pixelVal_in_0_4;
      end else if (10'h129 == _T_25[9:0]) begin
        image_0_297 <= io_pixelVal_in_0_3;
      end else if (10'h129 == _T_22[9:0]) begin
        image_0_297 <= io_pixelVal_in_0_2;
      end else if (10'h129 == _T_19[9:0]) begin
        image_0_297 <= io_pixelVal_in_0_1;
      end else if (10'h129 == _T_15[9:0]) begin
        image_0_297 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_298 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h12a == _T_37[9:0]) begin
        image_0_298 <= io_pixelVal_in_0_7;
      end else if (10'h12a == _T_34[9:0]) begin
        image_0_298 <= io_pixelVal_in_0_6;
      end else if (10'h12a == _T_31[9:0]) begin
        image_0_298 <= io_pixelVal_in_0_5;
      end else if (10'h12a == _T_28[9:0]) begin
        image_0_298 <= io_pixelVal_in_0_4;
      end else if (10'h12a == _T_25[9:0]) begin
        image_0_298 <= io_pixelVal_in_0_3;
      end else if (10'h12a == _T_22[9:0]) begin
        image_0_298 <= io_pixelVal_in_0_2;
      end else if (10'h12a == _T_19[9:0]) begin
        image_0_298 <= io_pixelVal_in_0_1;
      end else if (10'h12a == _T_15[9:0]) begin
        image_0_298 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_299 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h12b == _T_37[9:0]) begin
        image_0_299 <= io_pixelVal_in_0_7;
      end else if (10'h12b == _T_34[9:0]) begin
        image_0_299 <= io_pixelVal_in_0_6;
      end else if (10'h12b == _T_31[9:0]) begin
        image_0_299 <= io_pixelVal_in_0_5;
      end else if (10'h12b == _T_28[9:0]) begin
        image_0_299 <= io_pixelVal_in_0_4;
      end else if (10'h12b == _T_25[9:0]) begin
        image_0_299 <= io_pixelVal_in_0_3;
      end else if (10'h12b == _T_22[9:0]) begin
        image_0_299 <= io_pixelVal_in_0_2;
      end else if (10'h12b == _T_19[9:0]) begin
        image_0_299 <= io_pixelVal_in_0_1;
      end else if (10'h12b == _T_15[9:0]) begin
        image_0_299 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_300 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h12c == _T_37[9:0]) begin
        image_0_300 <= io_pixelVal_in_0_7;
      end else if (10'h12c == _T_34[9:0]) begin
        image_0_300 <= io_pixelVal_in_0_6;
      end else if (10'h12c == _T_31[9:0]) begin
        image_0_300 <= io_pixelVal_in_0_5;
      end else if (10'h12c == _T_28[9:0]) begin
        image_0_300 <= io_pixelVal_in_0_4;
      end else if (10'h12c == _T_25[9:0]) begin
        image_0_300 <= io_pixelVal_in_0_3;
      end else if (10'h12c == _T_22[9:0]) begin
        image_0_300 <= io_pixelVal_in_0_2;
      end else if (10'h12c == _T_19[9:0]) begin
        image_0_300 <= io_pixelVal_in_0_1;
      end else if (10'h12c == _T_15[9:0]) begin
        image_0_300 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_301 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h12d == _T_37[9:0]) begin
        image_0_301 <= io_pixelVal_in_0_7;
      end else if (10'h12d == _T_34[9:0]) begin
        image_0_301 <= io_pixelVal_in_0_6;
      end else if (10'h12d == _T_31[9:0]) begin
        image_0_301 <= io_pixelVal_in_0_5;
      end else if (10'h12d == _T_28[9:0]) begin
        image_0_301 <= io_pixelVal_in_0_4;
      end else if (10'h12d == _T_25[9:0]) begin
        image_0_301 <= io_pixelVal_in_0_3;
      end else if (10'h12d == _T_22[9:0]) begin
        image_0_301 <= io_pixelVal_in_0_2;
      end else if (10'h12d == _T_19[9:0]) begin
        image_0_301 <= io_pixelVal_in_0_1;
      end else if (10'h12d == _T_15[9:0]) begin
        image_0_301 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_302 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h12e == _T_37[9:0]) begin
        image_0_302 <= io_pixelVal_in_0_7;
      end else if (10'h12e == _T_34[9:0]) begin
        image_0_302 <= io_pixelVal_in_0_6;
      end else if (10'h12e == _T_31[9:0]) begin
        image_0_302 <= io_pixelVal_in_0_5;
      end else if (10'h12e == _T_28[9:0]) begin
        image_0_302 <= io_pixelVal_in_0_4;
      end else if (10'h12e == _T_25[9:0]) begin
        image_0_302 <= io_pixelVal_in_0_3;
      end else if (10'h12e == _T_22[9:0]) begin
        image_0_302 <= io_pixelVal_in_0_2;
      end else if (10'h12e == _T_19[9:0]) begin
        image_0_302 <= io_pixelVal_in_0_1;
      end else if (10'h12e == _T_15[9:0]) begin
        image_0_302 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_303 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h12f == _T_37[9:0]) begin
        image_0_303 <= io_pixelVal_in_0_7;
      end else if (10'h12f == _T_34[9:0]) begin
        image_0_303 <= io_pixelVal_in_0_6;
      end else if (10'h12f == _T_31[9:0]) begin
        image_0_303 <= io_pixelVal_in_0_5;
      end else if (10'h12f == _T_28[9:0]) begin
        image_0_303 <= io_pixelVal_in_0_4;
      end else if (10'h12f == _T_25[9:0]) begin
        image_0_303 <= io_pixelVal_in_0_3;
      end else if (10'h12f == _T_22[9:0]) begin
        image_0_303 <= io_pixelVal_in_0_2;
      end else if (10'h12f == _T_19[9:0]) begin
        image_0_303 <= io_pixelVal_in_0_1;
      end else if (10'h12f == _T_15[9:0]) begin
        image_0_303 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_304 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h130 == _T_37[9:0]) begin
        image_0_304 <= io_pixelVal_in_0_7;
      end else if (10'h130 == _T_34[9:0]) begin
        image_0_304 <= io_pixelVal_in_0_6;
      end else if (10'h130 == _T_31[9:0]) begin
        image_0_304 <= io_pixelVal_in_0_5;
      end else if (10'h130 == _T_28[9:0]) begin
        image_0_304 <= io_pixelVal_in_0_4;
      end else if (10'h130 == _T_25[9:0]) begin
        image_0_304 <= io_pixelVal_in_0_3;
      end else if (10'h130 == _T_22[9:0]) begin
        image_0_304 <= io_pixelVal_in_0_2;
      end else if (10'h130 == _T_19[9:0]) begin
        image_0_304 <= io_pixelVal_in_0_1;
      end else if (10'h130 == _T_15[9:0]) begin
        image_0_304 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_305 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h131 == _T_37[9:0]) begin
        image_0_305 <= io_pixelVal_in_0_7;
      end else if (10'h131 == _T_34[9:0]) begin
        image_0_305 <= io_pixelVal_in_0_6;
      end else if (10'h131 == _T_31[9:0]) begin
        image_0_305 <= io_pixelVal_in_0_5;
      end else if (10'h131 == _T_28[9:0]) begin
        image_0_305 <= io_pixelVal_in_0_4;
      end else if (10'h131 == _T_25[9:0]) begin
        image_0_305 <= io_pixelVal_in_0_3;
      end else if (10'h131 == _T_22[9:0]) begin
        image_0_305 <= io_pixelVal_in_0_2;
      end else if (10'h131 == _T_19[9:0]) begin
        image_0_305 <= io_pixelVal_in_0_1;
      end else if (10'h131 == _T_15[9:0]) begin
        image_0_305 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_306 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h132 == _T_37[9:0]) begin
        image_0_306 <= io_pixelVal_in_0_7;
      end else if (10'h132 == _T_34[9:0]) begin
        image_0_306 <= io_pixelVal_in_0_6;
      end else if (10'h132 == _T_31[9:0]) begin
        image_0_306 <= io_pixelVal_in_0_5;
      end else if (10'h132 == _T_28[9:0]) begin
        image_0_306 <= io_pixelVal_in_0_4;
      end else if (10'h132 == _T_25[9:0]) begin
        image_0_306 <= io_pixelVal_in_0_3;
      end else if (10'h132 == _T_22[9:0]) begin
        image_0_306 <= io_pixelVal_in_0_2;
      end else if (10'h132 == _T_19[9:0]) begin
        image_0_306 <= io_pixelVal_in_0_1;
      end else if (10'h132 == _T_15[9:0]) begin
        image_0_306 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_307 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h133 == _T_37[9:0]) begin
        image_0_307 <= io_pixelVal_in_0_7;
      end else if (10'h133 == _T_34[9:0]) begin
        image_0_307 <= io_pixelVal_in_0_6;
      end else if (10'h133 == _T_31[9:0]) begin
        image_0_307 <= io_pixelVal_in_0_5;
      end else if (10'h133 == _T_28[9:0]) begin
        image_0_307 <= io_pixelVal_in_0_4;
      end else if (10'h133 == _T_25[9:0]) begin
        image_0_307 <= io_pixelVal_in_0_3;
      end else if (10'h133 == _T_22[9:0]) begin
        image_0_307 <= io_pixelVal_in_0_2;
      end else if (10'h133 == _T_19[9:0]) begin
        image_0_307 <= io_pixelVal_in_0_1;
      end else if (10'h133 == _T_15[9:0]) begin
        image_0_307 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_308 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h134 == _T_37[9:0]) begin
        image_0_308 <= io_pixelVal_in_0_7;
      end else if (10'h134 == _T_34[9:0]) begin
        image_0_308 <= io_pixelVal_in_0_6;
      end else if (10'h134 == _T_31[9:0]) begin
        image_0_308 <= io_pixelVal_in_0_5;
      end else if (10'h134 == _T_28[9:0]) begin
        image_0_308 <= io_pixelVal_in_0_4;
      end else if (10'h134 == _T_25[9:0]) begin
        image_0_308 <= io_pixelVal_in_0_3;
      end else if (10'h134 == _T_22[9:0]) begin
        image_0_308 <= io_pixelVal_in_0_2;
      end else if (10'h134 == _T_19[9:0]) begin
        image_0_308 <= io_pixelVal_in_0_1;
      end else if (10'h134 == _T_15[9:0]) begin
        image_0_308 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_309 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h135 == _T_37[9:0]) begin
        image_0_309 <= io_pixelVal_in_0_7;
      end else if (10'h135 == _T_34[9:0]) begin
        image_0_309 <= io_pixelVal_in_0_6;
      end else if (10'h135 == _T_31[9:0]) begin
        image_0_309 <= io_pixelVal_in_0_5;
      end else if (10'h135 == _T_28[9:0]) begin
        image_0_309 <= io_pixelVal_in_0_4;
      end else if (10'h135 == _T_25[9:0]) begin
        image_0_309 <= io_pixelVal_in_0_3;
      end else if (10'h135 == _T_22[9:0]) begin
        image_0_309 <= io_pixelVal_in_0_2;
      end else if (10'h135 == _T_19[9:0]) begin
        image_0_309 <= io_pixelVal_in_0_1;
      end else if (10'h135 == _T_15[9:0]) begin
        image_0_309 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_310 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h136 == _T_37[9:0]) begin
        image_0_310 <= io_pixelVal_in_0_7;
      end else if (10'h136 == _T_34[9:0]) begin
        image_0_310 <= io_pixelVal_in_0_6;
      end else if (10'h136 == _T_31[9:0]) begin
        image_0_310 <= io_pixelVal_in_0_5;
      end else if (10'h136 == _T_28[9:0]) begin
        image_0_310 <= io_pixelVal_in_0_4;
      end else if (10'h136 == _T_25[9:0]) begin
        image_0_310 <= io_pixelVal_in_0_3;
      end else if (10'h136 == _T_22[9:0]) begin
        image_0_310 <= io_pixelVal_in_0_2;
      end else if (10'h136 == _T_19[9:0]) begin
        image_0_310 <= io_pixelVal_in_0_1;
      end else if (10'h136 == _T_15[9:0]) begin
        image_0_310 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_311 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h137 == _T_37[9:0]) begin
        image_0_311 <= io_pixelVal_in_0_7;
      end else if (10'h137 == _T_34[9:0]) begin
        image_0_311 <= io_pixelVal_in_0_6;
      end else if (10'h137 == _T_31[9:0]) begin
        image_0_311 <= io_pixelVal_in_0_5;
      end else if (10'h137 == _T_28[9:0]) begin
        image_0_311 <= io_pixelVal_in_0_4;
      end else if (10'h137 == _T_25[9:0]) begin
        image_0_311 <= io_pixelVal_in_0_3;
      end else if (10'h137 == _T_22[9:0]) begin
        image_0_311 <= io_pixelVal_in_0_2;
      end else if (10'h137 == _T_19[9:0]) begin
        image_0_311 <= io_pixelVal_in_0_1;
      end else if (10'h137 == _T_15[9:0]) begin
        image_0_311 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_312 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h138 == _T_37[9:0]) begin
        image_0_312 <= io_pixelVal_in_0_7;
      end else if (10'h138 == _T_34[9:0]) begin
        image_0_312 <= io_pixelVal_in_0_6;
      end else if (10'h138 == _T_31[9:0]) begin
        image_0_312 <= io_pixelVal_in_0_5;
      end else if (10'h138 == _T_28[9:0]) begin
        image_0_312 <= io_pixelVal_in_0_4;
      end else if (10'h138 == _T_25[9:0]) begin
        image_0_312 <= io_pixelVal_in_0_3;
      end else if (10'h138 == _T_22[9:0]) begin
        image_0_312 <= io_pixelVal_in_0_2;
      end else if (10'h138 == _T_19[9:0]) begin
        image_0_312 <= io_pixelVal_in_0_1;
      end else if (10'h138 == _T_15[9:0]) begin
        image_0_312 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_313 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h139 == _T_37[9:0]) begin
        image_0_313 <= io_pixelVal_in_0_7;
      end else if (10'h139 == _T_34[9:0]) begin
        image_0_313 <= io_pixelVal_in_0_6;
      end else if (10'h139 == _T_31[9:0]) begin
        image_0_313 <= io_pixelVal_in_0_5;
      end else if (10'h139 == _T_28[9:0]) begin
        image_0_313 <= io_pixelVal_in_0_4;
      end else if (10'h139 == _T_25[9:0]) begin
        image_0_313 <= io_pixelVal_in_0_3;
      end else if (10'h139 == _T_22[9:0]) begin
        image_0_313 <= io_pixelVal_in_0_2;
      end else if (10'h139 == _T_19[9:0]) begin
        image_0_313 <= io_pixelVal_in_0_1;
      end else if (10'h139 == _T_15[9:0]) begin
        image_0_313 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_314 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h13a == _T_37[9:0]) begin
        image_0_314 <= io_pixelVal_in_0_7;
      end else if (10'h13a == _T_34[9:0]) begin
        image_0_314 <= io_pixelVal_in_0_6;
      end else if (10'h13a == _T_31[9:0]) begin
        image_0_314 <= io_pixelVal_in_0_5;
      end else if (10'h13a == _T_28[9:0]) begin
        image_0_314 <= io_pixelVal_in_0_4;
      end else if (10'h13a == _T_25[9:0]) begin
        image_0_314 <= io_pixelVal_in_0_3;
      end else if (10'h13a == _T_22[9:0]) begin
        image_0_314 <= io_pixelVal_in_0_2;
      end else if (10'h13a == _T_19[9:0]) begin
        image_0_314 <= io_pixelVal_in_0_1;
      end else if (10'h13a == _T_15[9:0]) begin
        image_0_314 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_315 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h13b == _T_37[9:0]) begin
        image_0_315 <= io_pixelVal_in_0_7;
      end else if (10'h13b == _T_34[9:0]) begin
        image_0_315 <= io_pixelVal_in_0_6;
      end else if (10'h13b == _T_31[9:0]) begin
        image_0_315 <= io_pixelVal_in_0_5;
      end else if (10'h13b == _T_28[9:0]) begin
        image_0_315 <= io_pixelVal_in_0_4;
      end else if (10'h13b == _T_25[9:0]) begin
        image_0_315 <= io_pixelVal_in_0_3;
      end else if (10'h13b == _T_22[9:0]) begin
        image_0_315 <= io_pixelVal_in_0_2;
      end else if (10'h13b == _T_19[9:0]) begin
        image_0_315 <= io_pixelVal_in_0_1;
      end else if (10'h13b == _T_15[9:0]) begin
        image_0_315 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_316 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h13c == _T_37[9:0]) begin
        image_0_316 <= io_pixelVal_in_0_7;
      end else if (10'h13c == _T_34[9:0]) begin
        image_0_316 <= io_pixelVal_in_0_6;
      end else if (10'h13c == _T_31[9:0]) begin
        image_0_316 <= io_pixelVal_in_0_5;
      end else if (10'h13c == _T_28[9:0]) begin
        image_0_316 <= io_pixelVal_in_0_4;
      end else if (10'h13c == _T_25[9:0]) begin
        image_0_316 <= io_pixelVal_in_0_3;
      end else if (10'h13c == _T_22[9:0]) begin
        image_0_316 <= io_pixelVal_in_0_2;
      end else if (10'h13c == _T_19[9:0]) begin
        image_0_316 <= io_pixelVal_in_0_1;
      end else if (10'h13c == _T_15[9:0]) begin
        image_0_316 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_317 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h13d == _T_37[9:0]) begin
        image_0_317 <= io_pixelVal_in_0_7;
      end else if (10'h13d == _T_34[9:0]) begin
        image_0_317 <= io_pixelVal_in_0_6;
      end else if (10'h13d == _T_31[9:0]) begin
        image_0_317 <= io_pixelVal_in_0_5;
      end else if (10'h13d == _T_28[9:0]) begin
        image_0_317 <= io_pixelVal_in_0_4;
      end else if (10'h13d == _T_25[9:0]) begin
        image_0_317 <= io_pixelVal_in_0_3;
      end else if (10'h13d == _T_22[9:0]) begin
        image_0_317 <= io_pixelVal_in_0_2;
      end else if (10'h13d == _T_19[9:0]) begin
        image_0_317 <= io_pixelVal_in_0_1;
      end else if (10'h13d == _T_15[9:0]) begin
        image_0_317 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_318 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h13e == _T_37[9:0]) begin
        image_0_318 <= io_pixelVal_in_0_7;
      end else if (10'h13e == _T_34[9:0]) begin
        image_0_318 <= io_pixelVal_in_0_6;
      end else if (10'h13e == _T_31[9:0]) begin
        image_0_318 <= io_pixelVal_in_0_5;
      end else if (10'h13e == _T_28[9:0]) begin
        image_0_318 <= io_pixelVal_in_0_4;
      end else if (10'h13e == _T_25[9:0]) begin
        image_0_318 <= io_pixelVal_in_0_3;
      end else if (10'h13e == _T_22[9:0]) begin
        image_0_318 <= io_pixelVal_in_0_2;
      end else if (10'h13e == _T_19[9:0]) begin
        image_0_318 <= io_pixelVal_in_0_1;
      end else if (10'h13e == _T_15[9:0]) begin
        image_0_318 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_319 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h13f == _T_37[9:0]) begin
        image_0_319 <= io_pixelVal_in_0_7;
      end else if (10'h13f == _T_34[9:0]) begin
        image_0_319 <= io_pixelVal_in_0_6;
      end else if (10'h13f == _T_31[9:0]) begin
        image_0_319 <= io_pixelVal_in_0_5;
      end else if (10'h13f == _T_28[9:0]) begin
        image_0_319 <= io_pixelVal_in_0_4;
      end else if (10'h13f == _T_25[9:0]) begin
        image_0_319 <= io_pixelVal_in_0_3;
      end else if (10'h13f == _T_22[9:0]) begin
        image_0_319 <= io_pixelVal_in_0_2;
      end else if (10'h13f == _T_19[9:0]) begin
        image_0_319 <= io_pixelVal_in_0_1;
      end else if (10'h13f == _T_15[9:0]) begin
        image_0_319 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_320 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h140 == _T_37[9:0]) begin
        image_0_320 <= io_pixelVal_in_0_7;
      end else if (10'h140 == _T_34[9:0]) begin
        image_0_320 <= io_pixelVal_in_0_6;
      end else if (10'h140 == _T_31[9:0]) begin
        image_0_320 <= io_pixelVal_in_0_5;
      end else if (10'h140 == _T_28[9:0]) begin
        image_0_320 <= io_pixelVal_in_0_4;
      end else if (10'h140 == _T_25[9:0]) begin
        image_0_320 <= io_pixelVal_in_0_3;
      end else if (10'h140 == _T_22[9:0]) begin
        image_0_320 <= io_pixelVal_in_0_2;
      end else if (10'h140 == _T_19[9:0]) begin
        image_0_320 <= io_pixelVal_in_0_1;
      end else if (10'h140 == _T_15[9:0]) begin
        image_0_320 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_321 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h141 == _T_37[9:0]) begin
        image_0_321 <= io_pixelVal_in_0_7;
      end else if (10'h141 == _T_34[9:0]) begin
        image_0_321 <= io_pixelVal_in_0_6;
      end else if (10'h141 == _T_31[9:0]) begin
        image_0_321 <= io_pixelVal_in_0_5;
      end else if (10'h141 == _T_28[9:0]) begin
        image_0_321 <= io_pixelVal_in_0_4;
      end else if (10'h141 == _T_25[9:0]) begin
        image_0_321 <= io_pixelVal_in_0_3;
      end else if (10'h141 == _T_22[9:0]) begin
        image_0_321 <= io_pixelVal_in_0_2;
      end else if (10'h141 == _T_19[9:0]) begin
        image_0_321 <= io_pixelVal_in_0_1;
      end else if (10'h141 == _T_15[9:0]) begin
        image_0_321 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_322 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h142 == _T_37[9:0]) begin
        image_0_322 <= io_pixelVal_in_0_7;
      end else if (10'h142 == _T_34[9:0]) begin
        image_0_322 <= io_pixelVal_in_0_6;
      end else if (10'h142 == _T_31[9:0]) begin
        image_0_322 <= io_pixelVal_in_0_5;
      end else if (10'h142 == _T_28[9:0]) begin
        image_0_322 <= io_pixelVal_in_0_4;
      end else if (10'h142 == _T_25[9:0]) begin
        image_0_322 <= io_pixelVal_in_0_3;
      end else if (10'h142 == _T_22[9:0]) begin
        image_0_322 <= io_pixelVal_in_0_2;
      end else if (10'h142 == _T_19[9:0]) begin
        image_0_322 <= io_pixelVal_in_0_1;
      end else if (10'h142 == _T_15[9:0]) begin
        image_0_322 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_323 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h143 == _T_37[9:0]) begin
        image_0_323 <= io_pixelVal_in_0_7;
      end else if (10'h143 == _T_34[9:0]) begin
        image_0_323 <= io_pixelVal_in_0_6;
      end else if (10'h143 == _T_31[9:0]) begin
        image_0_323 <= io_pixelVal_in_0_5;
      end else if (10'h143 == _T_28[9:0]) begin
        image_0_323 <= io_pixelVal_in_0_4;
      end else if (10'h143 == _T_25[9:0]) begin
        image_0_323 <= io_pixelVal_in_0_3;
      end else if (10'h143 == _T_22[9:0]) begin
        image_0_323 <= io_pixelVal_in_0_2;
      end else if (10'h143 == _T_19[9:0]) begin
        image_0_323 <= io_pixelVal_in_0_1;
      end else if (10'h143 == _T_15[9:0]) begin
        image_0_323 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_324 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h144 == _T_37[9:0]) begin
        image_0_324 <= io_pixelVal_in_0_7;
      end else if (10'h144 == _T_34[9:0]) begin
        image_0_324 <= io_pixelVal_in_0_6;
      end else if (10'h144 == _T_31[9:0]) begin
        image_0_324 <= io_pixelVal_in_0_5;
      end else if (10'h144 == _T_28[9:0]) begin
        image_0_324 <= io_pixelVal_in_0_4;
      end else if (10'h144 == _T_25[9:0]) begin
        image_0_324 <= io_pixelVal_in_0_3;
      end else if (10'h144 == _T_22[9:0]) begin
        image_0_324 <= io_pixelVal_in_0_2;
      end else if (10'h144 == _T_19[9:0]) begin
        image_0_324 <= io_pixelVal_in_0_1;
      end else if (10'h144 == _T_15[9:0]) begin
        image_0_324 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_325 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h145 == _T_37[9:0]) begin
        image_0_325 <= io_pixelVal_in_0_7;
      end else if (10'h145 == _T_34[9:0]) begin
        image_0_325 <= io_pixelVal_in_0_6;
      end else if (10'h145 == _T_31[9:0]) begin
        image_0_325 <= io_pixelVal_in_0_5;
      end else if (10'h145 == _T_28[9:0]) begin
        image_0_325 <= io_pixelVal_in_0_4;
      end else if (10'h145 == _T_25[9:0]) begin
        image_0_325 <= io_pixelVal_in_0_3;
      end else if (10'h145 == _T_22[9:0]) begin
        image_0_325 <= io_pixelVal_in_0_2;
      end else if (10'h145 == _T_19[9:0]) begin
        image_0_325 <= io_pixelVal_in_0_1;
      end else if (10'h145 == _T_15[9:0]) begin
        image_0_325 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_326 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h146 == _T_37[9:0]) begin
        image_0_326 <= io_pixelVal_in_0_7;
      end else if (10'h146 == _T_34[9:0]) begin
        image_0_326 <= io_pixelVal_in_0_6;
      end else if (10'h146 == _T_31[9:0]) begin
        image_0_326 <= io_pixelVal_in_0_5;
      end else if (10'h146 == _T_28[9:0]) begin
        image_0_326 <= io_pixelVal_in_0_4;
      end else if (10'h146 == _T_25[9:0]) begin
        image_0_326 <= io_pixelVal_in_0_3;
      end else if (10'h146 == _T_22[9:0]) begin
        image_0_326 <= io_pixelVal_in_0_2;
      end else if (10'h146 == _T_19[9:0]) begin
        image_0_326 <= io_pixelVal_in_0_1;
      end else if (10'h146 == _T_15[9:0]) begin
        image_0_326 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_327 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h147 == _T_37[9:0]) begin
        image_0_327 <= io_pixelVal_in_0_7;
      end else if (10'h147 == _T_34[9:0]) begin
        image_0_327 <= io_pixelVal_in_0_6;
      end else if (10'h147 == _T_31[9:0]) begin
        image_0_327 <= io_pixelVal_in_0_5;
      end else if (10'h147 == _T_28[9:0]) begin
        image_0_327 <= io_pixelVal_in_0_4;
      end else if (10'h147 == _T_25[9:0]) begin
        image_0_327 <= io_pixelVal_in_0_3;
      end else if (10'h147 == _T_22[9:0]) begin
        image_0_327 <= io_pixelVal_in_0_2;
      end else if (10'h147 == _T_19[9:0]) begin
        image_0_327 <= io_pixelVal_in_0_1;
      end else if (10'h147 == _T_15[9:0]) begin
        image_0_327 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_328 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h148 == _T_37[9:0]) begin
        image_0_328 <= io_pixelVal_in_0_7;
      end else if (10'h148 == _T_34[9:0]) begin
        image_0_328 <= io_pixelVal_in_0_6;
      end else if (10'h148 == _T_31[9:0]) begin
        image_0_328 <= io_pixelVal_in_0_5;
      end else if (10'h148 == _T_28[9:0]) begin
        image_0_328 <= io_pixelVal_in_0_4;
      end else if (10'h148 == _T_25[9:0]) begin
        image_0_328 <= io_pixelVal_in_0_3;
      end else if (10'h148 == _T_22[9:0]) begin
        image_0_328 <= io_pixelVal_in_0_2;
      end else if (10'h148 == _T_19[9:0]) begin
        image_0_328 <= io_pixelVal_in_0_1;
      end else if (10'h148 == _T_15[9:0]) begin
        image_0_328 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_329 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h149 == _T_37[9:0]) begin
        image_0_329 <= io_pixelVal_in_0_7;
      end else if (10'h149 == _T_34[9:0]) begin
        image_0_329 <= io_pixelVal_in_0_6;
      end else if (10'h149 == _T_31[9:0]) begin
        image_0_329 <= io_pixelVal_in_0_5;
      end else if (10'h149 == _T_28[9:0]) begin
        image_0_329 <= io_pixelVal_in_0_4;
      end else if (10'h149 == _T_25[9:0]) begin
        image_0_329 <= io_pixelVal_in_0_3;
      end else if (10'h149 == _T_22[9:0]) begin
        image_0_329 <= io_pixelVal_in_0_2;
      end else if (10'h149 == _T_19[9:0]) begin
        image_0_329 <= io_pixelVal_in_0_1;
      end else if (10'h149 == _T_15[9:0]) begin
        image_0_329 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_330 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h14a == _T_37[9:0]) begin
        image_0_330 <= io_pixelVal_in_0_7;
      end else if (10'h14a == _T_34[9:0]) begin
        image_0_330 <= io_pixelVal_in_0_6;
      end else if (10'h14a == _T_31[9:0]) begin
        image_0_330 <= io_pixelVal_in_0_5;
      end else if (10'h14a == _T_28[9:0]) begin
        image_0_330 <= io_pixelVal_in_0_4;
      end else if (10'h14a == _T_25[9:0]) begin
        image_0_330 <= io_pixelVal_in_0_3;
      end else if (10'h14a == _T_22[9:0]) begin
        image_0_330 <= io_pixelVal_in_0_2;
      end else if (10'h14a == _T_19[9:0]) begin
        image_0_330 <= io_pixelVal_in_0_1;
      end else if (10'h14a == _T_15[9:0]) begin
        image_0_330 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_331 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h14b == _T_37[9:0]) begin
        image_0_331 <= io_pixelVal_in_0_7;
      end else if (10'h14b == _T_34[9:0]) begin
        image_0_331 <= io_pixelVal_in_0_6;
      end else if (10'h14b == _T_31[9:0]) begin
        image_0_331 <= io_pixelVal_in_0_5;
      end else if (10'h14b == _T_28[9:0]) begin
        image_0_331 <= io_pixelVal_in_0_4;
      end else if (10'h14b == _T_25[9:0]) begin
        image_0_331 <= io_pixelVal_in_0_3;
      end else if (10'h14b == _T_22[9:0]) begin
        image_0_331 <= io_pixelVal_in_0_2;
      end else if (10'h14b == _T_19[9:0]) begin
        image_0_331 <= io_pixelVal_in_0_1;
      end else if (10'h14b == _T_15[9:0]) begin
        image_0_331 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_332 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h14c == _T_37[9:0]) begin
        image_0_332 <= io_pixelVal_in_0_7;
      end else if (10'h14c == _T_34[9:0]) begin
        image_0_332 <= io_pixelVal_in_0_6;
      end else if (10'h14c == _T_31[9:0]) begin
        image_0_332 <= io_pixelVal_in_0_5;
      end else if (10'h14c == _T_28[9:0]) begin
        image_0_332 <= io_pixelVal_in_0_4;
      end else if (10'h14c == _T_25[9:0]) begin
        image_0_332 <= io_pixelVal_in_0_3;
      end else if (10'h14c == _T_22[9:0]) begin
        image_0_332 <= io_pixelVal_in_0_2;
      end else if (10'h14c == _T_19[9:0]) begin
        image_0_332 <= io_pixelVal_in_0_1;
      end else if (10'h14c == _T_15[9:0]) begin
        image_0_332 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_333 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h14d == _T_37[9:0]) begin
        image_0_333 <= io_pixelVal_in_0_7;
      end else if (10'h14d == _T_34[9:0]) begin
        image_0_333 <= io_pixelVal_in_0_6;
      end else if (10'h14d == _T_31[9:0]) begin
        image_0_333 <= io_pixelVal_in_0_5;
      end else if (10'h14d == _T_28[9:0]) begin
        image_0_333 <= io_pixelVal_in_0_4;
      end else if (10'h14d == _T_25[9:0]) begin
        image_0_333 <= io_pixelVal_in_0_3;
      end else if (10'h14d == _T_22[9:0]) begin
        image_0_333 <= io_pixelVal_in_0_2;
      end else if (10'h14d == _T_19[9:0]) begin
        image_0_333 <= io_pixelVal_in_0_1;
      end else if (10'h14d == _T_15[9:0]) begin
        image_0_333 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_334 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h14e == _T_37[9:0]) begin
        image_0_334 <= io_pixelVal_in_0_7;
      end else if (10'h14e == _T_34[9:0]) begin
        image_0_334 <= io_pixelVal_in_0_6;
      end else if (10'h14e == _T_31[9:0]) begin
        image_0_334 <= io_pixelVal_in_0_5;
      end else if (10'h14e == _T_28[9:0]) begin
        image_0_334 <= io_pixelVal_in_0_4;
      end else if (10'h14e == _T_25[9:0]) begin
        image_0_334 <= io_pixelVal_in_0_3;
      end else if (10'h14e == _T_22[9:0]) begin
        image_0_334 <= io_pixelVal_in_0_2;
      end else if (10'h14e == _T_19[9:0]) begin
        image_0_334 <= io_pixelVal_in_0_1;
      end else if (10'h14e == _T_15[9:0]) begin
        image_0_334 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_335 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h14f == _T_37[9:0]) begin
        image_0_335 <= io_pixelVal_in_0_7;
      end else if (10'h14f == _T_34[9:0]) begin
        image_0_335 <= io_pixelVal_in_0_6;
      end else if (10'h14f == _T_31[9:0]) begin
        image_0_335 <= io_pixelVal_in_0_5;
      end else if (10'h14f == _T_28[9:0]) begin
        image_0_335 <= io_pixelVal_in_0_4;
      end else if (10'h14f == _T_25[9:0]) begin
        image_0_335 <= io_pixelVal_in_0_3;
      end else if (10'h14f == _T_22[9:0]) begin
        image_0_335 <= io_pixelVal_in_0_2;
      end else if (10'h14f == _T_19[9:0]) begin
        image_0_335 <= io_pixelVal_in_0_1;
      end else if (10'h14f == _T_15[9:0]) begin
        image_0_335 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_336 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h150 == _T_37[9:0]) begin
        image_0_336 <= io_pixelVal_in_0_7;
      end else if (10'h150 == _T_34[9:0]) begin
        image_0_336 <= io_pixelVal_in_0_6;
      end else if (10'h150 == _T_31[9:0]) begin
        image_0_336 <= io_pixelVal_in_0_5;
      end else if (10'h150 == _T_28[9:0]) begin
        image_0_336 <= io_pixelVal_in_0_4;
      end else if (10'h150 == _T_25[9:0]) begin
        image_0_336 <= io_pixelVal_in_0_3;
      end else if (10'h150 == _T_22[9:0]) begin
        image_0_336 <= io_pixelVal_in_0_2;
      end else if (10'h150 == _T_19[9:0]) begin
        image_0_336 <= io_pixelVal_in_0_1;
      end else if (10'h150 == _T_15[9:0]) begin
        image_0_336 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_337 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h151 == _T_37[9:0]) begin
        image_0_337 <= io_pixelVal_in_0_7;
      end else if (10'h151 == _T_34[9:0]) begin
        image_0_337 <= io_pixelVal_in_0_6;
      end else if (10'h151 == _T_31[9:0]) begin
        image_0_337 <= io_pixelVal_in_0_5;
      end else if (10'h151 == _T_28[9:0]) begin
        image_0_337 <= io_pixelVal_in_0_4;
      end else if (10'h151 == _T_25[9:0]) begin
        image_0_337 <= io_pixelVal_in_0_3;
      end else if (10'h151 == _T_22[9:0]) begin
        image_0_337 <= io_pixelVal_in_0_2;
      end else if (10'h151 == _T_19[9:0]) begin
        image_0_337 <= io_pixelVal_in_0_1;
      end else if (10'h151 == _T_15[9:0]) begin
        image_0_337 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_338 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h152 == _T_37[9:0]) begin
        image_0_338 <= io_pixelVal_in_0_7;
      end else if (10'h152 == _T_34[9:0]) begin
        image_0_338 <= io_pixelVal_in_0_6;
      end else if (10'h152 == _T_31[9:0]) begin
        image_0_338 <= io_pixelVal_in_0_5;
      end else if (10'h152 == _T_28[9:0]) begin
        image_0_338 <= io_pixelVal_in_0_4;
      end else if (10'h152 == _T_25[9:0]) begin
        image_0_338 <= io_pixelVal_in_0_3;
      end else if (10'h152 == _T_22[9:0]) begin
        image_0_338 <= io_pixelVal_in_0_2;
      end else if (10'h152 == _T_19[9:0]) begin
        image_0_338 <= io_pixelVal_in_0_1;
      end else if (10'h152 == _T_15[9:0]) begin
        image_0_338 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_339 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h153 == _T_37[9:0]) begin
        image_0_339 <= io_pixelVal_in_0_7;
      end else if (10'h153 == _T_34[9:0]) begin
        image_0_339 <= io_pixelVal_in_0_6;
      end else if (10'h153 == _T_31[9:0]) begin
        image_0_339 <= io_pixelVal_in_0_5;
      end else if (10'h153 == _T_28[9:0]) begin
        image_0_339 <= io_pixelVal_in_0_4;
      end else if (10'h153 == _T_25[9:0]) begin
        image_0_339 <= io_pixelVal_in_0_3;
      end else if (10'h153 == _T_22[9:0]) begin
        image_0_339 <= io_pixelVal_in_0_2;
      end else if (10'h153 == _T_19[9:0]) begin
        image_0_339 <= io_pixelVal_in_0_1;
      end else if (10'h153 == _T_15[9:0]) begin
        image_0_339 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_340 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h154 == _T_37[9:0]) begin
        image_0_340 <= io_pixelVal_in_0_7;
      end else if (10'h154 == _T_34[9:0]) begin
        image_0_340 <= io_pixelVal_in_0_6;
      end else if (10'h154 == _T_31[9:0]) begin
        image_0_340 <= io_pixelVal_in_0_5;
      end else if (10'h154 == _T_28[9:0]) begin
        image_0_340 <= io_pixelVal_in_0_4;
      end else if (10'h154 == _T_25[9:0]) begin
        image_0_340 <= io_pixelVal_in_0_3;
      end else if (10'h154 == _T_22[9:0]) begin
        image_0_340 <= io_pixelVal_in_0_2;
      end else if (10'h154 == _T_19[9:0]) begin
        image_0_340 <= io_pixelVal_in_0_1;
      end else if (10'h154 == _T_15[9:0]) begin
        image_0_340 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_341 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h155 == _T_37[9:0]) begin
        image_0_341 <= io_pixelVal_in_0_7;
      end else if (10'h155 == _T_34[9:0]) begin
        image_0_341 <= io_pixelVal_in_0_6;
      end else if (10'h155 == _T_31[9:0]) begin
        image_0_341 <= io_pixelVal_in_0_5;
      end else if (10'h155 == _T_28[9:0]) begin
        image_0_341 <= io_pixelVal_in_0_4;
      end else if (10'h155 == _T_25[9:0]) begin
        image_0_341 <= io_pixelVal_in_0_3;
      end else if (10'h155 == _T_22[9:0]) begin
        image_0_341 <= io_pixelVal_in_0_2;
      end else if (10'h155 == _T_19[9:0]) begin
        image_0_341 <= io_pixelVal_in_0_1;
      end else if (10'h155 == _T_15[9:0]) begin
        image_0_341 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_342 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h156 == _T_37[9:0]) begin
        image_0_342 <= io_pixelVal_in_0_7;
      end else if (10'h156 == _T_34[9:0]) begin
        image_0_342 <= io_pixelVal_in_0_6;
      end else if (10'h156 == _T_31[9:0]) begin
        image_0_342 <= io_pixelVal_in_0_5;
      end else if (10'h156 == _T_28[9:0]) begin
        image_0_342 <= io_pixelVal_in_0_4;
      end else if (10'h156 == _T_25[9:0]) begin
        image_0_342 <= io_pixelVal_in_0_3;
      end else if (10'h156 == _T_22[9:0]) begin
        image_0_342 <= io_pixelVal_in_0_2;
      end else if (10'h156 == _T_19[9:0]) begin
        image_0_342 <= io_pixelVal_in_0_1;
      end else if (10'h156 == _T_15[9:0]) begin
        image_0_342 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_343 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h157 == _T_37[9:0]) begin
        image_0_343 <= io_pixelVal_in_0_7;
      end else if (10'h157 == _T_34[9:0]) begin
        image_0_343 <= io_pixelVal_in_0_6;
      end else if (10'h157 == _T_31[9:0]) begin
        image_0_343 <= io_pixelVal_in_0_5;
      end else if (10'h157 == _T_28[9:0]) begin
        image_0_343 <= io_pixelVal_in_0_4;
      end else if (10'h157 == _T_25[9:0]) begin
        image_0_343 <= io_pixelVal_in_0_3;
      end else if (10'h157 == _T_22[9:0]) begin
        image_0_343 <= io_pixelVal_in_0_2;
      end else if (10'h157 == _T_19[9:0]) begin
        image_0_343 <= io_pixelVal_in_0_1;
      end else if (10'h157 == _T_15[9:0]) begin
        image_0_343 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_344 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h158 == _T_37[9:0]) begin
        image_0_344 <= io_pixelVal_in_0_7;
      end else if (10'h158 == _T_34[9:0]) begin
        image_0_344 <= io_pixelVal_in_0_6;
      end else if (10'h158 == _T_31[9:0]) begin
        image_0_344 <= io_pixelVal_in_0_5;
      end else if (10'h158 == _T_28[9:0]) begin
        image_0_344 <= io_pixelVal_in_0_4;
      end else if (10'h158 == _T_25[9:0]) begin
        image_0_344 <= io_pixelVal_in_0_3;
      end else if (10'h158 == _T_22[9:0]) begin
        image_0_344 <= io_pixelVal_in_0_2;
      end else if (10'h158 == _T_19[9:0]) begin
        image_0_344 <= io_pixelVal_in_0_1;
      end else if (10'h158 == _T_15[9:0]) begin
        image_0_344 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_345 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h159 == _T_37[9:0]) begin
        image_0_345 <= io_pixelVal_in_0_7;
      end else if (10'h159 == _T_34[9:0]) begin
        image_0_345 <= io_pixelVal_in_0_6;
      end else if (10'h159 == _T_31[9:0]) begin
        image_0_345 <= io_pixelVal_in_0_5;
      end else if (10'h159 == _T_28[9:0]) begin
        image_0_345 <= io_pixelVal_in_0_4;
      end else if (10'h159 == _T_25[9:0]) begin
        image_0_345 <= io_pixelVal_in_0_3;
      end else if (10'h159 == _T_22[9:0]) begin
        image_0_345 <= io_pixelVal_in_0_2;
      end else if (10'h159 == _T_19[9:0]) begin
        image_0_345 <= io_pixelVal_in_0_1;
      end else if (10'h159 == _T_15[9:0]) begin
        image_0_345 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_346 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h15a == _T_37[9:0]) begin
        image_0_346 <= io_pixelVal_in_0_7;
      end else if (10'h15a == _T_34[9:0]) begin
        image_0_346 <= io_pixelVal_in_0_6;
      end else if (10'h15a == _T_31[9:0]) begin
        image_0_346 <= io_pixelVal_in_0_5;
      end else if (10'h15a == _T_28[9:0]) begin
        image_0_346 <= io_pixelVal_in_0_4;
      end else if (10'h15a == _T_25[9:0]) begin
        image_0_346 <= io_pixelVal_in_0_3;
      end else if (10'h15a == _T_22[9:0]) begin
        image_0_346 <= io_pixelVal_in_0_2;
      end else if (10'h15a == _T_19[9:0]) begin
        image_0_346 <= io_pixelVal_in_0_1;
      end else if (10'h15a == _T_15[9:0]) begin
        image_0_346 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_347 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h15b == _T_37[9:0]) begin
        image_0_347 <= io_pixelVal_in_0_7;
      end else if (10'h15b == _T_34[9:0]) begin
        image_0_347 <= io_pixelVal_in_0_6;
      end else if (10'h15b == _T_31[9:0]) begin
        image_0_347 <= io_pixelVal_in_0_5;
      end else if (10'h15b == _T_28[9:0]) begin
        image_0_347 <= io_pixelVal_in_0_4;
      end else if (10'h15b == _T_25[9:0]) begin
        image_0_347 <= io_pixelVal_in_0_3;
      end else if (10'h15b == _T_22[9:0]) begin
        image_0_347 <= io_pixelVal_in_0_2;
      end else if (10'h15b == _T_19[9:0]) begin
        image_0_347 <= io_pixelVal_in_0_1;
      end else if (10'h15b == _T_15[9:0]) begin
        image_0_347 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_348 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h15c == _T_37[9:0]) begin
        image_0_348 <= io_pixelVal_in_0_7;
      end else if (10'h15c == _T_34[9:0]) begin
        image_0_348 <= io_pixelVal_in_0_6;
      end else if (10'h15c == _T_31[9:0]) begin
        image_0_348 <= io_pixelVal_in_0_5;
      end else if (10'h15c == _T_28[9:0]) begin
        image_0_348 <= io_pixelVal_in_0_4;
      end else if (10'h15c == _T_25[9:0]) begin
        image_0_348 <= io_pixelVal_in_0_3;
      end else if (10'h15c == _T_22[9:0]) begin
        image_0_348 <= io_pixelVal_in_0_2;
      end else if (10'h15c == _T_19[9:0]) begin
        image_0_348 <= io_pixelVal_in_0_1;
      end else if (10'h15c == _T_15[9:0]) begin
        image_0_348 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_349 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h15d == _T_37[9:0]) begin
        image_0_349 <= io_pixelVal_in_0_7;
      end else if (10'h15d == _T_34[9:0]) begin
        image_0_349 <= io_pixelVal_in_0_6;
      end else if (10'h15d == _T_31[9:0]) begin
        image_0_349 <= io_pixelVal_in_0_5;
      end else if (10'h15d == _T_28[9:0]) begin
        image_0_349 <= io_pixelVal_in_0_4;
      end else if (10'h15d == _T_25[9:0]) begin
        image_0_349 <= io_pixelVal_in_0_3;
      end else if (10'h15d == _T_22[9:0]) begin
        image_0_349 <= io_pixelVal_in_0_2;
      end else if (10'h15d == _T_19[9:0]) begin
        image_0_349 <= io_pixelVal_in_0_1;
      end else if (10'h15d == _T_15[9:0]) begin
        image_0_349 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_350 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h15e == _T_37[9:0]) begin
        image_0_350 <= io_pixelVal_in_0_7;
      end else if (10'h15e == _T_34[9:0]) begin
        image_0_350 <= io_pixelVal_in_0_6;
      end else if (10'h15e == _T_31[9:0]) begin
        image_0_350 <= io_pixelVal_in_0_5;
      end else if (10'h15e == _T_28[9:0]) begin
        image_0_350 <= io_pixelVal_in_0_4;
      end else if (10'h15e == _T_25[9:0]) begin
        image_0_350 <= io_pixelVal_in_0_3;
      end else if (10'h15e == _T_22[9:0]) begin
        image_0_350 <= io_pixelVal_in_0_2;
      end else if (10'h15e == _T_19[9:0]) begin
        image_0_350 <= io_pixelVal_in_0_1;
      end else if (10'h15e == _T_15[9:0]) begin
        image_0_350 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_351 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h15f == _T_37[9:0]) begin
        image_0_351 <= io_pixelVal_in_0_7;
      end else if (10'h15f == _T_34[9:0]) begin
        image_0_351 <= io_pixelVal_in_0_6;
      end else if (10'h15f == _T_31[9:0]) begin
        image_0_351 <= io_pixelVal_in_0_5;
      end else if (10'h15f == _T_28[9:0]) begin
        image_0_351 <= io_pixelVal_in_0_4;
      end else if (10'h15f == _T_25[9:0]) begin
        image_0_351 <= io_pixelVal_in_0_3;
      end else if (10'h15f == _T_22[9:0]) begin
        image_0_351 <= io_pixelVal_in_0_2;
      end else if (10'h15f == _T_19[9:0]) begin
        image_0_351 <= io_pixelVal_in_0_1;
      end else if (10'h15f == _T_15[9:0]) begin
        image_0_351 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_352 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h160 == _T_37[9:0]) begin
        image_0_352 <= io_pixelVal_in_0_7;
      end else if (10'h160 == _T_34[9:0]) begin
        image_0_352 <= io_pixelVal_in_0_6;
      end else if (10'h160 == _T_31[9:0]) begin
        image_0_352 <= io_pixelVal_in_0_5;
      end else if (10'h160 == _T_28[9:0]) begin
        image_0_352 <= io_pixelVal_in_0_4;
      end else if (10'h160 == _T_25[9:0]) begin
        image_0_352 <= io_pixelVal_in_0_3;
      end else if (10'h160 == _T_22[9:0]) begin
        image_0_352 <= io_pixelVal_in_0_2;
      end else if (10'h160 == _T_19[9:0]) begin
        image_0_352 <= io_pixelVal_in_0_1;
      end else if (10'h160 == _T_15[9:0]) begin
        image_0_352 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_353 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h161 == _T_37[9:0]) begin
        image_0_353 <= io_pixelVal_in_0_7;
      end else if (10'h161 == _T_34[9:0]) begin
        image_0_353 <= io_pixelVal_in_0_6;
      end else if (10'h161 == _T_31[9:0]) begin
        image_0_353 <= io_pixelVal_in_0_5;
      end else if (10'h161 == _T_28[9:0]) begin
        image_0_353 <= io_pixelVal_in_0_4;
      end else if (10'h161 == _T_25[9:0]) begin
        image_0_353 <= io_pixelVal_in_0_3;
      end else if (10'h161 == _T_22[9:0]) begin
        image_0_353 <= io_pixelVal_in_0_2;
      end else if (10'h161 == _T_19[9:0]) begin
        image_0_353 <= io_pixelVal_in_0_1;
      end else if (10'h161 == _T_15[9:0]) begin
        image_0_353 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_354 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h162 == _T_37[9:0]) begin
        image_0_354 <= io_pixelVal_in_0_7;
      end else if (10'h162 == _T_34[9:0]) begin
        image_0_354 <= io_pixelVal_in_0_6;
      end else if (10'h162 == _T_31[9:0]) begin
        image_0_354 <= io_pixelVal_in_0_5;
      end else if (10'h162 == _T_28[9:0]) begin
        image_0_354 <= io_pixelVal_in_0_4;
      end else if (10'h162 == _T_25[9:0]) begin
        image_0_354 <= io_pixelVal_in_0_3;
      end else if (10'h162 == _T_22[9:0]) begin
        image_0_354 <= io_pixelVal_in_0_2;
      end else if (10'h162 == _T_19[9:0]) begin
        image_0_354 <= io_pixelVal_in_0_1;
      end else if (10'h162 == _T_15[9:0]) begin
        image_0_354 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_355 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h163 == _T_37[9:0]) begin
        image_0_355 <= io_pixelVal_in_0_7;
      end else if (10'h163 == _T_34[9:0]) begin
        image_0_355 <= io_pixelVal_in_0_6;
      end else if (10'h163 == _T_31[9:0]) begin
        image_0_355 <= io_pixelVal_in_0_5;
      end else if (10'h163 == _T_28[9:0]) begin
        image_0_355 <= io_pixelVal_in_0_4;
      end else if (10'h163 == _T_25[9:0]) begin
        image_0_355 <= io_pixelVal_in_0_3;
      end else if (10'h163 == _T_22[9:0]) begin
        image_0_355 <= io_pixelVal_in_0_2;
      end else if (10'h163 == _T_19[9:0]) begin
        image_0_355 <= io_pixelVal_in_0_1;
      end else if (10'h163 == _T_15[9:0]) begin
        image_0_355 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_356 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h164 == _T_37[9:0]) begin
        image_0_356 <= io_pixelVal_in_0_7;
      end else if (10'h164 == _T_34[9:0]) begin
        image_0_356 <= io_pixelVal_in_0_6;
      end else if (10'h164 == _T_31[9:0]) begin
        image_0_356 <= io_pixelVal_in_0_5;
      end else if (10'h164 == _T_28[9:0]) begin
        image_0_356 <= io_pixelVal_in_0_4;
      end else if (10'h164 == _T_25[9:0]) begin
        image_0_356 <= io_pixelVal_in_0_3;
      end else if (10'h164 == _T_22[9:0]) begin
        image_0_356 <= io_pixelVal_in_0_2;
      end else if (10'h164 == _T_19[9:0]) begin
        image_0_356 <= io_pixelVal_in_0_1;
      end else if (10'h164 == _T_15[9:0]) begin
        image_0_356 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_357 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h165 == _T_37[9:0]) begin
        image_0_357 <= io_pixelVal_in_0_7;
      end else if (10'h165 == _T_34[9:0]) begin
        image_0_357 <= io_pixelVal_in_0_6;
      end else if (10'h165 == _T_31[9:0]) begin
        image_0_357 <= io_pixelVal_in_0_5;
      end else if (10'h165 == _T_28[9:0]) begin
        image_0_357 <= io_pixelVal_in_0_4;
      end else if (10'h165 == _T_25[9:0]) begin
        image_0_357 <= io_pixelVal_in_0_3;
      end else if (10'h165 == _T_22[9:0]) begin
        image_0_357 <= io_pixelVal_in_0_2;
      end else if (10'h165 == _T_19[9:0]) begin
        image_0_357 <= io_pixelVal_in_0_1;
      end else if (10'h165 == _T_15[9:0]) begin
        image_0_357 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_358 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h166 == _T_37[9:0]) begin
        image_0_358 <= io_pixelVal_in_0_7;
      end else if (10'h166 == _T_34[9:0]) begin
        image_0_358 <= io_pixelVal_in_0_6;
      end else if (10'h166 == _T_31[9:0]) begin
        image_0_358 <= io_pixelVal_in_0_5;
      end else if (10'h166 == _T_28[9:0]) begin
        image_0_358 <= io_pixelVal_in_0_4;
      end else if (10'h166 == _T_25[9:0]) begin
        image_0_358 <= io_pixelVal_in_0_3;
      end else if (10'h166 == _T_22[9:0]) begin
        image_0_358 <= io_pixelVal_in_0_2;
      end else if (10'h166 == _T_19[9:0]) begin
        image_0_358 <= io_pixelVal_in_0_1;
      end else if (10'h166 == _T_15[9:0]) begin
        image_0_358 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_359 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h167 == _T_37[9:0]) begin
        image_0_359 <= io_pixelVal_in_0_7;
      end else if (10'h167 == _T_34[9:0]) begin
        image_0_359 <= io_pixelVal_in_0_6;
      end else if (10'h167 == _T_31[9:0]) begin
        image_0_359 <= io_pixelVal_in_0_5;
      end else if (10'h167 == _T_28[9:0]) begin
        image_0_359 <= io_pixelVal_in_0_4;
      end else if (10'h167 == _T_25[9:0]) begin
        image_0_359 <= io_pixelVal_in_0_3;
      end else if (10'h167 == _T_22[9:0]) begin
        image_0_359 <= io_pixelVal_in_0_2;
      end else if (10'h167 == _T_19[9:0]) begin
        image_0_359 <= io_pixelVal_in_0_1;
      end else if (10'h167 == _T_15[9:0]) begin
        image_0_359 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_360 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h168 == _T_37[9:0]) begin
        image_0_360 <= io_pixelVal_in_0_7;
      end else if (10'h168 == _T_34[9:0]) begin
        image_0_360 <= io_pixelVal_in_0_6;
      end else if (10'h168 == _T_31[9:0]) begin
        image_0_360 <= io_pixelVal_in_0_5;
      end else if (10'h168 == _T_28[9:0]) begin
        image_0_360 <= io_pixelVal_in_0_4;
      end else if (10'h168 == _T_25[9:0]) begin
        image_0_360 <= io_pixelVal_in_0_3;
      end else if (10'h168 == _T_22[9:0]) begin
        image_0_360 <= io_pixelVal_in_0_2;
      end else if (10'h168 == _T_19[9:0]) begin
        image_0_360 <= io_pixelVal_in_0_1;
      end else if (10'h168 == _T_15[9:0]) begin
        image_0_360 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_361 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h169 == _T_37[9:0]) begin
        image_0_361 <= io_pixelVal_in_0_7;
      end else if (10'h169 == _T_34[9:0]) begin
        image_0_361 <= io_pixelVal_in_0_6;
      end else if (10'h169 == _T_31[9:0]) begin
        image_0_361 <= io_pixelVal_in_0_5;
      end else if (10'h169 == _T_28[9:0]) begin
        image_0_361 <= io_pixelVal_in_0_4;
      end else if (10'h169 == _T_25[9:0]) begin
        image_0_361 <= io_pixelVal_in_0_3;
      end else if (10'h169 == _T_22[9:0]) begin
        image_0_361 <= io_pixelVal_in_0_2;
      end else if (10'h169 == _T_19[9:0]) begin
        image_0_361 <= io_pixelVal_in_0_1;
      end else if (10'h169 == _T_15[9:0]) begin
        image_0_361 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_362 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h16a == _T_37[9:0]) begin
        image_0_362 <= io_pixelVal_in_0_7;
      end else if (10'h16a == _T_34[9:0]) begin
        image_0_362 <= io_pixelVal_in_0_6;
      end else if (10'h16a == _T_31[9:0]) begin
        image_0_362 <= io_pixelVal_in_0_5;
      end else if (10'h16a == _T_28[9:0]) begin
        image_0_362 <= io_pixelVal_in_0_4;
      end else if (10'h16a == _T_25[9:0]) begin
        image_0_362 <= io_pixelVal_in_0_3;
      end else if (10'h16a == _T_22[9:0]) begin
        image_0_362 <= io_pixelVal_in_0_2;
      end else if (10'h16a == _T_19[9:0]) begin
        image_0_362 <= io_pixelVal_in_0_1;
      end else if (10'h16a == _T_15[9:0]) begin
        image_0_362 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_363 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h16b == _T_37[9:0]) begin
        image_0_363 <= io_pixelVal_in_0_7;
      end else if (10'h16b == _T_34[9:0]) begin
        image_0_363 <= io_pixelVal_in_0_6;
      end else if (10'h16b == _T_31[9:0]) begin
        image_0_363 <= io_pixelVal_in_0_5;
      end else if (10'h16b == _T_28[9:0]) begin
        image_0_363 <= io_pixelVal_in_0_4;
      end else if (10'h16b == _T_25[9:0]) begin
        image_0_363 <= io_pixelVal_in_0_3;
      end else if (10'h16b == _T_22[9:0]) begin
        image_0_363 <= io_pixelVal_in_0_2;
      end else if (10'h16b == _T_19[9:0]) begin
        image_0_363 <= io_pixelVal_in_0_1;
      end else if (10'h16b == _T_15[9:0]) begin
        image_0_363 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_364 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h16c == _T_37[9:0]) begin
        image_0_364 <= io_pixelVal_in_0_7;
      end else if (10'h16c == _T_34[9:0]) begin
        image_0_364 <= io_pixelVal_in_0_6;
      end else if (10'h16c == _T_31[9:0]) begin
        image_0_364 <= io_pixelVal_in_0_5;
      end else if (10'h16c == _T_28[9:0]) begin
        image_0_364 <= io_pixelVal_in_0_4;
      end else if (10'h16c == _T_25[9:0]) begin
        image_0_364 <= io_pixelVal_in_0_3;
      end else if (10'h16c == _T_22[9:0]) begin
        image_0_364 <= io_pixelVal_in_0_2;
      end else if (10'h16c == _T_19[9:0]) begin
        image_0_364 <= io_pixelVal_in_0_1;
      end else if (10'h16c == _T_15[9:0]) begin
        image_0_364 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_365 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h16d == _T_37[9:0]) begin
        image_0_365 <= io_pixelVal_in_0_7;
      end else if (10'h16d == _T_34[9:0]) begin
        image_0_365 <= io_pixelVal_in_0_6;
      end else if (10'h16d == _T_31[9:0]) begin
        image_0_365 <= io_pixelVal_in_0_5;
      end else if (10'h16d == _T_28[9:0]) begin
        image_0_365 <= io_pixelVal_in_0_4;
      end else if (10'h16d == _T_25[9:0]) begin
        image_0_365 <= io_pixelVal_in_0_3;
      end else if (10'h16d == _T_22[9:0]) begin
        image_0_365 <= io_pixelVal_in_0_2;
      end else if (10'h16d == _T_19[9:0]) begin
        image_0_365 <= io_pixelVal_in_0_1;
      end else if (10'h16d == _T_15[9:0]) begin
        image_0_365 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_366 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h16e == _T_37[9:0]) begin
        image_0_366 <= io_pixelVal_in_0_7;
      end else if (10'h16e == _T_34[9:0]) begin
        image_0_366 <= io_pixelVal_in_0_6;
      end else if (10'h16e == _T_31[9:0]) begin
        image_0_366 <= io_pixelVal_in_0_5;
      end else if (10'h16e == _T_28[9:0]) begin
        image_0_366 <= io_pixelVal_in_0_4;
      end else if (10'h16e == _T_25[9:0]) begin
        image_0_366 <= io_pixelVal_in_0_3;
      end else if (10'h16e == _T_22[9:0]) begin
        image_0_366 <= io_pixelVal_in_0_2;
      end else if (10'h16e == _T_19[9:0]) begin
        image_0_366 <= io_pixelVal_in_0_1;
      end else if (10'h16e == _T_15[9:0]) begin
        image_0_366 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_367 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h16f == _T_37[9:0]) begin
        image_0_367 <= io_pixelVal_in_0_7;
      end else if (10'h16f == _T_34[9:0]) begin
        image_0_367 <= io_pixelVal_in_0_6;
      end else if (10'h16f == _T_31[9:0]) begin
        image_0_367 <= io_pixelVal_in_0_5;
      end else if (10'h16f == _T_28[9:0]) begin
        image_0_367 <= io_pixelVal_in_0_4;
      end else if (10'h16f == _T_25[9:0]) begin
        image_0_367 <= io_pixelVal_in_0_3;
      end else if (10'h16f == _T_22[9:0]) begin
        image_0_367 <= io_pixelVal_in_0_2;
      end else if (10'h16f == _T_19[9:0]) begin
        image_0_367 <= io_pixelVal_in_0_1;
      end else if (10'h16f == _T_15[9:0]) begin
        image_0_367 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_368 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h170 == _T_37[9:0]) begin
        image_0_368 <= io_pixelVal_in_0_7;
      end else if (10'h170 == _T_34[9:0]) begin
        image_0_368 <= io_pixelVal_in_0_6;
      end else if (10'h170 == _T_31[9:0]) begin
        image_0_368 <= io_pixelVal_in_0_5;
      end else if (10'h170 == _T_28[9:0]) begin
        image_0_368 <= io_pixelVal_in_0_4;
      end else if (10'h170 == _T_25[9:0]) begin
        image_0_368 <= io_pixelVal_in_0_3;
      end else if (10'h170 == _T_22[9:0]) begin
        image_0_368 <= io_pixelVal_in_0_2;
      end else if (10'h170 == _T_19[9:0]) begin
        image_0_368 <= io_pixelVal_in_0_1;
      end else if (10'h170 == _T_15[9:0]) begin
        image_0_368 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_369 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h171 == _T_37[9:0]) begin
        image_0_369 <= io_pixelVal_in_0_7;
      end else if (10'h171 == _T_34[9:0]) begin
        image_0_369 <= io_pixelVal_in_0_6;
      end else if (10'h171 == _T_31[9:0]) begin
        image_0_369 <= io_pixelVal_in_0_5;
      end else if (10'h171 == _T_28[9:0]) begin
        image_0_369 <= io_pixelVal_in_0_4;
      end else if (10'h171 == _T_25[9:0]) begin
        image_0_369 <= io_pixelVal_in_0_3;
      end else if (10'h171 == _T_22[9:0]) begin
        image_0_369 <= io_pixelVal_in_0_2;
      end else if (10'h171 == _T_19[9:0]) begin
        image_0_369 <= io_pixelVal_in_0_1;
      end else if (10'h171 == _T_15[9:0]) begin
        image_0_369 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_370 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h172 == _T_37[9:0]) begin
        image_0_370 <= io_pixelVal_in_0_7;
      end else if (10'h172 == _T_34[9:0]) begin
        image_0_370 <= io_pixelVal_in_0_6;
      end else if (10'h172 == _T_31[9:0]) begin
        image_0_370 <= io_pixelVal_in_0_5;
      end else if (10'h172 == _T_28[9:0]) begin
        image_0_370 <= io_pixelVal_in_0_4;
      end else if (10'h172 == _T_25[9:0]) begin
        image_0_370 <= io_pixelVal_in_0_3;
      end else if (10'h172 == _T_22[9:0]) begin
        image_0_370 <= io_pixelVal_in_0_2;
      end else if (10'h172 == _T_19[9:0]) begin
        image_0_370 <= io_pixelVal_in_0_1;
      end else if (10'h172 == _T_15[9:0]) begin
        image_0_370 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_371 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h173 == _T_37[9:0]) begin
        image_0_371 <= io_pixelVal_in_0_7;
      end else if (10'h173 == _T_34[9:0]) begin
        image_0_371 <= io_pixelVal_in_0_6;
      end else if (10'h173 == _T_31[9:0]) begin
        image_0_371 <= io_pixelVal_in_0_5;
      end else if (10'h173 == _T_28[9:0]) begin
        image_0_371 <= io_pixelVal_in_0_4;
      end else if (10'h173 == _T_25[9:0]) begin
        image_0_371 <= io_pixelVal_in_0_3;
      end else if (10'h173 == _T_22[9:0]) begin
        image_0_371 <= io_pixelVal_in_0_2;
      end else if (10'h173 == _T_19[9:0]) begin
        image_0_371 <= io_pixelVal_in_0_1;
      end else if (10'h173 == _T_15[9:0]) begin
        image_0_371 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_372 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h174 == _T_37[9:0]) begin
        image_0_372 <= io_pixelVal_in_0_7;
      end else if (10'h174 == _T_34[9:0]) begin
        image_0_372 <= io_pixelVal_in_0_6;
      end else if (10'h174 == _T_31[9:0]) begin
        image_0_372 <= io_pixelVal_in_0_5;
      end else if (10'h174 == _T_28[9:0]) begin
        image_0_372 <= io_pixelVal_in_0_4;
      end else if (10'h174 == _T_25[9:0]) begin
        image_0_372 <= io_pixelVal_in_0_3;
      end else if (10'h174 == _T_22[9:0]) begin
        image_0_372 <= io_pixelVal_in_0_2;
      end else if (10'h174 == _T_19[9:0]) begin
        image_0_372 <= io_pixelVal_in_0_1;
      end else if (10'h174 == _T_15[9:0]) begin
        image_0_372 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_373 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h175 == _T_37[9:0]) begin
        image_0_373 <= io_pixelVal_in_0_7;
      end else if (10'h175 == _T_34[9:0]) begin
        image_0_373 <= io_pixelVal_in_0_6;
      end else if (10'h175 == _T_31[9:0]) begin
        image_0_373 <= io_pixelVal_in_0_5;
      end else if (10'h175 == _T_28[9:0]) begin
        image_0_373 <= io_pixelVal_in_0_4;
      end else if (10'h175 == _T_25[9:0]) begin
        image_0_373 <= io_pixelVal_in_0_3;
      end else if (10'h175 == _T_22[9:0]) begin
        image_0_373 <= io_pixelVal_in_0_2;
      end else if (10'h175 == _T_19[9:0]) begin
        image_0_373 <= io_pixelVal_in_0_1;
      end else if (10'h175 == _T_15[9:0]) begin
        image_0_373 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_374 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h176 == _T_37[9:0]) begin
        image_0_374 <= io_pixelVal_in_0_7;
      end else if (10'h176 == _T_34[9:0]) begin
        image_0_374 <= io_pixelVal_in_0_6;
      end else if (10'h176 == _T_31[9:0]) begin
        image_0_374 <= io_pixelVal_in_0_5;
      end else if (10'h176 == _T_28[9:0]) begin
        image_0_374 <= io_pixelVal_in_0_4;
      end else if (10'h176 == _T_25[9:0]) begin
        image_0_374 <= io_pixelVal_in_0_3;
      end else if (10'h176 == _T_22[9:0]) begin
        image_0_374 <= io_pixelVal_in_0_2;
      end else if (10'h176 == _T_19[9:0]) begin
        image_0_374 <= io_pixelVal_in_0_1;
      end else if (10'h176 == _T_15[9:0]) begin
        image_0_374 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_375 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h177 == _T_37[9:0]) begin
        image_0_375 <= io_pixelVal_in_0_7;
      end else if (10'h177 == _T_34[9:0]) begin
        image_0_375 <= io_pixelVal_in_0_6;
      end else if (10'h177 == _T_31[9:0]) begin
        image_0_375 <= io_pixelVal_in_0_5;
      end else if (10'h177 == _T_28[9:0]) begin
        image_0_375 <= io_pixelVal_in_0_4;
      end else if (10'h177 == _T_25[9:0]) begin
        image_0_375 <= io_pixelVal_in_0_3;
      end else if (10'h177 == _T_22[9:0]) begin
        image_0_375 <= io_pixelVal_in_0_2;
      end else if (10'h177 == _T_19[9:0]) begin
        image_0_375 <= io_pixelVal_in_0_1;
      end else if (10'h177 == _T_15[9:0]) begin
        image_0_375 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_376 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h178 == _T_37[9:0]) begin
        image_0_376 <= io_pixelVal_in_0_7;
      end else if (10'h178 == _T_34[9:0]) begin
        image_0_376 <= io_pixelVal_in_0_6;
      end else if (10'h178 == _T_31[9:0]) begin
        image_0_376 <= io_pixelVal_in_0_5;
      end else if (10'h178 == _T_28[9:0]) begin
        image_0_376 <= io_pixelVal_in_0_4;
      end else if (10'h178 == _T_25[9:0]) begin
        image_0_376 <= io_pixelVal_in_0_3;
      end else if (10'h178 == _T_22[9:0]) begin
        image_0_376 <= io_pixelVal_in_0_2;
      end else if (10'h178 == _T_19[9:0]) begin
        image_0_376 <= io_pixelVal_in_0_1;
      end else if (10'h178 == _T_15[9:0]) begin
        image_0_376 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_377 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h179 == _T_37[9:0]) begin
        image_0_377 <= io_pixelVal_in_0_7;
      end else if (10'h179 == _T_34[9:0]) begin
        image_0_377 <= io_pixelVal_in_0_6;
      end else if (10'h179 == _T_31[9:0]) begin
        image_0_377 <= io_pixelVal_in_0_5;
      end else if (10'h179 == _T_28[9:0]) begin
        image_0_377 <= io_pixelVal_in_0_4;
      end else if (10'h179 == _T_25[9:0]) begin
        image_0_377 <= io_pixelVal_in_0_3;
      end else if (10'h179 == _T_22[9:0]) begin
        image_0_377 <= io_pixelVal_in_0_2;
      end else if (10'h179 == _T_19[9:0]) begin
        image_0_377 <= io_pixelVal_in_0_1;
      end else if (10'h179 == _T_15[9:0]) begin
        image_0_377 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_378 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h17a == _T_37[9:0]) begin
        image_0_378 <= io_pixelVal_in_0_7;
      end else if (10'h17a == _T_34[9:0]) begin
        image_0_378 <= io_pixelVal_in_0_6;
      end else if (10'h17a == _T_31[9:0]) begin
        image_0_378 <= io_pixelVal_in_0_5;
      end else if (10'h17a == _T_28[9:0]) begin
        image_0_378 <= io_pixelVal_in_0_4;
      end else if (10'h17a == _T_25[9:0]) begin
        image_0_378 <= io_pixelVal_in_0_3;
      end else if (10'h17a == _T_22[9:0]) begin
        image_0_378 <= io_pixelVal_in_0_2;
      end else if (10'h17a == _T_19[9:0]) begin
        image_0_378 <= io_pixelVal_in_0_1;
      end else if (10'h17a == _T_15[9:0]) begin
        image_0_378 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_379 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h17b == _T_37[9:0]) begin
        image_0_379 <= io_pixelVal_in_0_7;
      end else if (10'h17b == _T_34[9:0]) begin
        image_0_379 <= io_pixelVal_in_0_6;
      end else if (10'h17b == _T_31[9:0]) begin
        image_0_379 <= io_pixelVal_in_0_5;
      end else if (10'h17b == _T_28[9:0]) begin
        image_0_379 <= io_pixelVal_in_0_4;
      end else if (10'h17b == _T_25[9:0]) begin
        image_0_379 <= io_pixelVal_in_0_3;
      end else if (10'h17b == _T_22[9:0]) begin
        image_0_379 <= io_pixelVal_in_0_2;
      end else if (10'h17b == _T_19[9:0]) begin
        image_0_379 <= io_pixelVal_in_0_1;
      end else if (10'h17b == _T_15[9:0]) begin
        image_0_379 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_380 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h17c == _T_37[9:0]) begin
        image_0_380 <= io_pixelVal_in_0_7;
      end else if (10'h17c == _T_34[9:0]) begin
        image_0_380 <= io_pixelVal_in_0_6;
      end else if (10'h17c == _T_31[9:0]) begin
        image_0_380 <= io_pixelVal_in_0_5;
      end else if (10'h17c == _T_28[9:0]) begin
        image_0_380 <= io_pixelVal_in_0_4;
      end else if (10'h17c == _T_25[9:0]) begin
        image_0_380 <= io_pixelVal_in_0_3;
      end else if (10'h17c == _T_22[9:0]) begin
        image_0_380 <= io_pixelVal_in_0_2;
      end else if (10'h17c == _T_19[9:0]) begin
        image_0_380 <= io_pixelVal_in_0_1;
      end else if (10'h17c == _T_15[9:0]) begin
        image_0_380 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_381 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h17d == _T_37[9:0]) begin
        image_0_381 <= io_pixelVal_in_0_7;
      end else if (10'h17d == _T_34[9:0]) begin
        image_0_381 <= io_pixelVal_in_0_6;
      end else if (10'h17d == _T_31[9:0]) begin
        image_0_381 <= io_pixelVal_in_0_5;
      end else if (10'h17d == _T_28[9:0]) begin
        image_0_381 <= io_pixelVal_in_0_4;
      end else if (10'h17d == _T_25[9:0]) begin
        image_0_381 <= io_pixelVal_in_0_3;
      end else if (10'h17d == _T_22[9:0]) begin
        image_0_381 <= io_pixelVal_in_0_2;
      end else if (10'h17d == _T_19[9:0]) begin
        image_0_381 <= io_pixelVal_in_0_1;
      end else if (10'h17d == _T_15[9:0]) begin
        image_0_381 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_382 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h17e == _T_37[9:0]) begin
        image_0_382 <= io_pixelVal_in_0_7;
      end else if (10'h17e == _T_34[9:0]) begin
        image_0_382 <= io_pixelVal_in_0_6;
      end else if (10'h17e == _T_31[9:0]) begin
        image_0_382 <= io_pixelVal_in_0_5;
      end else if (10'h17e == _T_28[9:0]) begin
        image_0_382 <= io_pixelVal_in_0_4;
      end else if (10'h17e == _T_25[9:0]) begin
        image_0_382 <= io_pixelVal_in_0_3;
      end else if (10'h17e == _T_22[9:0]) begin
        image_0_382 <= io_pixelVal_in_0_2;
      end else if (10'h17e == _T_19[9:0]) begin
        image_0_382 <= io_pixelVal_in_0_1;
      end else if (10'h17e == _T_15[9:0]) begin
        image_0_382 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_383 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h17f == _T_37[9:0]) begin
        image_0_383 <= io_pixelVal_in_0_7;
      end else if (10'h17f == _T_34[9:0]) begin
        image_0_383 <= io_pixelVal_in_0_6;
      end else if (10'h17f == _T_31[9:0]) begin
        image_0_383 <= io_pixelVal_in_0_5;
      end else if (10'h17f == _T_28[9:0]) begin
        image_0_383 <= io_pixelVal_in_0_4;
      end else if (10'h17f == _T_25[9:0]) begin
        image_0_383 <= io_pixelVal_in_0_3;
      end else if (10'h17f == _T_22[9:0]) begin
        image_0_383 <= io_pixelVal_in_0_2;
      end else if (10'h17f == _T_19[9:0]) begin
        image_0_383 <= io_pixelVal_in_0_1;
      end else if (10'h17f == _T_15[9:0]) begin
        image_0_383 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_384 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h180 == _T_37[9:0]) begin
        image_0_384 <= io_pixelVal_in_0_7;
      end else if (10'h180 == _T_34[9:0]) begin
        image_0_384 <= io_pixelVal_in_0_6;
      end else if (10'h180 == _T_31[9:0]) begin
        image_0_384 <= io_pixelVal_in_0_5;
      end else if (10'h180 == _T_28[9:0]) begin
        image_0_384 <= io_pixelVal_in_0_4;
      end else if (10'h180 == _T_25[9:0]) begin
        image_0_384 <= io_pixelVal_in_0_3;
      end else if (10'h180 == _T_22[9:0]) begin
        image_0_384 <= io_pixelVal_in_0_2;
      end else if (10'h180 == _T_19[9:0]) begin
        image_0_384 <= io_pixelVal_in_0_1;
      end else if (10'h180 == _T_15[9:0]) begin
        image_0_384 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_385 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h181 == _T_37[9:0]) begin
        image_0_385 <= io_pixelVal_in_0_7;
      end else if (10'h181 == _T_34[9:0]) begin
        image_0_385 <= io_pixelVal_in_0_6;
      end else if (10'h181 == _T_31[9:0]) begin
        image_0_385 <= io_pixelVal_in_0_5;
      end else if (10'h181 == _T_28[9:0]) begin
        image_0_385 <= io_pixelVal_in_0_4;
      end else if (10'h181 == _T_25[9:0]) begin
        image_0_385 <= io_pixelVal_in_0_3;
      end else if (10'h181 == _T_22[9:0]) begin
        image_0_385 <= io_pixelVal_in_0_2;
      end else if (10'h181 == _T_19[9:0]) begin
        image_0_385 <= io_pixelVal_in_0_1;
      end else if (10'h181 == _T_15[9:0]) begin
        image_0_385 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_386 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h182 == _T_37[9:0]) begin
        image_0_386 <= io_pixelVal_in_0_7;
      end else if (10'h182 == _T_34[9:0]) begin
        image_0_386 <= io_pixelVal_in_0_6;
      end else if (10'h182 == _T_31[9:0]) begin
        image_0_386 <= io_pixelVal_in_0_5;
      end else if (10'h182 == _T_28[9:0]) begin
        image_0_386 <= io_pixelVal_in_0_4;
      end else if (10'h182 == _T_25[9:0]) begin
        image_0_386 <= io_pixelVal_in_0_3;
      end else if (10'h182 == _T_22[9:0]) begin
        image_0_386 <= io_pixelVal_in_0_2;
      end else if (10'h182 == _T_19[9:0]) begin
        image_0_386 <= io_pixelVal_in_0_1;
      end else if (10'h182 == _T_15[9:0]) begin
        image_0_386 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_387 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h183 == _T_37[9:0]) begin
        image_0_387 <= io_pixelVal_in_0_7;
      end else if (10'h183 == _T_34[9:0]) begin
        image_0_387 <= io_pixelVal_in_0_6;
      end else if (10'h183 == _T_31[9:0]) begin
        image_0_387 <= io_pixelVal_in_0_5;
      end else if (10'h183 == _T_28[9:0]) begin
        image_0_387 <= io_pixelVal_in_0_4;
      end else if (10'h183 == _T_25[9:0]) begin
        image_0_387 <= io_pixelVal_in_0_3;
      end else if (10'h183 == _T_22[9:0]) begin
        image_0_387 <= io_pixelVal_in_0_2;
      end else if (10'h183 == _T_19[9:0]) begin
        image_0_387 <= io_pixelVal_in_0_1;
      end else if (10'h183 == _T_15[9:0]) begin
        image_0_387 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_388 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h184 == _T_37[9:0]) begin
        image_0_388 <= io_pixelVal_in_0_7;
      end else if (10'h184 == _T_34[9:0]) begin
        image_0_388 <= io_pixelVal_in_0_6;
      end else if (10'h184 == _T_31[9:0]) begin
        image_0_388 <= io_pixelVal_in_0_5;
      end else if (10'h184 == _T_28[9:0]) begin
        image_0_388 <= io_pixelVal_in_0_4;
      end else if (10'h184 == _T_25[9:0]) begin
        image_0_388 <= io_pixelVal_in_0_3;
      end else if (10'h184 == _T_22[9:0]) begin
        image_0_388 <= io_pixelVal_in_0_2;
      end else if (10'h184 == _T_19[9:0]) begin
        image_0_388 <= io_pixelVal_in_0_1;
      end else if (10'h184 == _T_15[9:0]) begin
        image_0_388 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_389 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h185 == _T_37[9:0]) begin
        image_0_389 <= io_pixelVal_in_0_7;
      end else if (10'h185 == _T_34[9:0]) begin
        image_0_389 <= io_pixelVal_in_0_6;
      end else if (10'h185 == _T_31[9:0]) begin
        image_0_389 <= io_pixelVal_in_0_5;
      end else if (10'h185 == _T_28[9:0]) begin
        image_0_389 <= io_pixelVal_in_0_4;
      end else if (10'h185 == _T_25[9:0]) begin
        image_0_389 <= io_pixelVal_in_0_3;
      end else if (10'h185 == _T_22[9:0]) begin
        image_0_389 <= io_pixelVal_in_0_2;
      end else if (10'h185 == _T_19[9:0]) begin
        image_0_389 <= io_pixelVal_in_0_1;
      end else if (10'h185 == _T_15[9:0]) begin
        image_0_389 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_390 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h186 == _T_37[9:0]) begin
        image_0_390 <= io_pixelVal_in_0_7;
      end else if (10'h186 == _T_34[9:0]) begin
        image_0_390 <= io_pixelVal_in_0_6;
      end else if (10'h186 == _T_31[9:0]) begin
        image_0_390 <= io_pixelVal_in_0_5;
      end else if (10'h186 == _T_28[9:0]) begin
        image_0_390 <= io_pixelVal_in_0_4;
      end else if (10'h186 == _T_25[9:0]) begin
        image_0_390 <= io_pixelVal_in_0_3;
      end else if (10'h186 == _T_22[9:0]) begin
        image_0_390 <= io_pixelVal_in_0_2;
      end else if (10'h186 == _T_19[9:0]) begin
        image_0_390 <= io_pixelVal_in_0_1;
      end else if (10'h186 == _T_15[9:0]) begin
        image_0_390 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_391 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h187 == _T_37[9:0]) begin
        image_0_391 <= io_pixelVal_in_0_7;
      end else if (10'h187 == _T_34[9:0]) begin
        image_0_391 <= io_pixelVal_in_0_6;
      end else if (10'h187 == _T_31[9:0]) begin
        image_0_391 <= io_pixelVal_in_0_5;
      end else if (10'h187 == _T_28[9:0]) begin
        image_0_391 <= io_pixelVal_in_0_4;
      end else if (10'h187 == _T_25[9:0]) begin
        image_0_391 <= io_pixelVal_in_0_3;
      end else if (10'h187 == _T_22[9:0]) begin
        image_0_391 <= io_pixelVal_in_0_2;
      end else if (10'h187 == _T_19[9:0]) begin
        image_0_391 <= io_pixelVal_in_0_1;
      end else if (10'h187 == _T_15[9:0]) begin
        image_0_391 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_392 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h188 == _T_37[9:0]) begin
        image_0_392 <= io_pixelVal_in_0_7;
      end else if (10'h188 == _T_34[9:0]) begin
        image_0_392 <= io_pixelVal_in_0_6;
      end else if (10'h188 == _T_31[9:0]) begin
        image_0_392 <= io_pixelVal_in_0_5;
      end else if (10'h188 == _T_28[9:0]) begin
        image_0_392 <= io_pixelVal_in_0_4;
      end else if (10'h188 == _T_25[9:0]) begin
        image_0_392 <= io_pixelVal_in_0_3;
      end else if (10'h188 == _T_22[9:0]) begin
        image_0_392 <= io_pixelVal_in_0_2;
      end else if (10'h188 == _T_19[9:0]) begin
        image_0_392 <= io_pixelVal_in_0_1;
      end else if (10'h188 == _T_15[9:0]) begin
        image_0_392 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_393 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h189 == _T_37[9:0]) begin
        image_0_393 <= io_pixelVal_in_0_7;
      end else if (10'h189 == _T_34[9:0]) begin
        image_0_393 <= io_pixelVal_in_0_6;
      end else if (10'h189 == _T_31[9:0]) begin
        image_0_393 <= io_pixelVal_in_0_5;
      end else if (10'h189 == _T_28[9:0]) begin
        image_0_393 <= io_pixelVal_in_0_4;
      end else if (10'h189 == _T_25[9:0]) begin
        image_0_393 <= io_pixelVal_in_0_3;
      end else if (10'h189 == _T_22[9:0]) begin
        image_0_393 <= io_pixelVal_in_0_2;
      end else if (10'h189 == _T_19[9:0]) begin
        image_0_393 <= io_pixelVal_in_0_1;
      end else if (10'h189 == _T_15[9:0]) begin
        image_0_393 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_394 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h18a == _T_37[9:0]) begin
        image_0_394 <= io_pixelVal_in_0_7;
      end else if (10'h18a == _T_34[9:0]) begin
        image_0_394 <= io_pixelVal_in_0_6;
      end else if (10'h18a == _T_31[9:0]) begin
        image_0_394 <= io_pixelVal_in_0_5;
      end else if (10'h18a == _T_28[9:0]) begin
        image_0_394 <= io_pixelVal_in_0_4;
      end else if (10'h18a == _T_25[9:0]) begin
        image_0_394 <= io_pixelVal_in_0_3;
      end else if (10'h18a == _T_22[9:0]) begin
        image_0_394 <= io_pixelVal_in_0_2;
      end else if (10'h18a == _T_19[9:0]) begin
        image_0_394 <= io_pixelVal_in_0_1;
      end else if (10'h18a == _T_15[9:0]) begin
        image_0_394 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_395 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h18b == _T_37[9:0]) begin
        image_0_395 <= io_pixelVal_in_0_7;
      end else if (10'h18b == _T_34[9:0]) begin
        image_0_395 <= io_pixelVal_in_0_6;
      end else if (10'h18b == _T_31[9:0]) begin
        image_0_395 <= io_pixelVal_in_0_5;
      end else if (10'h18b == _T_28[9:0]) begin
        image_0_395 <= io_pixelVal_in_0_4;
      end else if (10'h18b == _T_25[9:0]) begin
        image_0_395 <= io_pixelVal_in_0_3;
      end else if (10'h18b == _T_22[9:0]) begin
        image_0_395 <= io_pixelVal_in_0_2;
      end else if (10'h18b == _T_19[9:0]) begin
        image_0_395 <= io_pixelVal_in_0_1;
      end else if (10'h18b == _T_15[9:0]) begin
        image_0_395 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_396 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h18c == _T_37[9:0]) begin
        image_0_396 <= io_pixelVal_in_0_7;
      end else if (10'h18c == _T_34[9:0]) begin
        image_0_396 <= io_pixelVal_in_0_6;
      end else if (10'h18c == _T_31[9:0]) begin
        image_0_396 <= io_pixelVal_in_0_5;
      end else if (10'h18c == _T_28[9:0]) begin
        image_0_396 <= io_pixelVal_in_0_4;
      end else if (10'h18c == _T_25[9:0]) begin
        image_0_396 <= io_pixelVal_in_0_3;
      end else if (10'h18c == _T_22[9:0]) begin
        image_0_396 <= io_pixelVal_in_0_2;
      end else if (10'h18c == _T_19[9:0]) begin
        image_0_396 <= io_pixelVal_in_0_1;
      end else if (10'h18c == _T_15[9:0]) begin
        image_0_396 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_397 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h18d == _T_37[9:0]) begin
        image_0_397 <= io_pixelVal_in_0_7;
      end else if (10'h18d == _T_34[9:0]) begin
        image_0_397 <= io_pixelVal_in_0_6;
      end else if (10'h18d == _T_31[9:0]) begin
        image_0_397 <= io_pixelVal_in_0_5;
      end else if (10'h18d == _T_28[9:0]) begin
        image_0_397 <= io_pixelVal_in_0_4;
      end else if (10'h18d == _T_25[9:0]) begin
        image_0_397 <= io_pixelVal_in_0_3;
      end else if (10'h18d == _T_22[9:0]) begin
        image_0_397 <= io_pixelVal_in_0_2;
      end else if (10'h18d == _T_19[9:0]) begin
        image_0_397 <= io_pixelVal_in_0_1;
      end else if (10'h18d == _T_15[9:0]) begin
        image_0_397 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_398 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h18e == _T_37[9:0]) begin
        image_0_398 <= io_pixelVal_in_0_7;
      end else if (10'h18e == _T_34[9:0]) begin
        image_0_398 <= io_pixelVal_in_0_6;
      end else if (10'h18e == _T_31[9:0]) begin
        image_0_398 <= io_pixelVal_in_0_5;
      end else if (10'h18e == _T_28[9:0]) begin
        image_0_398 <= io_pixelVal_in_0_4;
      end else if (10'h18e == _T_25[9:0]) begin
        image_0_398 <= io_pixelVal_in_0_3;
      end else if (10'h18e == _T_22[9:0]) begin
        image_0_398 <= io_pixelVal_in_0_2;
      end else if (10'h18e == _T_19[9:0]) begin
        image_0_398 <= io_pixelVal_in_0_1;
      end else if (10'h18e == _T_15[9:0]) begin
        image_0_398 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_399 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h18f == _T_37[9:0]) begin
        image_0_399 <= io_pixelVal_in_0_7;
      end else if (10'h18f == _T_34[9:0]) begin
        image_0_399 <= io_pixelVal_in_0_6;
      end else if (10'h18f == _T_31[9:0]) begin
        image_0_399 <= io_pixelVal_in_0_5;
      end else if (10'h18f == _T_28[9:0]) begin
        image_0_399 <= io_pixelVal_in_0_4;
      end else if (10'h18f == _T_25[9:0]) begin
        image_0_399 <= io_pixelVal_in_0_3;
      end else if (10'h18f == _T_22[9:0]) begin
        image_0_399 <= io_pixelVal_in_0_2;
      end else if (10'h18f == _T_19[9:0]) begin
        image_0_399 <= io_pixelVal_in_0_1;
      end else if (10'h18f == _T_15[9:0]) begin
        image_0_399 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_400 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h190 == _T_37[9:0]) begin
        image_0_400 <= io_pixelVal_in_0_7;
      end else if (10'h190 == _T_34[9:0]) begin
        image_0_400 <= io_pixelVal_in_0_6;
      end else if (10'h190 == _T_31[9:0]) begin
        image_0_400 <= io_pixelVal_in_0_5;
      end else if (10'h190 == _T_28[9:0]) begin
        image_0_400 <= io_pixelVal_in_0_4;
      end else if (10'h190 == _T_25[9:0]) begin
        image_0_400 <= io_pixelVal_in_0_3;
      end else if (10'h190 == _T_22[9:0]) begin
        image_0_400 <= io_pixelVal_in_0_2;
      end else if (10'h190 == _T_19[9:0]) begin
        image_0_400 <= io_pixelVal_in_0_1;
      end else if (10'h190 == _T_15[9:0]) begin
        image_0_400 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_401 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h191 == _T_37[9:0]) begin
        image_0_401 <= io_pixelVal_in_0_7;
      end else if (10'h191 == _T_34[9:0]) begin
        image_0_401 <= io_pixelVal_in_0_6;
      end else if (10'h191 == _T_31[9:0]) begin
        image_0_401 <= io_pixelVal_in_0_5;
      end else if (10'h191 == _T_28[9:0]) begin
        image_0_401 <= io_pixelVal_in_0_4;
      end else if (10'h191 == _T_25[9:0]) begin
        image_0_401 <= io_pixelVal_in_0_3;
      end else if (10'h191 == _T_22[9:0]) begin
        image_0_401 <= io_pixelVal_in_0_2;
      end else if (10'h191 == _T_19[9:0]) begin
        image_0_401 <= io_pixelVal_in_0_1;
      end else if (10'h191 == _T_15[9:0]) begin
        image_0_401 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_402 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h192 == _T_37[9:0]) begin
        image_0_402 <= io_pixelVal_in_0_7;
      end else if (10'h192 == _T_34[9:0]) begin
        image_0_402 <= io_pixelVal_in_0_6;
      end else if (10'h192 == _T_31[9:0]) begin
        image_0_402 <= io_pixelVal_in_0_5;
      end else if (10'h192 == _T_28[9:0]) begin
        image_0_402 <= io_pixelVal_in_0_4;
      end else if (10'h192 == _T_25[9:0]) begin
        image_0_402 <= io_pixelVal_in_0_3;
      end else if (10'h192 == _T_22[9:0]) begin
        image_0_402 <= io_pixelVal_in_0_2;
      end else if (10'h192 == _T_19[9:0]) begin
        image_0_402 <= io_pixelVal_in_0_1;
      end else if (10'h192 == _T_15[9:0]) begin
        image_0_402 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_403 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h193 == _T_37[9:0]) begin
        image_0_403 <= io_pixelVal_in_0_7;
      end else if (10'h193 == _T_34[9:0]) begin
        image_0_403 <= io_pixelVal_in_0_6;
      end else if (10'h193 == _T_31[9:0]) begin
        image_0_403 <= io_pixelVal_in_0_5;
      end else if (10'h193 == _T_28[9:0]) begin
        image_0_403 <= io_pixelVal_in_0_4;
      end else if (10'h193 == _T_25[9:0]) begin
        image_0_403 <= io_pixelVal_in_0_3;
      end else if (10'h193 == _T_22[9:0]) begin
        image_0_403 <= io_pixelVal_in_0_2;
      end else if (10'h193 == _T_19[9:0]) begin
        image_0_403 <= io_pixelVal_in_0_1;
      end else if (10'h193 == _T_15[9:0]) begin
        image_0_403 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_404 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h194 == _T_37[9:0]) begin
        image_0_404 <= io_pixelVal_in_0_7;
      end else if (10'h194 == _T_34[9:0]) begin
        image_0_404 <= io_pixelVal_in_0_6;
      end else if (10'h194 == _T_31[9:0]) begin
        image_0_404 <= io_pixelVal_in_0_5;
      end else if (10'h194 == _T_28[9:0]) begin
        image_0_404 <= io_pixelVal_in_0_4;
      end else if (10'h194 == _T_25[9:0]) begin
        image_0_404 <= io_pixelVal_in_0_3;
      end else if (10'h194 == _T_22[9:0]) begin
        image_0_404 <= io_pixelVal_in_0_2;
      end else if (10'h194 == _T_19[9:0]) begin
        image_0_404 <= io_pixelVal_in_0_1;
      end else if (10'h194 == _T_15[9:0]) begin
        image_0_404 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_405 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h195 == _T_37[9:0]) begin
        image_0_405 <= io_pixelVal_in_0_7;
      end else if (10'h195 == _T_34[9:0]) begin
        image_0_405 <= io_pixelVal_in_0_6;
      end else if (10'h195 == _T_31[9:0]) begin
        image_0_405 <= io_pixelVal_in_0_5;
      end else if (10'h195 == _T_28[9:0]) begin
        image_0_405 <= io_pixelVal_in_0_4;
      end else if (10'h195 == _T_25[9:0]) begin
        image_0_405 <= io_pixelVal_in_0_3;
      end else if (10'h195 == _T_22[9:0]) begin
        image_0_405 <= io_pixelVal_in_0_2;
      end else if (10'h195 == _T_19[9:0]) begin
        image_0_405 <= io_pixelVal_in_0_1;
      end else if (10'h195 == _T_15[9:0]) begin
        image_0_405 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_406 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h196 == _T_37[9:0]) begin
        image_0_406 <= io_pixelVal_in_0_7;
      end else if (10'h196 == _T_34[9:0]) begin
        image_0_406 <= io_pixelVal_in_0_6;
      end else if (10'h196 == _T_31[9:0]) begin
        image_0_406 <= io_pixelVal_in_0_5;
      end else if (10'h196 == _T_28[9:0]) begin
        image_0_406 <= io_pixelVal_in_0_4;
      end else if (10'h196 == _T_25[9:0]) begin
        image_0_406 <= io_pixelVal_in_0_3;
      end else if (10'h196 == _T_22[9:0]) begin
        image_0_406 <= io_pixelVal_in_0_2;
      end else if (10'h196 == _T_19[9:0]) begin
        image_0_406 <= io_pixelVal_in_0_1;
      end else if (10'h196 == _T_15[9:0]) begin
        image_0_406 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_407 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h197 == _T_37[9:0]) begin
        image_0_407 <= io_pixelVal_in_0_7;
      end else if (10'h197 == _T_34[9:0]) begin
        image_0_407 <= io_pixelVal_in_0_6;
      end else if (10'h197 == _T_31[9:0]) begin
        image_0_407 <= io_pixelVal_in_0_5;
      end else if (10'h197 == _T_28[9:0]) begin
        image_0_407 <= io_pixelVal_in_0_4;
      end else if (10'h197 == _T_25[9:0]) begin
        image_0_407 <= io_pixelVal_in_0_3;
      end else if (10'h197 == _T_22[9:0]) begin
        image_0_407 <= io_pixelVal_in_0_2;
      end else if (10'h197 == _T_19[9:0]) begin
        image_0_407 <= io_pixelVal_in_0_1;
      end else if (10'h197 == _T_15[9:0]) begin
        image_0_407 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_408 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h198 == _T_37[9:0]) begin
        image_0_408 <= io_pixelVal_in_0_7;
      end else if (10'h198 == _T_34[9:0]) begin
        image_0_408 <= io_pixelVal_in_0_6;
      end else if (10'h198 == _T_31[9:0]) begin
        image_0_408 <= io_pixelVal_in_0_5;
      end else if (10'h198 == _T_28[9:0]) begin
        image_0_408 <= io_pixelVal_in_0_4;
      end else if (10'h198 == _T_25[9:0]) begin
        image_0_408 <= io_pixelVal_in_0_3;
      end else if (10'h198 == _T_22[9:0]) begin
        image_0_408 <= io_pixelVal_in_0_2;
      end else if (10'h198 == _T_19[9:0]) begin
        image_0_408 <= io_pixelVal_in_0_1;
      end else if (10'h198 == _T_15[9:0]) begin
        image_0_408 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_409 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h199 == _T_37[9:0]) begin
        image_0_409 <= io_pixelVal_in_0_7;
      end else if (10'h199 == _T_34[9:0]) begin
        image_0_409 <= io_pixelVal_in_0_6;
      end else if (10'h199 == _T_31[9:0]) begin
        image_0_409 <= io_pixelVal_in_0_5;
      end else if (10'h199 == _T_28[9:0]) begin
        image_0_409 <= io_pixelVal_in_0_4;
      end else if (10'h199 == _T_25[9:0]) begin
        image_0_409 <= io_pixelVal_in_0_3;
      end else if (10'h199 == _T_22[9:0]) begin
        image_0_409 <= io_pixelVal_in_0_2;
      end else if (10'h199 == _T_19[9:0]) begin
        image_0_409 <= io_pixelVal_in_0_1;
      end else if (10'h199 == _T_15[9:0]) begin
        image_0_409 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_410 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h19a == _T_37[9:0]) begin
        image_0_410 <= io_pixelVal_in_0_7;
      end else if (10'h19a == _T_34[9:0]) begin
        image_0_410 <= io_pixelVal_in_0_6;
      end else if (10'h19a == _T_31[9:0]) begin
        image_0_410 <= io_pixelVal_in_0_5;
      end else if (10'h19a == _T_28[9:0]) begin
        image_0_410 <= io_pixelVal_in_0_4;
      end else if (10'h19a == _T_25[9:0]) begin
        image_0_410 <= io_pixelVal_in_0_3;
      end else if (10'h19a == _T_22[9:0]) begin
        image_0_410 <= io_pixelVal_in_0_2;
      end else if (10'h19a == _T_19[9:0]) begin
        image_0_410 <= io_pixelVal_in_0_1;
      end else if (10'h19a == _T_15[9:0]) begin
        image_0_410 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_411 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h19b == _T_37[9:0]) begin
        image_0_411 <= io_pixelVal_in_0_7;
      end else if (10'h19b == _T_34[9:0]) begin
        image_0_411 <= io_pixelVal_in_0_6;
      end else if (10'h19b == _T_31[9:0]) begin
        image_0_411 <= io_pixelVal_in_0_5;
      end else if (10'h19b == _T_28[9:0]) begin
        image_0_411 <= io_pixelVal_in_0_4;
      end else if (10'h19b == _T_25[9:0]) begin
        image_0_411 <= io_pixelVal_in_0_3;
      end else if (10'h19b == _T_22[9:0]) begin
        image_0_411 <= io_pixelVal_in_0_2;
      end else if (10'h19b == _T_19[9:0]) begin
        image_0_411 <= io_pixelVal_in_0_1;
      end else if (10'h19b == _T_15[9:0]) begin
        image_0_411 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_412 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h19c == _T_37[9:0]) begin
        image_0_412 <= io_pixelVal_in_0_7;
      end else if (10'h19c == _T_34[9:0]) begin
        image_0_412 <= io_pixelVal_in_0_6;
      end else if (10'h19c == _T_31[9:0]) begin
        image_0_412 <= io_pixelVal_in_0_5;
      end else if (10'h19c == _T_28[9:0]) begin
        image_0_412 <= io_pixelVal_in_0_4;
      end else if (10'h19c == _T_25[9:0]) begin
        image_0_412 <= io_pixelVal_in_0_3;
      end else if (10'h19c == _T_22[9:0]) begin
        image_0_412 <= io_pixelVal_in_0_2;
      end else if (10'h19c == _T_19[9:0]) begin
        image_0_412 <= io_pixelVal_in_0_1;
      end else if (10'h19c == _T_15[9:0]) begin
        image_0_412 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_413 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h19d == _T_37[9:0]) begin
        image_0_413 <= io_pixelVal_in_0_7;
      end else if (10'h19d == _T_34[9:0]) begin
        image_0_413 <= io_pixelVal_in_0_6;
      end else if (10'h19d == _T_31[9:0]) begin
        image_0_413 <= io_pixelVal_in_0_5;
      end else if (10'h19d == _T_28[9:0]) begin
        image_0_413 <= io_pixelVal_in_0_4;
      end else if (10'h19d == _T_25[9:0]) begin
        image_0_413 <= io_pixelVal_in_0_3;
      end else if (10'h19d == _T_22[9:0]) begin
        image_0_413 <= io_pixelVal_in_0_2;
      end else if (10'h19d == _T_19[9:0]) begin
        image_0_413 <= io_pixelVal_in_0_1;
      end else if (10'h19d == _T_15[9:0]) begin
        image_0_413 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_414 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h19e == _T_37[9:0]) begin
        image_0_414 <= io_pixelVal_in_0_7;
      end else if (10'h19e == _T_34[9:0]) begin
        image_0_414 <= io_pixelVal_in_0_6;
      end else if (10'h19e == _T_31[9:0]) begin
        image_0_414 <= io_pixelVal_in_0_5;
      end else if (10'h19e == _T_28[9:0]) begin
        image_0_414 <= io_pixelVal_in_0_4;
      end else if (10'h19e == _T_25[9:0]) begin
        image_0_414 <= io_pixelVal_in_0_3;
      end else if (10'h19e == _T_22[9:0]) begin
        image_0_414 <= io_pixelVal_in_0_2;
      end else if (10'h19e == _T_19[9:0]) begin
        image_0_414 <= io_pixelVal_in_0_1;
      end else if (10'h19e == _T_15[9:0]) begin
        image_0_414 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_415 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h19f == _T_37[9:0]) begin
        image_0_415 <= io_pixelVal_in_0_7;
      end else if (10'h19f == _T_34[9:0]) begin
        image_0_415 <= io_pixelVal_in_0_6;
      end else if (10'h19f == _T_31[9:0]) begin
        image_0_415 <= io_pixelVal_in_0_5;
      end else if (10'h19f == _T_28[9:0]) begin
        image_0_415 <= io_pixelVal_in_0_4;
      end else if (10'h19f == _T_25[9:0]) begin
        image_0_415 <= io_pixelVal_in_0_3;
      end else if (10'h19f == _T_22[9:0]) begin
        image_0_415 <= io_pixelVal_in_0_2;
      end else if (10'h19f == _T_19[9:0]) begin
        image_0_415 <= io_pixelVal_in_0_1;
      end else if (10'h19f == _T_15[9:0]) begin
        image_0_415 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_416 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1a0 == _T_37[9:0]) begin
        image_0_416 <= io_pixelVal_in_0_7;
      end else if (10'h1a0 == _T_34[9:0]) begin
        image_0_416 <= io_pixelVal_in_0_6;
      end else if (10'h1a0 == _T_31[9:0]) begin
        image_0_416 <= io_pixelVal_in_0_5;
      end else if (10'h1a0 == _T_28[9:0]) begin
        image_0_416 <= io_pixelVal_in_0_4;
      end else if (10'h1a0 == _T_25[9:0]) begin
        image_0_416 <= io_pixelVal_in_0_3;
      end else if (10'h1a0 == _T_22[9:0]) begin
        image_0_416 <= io_pixelVal_in_0_2;
      end else if (10'h1a0 == _T_19[9:0]) begin
        image_0_416 <= io_pixelVal_in_0_1;
      end else if (10'h1a0 == _T_15[9:0]) begin
        image_0_416 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_417 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1a1 == _T_37[9:0]) begin
        image_0_417 <= io_pixelVal_in_0_7;
      end else if (10'h1a1 == _T_34[9:0]) begin
        image_0_417 <= io_pixelVal_in_0_6;
      end else if (10'h1a1 == _T_31[9:0]) begin
        image_0_417 <= io_pixelVal_in_0_5;
      end else if (10'h1a1 == _T_28[9:0]) begin
        image_0_417 <= io_pixelVal_in_0_4;
      end else if (10'h1a1 == _T_25[9:0]) begin
        image_0_417 <= io_pixelVal_in_0_3;
      end else if (10'h1a1 == _T_22[9:0]) begin
        image_0_417 <= io_pixelVal_in_0_2;
      end else if (10'h1a1 == _T_19[9:0]) begin
        image_0_417 <= io_pixelVal_in_0_1;
      end else if (10'h1a1 == _T_15[9:0]) begin
        image_0_417 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_418 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1a2 == _T_37[9:0]) begin
        image_0_418 <= io_pixelVal_in_0_7;
      end else if (10'h1a2 == _T_34[9:0]) begin
        image_0_418 <= io_pixelVal_in_0_6;
      end else if (10'h1a2 == _T_31[9:0]) begin
        image_0_418 <= io_pixelVal_in_0_5;
      end else if (10'h1a2 == _T_28[9:0]) begin
        image_0_418 <= io_pixelVal_in_0_4;
      end else if (10'h1a2 == _T_25[9:0]) begin
        image_0_418 <= io_pixelVal_in_0_3;
      end else if (10'h1a2 == _T_22[9:0]) begin
        image_0_418 <= io_pixelVal_in_0_2;
      end else if (10'h1a2 == _T_19[9:0]) begin
        image_0_418 <= io_pixelVal_in_0_1;
      end else if (10'h1a2 == _T_15[9:0]) begin
        image_0_418 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_419 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1a3 == _T_37[9:0]) begin
        image_0_419 <= io_pixelVal_in_0_7;
      end else if (10'h1a3 == _T_34[9:0]) begin
        image_0_419 <= io_pixelVal_in_0_6;
      end else if (10'h1a3 == _T_31[9:0]) begin
        image_0_419 <= io_pixelVal_in_0_5;
      end else if (10'h1a3 == _T_28[9:0]) begin
        image_0_419 <= io_pixelVal_in_0_4;
      end else if (10'h1a3 == _T_25[9:0]) begin
        image_0_419 <= io_pixelVal_in_0_3;
      end else if (10'h1a3 == _T_22[9:0]) begin
        image_0_419 <= io_pixelVal_in_0_2;
      end else if (10'h1a3 == _T_19[9:0]) begin
        image_0_419 <= io_pixelVal_in_0_1;
      end else if (10'h1a3 == _T_15[9:0]) begin
        image_0_419 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_420 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1a4 == _T_37[9:0]) begin
        image_0_420 <= io_pixelVal_in_0_7;
      end else if (10'h1a4 == _T_34[9:0]) begin
        image_0_420 <= io_pixelVal_in_0_6;
      end else if (10'h1a4 == _T_31[9:0]) begin
        image_0_420 <= io_pixelVal_in_0_5;
      end else if (10'h1a4 == _T_28[9:0]) begin
        image_0_420 <= io_pixelVal_in_0_4;
      end else if (10'h1a4 == _T_25[9:0]) begin
        image_0_420 <= io_pixelVal_in_0_3;
      end else if (10'h1a4 == _T_22[9:0]) begin
        image_0_420 <= io_pixelVal_in_0_2;
      end else if (10'h1a4 == _T_19[9:0]) begin
        image_0_420 <= io_pixelVal_in_0_1;
      end else if (10'h1a4 == _T_15[9:0]) begin
        image_0_420 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_421 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1a5 == _T_37[9:0]) begin
        image_0_421 <= io_pixelVal_in_0_7;
      end else if (10'h1a5 == _T_34[9:0]) begin
        image_0_421 <= io_pixelVal_in_0_6;
      end else if (10'h1a5 == _T_31[9:0]) begin
        image_0_421 <= io_pixelVal_in_0_5;
      end else if (10'h1a5 == _T_28[9:0]) begin
        image_0_421 <= io_pixelVal_in_0_4;
      end else if (10'h1a5 == _T_25[9:0]) begin
        image_0_421 <= io_pixelVal_in_0_3;
      end else if (10'h1a5 == _T_22[9:0]) begin
        image_0_421 <= io_pixelVal_in_0_2;
      end else if (10'h1a5 == _T_19[9:0]) begin
        image_0_421 <= io_pixelVal_in_0_1;
      end else if (10'h1a5 == _T_15[9:0]) begin
        image_0_421 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_422 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1a6 == _T_37[9:0]) begin
        image_0_422 <= io_pixelVal_in_0_7;
      end else if (10'h1a6 == _T_34[9:0]) begin
        image_0_422 <= io_pixelVal_in_0_6;
      end else if (10'h1a6 == _T_31[9:0]) begin
        image_0_422 <= io_pixelVal_in_0_5;
      end else if (10'h1a6 == _T_28[9:0]) begin
        image_0_422 <= io_pixelVal_in_0_4;
      end else if (10'h1a6 == _T_25[9:0]) begin
        image_0_422 <= io_pixelVal_in_0_3;
      end else if (10'h1a6 == _T_22[9:0]) begin
        image_0_422 <= io_pixelVal_in_0_2;
      end else if (10'h1a6 == _T_19[9:0]) begin
        image_0_422 <= io_pixelVal_in_0_1;
      end else if (10'h1a6 == _T_15[9:0]) begin
        image_0_422 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_423 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1a7 == _T_37[9:0]) begin
        image_0_423 <= io_pixelVal_in_0_7;
      end else if (10'h1a7 == _T_34[9:0]) begin
        image_0_423 <= io_pixelVal_in_0_6;
      end else if (10'h1a7 == _T_31[9:0]) begin
        image_0_423 <= io_pixelVal_in_0_5;
      end else if (10'h1a7 == _T_28[9:0]) begin
        image_0_423 <= io_pixelVal_in_0_4;
      end else if (10'h1a7 == _T_25[9:0]) begin
        image_0_423 <= io_pixelVal_in_0_3;
      end else if (10'h1a7 == _T_22[9:0]) begin
        image_0_423 <= io_pixelVal_in_0_2;
      end else if (10'h1a7 == _T_19[9:0]) begin
        image_0_423 <= io_pixelVal_in_0_1;
      end else if (10'h1a7 == _T_15[9:0]) begin
        image_0_423 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_424 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1a8 == _T_37[9:0]) begin
        image_0_424 <= io_pixelVal_in_0_7;
      end else if (10'h1a8 == _T_34[9:0]) begin
        image_0_424 <= io_pixelVal_in_0_6;
      end else if (10'h1a8 == _T_31[9:0]) begin
        image_0_424 <= io_pixelVal_in_0_5;
      end else if (10'h1a8 == _T_28[9:0]) begin
        image_0_424 <= io_pixelVal_in_0_4;
      end else if (10'h1a8 == _T_25[9:0]) begin
        image_0_424 <= io_pixelVal_in_0_3;
      end else if (10'h1a8 == _T_22[9:0]) begin
        image_0_424 <= io_pixelVal_in_0_2;
      end else if (10'h1a8 == _T_19[9:0]) begin
        image_0_424 <= io_pixelVal_in_0_1;
      end else if (10'h1a8 == _T_15[9:0]) begin
        image_0_424 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_425 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1a9 == _T_37[9:0]) begin
        image_0_425 <= io_pixelVal_in_0_7;
      end else if (10'h1a9 == _T_34[9:0]) begin
        image_0_425 <= io_pixelVal_in_0_6;
      end else if (10'h1a9 == _T_31[9:0]) begin
        image_0_425 <= io_pixelVal_in_0_5;
      end else if (10'h1a9 == _T_28[9:0]) begin
        image_0_425 <= io_pixelVal_in_0_4;
      end else if (10'h1a9 == _T_25[9:0]) begin
        image_0_425 <= io_pixelVal_in_0_3;
      end else if (10'h1a9 == _T_22[9:0]) begin
        image_0_425 <= io_pixelVal_in_0_2;
      end else if (10'h1a9 == _T_19[9:0]) begin
        image_0_425 <= io_pixelVal_in_0_1;
      end else if (10'h1a9 == _T_15[9:0]) begin
        image_0_425 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_426 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1aa == _T_37[9:0]) begin
        image_0_426 <= io_pixelVal_in_0_7;
      end else if (10'h1aa == _T_34[9:0]) begin
        image_0_426 <= io_pixelVal_in_0_6;
      end else if (10'h1aa == _T_31[9:0]) begin
        image_0_426 <= io_pixelVal_in_0_5;
      end else if (10'h1aa == _T_28[9:0]) begin
        image_0_426 <= io_pixelVal_in_0_4;
      end else if (10'h1aa == _T_25[9:0]) begin
        image_0_426 <= io_pixelVal_in_0_3;
      end else if (10'h1aa == _T_22[9:0]) begin
        image_0_426 <= io_pixelVal_in_0_2;
      end else if (10'h1aa == _T_19[9:0]) begin
        image_0_426 <= io_pixelVal_in_0_1;
      end else if (10'h1aa == _T_15[9:0]) begin
        image_0_426 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_427 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1ab == _T_37[9:0]) begin
        image_0_427 <= io_pixelVal_in_0_7;
      end else if (10'h1ab == _T_34[9:0]) begin
        image_0_427 <= io_pixelVal_in_0_6;
      end else if (10'h1ab == _T_31[9:0]) begin
        image_0_427 <= io_pixelVal_in_0_5;
      end else if (10'h1ab == _T_28[9:0]) begin
        image_0_427 <= io_pixelVal_in_0_4;
      end else if (10'h1ab == _T_25[9:0]) begin
        image_0_427 <= io_pixelVal_in_0_3;
      end else if (10'h1ab == _T_22[9:0]) begin
        image_0_427 <= io_pixelVal_in_0_2;
      end else if (10'h1ab == _T_19[9:0]) begin
        image_0_427 <= io_pixelVal_in_0_1;
      end else if (10'h1ab == _T_15[9:0]) begin
        image_0_427 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_428 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1ac == _T_37[9:0]) begin
        image_0_428 <= io_pixelVal_in_0_7;
      end else if (10'h1ac == _T_34[9:0]) begin
        image_0_428 <= io_pixelVal_in_0_6;
      end else if (10'h1ac == _T_31[9:0]) begin
        image_0_428 <= io_pixelVal_in_0_5;
      end else if (10'h1ac == _T_28[9:0]) begin
        image_0_428 <= io_pixelVal_in_0_4;
      end else if (10'h1ac == _T_25[9:0]) begin
        image_0_428 <= io_pixelVal_in_0_3;
      end else if (10'h1ac == _T_22[9:0]) begin
        image_0_428 <= io_pixelVal_in_0_2;
      end else if (10'h1ac == _T_19[9:0]) begin
        image_0_428 <= io_pixelVal_in_0_1;
      end else if (10'h1ac == _T_15[9:0]) begin
        image_0_428 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_429 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1ad == _T_37[9:0]) begin
        image_0_429 <= io_pixelVal_in_0_7;
      end else if (10'h1ad == _T_34[9:0]) begin
        image_0_429 <= io_pixelVal_in_0_6;
      end else if (10'h1ad == _T_31[9:0]) begin
        image_0_429 <= io_pixelVal_in_0_5;
      end else if (10'h1ad == _T_28[9:0]) begin
        image_0_429 <= io_pixelVal_in_0_4;
      end else if (10'h1ad == _T_25[9:0]) begin
        image_0_429 <= io_pixelVal_in_0_3;
      end else if (10'h1ad == _T_22[9:0]) begin
        image_0_429 <= io_pixelVal_in_0_2;
      end else if (10'h1ad == _T_19[9:0]) begin
        image_0_429 <= io_pixelVal_in_0_1;
      end else if (10'h1ad == _T_15[9:0]) begin
        image_0_429 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_430 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1ae == _T_37[9:0]) begin
        image_0_430 <= io_pixelVal_in_0_7;
      end else if (10'h1ae == _T_34[9:0]) begin
        image_0_430 <= io_pixelVal_in_0_6;
      end else if (10'h1ae == _T_31[9:0]) begin
        image_0_430 <= io_pixelVal_in_0_5;
      end else if (10'h1ae == _T_28[9:0]) begin
        image_0_430 <= io_pixelVal_in_0_4;
      end else if (10'h1ae == _T_25[9:0]) begin
        image_0_430 <= io_pixelVal_in_0_3;
      end else if (10'h1ae == _T_22[9:0]) begin
        image_0_430 <= io_pixelVal_in_0_2;
      end else if (10'h1ae == _T_19[9:0]) begin
        image_0_430 <= io_pixelVal_in_0_1;
      end else if (10'h1ae == _T_15[9:0]) begin
        image_0_430 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_431 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1af == _T_37[9:0]) begin
        image_0_431 <= io_pixelVal_in_0_7;
      end else if (10'h1af == _T_34[9:0]) begin
        image_0_431 <= io_pixelVal_in_0_6;
      end else if (10'h1af == _T_31[9:0]) begin
        image_0_431 <= io_pixelVal_in_0_5;
      end else if (10'h1af == _T_28[9:0]) begin
        image_0_431 <= io_pixelVal_in_0_4;
      end else if (10'h1af == _T_25[9:0]) begin
        image_0_431 <= io_pixelVal_in_0_3;
      end else if (10'h1af == _T_22[9:0]) begin
        image_0_431 <= io_pixelVal_in_0_2;
      end else if (10'h1af == _T_19[9:0]) begin
        image_0_431 <= io_pixelVal_in_0_1;
      end else if (10'h1af == _T_15[9:0]) begin
        image_0_431 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_432 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1b0 == _T_37[9:0]) begin
        image_0_432 <= io_pixelVal_in_0_7;
      end else if (10'h1b0 == _T_34[9:0]) begin
        image_0_432 <= io_pixelVal_in_0_6;
      end else if (10'h1b0 == _T_31[9:0]) begin
        image_0_432 <= io_pixelVal_in_0_5;
      end else if (10'h1b0 == _T_28[9:0]) begin
        image_0_432 <= io_pixelVal_in_0_4;
      end else if (10'h1b0 == _T_25[9:0]) begin
        image_0_432 <= io_pixelVal_in_0_3;
      end else if (10'h1b0 == _T_22[9:0]) begin
        image_0_432 <= io_pixelVal_in_0_2;
      end else if (10'h1b0 == _T_19[9:0]) begin
        image_0_432 <= io_pixelVal_in_0_1;
      end else if (10'h1b0 == _T_15[9:0]) begin
        image_0_432 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_433 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1b1 == _T_37[9:0]) begin
        image_0_433 <= io_pixelVal_in_0_7;
      end else if (10'h1b1 == _T_34[9:0]) begin
        image_0_433 <= io_pixelVal_in_0_6;
      end else if (10'h1b1 == _T_31[9:0]) begin
        image_0_433 <= io_pixelVal_in_0_5;
      end else if (10'h1b1 == _T_28[9:0]) begin
        image_0_433 <= io_pixelVal_in_0_4;
      end else if (10'h1b1 == _T_25[9:0]) begin
        image_0_433 <= io_pixelVal_in_0_3;
      end else if (10'h1b1 == _T_22[9:0]) begin
        image_0_433 <= io_pixelVal_in_0_2;
      end else if (10'h1b1 == _T_19[9:0]) begin
        image_0_433 <= io_pixelVal_in_0_1;
      end else if (10'h1b1 == _T_15[9:0]) begin
        image_0_433 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_434 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1b2 == _T_37[9:0]) begin
        image_0_434 <= io_pixelVal_in_0_7;
      end else if (10'h1b2 == _T_34[9:0]) begin
        image_0_434 <= io_pixelVal_in_0_6;
      end else if (10'h1b2 == _T_31[9:0]) begin
        image_0_434 <= io_pixelVal_in_0_5;
      end else if (10'h1b2 == _T_28[9:0]) begin
        image_0_434 <= io_pixelVal_in_0_4;
      end else if (10'h1b2 == _T_25[9:0]) begin
        image_0_434 <= io_pixelVal_in_0_3;
      end else if (10'h1b2 == _T_22[9:0]) begin
        image_0_434 <= io_pixelVal_in_0_2;
      end else if (10'h1b2 == _T_19[9:0]) begin
        image_0_434 <= io_pixelVal_in_0_1;
      end else if (10'h1b2 == _T_15[9:0]) begin
        image_0_434 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_435 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1b3 == _T_37[9:0]) begin
        image_0_435 <= io_pixelVal_in_0_7;
      end else if (10'h1b3 == _T_34[9:0]) begin
        image_0_435 <= io_pixelVal_in_0_6;
      end else if (10'h1b3 == _T_31[9:0]) begin
        image_0_435 <= io_pixelVal_in_0_5;
      end else if (10'h1b3 == _T_28[9:0]) begin
        image_0_435 <= io_pixelVal_in_0_4;
      end else if (10'h1b3 == _T_25[9:0]) begin
        image_0_435 <= io_pixelVal_in_0_3;
      end else if (10'h1b3 == _T_22[9:0]) begin
        image_0_435 <= io_pixelVal_in_0_2;
      end else if (10'h1b3 == _T_19[9:0]) begin
        image_0_435 <= io_pixelVal_in_0_1;
      end else if (10'h1b3 == _T_15[9:0]) begin
        image_0_435 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_436 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1b4 == _T_37[9:0]) begin
        image_0_436 <= io_pixelVal_in_0_7;
      end else if (10'h1b4 == _T_34[9:0]) begin
        image_0_436 <= io_pixelVal_in_0_6;
      end else if (10'h1b4 == _T_31[9:0]) begin
        image_0_436 <= io_pixelVal_in_0_5;
      end else if (10'h1b4 == _T_28[9:0]) begin
        image_0_436 <= io_pixelVal_in_0_4;
      end else if (10'h1b4 == _T_25[9:0]) begin
        image_0_436 <= io_pixelVal_in_0_3;
      end else if (10'h1b4 == _T_22[9:0]) begin
        image_0_436 <= io_pixelVal_in_0_2;
      end else if (10'h1b4 == _T_19[9:0]) begin
        image_0_436 <= io_pixelVal_in_0_1;
      end else if (10'h1b4 == _T_15[9:0]) begin
        image_0_436 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_437 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1b5 == _T_37[9:0]) begin
        image_0_437 <= io_pixelVal_in_0_7;
      end else if (10'h1b5 == _T_34[9:0]) begin
        image_0_437 <= io_pixelVal_in_0_6;
      end else if (10'h1b5 == _T_31[9:0]) begin
        image_0_437 <= io_pixelVal_in_0_5;
      end else if (10'h1b5 == _T_28[9:0]) begin
        image_0_437 <= io_pixelVal_in_0_4;
      end else if (10'h1b5 == _T_25[9:0]) begin
        image_0_437 <= io_pixelVal_in_0_3;
      end else if (10'h1b5 == _T_22[9:0]) begin
        image_0_437 <= io_pixelVal_in_0_2;
      end else if (10'h1b5 == _T_19[9:0]) begin
        image_0_437 <= io_pixelVal_in_0_1;
      end else if (10'h1b5 == _T_15[9:0]) begin
        image_0_437 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_438 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1b6 == _T_37[9:0]) begin
        image_0_438 <= io_pixelVal_in_0_7;
      end else if (10'h1b6 == _T_34[9:0]) begin
        image_0_438 <= io_pixelVal_in_0_6;
      end else if (10'h1b6 == _T_31[9:0]) begin
        image_0_438 <= io_pixelVal_in_0_5;
      end else if (10'h1b6 == _T_28[9:0]) begin
        image_0_438 <= io_pixelVal_in_0_4;
      end else if (10'h1b6 == _T_25[9:0]) begin
        image_0_438 <= io_pixelVal_in_0_3;
      end else if (10'h1b6 == _T_22[9:0]) begin
        image_0_438 <= io_pixelVal_in_0_2;
      end else if (10'h1b6 == _T_19[9:0]) begin
        image_0_438 <= io_pixelVal_in_0_1;
      end else if (10'h1b6 == _T_15[9:0]) begin
        image_0_438 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_439 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1b7 == _T_37[9:0]) begin
        image_0_439 <= io_pixelVal_in_0_7;
      end else if (10'h1b7 == _T_34[9:0]) begin
        image_0_439 <= io_pixelVal_in_0_6;
      end else if (10'h1b7 == _T_31[9:0]) begin
        image_0_439 <= io_pixelVal_in_0_5;
      end else if (10'h1b7 == _T_28[9:0]) begin
        image_0_439 <= io_pixelVal_in_0_4;
      end else if (10'h1b7 == _T_25[9:0]) begin
        image_0_439 <= io_pixelVal_in_0_3;
      end else if (10'h1b7 == _T_22[9:0]) begin
        image_0_439 <= io_pixelVal_in_0_2;
      end else if (10'h1b7 == _T_19[9:0]) begin
        image_0_439 <= io_pixelVal_in_0_1;
      end else if (10'h1b7 == _T_15[9:0]) begin
        image_0_439 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_440 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1b8 == _T_37[9:0]) begin
        image_0_440 <= io_pixelVal_in_0_7;
      end else if (10'h1b8 == _T_34[9:0]) begin
        image_0_440 <= io_pixelVal_in_0_6;
      end else if (10'h1b8 == _T_31[9:0]) begin
        image_0_440 <= io_pixelVal_in_0_5;
      end else if (10'h1b8 == _T_28[9:0]) begin
        image_0_440 <= io_pixelVal_in_0_4;
      end else if (10'h1b8 == _T_25[9:0]) begin
        image_0_440 <= io_pixelVal_in_0_3;
      end else if (10'h1b8 == _T_22[9:0]) begin
        image_0_440 <= io_pixelVal_in_0_2;
      end else if (10'h1b8 == _T_19[9:0]) begin
        image_0_440 <= io_pixelVal_in_0_1;
      end else if (10'h1b8 == _T_15[9:0]) begin
        image_0_440 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_441 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1b9 == _T_37[9:0]) begin
        image_0_441 <= io_pixelVal_in_0_7;
      end else if (10'h1b9 == _T_34[9:0]) begin
        image_0_441 <= io_pixelVal_in_0_6;
      end else if (10'h1b9 == _T_31[9:0]) begin
        image_0_441 <= io_pixelVal_in_0_5;
      end else if (10'h1b9 == _T_28[9:0]) begin
        image_0_441 <= io_pixelVal_in_0_4;
      end else if (10'h1b9 == _T_25[9:0]) begin
        image_0_441 <= io_pixelVal_in_0_3;
      end else if (10'h1b9 == _T_22[9:0]) begin
        image_0_441 <= io_pixelVal_in_0_2;
      end else if (10'h1b9 == _T_19[9:0]) begin
        image_0_441 <= io_pixelVal_in_0_1;
      end else if (10'h1b9 == _T_15[9:0]) begin
        image_0_441 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_442 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1ba == _T_37[9:0]) begin
        image_0_442 <= io_pixelVal_in_0_7;
      end else if (10'h1ba == _T_34[9:0]) begin
        image_0_442 <= io_pixelVal_in_0_6;
      end else if (10'h1ba == _T_31[9:0]) begin
        image_0_442 <= io_pixelVal_in_0_5;
      end else if (10'h1ba == _T_28[9:0]) begin
        image_0_442 <= io_pixelVal_in_0_4;
      end else if (10'h1ba == _T_25[9:0]) begin
        image_0_442 <= io_pixelVal_in_0_3;
      end else if (10'h1ba == _T_22[9:0]) begin
        image_0_442 <= io_pixelVal_in_0_2;
      end else if (10'h1ba == _T_19[9:0]) begin
        image_0_442 <= io_pixelVal_in_0_1;
      end else if (10'h1ba == _T_15[9:0]) begin
        image_0_442 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_443 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1bb == _T_37[9:0]) begin
        image_0_443 <= io_pixelVal_in_0_7;
      end else if (10'h1bb == _T_34[9:0]) begin
        image_0_443 <= io_pixelVal_in_0_6;
      end else if (10'h1bb == _T_31[9:0]) begin
        image_0_443 <= io_pixelVal_in_0_5;
      end else if (10'h1bb == _T_28[9:0]) begin
        image_0_443 <= io_pixelVal_in_0_4;
      end else if (10'h1bb == _T_25[9:0]) begin
        image_0_443 <= io_pixelVal_in_0_3;
      end else if (10'h1bb == _T_22[9:0]) begin
        image_0_443 <= io_pixelVal_in_0_2;
      end else if (10'h1bb == _T_19[9:0]) begin
        image_0_443 <= io_pixelVal_in_0_1;
      end else if (10'h1bb == _T_15[9:0]) begin
        image_0_443 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_444 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1bc == _T_37[9:0]) begin
        image_0_444 <= io_pixelVal_in_0_7;
      end else if (10'h1bc == _T_34[9:0]) begin
        image_0_444 <= io_pixelVal_in_0_6;
      end else if (10'h1bc == _T_31[9:0]) begin
        image_0_444 <= io_pixelVal_in_0_5;
      end else if (10'h1bc == _T_28[9:0]) begin
        image_0_444 <= io_pixelVal_in_0_4;
      end else if (10'h1bc == _T_25[9:0]) begin
        image_0_444 <= io_pixelVal_in_0_3;
      end else if (10'h1bc == _T_22[9:0]) begin
        image_0_444 <= io_pixelVal_in_0_2;
      end else if (10'h1bc == _T_19[9:0]) begin
        image_0_444 <= io_pixelVal_in_0_1;
      end else if (10'h1bc == _T_15[9:0]) begin
        image_0_444 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_445 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1bd == _T_37[9:0]) begin
        image_0_445 <= io_pixelVal_in_0_7;
      end else if (10'h1bd == _T_34[9:0]) begin
        image_0_445 <= io_pixelVal_in_0_6;
      end else if (10'h1bd == _T_31[9:0]) begin
        image_0_445 <= io_pixelVal_in_0_5;
      end else if (10'h1bd == _T_28[9:0]) begin
        image_0_445 <= io_pixelVal_in_0_4;
      end else if (10'h1bd == _T_25[9:0]) begin
        image_0_445 <= io_pixelVal_in_0_3;
      end else if (10'h1bd == _T_22[9:0]) begin
        image_0_445 <= io_pixelVal_in_0_2;
      end else if (10'h1bd == _T_19[9:0]) begin
        image_0_445 <= io_pixelVal_in_0_1;
      end else if (10'h1bd == _T_15[9:0]) begin
        image_0_445 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_446 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1be == _T_37[9:0]) begin
        image_0_446 <= io_pixelVal_in_0_7;
      end else if (10'h1be == _T_34[9:0]) begin
        image_0_446 <= io_pixelVal_in_0_6;
      end else if (10'h1be == _T_31[9:0]) begin
        image_0_446 <= io_pixelVal_in_0_5;
      end else if (10'h1be == _T_28[9:0]) begin
        image_0_446 <= io_pixelVal_in_0_4;
      end else if (10'h1be == _T_25[9:0]) begin
        image_0_446 <= io_pixelVal_in_0_3;
      end else if (10'h1be == _T_22[9:0]) begin
        image_0_446 <= io_pixelVal_in_0_2;
      end else if (10'h1be == _T_19[9:0]) begin
        image_0_446 <= io_pixelVal_in_0_1;
      end else if (10'h1be == _T_15[9:0]) begin
        image_0_446 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_447 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1bf == _T_37[9:0]) begin
        image_0_447 <= io_pixelVal_in_0_7;
      end else if (10'h1bf == _T_34[9:0]) begin
        image_0_447 <= io_pixelVal_in_0_6;
      end else if (10'h1bf == _T_31[9:0]) begin
        image_0_447 <= io_pixelVal_in_0_5;
      end else if (10'h1bf == _T_28[9:0]) begin
        image_0_447 <= io_pixelVal_in_0_4;
      end else if (10'h1bf == _T_25[9:0]) begin
        image_0_447 <= io_pixelVal_in_0_3;
      end else if (10'h1bf == _T_22[9:0]) begin
        image_0_447 <= io_pixelVal_in_0_2;
      end else if (10'h1bf == _T_19[9:0]) begin
        image_0_447 <= io_pixelVal_in_0_1;
      end else if (10'h1bf == _T_15[9:0]) begin
        image_0_447 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_448 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1c0 == _T_37[9:0]) begin
        image_0_448 <= io_pixelVal_in_0_7;
      end else if (10'h1c0 == _T_34[9:0]) begin
        image_0_448 <= io_pixelVal_in_0_6;
      end else if (10'h1c0 == _T_31[9:0]) begin
        image_0_448 <= io_pixelVal_in_0_5;
      end else if (10'h1c0 == _T_28[9:0]) begin
        image_0_448 <= io_pixelVal_in_0_4;
      end else if (10'h1c0 == _T_25[9:0]) begin
        image_0_448 <= io_pixelVal_in_0_3;
      end else if (10'h1c0 == _T_22[9:0]) begin
        image_0_448 <= io_pixelVal_in_0_2;
      end else if (10'h1c0 == _T_19[9:0]) begin
        image_0_448 <= io_pixelVal_in_0_1;
      end else if (10'h1c0 == _T_15[9:0]) begin
        image_0_448 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_449 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1c1 == _T_37[9:0]) begin
        image_0_449 <= io_pixelVal_in_0_7;
      end else if (10'h1c1 == _T_34[9:0]) begin
        image_0_449 <= io_pixelVal_in_0_6;
      end else if (10'h1c1 == _T_31[9:0]) begin
        image_0_449 <= io_pixelVal_in_0_5;
      end else if (10'h1c1 == _T_28[9:0]) begin
        image_0_449 <= io_pixelVal_in_0_4;
      end else if (10'h1c1 == _T_25[9:0]) begin
        image_0_449 <= io_pixelVal_in_0_3;
      end else if (10'h1c1 == _T_22[9:0]) begin
        image_0_449 <= io_pixelVal_in_0_2;
      end else if (10'h1c1 == _T_19[9:0]) begin
        image_0_449 <= io_pixelVal_in_0_1;
      end else if (10'h1c1 == _T_15[9:0]) begin
        image_0_449 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_450 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1c2 == _T_37[9:0]) begin
        image_0_450 <= io_pixelVal_in_0_7;
      end else if (10'h1c2 == _T_34[9:0]) begin
        image_0_450 <= io_pixelVal_in_0_6;
      end else if (10'h1c2 == _T_31[9:0]) begin
        image_0_450 <= io_pixelVal_in_0_5;
      end else if (10'h1c2 == _T_28[9:0]) begin
        image_0_450 <= io_pixelVal_in_0_4;
      end else if (10'h1c2 == _T_25[9:0]) begin
        image_0_450 <= io_pixelVal_in_0_3;
      end else if (10'h1c2 == _T_22[9:0]) begin
        image_0_450 <= io_pixelVal_in_0_2;
      end else if (10'h1c2 == _T_19[9:0]) begin
        image_0_450 <= io_pixelVal_in_0_1;
      end else if (10'h1c2 == _T_15[9:0]) begin
        image_0_450 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_451 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1c3 == _T_37[9:0]) begin
        image_0_451 <= io_pixelVal_in_0_7;
      end else if (10'h1c3 == _T_34[9:0]) begin
        image_0_451 <= io_pixelVal_in_0_6;
      end else if (10'h1c3 == _T_31[9:0]) begin
        image_0_451 <= io_pixelVal_in_0_5;
      end else if (10'h1c3 == _T_28[9:0]) begin
        image_0_451 <= io_pixelVal_in_0_4;
      end else if (10'h1c3 == _T_25[9:0]) begin
        image_0_451 <= io_pixelVal_in_0_3;
      end else if (10'h1c3 == _T_22[9:0]) begin
        image_0_451 <= io_pixelVal_in_0_2;
      end else if (10'h1c3 == _T_19[9:0]) begin
        image_0_451 <= io_pixelVal_in_0_1;
      end else if (10'h1c3 == _T_15[9:0]) begin
        image_0_451 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_452 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1c4 == _T_37[9:0]) begin
        image_0_452 <= io_pixelVal_in_0_7;
      end else if (10'h1c4 == _T_34[9:0]) begin
        image_0_452 <= io_pixelVal_in_0_6;
      end else if (10'h1c4 == _T_31[9:0]) begin
        image_0_452 <= io_pixelVal_in_0_5;
      end else if (10'h1c4 == _T_28[9:0]) begin
        image_0_452 <= io_pixelVal_in_0_4;
      end else if (10'h1c4 == _T_25[9:0]) begin
        image_0_452 <= io_pixelVal_in_0_3;
      end else if (10'h1c4 == _T_22[9:0]) begin
        image_0_452 <= io_pixelVal_in_0_2;
      end else if (10'h1c4 == _T_19[9:0]) begin
        image_0_452 <= io_pixelVal_in_0_1;
      end else if (10'h1c4 == _T_15[9:0]) begin
        image_0_452 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_453 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1c5 == _T_37[9:0]) begin
        image_0_453 <= io_pixelVal_in_0_7;
      end else if (10'h1c5 == _T_34[9:0]) begin
        image_0_453 <= io_pixelVal_in_0_6;
      end else if (10'h1c5 == _T_31[9:0]) begin
        image_0_453 <= io_pixelVal_in_0_5;
      end else if (10'h1c5 == _T_28[9:0]) begin
        image_0_453 <= io_pixelVal_in_0_4;
      end else if (10'h1c5 == _T_25[9:0]) begin
        image_0_453 <= io_pixelVal_in_0_3;
      end else if (10'h1c5 == _T_22[9:0]) begin
        image_0_453 <= io_pixelVal_in_0_2;
      end else if (10'h1c5 == _T_19[9:0]) begin
        image_0_453 <= io_pixelVal_in_0_1;
      end else if (10'h1c5 == _T_15[9:0]) begin
        image_0_453 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_454 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1c6 == _T_37[9:0]) begin
        image_0_454 <= io_pixelVal_in_0_7;
      end else if (10'h1c6 == _T_34[9:0]) begin
        image_0_454 <= io_pixelVal_in_0_6;
      end else if (10'h1c6 == _T_31[9:0]) begin
        image_0_454 <= io_pixelVal_in_0_5;
      end else if (10'h1c6 == _T_28[9:0]) begin
        image_0_454 <= io_pixelVal_in_0_4;
      end else if (10'h1c6 == _T_25[9:0]) begin
        image_0_454 <= io_pixelVal_in_0_3;
      end else if (10'h1c6 == _T_22[9:0]) begin
        image_0_454 <= io_pixelVal_in_0_2;
      end else if (10'h1c6 == _T_19[9:0]) begin
        image_0_454 <= io_pixelVal_in_0_1;
      end else if (10'h1c6 == _T_15[9:0]) begin
        image_0_454 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_455 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1c7 == _T_37[9:0]) begin
        image_0_455 <= io_pixelVal_in_0_7;
      end else if (10'h1c7 == _T_34[9:0]) begin
        image_0_455 <= io_pixelVal_in_0_6;
      end else if (10'h1c7 == _T_31[9:0]) begin
        image_0_455 <= io_pixelVal_in_0_5;
      end else if (10'h1c7 == _T_28[9:0]) begin
        image_0_455 <= io_pixelVal_in_0_4;
      end else if (10'h1c7 == _T_25[9:0]) begin
        image_0_455 <= io_pixelVal_in_0_3;
      end else if (10'h1c7 == _T_22[9:0]) begin
        image_0_455 <= io_pixelVal_in_0_2;
      end else if (10'h1c7 == _T_19[9:0]) begin
        image_0_455 <= io_pixelVal_in_0_1;
      end else if (10'h1c7 == _T_15[9:0]) begin
        image_0_455 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_456 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1c8 == _T_37[9:0]) begin
        image_0_456 <= io_pixelVal_in_0_7;
      end else if (10'h1c8 == _T_34[9:0]) begin
        image_0_456 <= io_pixelVal_in_0_6;
      end else if (10'h1c8 == _T_31[9:0]) begin
        image_0_456 <= io_pixelVal_in_0_5;
      end else if (10'h1c8 == _T_28[9:0]) begin
        image_0_456 <= io_pixelVal_in_0_4;
      end else if (10'h1c8 == _T_25[9:0]) begin
        image_0_456 <= io_pixelVal_in_0_3;
      end else if (10'h1c8 == _T_22[9:0]) begin
        image_0_456 <= io_pixelVal_in_0_2;
      end else if (10'h1c8 == _T_19[9:0]) begin
        image_0_456 <= io_pixelVal_in_0_1;
      end else if (10'h1c8 == _T_15[9:0]) begin
        image_0_456 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_457 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1c9 == _T_37[9:0]) begin
        image_0_457 <= io_pixelVal_in_0_7;
      end else if (10'h1c9 == _T_34[9:0]) begin
        image_0_457 <= io_pixelVal_in_0_6;
      end else if (10'h1c9 == _T_31[9:0]) begin
        image_0_457 <= io_pixelVal_in_0_5;
      end else if (10'h1c9 == _T_28[9:0]) begin
        image_0_457 <= io_pixelVal_in_0_4;
      end else if (10'h1c9 == _T_25[9:0]) begin
        image_0_457 <= io_pixelVal_in_0_3;
      end else if (10'h1c9 == _T_22[9:0]) begin
        image_0_457 <= io_pixelVal_in_0_2;
      end else if (10'h1c9 == _T_19[9:0]) begin
        image_0_457 <= io_pixelVal_in_0_1;
      end else if (10'h1c9 == _T_15[9:0]) begin
        image_0_457 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_458 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1ca == _T_37[9:0]) begin
        image_0_458 <= io_pixelVal_in_0_7;
      end else if (10'h1ca == _T_34[9:0]) begin
        image_0_458 <= io_pixelVal_in_0_6;
      end else if (10'h1ca == _T_31[9:0]) begin
        image_0_458 <= io_pixelVal_in_0_5;
      end else if (10'h1ca == _T_28[9:0]) begin
        image_0_458 <= io_pixelVal_in_0_4;
      end else if (10'h1ca == _T_25[9:0]) begin
        image_0_458 <= io_pixelVal_in_0_3;
      end else if (10'h1ca == _T_22[9:0]) begin
        image_0_458 <= io_pixelVal_in_0_2;
      end else if (10'h1ca == _T_19[9:0]) begin
        image_0_458 <= io_pixelVal_in_0_1;
      end else if (10'h1ca == _T_15[9:0]) begin
        image_0_458 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_459 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1cb == _T_37[9:0]) begin
        image_0_459 <= io_pixelVal_in_0_7;
      end else if (10'h1cb == _T_34[9:0]) begin
        image_0_459 <= io_pixelVal_in_0_6;
      end else if (10'h1cb == _T_31[9:0]) begin
        image_0_459 <= io_pixelVal_in_0_5;
      end else if (10'h1cb == _T_28[9:0]) begin
        image_0_459 <= io_pixelVal_in_0_4;
      end else if (10'h1cb == _T_25[9:0]) begin
        image_0_459 <= io_pixelVal_in_0_3;
      end else if (10'h1cb == _T_22[9:0]) begin
        image_0_459 <= io_pixelVal_in_0_2;
      end else if (10'h1cb == _T_19[9:0]) begin
        image_0_459 <= io_pixelVal_in_0_1;
      end else if (10'h1cb == _T_15[9:0]) begin
        image_0_459 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_460 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1cc == _T_37[9:0]) begin
        image_0_460 <= io_pixelVal_in_0_7;
      end else if (10'h1cc == _T_34[9:0]) begin
        image_0_460 <= io_pixelVal_in_0_6;
      end else if (10'h1cc == _T_31[9:0]) begin
        image_0_460 <= io_pixelVal_in_0_5;
      end else if (10'h1cc == _T_28[9:0]) begin
        image_0_460 <= io_pixelVal_in_0_4;
      end else if (10'h1cc == _T_25[9:0]) begin
        image_0_460 <= io_pixelVal_in_0_3;
      end else if (10'h1cc == _T_22[9:0]) begin
        image_0_460 <= io_pixelVal_in_0_2;
      end else if (10'h1cc == _T_19[9:0]) begin
        image_0_460 <= io_pixelVal_in_0_1;
      end else if (10'h1cc == _T_15[9:0]) begin
        image_0_460 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_461 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1cd == _T_37[9:0]) begin
        image_0_461 <= io_pixelVal_in_0_7;
      end else if (10'h1cd == _T_34[9:0]) begin
        image_0_461 <= io_pixelVal_in_0_6;
      end else if (10'h1cd == _T_31[9:0]) begin
        image_0_461 <= io_pixelVal_in_0_5;
      end else if (10'h1cd == _T_28[9:0]) begin
        image_0_461 <= io_pixelVal_in_0_4;
      end else if (10'h1cd == _T_25[9:0]) begin
        image_0_461 <= io_pixelVal_in_0_3;
      end else if (10'h1cd == _T_22[9:0]) begin
        image_0_461 <= io_pixelVal_in_0_2;
      end else if (10'h1cd == _T_19[9:0]) begin
        image_0_461 <= io_pixelVal_in_0_1;
      end else if (10'h1cd == _T_15[9:0]) begin
        image_0_461 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_462 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1ce == _T_37[9:0]) begin
        image_0_462 <= io_pixelVal_in_0_7;
      end else if (10'h1ce == _T_34[9:0]) begin
        image_0_462 <= io_pixelVal_in_0_6;
      end else if (10'h1ce == _T_31[9:0]) begin
        image_0_462 <= io_pixelVal_in_0_5;
      end else if (10'h1ce == _T_28[9:0]) begin
        image_0_462 <= io_pixelVal_in_0_4;
      end else if (10'h1ce == _T_25[9:0]) begin
        image_0_462 <= io_pixelVal_in_0_3;
      end else if (10'h1ce == _T_22[9:0]) begin
        image_0_462 <= io_pixelVal_in_0_2;
      end else if (10'h1ce == _T_19[9:0]) begin
        image_0_462 <= io_pixelVal_in_0_1;
      end else if (10'h1ce == _T_15[9:0]) begin
        image_0_462 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_463 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1cf == _T_37[9:0]) begin
        image_0_463 <= io_pixelVal_in_0_7;
      end else if (10'h1cf == _T_34[9:0]) begin
        image_0_463 <= io_pixelVal_in_0_6;
      end else if (10'h1cf == _T_31[9:0]) begin
        image_0_463 <= io_pixelVal_in_0_5;
      end else if (10'h1cf == _T_28[9:0]) begin
        image_0_463 <= io_pixelVal_in_0_4;
      end else if (10'h1cf == _T_25[9:0]) begin
        image_0_463 <= io_pixelVal_in_0_3;
      end else if (10'h1cf == _T_22[9:0]) begin
        image_0_463 <= io_pixelVal_in_0_2;
      end else if (10'h1cf == _T_19[9:0]) begin
        image_0_463 <= io_pixelVal_in_0_1;
      end else if (10'h1cf == _T_15[9:0]) begin
        image_0_463 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_464 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1d0 == _T_37[9:0]) begin
        image_0_464 <= io_pixelVal_in_0_7;
      end else if (10'h1d0 == _T_34[9:0]) begin
        image_0_464 <= io_pixelVal_in_0_6;
      end else if (10'h1d0 == _T_31[9:0]) begin
        image_0_464 <= io_pixelVal_in_0_5;
      end else if (10'h1d0 == _T_28[9:0]) begin
        image_0_464 <= io_pixelVal_in_0_4;
      end else if (10'h1d0 == _T_25[9:0]) begin
        image_0_464 <= io_pixelVal_in_0_3;
      end else if (10'h1d0 == _T_22[9:0]) begin
        image_0_464 <= io_pixelVal_in_0_2;
      end else if (10'h1d0 == _T_19[9:0]) begin
        image_0_464 <= io_pixelVal_in_0_1;
      end else if (10'h1d0 == _T_15[9:0]) begin
        image_0_464 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_465 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1d1 == _T_37[9:0]) begin
        image_0_465 <= io_pixelVal_in_0_7;
      end else if (10'h1d1 == _T_34[9:0]) begin
        image_0_465 <= io_pixelVal_in_0_6;
      end else if (10'h1d1 == _T_31[9:0]) begin
        image_0_465 <= io_pixelVal_in_0_5;
      end else if (10'h1d1 == _T_28[9:0]) begin
        image_0_465 <= io_pixelVal_in_0_4;
      end else if (10'h1d1 == _T_25[9:0]) begin
        image_0_465 <= io_pixelVal_in_0_3;
      end else if (10'h1d1 == _T_22[9:0]) begin
        image_0_465 <= io_pixelVal_in_0_2;
      end else if (10'h1d1 == _T_19[9:0]) begin
        image_0_465 <= io_pixelVal_in_0_1;
      end else if (10'h1d1 == _T_15[9:0]) begin
        image_0_465 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_466 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1d2 == _T_37[9:0]) begin
        image_0_466 <= io_pixelVal_in_0_7;
      end else if (10'h1d2 == _T_34[9:0]) begin
        image_0_466 <= io_pixelVal_in_0_6;
      end else if (10'h1d2 == _T_31[9:0]) begin
        image_0_466 <= io_pixelVal_in_0_5;
      end else if (10'h1d2 == _T_28[9:0]) begin
        image_0_466 <= io_pixelVal_in_0_4;
      end else if (10'h1d2 == _T_25[9:0]) begin
        image_0_466 <= io_pixelVal_in_0_3;
      end else if (10'h1d2 == _T_22[9:0]) begin
        image_0_466 <= io_pixelVal_in_0_2;
      end else if (10'h1d2 == _T_19[9:0]) begin
        image_0_466 <= io_pixelVal_in_0_1;
      end else if (10'h1d2 == _T_15[9:0]) begin
        image_0_466 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_467 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1d3 == _T_37[9:0]) begin
        image_0_467 <= io_pixelVal_in_0_7;
      end else if (10'h1d3 == _T_34[9:0]) begin
        image_0_467 <= io_pixelVal_in_0_6;
      end else if (10'h1d3 == _T_31[9:0]) begin
        image_0_467 <= io_pixelVal_in_0_5;
      end else if (10'h1d3 == _T_28[9:0]) begin
        image_0_467 <= io_pixelVal_in_0_4;
      end else if (10'h1d3 == _T_25[9:0]) begin
        image_0_467 <= io_pixelVal_in_0_3;
      end else if (10'h1d3 == _T_22[9:0]) begin
        image_0_467 <= io_pixelVal_in_0_2;
      end else if (10'h1d3 == _T_19[9:0]) begin
        image_0_467 <= io_pixelVal_in_0_1;
      end else if (10'h1d3 == _T_15[9:0]) begin
        image_0_467 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_468 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1d4 == _T_37[9:0]) begin
        image_0_468 <= io_pixelVal_in_0_7;
      end else if (10'h1d4 == _T_34[9:0]) begin
        image_0_468 <= io_pixelVal_in_0_6;
      end else if (10'h1d4 == _T_31[9:0]) begin
        image_0_468 <= io_pixelVal_in_0_5;
      end else if (10'h1d4 == _T_28[9:0]) begin
        image_0_468 <= io_pixelVal_in_0_4;
      end else if (10'h1d4 == _T_25[9:0]) begin
        image_0_468 <= io_pixelVal_in_0_3;
      end else if (10'h1d4 == _T_22[9:0]) begin
        image_0_468 <= io_pixelVal_in_0_2;
      end else if (10'h1d4 == _T_19[9:0]) begin
        image_0_468 <= io_pixelVal_in_0_1;
      end else if (10'h1d4 == _T_15[9:0]) begin
        image_0_468 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_469 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1d5 == _T_37[9:0]) begin
        image_0_469 <= io_pixelVal_in_0_7;
      end else if (10'h1d5 == _T_34[9:0]) begin
        image_0_469 <= io_pixelVal_in_0_6;
      end else if (10'h1d5 == _T_31[9:0]) begin
        image_0_469 <= io_pixelVal_in_0_5;
      end else if (10'h1d5 == _T_28[9:0]) begin
        image_0_469 <= io_pixelVal_in_0_4;
      end else if (10'h1d5 == _T_25[9:0]) begin
        image_0_469 <= io_pixelVal_in_0_3;
      end else if (10'h1d5 == _T_22[9:0]) begin
        image_0_469 <= io_pixelVal_in_0_2;
      end else if (10'h1d5 == _T_19[9:0]) begin
        image_0_469 <= io_pixelVal_in_0_1;
      end else if (10'h1d5 == _T_15[9:0]) begin
        image_0_469 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_470 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1d6 == _T_37[9:0]) begin
        image_0_470 <= io_pixelVal_in_0_7;
      end else if (10'h1d6 == _T_34[9:0]) begin
        image_0_470 <= io_pixelVal_in_0_6;
      end else if (10'h1d6 == _T_31[9:0]) begin
        image_0_470 <= io_pixelVal_in_0_5;
      end else if (10'h1d6 == _T_28[9:0]) begin
        image_0_470 <= io_pixelVal_in_0_4;
      end else if (10'h1d6 == _T_25[9:0]) begin
        image_0_470 <= io_pixelVal_in_0_3;
      end else if (10'h1d6 == _T_22[9:0]) begin
        image_0_470 <= io_pixelVal_in_0_2;
      end else if (10'h1d6 == _T_19[9:0]) begin
        image_0_470 <= io_pixelVal_in_0_1;
      end else if (10'h1d6 == _T_15[9:0]) begin
        image_0_470 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_471 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1d7 == _T_37[9:0]) begin
        image_0_471 <= io_pixelVal_in_0_7;
      end else if (10'h1d7 == _T_34[9:0]) begin
        image_0_471 <= io_pixelVal_in_0_6;
      end else if (10'h1d7 == _T_31[9:0]) begin
        image_0_471 <= io_pixelVal_in_0_5;
      end else if (10'h1d7 == _T_28[9:0]) begin
        image_0_471 <= io_pixelVal_in_0_4;
      end else if (10'h1d7 == _T_25[9:0]) begin
        image_0_471 <= io_pixelVal_in_0_3;
      end else if (10'h1d7 == _T_22[9:0]) begin
        image_0_471 <= io_pixelVal_in_0_2;
      end else if (10'h1d7 == _T_19[9:0]) begin
        image_0_471 <= io_pixelVal_in_0_1;
      end else if (10'h1d7 == _T_15[9:0]) begin
        image_0_471 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_472 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1d8 == _T_37[9:0]) begin
        image_0_472 <= io_pixelVal_in_0_7;
      end else if (10'h1d8 == _T_34[9:0]) begin
        image_0_472 <= io_pixelVal_in_0_6;
      end else if (10'h1d8 == _T_31[9:0]) begin
        image_0_472 <= io_pixelVal_in_0_5;
      end else if (10'h1d8 == _T_28[9:0]) begin
        image_0_472 <= io_pixelVal_in_0_4;
      end else if (10'h1d8 == _T_25[9:0]) begin
        image_0_472 <= io_pixelVal_in_0_3;
      end else if (10'h1d8 == _T_22[9:0]) begin
        image_0_472 <= io_pixelVal_in_0_2;
      end else if (10'h1d8 == _T_19[9:0]) begin
        image_0_472 <= io_pixelVal_in_0_1;
      end else if (10'h1d8 == _T_15[9:0]) begin
        image_0_472 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_473 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1d9 == _T_37[9:0]) begin
        image_0_473 <= io_pixelVal_in_0_7;
      end else if (10'h1d9 == _T_34[9:0]) begin
        image_0_473 <= io_pixelVal_in_0_6;
      end else if (10'h1d9 == _T_31[9:0]) begin
        image_0_473 <= io_pixelVal_in_0_5;
      end else if (10'h1d9 == _T_28[9:0]) begin
        image_0_473 <= io_pixelVal_in_0_4;
      end else if (10'h1d9 == _T_25[9:0]) begin
        image_0_473 <= io_pixelVal_in_0_3;
      end else if (10'h1d9 == _T_22[9:0]) begin
        image_0_473 <= io_pixelVal_in_0_2;
      end else if (10'h1d9 == _T_19[9:0]) begin
        image_0_473 <= io_pixelVal_in_0_1;
      end else if (10'h1d9 == _T_15[9:0]) begin
        image_0_473 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_474 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1da == _T_37[9:0]) begin
        image_0_474 <= io_pixelVal_in_0_7;
      end else if (10'h1da == _T_34[9:0]) begin
        image_0_474 <= io_pixelVal_in_0_6;
      end else if (10'h1da == _T_31[9:0]) begin
        image_0_474 <= io_pixelVal_in_0_5;
      end else if (10'h1da == _T_28[9:0]) begin
        image_0_474 <= io_pixelVal_in_0_4;
      end else if (10'h1da == _T_25[9:0]) begin
        image_0_474 <= io_pixelVal_in_0_3;
      end else if (10'h1da == _T_22[9:0]) begin
        image_0_474 <= io_pixelVal_in_0_2;
      end else if (10'h1da == _T_19[9:0]) begin
        image_0_474 <= io_pixelVal_in_0_1;
      end else if (10'h1da == _T_15[9:0]) begin
        image_0_474 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_475 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1db == _T_37[9:0]) begin
        image_0_475 <= io_pixelVal_in_0_7;
      end else if (10'h1db == _T_34[9:0]) begin
        image_0_475 <= io_pixelVal_in_0_6;
      end else if (10'h1db == _T_31[9:0]) begin
        image_0_475 <= io_pixelVal_in_0_5;
      end else if (10'h1db == _T_28[9:0]) begin
        image_0_475 <= io_pixelVal_in_0_4;
      end else if (10'h1db == _T_25[9:0]) begin
        image_0_475 <= io_pixelVal_in_0_3;
      end else if (10'h1db == _T_22[9:0]) begin
        image_0_475 <= io_pixelVal_in_0_2;
      end else if (10'h1db == _T_19[9:0]) begin
        image_0_475 <= io_pixelVal_in_0_1;
      end else if (10'h1db == _T_15[9:0]) begin
        image_0_475 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_476 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1dc == _T_37[9:0]) begin
        image_0_476 <= io_pixelVal_in_0_7;
      end else if (10'h1dc == _T_34[9:0]) begin
        image_0_476 <= io_pixelVal_in_0_6;
      end else if (10'h1dc == _T_31[9:0]) begin
        image_0_476 <= io_pixelVal_in_0_5;
      end else if (10'h1dc == _T_28[9:0]) begin
        image_0_476 <= io_pixelVal_in_0_4;
      end else if (10'h1dc == _T_25[9:0]) begin
        image_0_476 <= io_pixelVal_in_0_3;
      end else if (10'h1dc == _T_22[9:0]) begin
        image_0_476 <= io_pixelVal_in_0_2;
      end else if (10'h1dc == _T_19[9:0]) begin
        image_0_476 <= io_pixelVal_in_0_1;
      end else if (10'h1dc == _T_15[9:0]) begin
        image_0_476 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_477 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1dd == _T_37[9:0]) begin
        image_0_477 <= io_pixelVal_in_0_7;
      end else if (10'h1dd == _T_34[9:0]) begin
        image_0_477 <= io_pixelVal_in_0_6;
      end else if (10'h1dd == _T_31[9:0]) begin
        image_0_477 <= io_pixelVal_in_0_5;
      end else if (10'h1dd == _T_28[9:0]) begin
        image_0_477 <= io_pixelVal_in_0_4;
      end else if (10'h1dd == _T_25[9:0]) begin
        image_0_477 <= io_pixelVal_in_0_3;
      end else if (10'h1dd == _T_22[9:0]) begin
        image_0_477 <= io_pixelVal_in_0_2;
      end else if (10'h1dd == _T_19[9:0]) begin
        image_0_477 <= io_pixelVal_in_0_1;
      end else if (10'h1dd == _T_15[9:0]) begin
        image_0_477 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_478 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1de == _T_37[9:0]) begin
        image_0_478 <= io_pixelVal_in_0_7;
      end else if (10'h1de == _T_34[9:0]) begin
        image_0_478 <= io_pixelVal_in_0_6;
      end else if (10'h1de == _T_31[9:0]) begin
        image_0_478 <= io_pixelVal_in_0_5;
      end else if (10'h1de == _T_28[9:0]) begin
        image_0_478 <= io_pixelVal_in_0_4;
      end else if (10'h1de == _T_25[9:0]) begin
        image_0_478 <= io_pixelVal_in_0_3;
      end else if (10'h1de == _T_22[9:0]) begin
        image_0_478 <= io_pixelVal_in_0_2;
      end else if (10'h1de == _T_19[9:0]) begin
        image_0_478 <= io_pixelVal_in_0_1;
      end else if (10'h1de == _T_15[9:0]) begin
        image_0_478 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_479 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1df == _T_37[9:0]) begin
        image_0_479 <= io_pixelVal_in_0_7;
      end else if (10'h1df == _T_34[9:0]) begin
        image_0_479 <= io_pixelVal_in_0_6;
      end else if (10'h1df == _T_31[9:0]) begin
        image_0_479 <= io_pixelVal_in_0_5;
      end else if (10'h1df == _T_28[9:0]) begin
        image_0_479 <= io_pixelVal_in_0_4;
      end else if (10'h1df == _T_25[9:0]) begin
        image_0_479 <= io_pixelVal_in_0_3;
      end else if (10'h1df == _T_22[9:0]) begin
        image_0_479 <= io_pixelVal_in_0_2;
      end else if (10'h1df == _T_19[9:0]) begin
        image_0_479 <= io_pixelVal_in_0_1;
      end else if (10'h1df == _T_15[9:0]) begin
        image_0_479 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_480 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1e0 == _T_37[9:0]) begin
        image_0_480 <= io_pixelVal_in_0_7;
      end else if (10'h1e0 == _T_34[9:0]) begin
        image_0_480 <= io_pixelVal_in_0_6;
      end else if (10'h1e0 == _T_31[9:0]) begin
        image_0_480 <= io_pixelVal_in_0_5;
      end else if (10'h1e0 == _T_28[9:0]) begin
        image_0_480 <= io_pixelVal_in_0_4;
      end else if (10'h1e0 == _T_25[9:0]) begin
        image_0_480 <= io_pixelVal_in_0_3;
      end else if (10'h1e0 == _T_22[9:0]) begin
        image_0_480 <= io_pixelVal_in_0_2;
      end else if (10'h1e0 == _T_19[9:0]) begin
        image_0_480 <= io_pixelVal_in_0_1;
      end else if (10'h1e0 == _T_15[9:0]) begin
        image_0_480 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_481 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1e1 == _T_37[9:0]) begin
        image_0_481 <= io_pixelVal_in_0_7;
      end else if (10'h1e1 == _T_34[9:0]) begin
        image_0_481 <= io_pixelVal_in_0_6;
      end else if (10'h1e1 == _T_31[9:0]) begin
        image_0_481 <= io_pixelVal_in_0_5;
      end else if (10'h1e1 == _T_28[9:0]) begin
        image_0_481 <= io_pixelVal_in_0_4;
      end else if (10'h1e1 == _T_25[9:0]) begin
        image_0_481 <= io_pixelVal_in_0_3;
      end else if (10'h1e1 == _T_22[9:0]) begin
        image_0_481 <= io_pixelVal_in_0_2;
      end else if (10'h1e1 == _T_19[9:0]) begin
        image_0_481 <= io_pixelVal_in_0_1;
      end else if (10'h1e1 == _T_15[9:0]) begin
        image_0_481 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_482 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1e2 == _T_37[9:0]) begin
        image_0_482 <= io_pixelVal_in_0_7;
      end else if (10'h1e2 == _T_34[9:0]) begin
        image_0_482 <= io_pixelVal_in_0_6;
      end else if (10'h1e2 == _T_31[9:0]) begin
        image_0_482 <= io_pixelVal_in_0_5;
      end else if (10'h1e2 == _T_28[9:0]) begin
        image_0_482 <= io_pixelVal_in_0_4;
      end else if (10'h1e2 == _T_25[9:0]) begin
        image_0_482 <= io_pixelVal_in_0_3;
      end else if (10'h1e2 == _T_22[9:0]) begin
        image_0_482 <= io_pixelVal_in_0_2;
      end else if (10'h1e2 == _T_19[9:0]) begin
        image_0_482 <= io_pixelVal_in_0_1;
      end else if (10'h1e2 == _T_15[9:0]) begin
        image_0_482 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_483 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1e3 == _T_37[9:0]) begin
        image_0_483 <= io_pixelVal_in_0_7;
      end else if (10'h1e3 == _T_34[9:0]) begin
        image_0_483 <= io_pixelVal_in_0_6;
      end else if (10'h1e3 == _T_31[9:0]) begin
        image_0_483 <= io_pixelVal_in_0_5;
      end else if (10'h1e3 == _T_28[9:0]) begin
        image_0_483 <= io_pixelVal_in_0_4;
      end else if (10'h1e3 == _T_25[9:0]) begin
        image_0_483 <= io_pixelVal_in_0_3;
      end else if (10'h1e3 == _T_22[9:0]) begin
        image_0_483 <= io_pixelVal_in_0_2;
      end else if (10'h1e3 == _T_19[9:0]) begin
        image_0_483 <= io_pixelVal_in_0_1;
      end else if (10'h1e3 == _T_15[9:0]) begin
        image_0_483 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_484 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1e4 == _T_37[9:0]) begin
        image_0_484 <= io_pixelVal_in_0_7;
      end else if (10'h1e4 == _T_34[9:0]) begin
        image_0_484 <= io_pixelVal_in_0_6;
      end else if (10'h1e4 == _T_31[9:0]) begin
        image_0_484 <= io_pixelVal_in_0_5;
      end else if (10'h1e4 == _T_28[9:0]) begin
        image_0_484 <= io_pixelVal_in_0_4;
      end else if (10'h1e4 == _T_25[9:0]) begin
        image_0_484 <= io_pixelVal_in_0_3;
      end else if (10'h1e4 == _T_22[9:0]) begin
        image_0_484 <= io_pixelVal_in_0_2;
      end else if (10'h1e4 == _T_19[9:0]) begin
        image_0_484 <= io_pixelVal_in_0_1;
      end else if (10'h1e4 == _T_15[9:0]) begin
        image_0_484 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_485 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1e5 == _T_37[9:0]) begin
        image_0_485 <= io_pixelVal_in_0_7;
      end else if (10'h1e5 == _T_34[9:0]) begin
        image_0_485 <= io_pixelVal_in_0_6;
      end else if (10'h1e5 == _T_31[9:0]) begin
        image_0_485 <= io_pixelVal_in_0_5;
      end else if (10'h1e5 == _T_28[9:0]) begin
        image_0_485 <= io_pixelVal_in_0_4;
      end else if (10'h1e5 == _T_25[9:0]) begin
        image_0_485 <= io_pixelVal_in_0_3;
      end else if (10'h1e5 == _T_22[9:0]) begin
        image_0_485 <= io_pixelVal_in_0_2;
      end else if (10'h1e5 == _T_19[9:0]) begin
        image_0_485 <= io_pixelVal_in_0_1;
      end else if (10'h1e5 == _T_15[9:0]) begin
        image_0_485 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_486 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1e6 == _T_37[9:0]) begin
        image_0_486 <= io_pixelVal_in_0_7;
      end else if (10'h1e6 == _T_34[9:0]) begin
        image_0_486 <= io_pixelVal_in_0_6;
      end else if (10'h1e6 == _T_31[9:0]) begin
        image_0_486 <= io_pixelVal_in_0_5;
      end else if (10'h1e6 == _T_28[9:0]) begin
        image_0_486 <= io_pixelVal_in_0_4;
      end else if (10'h1e6 == _T_25[9:0]) begin
        image_0_486 <= io_pixelVal_in_0_3;
      end else if (10'h1e6 == _T_22[9:0]) begin
        image_0_486 <= io_pixelVal_in_0_2;
      end else if (10'h1e6 == _T_19[9:0]) begin
        image_0_486 <= io_pixelVal_in_0_1;
      end else if (10'h1e6 == _T_15[9:0]) begin
        image_0_486 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_487 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1e7 == _T_37[9:0]) begin
        image_0_487 <= io_pixelVal_in_0_7;
      end else if (10'h1e7 == _T_34[9:0]) begin
        image_0_487 <= io_pixelVal_in_0_6;
      end else if (10'h1e7 == _T_31[9:0]) begin
        image_0_487 <= io_pixelVal_in_0_5;
      end else if (10'h1e7 == _T_28[9:0]) begin
        image_0_487 <= io_pixelVal_in_0_4;
      end else if (10'h1e7 == _T_25[9:0]) begin
        image_0_487 <= io_pixelVal_in_0_3;
      end else if (10'h1e7 == _T_22[9:0]) begin
        image_0_487 <= io_pixelVal_in_0_2;
      end else if (10'h1e7 == _T_19[9:0]) begin
        image_0_487 <= io_pixelVal_in_0_1;
      end else if (10'h1e7 == _T_15[9:0]) begin
        image_0_487 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_488 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1e8 == _T_37[9:0]) begin
        image_0_488 <= io_pixelVal_in_0_7;
      end else if (10'h1e8 == _T_34[9:0]) begin
        image_0_488 <= io_pixelVal_in_0_6;
      end else if (10'h1e8 == _T_31[9:0]) begin
        image_0_488 <= io_pixelVal_in_0_5;
      end else if (10'h1e8 == _T_28[9:0]) begin
        image_0_488 <= io_pixelVal_in_0_4;
      end else if (10'h1e8 == _T_25[9:0]) begin
        image_0_488 <= io_pixelVal_in_0_3;
      end else if (10'h1e8 == _T_22[9:0]) begin
        image_0_488 <= io_pixelVal_in_0_2;
      end else if (10'h1e8 == _T_19[9:0]) begin
        image_0_488 <= io_pixelVal_in_0_1;
      end else if (10'h1e8 == _T_15[9:0]) begin
        image_0_488 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_489 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1e9 == _T_37[9:0]) begin
        image_0_489 <= io_pixelVal_in_0_7;
      end else if (10'h1e9 == _T_34[9:0]) begin
        image_0_489 <= io_pixelVal_in_0_6;
      end else if (10'h1e9 == _T_31[9:0]) begin
        image_0_489 <= io_pixelVal_in_0_5;
      end else if (10'h1e9 == _T_28[9:0]) begin
        image_0_489 <= io_pixelVal_in_0_4;
      end else if (10'h1e9 == _T_25[9:0]) begin
        image_0_489 <= io_pixelVal_in_0_3;
      end else if (10'h1e9 == _T_22[9:0]) begin
        image_0_489 <= io_pixelVal_in_0_2;
      end else if (10'h1e9 == _T_19[9:0]) begin
        image_0_489 <= io_pixelVal_in_0_1;
      end else if (10'h1e9 == _T_15[9:0]) begin
        image_0_489 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_490 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1ea == _T_37[9:0]) begin
        image_0_490 <= io_pixelVal_in_0_7;
      end else if (10'h1ea == _T_34[9:0]) begin
        image_0_490 <= io_pixelVal_in_0_6;
      end else if (10'h1ea == _T_31[9:0]) begin
        image_0_490 <= io_pixelVal_in_0_5;
      end else if (10'h1ea == _T_28[9:0]) begin
        image_0_490 <= io_pixelVal_in_0_4;
      end else if (10'h1ea == _T_25[9:0]) begin
        image_0_490 <= io_pixelVal_in_0_3;
      end else if (10'h1ea == _T_22[9:0]) begin
        image_0_490 <= io_pixelVal_in_0_2;
      end else if (10'h1ea == _T_19[9:0]) begin
        image_0_490 <= io_pixelVal_in_0_1;
      end else if (10'h1ea == _T_15[9:0]) begin
        image_0_490 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_491 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1eb == _T_37[9:0]) begin
        image_0_491 <= io_pixelVal_in_0_7;
      end else if (10'h1eb == _T_34[9:0]) begin
        image_0_491 <= io_pixelVal_in_0_6;
      end else if (10'h1eb == _T_31[9:0]) begin
        image_0_491 <= io_pixelVal_in_0_5;
      end else if (10'h1eb == _T_28[9:0]) begin
        image_0_491 <= io_pixelVal_in_0_4;
      end else if (10'h1eb == _T_25[9:0]) begin
        image_0_491 <= io_pixelVal_in_0_3;
      end else if (10'h1eb == _T_22[9:0]) begin
        image_0_491 <= io_pixelVal_in_0_2;
      end else if (10'h1eb == _T_19[9:0]) begin
        image_0_491 <= io_pixelVal_in_0_1;
      end else if (10'h1eb == _T_15[9:0]) begin
        image_0_491 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_492 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1ec == _T_37[9:0]) begin
        image_0_492 <= io_pixelVal_in_0_7;
      end else if (10'h1ec == _T_34[9:0]) begin
        image_0_492 <= io_pixelVal_in_0_6;
      end else if (10'h1ec == _T_31[9:0]) begin
        image_0_492 <= io_pixelVal_in_0_5;
      end else if (10'h1ec == _T_28[9:0]) begin
        image_0_492 <= io_pixelVal_in_0_4;
      end else if (10'h1ec == _T_25[9:0]) begin
        image_0_492 <= io_pixelVal_in_0_3;
      end else if (10'h1ec == _T_22[9:0]) begin
        image_0_492 <= io_pixelVal_in_0_2;
      end else if (10'h1ec == _T_19[9:0]) begin
        image_0_492 <= io_pixelVal_in_0_1;
      end else if (10'h1ec == _T_15[9:0]) begin
        image_0_492 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_493 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1ed == _T_37[9:0]) begin
        image_0_493 <= io_pixelVal_in_0_7;
      end else if (10'h1ed == _T_34[9:0]) begin
        image_0_493 <= io_pixelVal_in_0_6;
      end else if (10'h1ed == _T_31[9:0]) begin
        image_0_493 <= io_pixelVal_in_0_5;
      end else if (10'h1ed == _T_28[9:0]) begin
        image_0_493 <= io_pixelVal_in_0_4;
      end else if (10'h1ed == _T_25[9:0]) begin
        image_0_493 <= io_pixelVal_in_0_3;
      end else if (10'h1ed == _T_22[9:0]) begin
        image_0_493 <= io_pixelVal_in_0_2;
      end else if (10'h1ed == _T_19[9:0]) begin
        image_0_493 <= io_pixelVal_in_0_1;
      end else if (10'h1ed == _T_15[9:0]) begin
        image_0_493 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_494 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1ee == _T_37[9:0]) begin
        image_0_494 <= io_pixelVal_in_0_7;
      end else if (10'h1ee == _T_34[9:0]) begin
        image_0_494 <= io_pixelVal_in_0_6;
      end else if (10'h1ee == _T_31[9:0]) begin
        image_0_494 <= io_pixelVal_in_0_5;
      end else if (10'h1ee == _T_28[9:0]) begin
        image_0_494 <= io_pixelVal_in_0_4;
      end else if (10'h1ee == _T_25[9:0]) begin
        image_0_494 <= io_pixelVal_in_0_3;
      end else if (10'h1ee == _T_22[9:0]) begin
        image_0_494 <= io_pixelVal_in_0_2;
      end else if (10'h1ee == _T_19[9:0]) begin
        image_0_494 <= io_pixelVal_in_0_1;
      end else if (10'h1ee == _T_15[9:0]) begin
        image_0_494 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_495 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1ef == _T_37[9:0]) begin
        image_0_495 <= io_pixelVal_in_0_7;
      end else if (10'h1ef == _T_34[9:0]) begin
        image_0_495 <= io_pixelVal_in_0_6;
      end else if (10'h1ef == _T_31[9:0]) begin
        image_0_495 <= io_pixelVal_in_0_5;
      end else if (10'h1ef == _T_28[9:0]) begin
        image_0_495 <= io_pixelVal_in_0_4;
      end else if (10'h1ef == _T_25[9:0]) begin
        image_0_495 <= io_pixelVal_in_0_3;
      end else if (10'h1ef == _T_22[9:0]) begin
        image_0_495 <= io_pixelVal_in_0_2;
      end else if (10'h1ef == _T_19[9:0]) begin
        image_0_495 <= io_pixelVal_in_0_1;
      end else if (10'h1ef == _T_15[9:0]) begin
        image_0_495 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_496 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1f0 == _T_37[9:0]) begin
        image_0_496 <= io_pixelVal_in_0_7;
      end else if (10'h1f0 == _T_34[9:0]) begin
        image_0_496 <= io_pixelVal_in_0_6;
      end else if (10'h1f0 == _T_31[9:0]) begin
        image_0_496 <= io_pixelVal_in_0_5;
      end else if (10'h1f0 == _T_28[9:0]) begin
        image_0_496 <= io_pixelVal_in_0_4;
      end else if (10'h1f0 == _T_25[9:0]) begin
        image_0_496 <= io_pixelVal_in_0_3;
      end else if (10'h1f0 == _T_22[9:0]) begin
        image_0_496 <= io_pixelVal_in_0_2;
      end else if (10'h1f0 == _T_19[9:0]) begin
        image_0_496 <= io_pixelVal_in_0_1;
      end else if (10'h1f0 == _T_15[9:0]) begin
        image_0_496 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_497 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1f1 == _T_37[9:0]) begin
        image_0_497 <= io_pixelVal_in_0_7;
      end else if (10'h1f1 == _T_34[9:0]) begin
        image_0_497 <= io_pixelVal_in_0_6;
      end else if (10'h1f1 == _T_31[9:0]) begin
        image_0_497 <= io_pixelVal_in_0_5;
      end else if (10'h1f1 == _T_28[9:0]) begin
        image_0_497 <= io_pixelVal_in_0_4;
      end else if (10'h1f1 == _T_25[9:0]) begin
        image_0_497 <= io_pixelVal_in_0_3;
      end else if (10'h1f1 == _T_22[9:0]) begin
        image_0_497 <= io_pixelVal_in_0_2;
      end else if (10'h1f1 == _T_19[9:0]) begin
        image_0_497 <= io_pixelVal_in_0_1;
      end else if (10'h1f1 == _T_15[9:0]) begin
        image_0_497 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_498 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1f2 == _T_37[9:0]) begin
        image_0_498 <= io_pixelVal_in_0_7;
      end else if (10'h1f2 == _T_34[9:0]) begin
        image_0_498 <= io_pixelVal_in_0_6;
      end else if (10'h1f2 == _T_31[9:0]) begin
        image_0_498 <= io_pixelVal_in_0_5;
      end else if (10'h1f2 == _T_28[9:0]) begin
        image_0_498 <= io_pixelVal_in_0_4;
      end else if (10'h1f2 == _T_25[9:0]) begin
        image_0_498 <= io_pixelVal_in_0_3;
      end else if (10'h1f2 == _T_22[9:0]) begin
        image_0_498 <= io_pixelVal_in_0_2;
      end else if (10'h1f2 == _T_19[9:0]) begin
        image_0_498 <= io_pixelVal_in_0_1;
      end else if (10'h1f2 == _T_15[9:0]) begin
        image_0_498 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_499 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1f3 == _T_37[9:0]) begin
        image_0_499 <= io_pixelVal_in_0_7;
      end else if (10'h1f3 == _T_34[9:0]) begin
        image_0_499 <= io_pixelVal_in_0_6;
      end else if (10'h1f3 == _T_31[9:0]) begin
        image_0_499 <= io_pixelVal_in_0_5;
      end else if (10'h1f3 == _T_28[9:0]) begin
        image_0_499 <= io_pixelVal_in_0_4;
      end else if (10'h1f3 == _T_25[9:0]) begin
        image_0_499 <= io_pixelVal_in_0_3;
      end else if (10'h1f3 == _T_22[9:0]) begin
        image_0_499 <= io_pixelVal_in_0_2;
      end else if (10'h1f3 == _T_19[9:0]) begin
        image_0_499 <= io_pixelVal_in_0_1;
      end else if (10'h1f3 == _T_15[9:0]) begin
        image_0_499 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_500 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1f4 == _T_37[9:0]) begin
        image_0_500 <= io_pixelVal_in_0_7;
      end else if (10'h1f4 == _T_34[9:0]) begin
        image_0_500 <= io_pixelVal_in_0_6;
      end else if (10'h1f4 == _T_31[9:0]) begin
        image_0_500 <= io_pixelVal_in_0_5;
      end else if (10'h1f4 == _T_28[9:0]) begin
        image_0_500 <= io_pixelVal_in_0_4;
      end else if (10'h1f4 == _T_25[9:0]) begin
        image_0_500 <= io_pixelVal_in_0_3;
      end else if (10'h1f4 == _T_22[9:0]) begin
        image_0_500 <= io_pixelVal_in_0_2;
      end else if (10'h1f4 == _T_19[9:0]) begin
        image_0_500 <= io_pixelVal_in_0_1;
      end else if (10'h1f4 == _T_15[9:0]) begin
        image_0_500 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_501 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1f5 == _T_37[9:0]) begin
        image_0_501 <= io_pixelVal_in_0_7;
      end else if (10'h1f5 == _T_34[9:0]) begin
        image_0_501 <= io_pixelVal_in_0_6;
      end else if (10'h1f5 == _T_31[9:0]) begin
        image_0_501 <= io_pixelVal_in_0_5;
      end else if (10'h1f5 == _T_28[9:0]) begin
        image_0_501 <= io_pixelVal_in_0_4;
      end else if (10'h1f5 == _T_25[9:0]) begin
        image_0_501 <= io_pixelVal_in_0_3;
      end else if (10'h1f5 == _T_22[9:0]) begin
        image_0_501 <= io_pixelVal_in_0_2;
      end else if (10'h1f5 == _T_19[9:0]) begin
        image_0_501 <= io_pixelVal_in_0_1;
      end else if (10'h1f5 == _T_15[9:0]) begin
        image_0_501 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_502 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1f6 == _T_37[9:0]) begin
        image_0_502 <= io_pixelVal_in_0_7;
      end else if (10'h1f6 == _T_34[9:0]) begin
        image_0_502 <= io_pixelVal_in_0_6;
      end else if (10'h1f6 == _T_31[9:0]) begin
        image_0_502 <= io_pixelVal_in_0_5;
      end else if (10'h1f6 == _T_28[9:0]) begin
        image_0_502 <= io_pixelVal_in_0_4;
      end else if (10'h1f6 == _T_25[9:0]) begin
        image_0_502 <= io_pixelVal_in_0_3;
      end else if (10'h1f6 == _T_22[9:0]) begin
        image_0_502 <= io_pixelVal_in_0_2;
      end else if (10'h1f6 == _T_19[9:0]) begin
        image_0_502 <= io_pixelVal_in_0_1;
      end else if (10'h1f6 == _T_15[9:0]) begin
        image_0_502 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_503 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1f7 == _T_37[9:0]) begin
        image_0_503 <= io_pixelVal_in_0_7;
      end else if (10'h1f7 == _T_34[9:0]) begin
        image_0_503 <= io_pixelVal_in_0_6;
      end else if (10'h1f7 == _T_31[9:0]) begin
        image_0_503 <= io_pixelVal_in_0_5;
      end else if (10'h1f7 == _T_28[9:0]) begin
        image_0_503 <= io_pixelVal_in_0_4;
      end else if (10'h1f7 == _T_25[9:0]) begin
        image_0_503 <= io_pixelVal_in_0_3;
      end else if (10'h1f7 == _T_22[9:0]) begin
        image_0_503 <= io_pixelVal_in_0_2;
      end else if (10'h1f7 == _T_19[9:0]) begin
        image_0_503 <= io_pixelVal_in_0_1;
      end else if (10'h1f7 == _T_15[9:0]) begin
        image_0_503 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_504 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1f8 == _T_37[9:0]) begin
        image_0_504 <= io_pixelVal_in_0_7;
      end else if (10'h1f8 == _T_34[9:0]) begin
        image_0_504 <= io_pixelVal_in_0_6;
      end else if (10'h1f8 == _T_31[9:0]) begin
        image_0_504 <= io_pixelVal_in_0_5;
      end else if (10'h1f8 == _T_28[9:0]) begin
        image_0_504 <= io_pixelVal_in_0_4;
      end else if (10'h1f8 == _T_25[9:0]) begin
        image_0_504 <= io_pixelVal_in_0_3;
      end else if (10'h1f8 == _T_22[9:0]) begin
        image_0_504 <= io_pixelVal_in_0_2;
      end else if (10'h1f8 == _T_19[9:0]) begin
        image_0_504 <= io_pixelVal_in_0_1;
      end else if (10'h1f8 == _T_15[9:0]) begin
        image_0_504 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_505 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1f9 == _T_37[9:0]) begin
        image_0_505 <= io_pixelVal_in_0_7;
      end else if (10'h1f9 == _T_34[9:0]) begin
        image_0_505 <= io_pixelVal_in_0_6;
      end else if (10'h1f9 == _T_31[9:0]) begin
        image_0_505 <= io_pixelVal_in_0_5;
      end else if (10'h1f9 == _T_28[9:0]) begin
        image_0_505 <= io_pixelVal_in_0_4;
      end else if (10'h1f9 == _T_25[9:0]) begin
        image_0_505 <= io_pixelVal_in_0_3;
      end else if (10'h1f9 == _T_22[9:0]) begin
        image_0_505 <= io_pixelVal_in_0_2;
      end else if (10'h1f9 == _T_19[9:0]) begin
        image_0_505 <= io_pixelVal_in_0_1;
      end else if (10'h1f9 == _T_15[9:0]) begin
        image_0_505 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_506 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1fa == _T_37[9:0]) begin
        image_0_506 <= io_pixelVal_in_0_7;
      end else if (10'h1fa == _T_34[9:0]) begin
        image_0_506 <= io_pixelVal_in_0_6;
      end else if (10'h1fa == _T_31[9:0]) begin
        image_0_506 <= io_pixelVal_in_0_5;
      end else if (10'h1fa == _T_28[9:0]) begin
        image_0_506 <= io_pixelVal_in_0_4;
      end else if (10'h1fa == _T_25[9:0]) begin
        image_0_506 <= io_pixelVal_in_0_3;
      end else if (10'h1fa == _T_22[9:0]) begin
        image_0_506 <= io_pixelVal_in_0_2;
      end else if (10'h1fa == _T_19[9:0]) begin
        image_0_506 <= io_pixelVal_in_0_1;
      end else if (10'h1fa == _T_15[9:0]) begin
        image_0_506 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_507 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1fb == _T_37[9:0]) begin
        image_0_507 <= io_pixelVal_in_0_7;
      end else if (10'h1fb == _T_34[9:0]) begin
        image_0_507 <= io_pixelVal_in_0_6;
      end else if (10'h1fb == _T_31[9:0]) begin
        image_0_507 <= io_pixelVal_in_0_5;
      end else if (10'h1fb == _T_28[9:0]) begin
        image_0_507 <= io_pixelVal_in_0_4;
      end else if (10'h1fb == _T_25[9:0]) begin
        image_0_507 <= io_pixelVal_in_0_3;
      end else if (10'h1fb == _T_22[9:0]) begin
        image_0_507 <= io_pixelVal_in_0_2;
      end else if (10'h1fb == _T_19[9:0]) begin
        image_0_507 <= io_pixelVal_in_0_1;
      end else if (10'h1fb == _T_15[9:0]) begin
        image_0_507 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_508 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1fc == _T_37[9:0]) begin
        image_0_508 <= io_pixelVal_in_0_7;
      end else if (10'h1fc == _T_34[9:0]) begin
        image_0_508 <= io_pixelVal_in_0_6;
      end else if (10'h1fc == _T_31[9:0]) begin
        image_0_508 <= io_pixelVal_in_0_5;
      end else if (10'h1fc == _T_28[9:0]) begin
        image_0_508 <= io_pixelVal_in_0_4;
      end else if (10'h1fc == _T_25[9:0]) begin
        image_0_508 <= io_pixelVal_in_0_3;
      end else if (10'h1fc == _T_22[9:0]) begin
        image_0_508 <= io_pixelVal_in_0_2;
      end else if (10'h1fc == _T_19[9:0]) begin
        image_0_508 <= io_pixelVal_in_0_1;
      end else if (10'h1fc == _T_15[9:0]) begin
        image_0_508 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_509 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1fd == _T_37[9:0]) begin
        image_0_509 <= io_pixelVal_in_0_7;
      end else if (10'h1fd == _T_34[9:0]) begin
        image_0_509 <= io_pixelVal_in_0_6;
      end else if (10'h1fd == _T_31[9:0]) begin
        image_0_509 <= io_pixelVal_in_0_5;
      end else if (10'h1fd == _T_28[9:0]) begin
        image_0_509 <= io_pixelVal_in_0_4;
      end else if (10'h1fd == _T_25[9:0]) begin
        image_0_509 <= io_pixelVal_in_0_3;
      end else if (10'h1fd == _T_22[9:0]) begin
        image_0_509 <= io_pixelVal_in_0_2;
      end else if (10'h1fd == _T_19[9:0]) begin
        image_0_509 <= io_pixelVal_in_0_1;
      end else if (10'h1fd == _T_15[9:0]) begin
        image_0_509 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_510 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1fe == _T_37[9:0]) begin
        image_0_510 <= io_pixelVal_in_0_7;
      end else if (10'h1fe == _T_34[9:0]) begin
        image_0_510 <= io_pixelVal_in_0_6;
      end else if (10'h1fe == _T_31[9:0]) begin
        image_0_510 <= io_pixelVal_in_0_5;
      end else if (10'h1fe == _T_28[9:0]) begin
        image_0_510 <= io_pixelVal_in_0_4;
      end else if (10'h1fe == _T_25[9:0]) begin
        image_0_510 <= io_pixelVal_in_0_3;
      end else if (10'h1fe == _T_22[9:0]) begin
        image_0_510 <= io_pixelVal_in_0_2;
      end else if (10'h1fe == _T_19[9:0]) begin
        image_0_510 <= io_pixelVal_in_0_1;
      end else if (10'h1fe == _T_15[9:0]) begin
        image_0_510 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_511 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1ff == _T_37[9:0]) begin
        image_0_511 <= io_pixelVal_in_0_7;
      end else if (10'h1ff == _T_34[9:0]) begin
        image_0_511 <= io_pixelVal_in_0_6;
      end else if (10'h1ff == _T_31[9:0]) begin
        image_0_511 <= io_pixelVal_in_0_5;
      end else if (10'h1ff == _T_28[9:0]) begin
        image_0_511 <= io_pixelVal_in_0_4;
      end else if (10'h1ff == _T_25[9:0]) begin
        image_0_511 <= io_pixelVal_in_0_3;
      end else if (10'h1ff == _T_22[9:0]) begin
        image_0_511 <= io_pixelVal_in_0_2;
      end else if (10'h1ff == _T_19[9:0]) begin
        image_0_511 <= io_pixelVal_in_0_1;
      end else if (10'h1ff == _T_15[9:0]) begin
        image_0_511 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_512 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h200 == _T_37[9:0]) begin
        image_0_512 <= io_pixelVal_in_0_7;
      end else if (10'h200 == _T_34[9:0]) begin
        image_0_512 <= io_pixelVal_in_0_6;
      end else if (10'h200 == _T_31[9:0]) begin
        image_0_512 <= io_pixelVal_in_0_5;
      end else if (10'h200 == _T_28[9:0]) begin
        image_0_512 <= io_pixelVal_in_0_4;
      end else if (10'h200 == _T_25[9:0]) begin
        image_0_512 <= io_pixelVal_in_0_3;
      end else if (10'h200 == _T_22[9:0]) begin
        image_0_512 <= io_pixelVal_in_0_2;
      end else if (10'h200 == _T_19[9:0]) begin
        image_0_512 <= io_pixelVal_in_0_1;
      end else if (10'h200 == _T_15[9:0]) begin
        image_0_512 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_513 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h201 == _T_37[9:0]) begin
        image_0_513 <= io_pixelVal_in_0_7;
      end else if (10'h201 == _T_34[9:0]) begin
        image_0_513 <= io_pixelVal_in_0_6;
      end else if (10'h201 == _T_31[9:0]) begin
        image_0_513 <= io_pixelVal_in_0_5;
      end else if (10'h201 == _T_28[9:0]) begin
        image_0_513 <= io_pixelVal_in_0_4;
      end else if (10'h201 == _T_25[9:0]) begin
        image_0_513 <= io_pixelVal_in_0_3;
      end else if (10'h201 == _T_22[9:0]) begin
        image_0_513 <= io_pixelVal_in_0_2;
      end else if (10'h201 == _T_19[9:0]) begin
        image_0_513 <= io_pixelVal_in_0_1;
      end else if (10'h201 == _T_15[9:0]) begin
        image_0_513 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_514 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h202 == _T_37[9:0]) begin
        image_0_514 <= io_pixelVal_in_0_7;
      end else if (10'h202 == _T_34[9:0]) begin
        image_0_514 <= io_pixelVal_in_0_6;
      end else if (10'h202 == _T_31[9:0]) begin
        image_0_514 <= io_pixelVal_in_0_5;
      end else if (10'h202 == _T_28[9:0]) begin
        image_0_514 <= io_pixelVal_in_0_4;
      end else if (10'h202 == _T_25[9:0]) begin
        image_0_514 <= io_pixelVal_in_0_3;
      end else if (10'h202 == _T_22[9:0]) begin
        image_0_514 <= io_pixelVal_in_0_2;
      end else if (10'h202 == _T_19[9:0]) begin
        image_0_514 <= io_pixelVal_in_0_1;
      end else if (10'h202 == _T_15[9:0]) begin
        image_0_514 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_515 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h203 == _T_37[9:0]) begin
        image_0_515 <= io_pixelVal_in_0_7;
      end else if (10'h203 == _T_34[9:0]) begin
        image_0_515 <= io_pixelVal_in_0_6;
      end else if (10'h203 == _T_31[9:0]) begin
        image_0_515 <= io_pixelVal_in_0_5;
      end else if (10'h203 == _T_28[9:0]) begin
        image_0_515 <= io_pixelVal_in_0_4;
      end else if (10'h203 == _T_25[9:0]) begin
        image_0_515 <= io_pixelVal_in_0_3;
      end else if (10'h203 == _T_22[9:0]) begin
        image_0_515 <= io_pixelVal_in_0_2;
      end else if (10'h203 == _T_19[9:0]) begin
        image_0_515 <= io_pixelVal_in_0_1;
      end else if (10'h203 == _T_15[9:0]) begin
        image_0_515 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_516 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h204 == _T_37[9:0]) begin
        image_0_516 <= io_pixelVal_in_0_7;
      end else if (10'h204 == _T_34[9:0]) begin
        image_0_516 <= io_pixelVal_in_0_6;
      end else if (10'h204 == _T_31[9:0]) begin
        image_0_516 <= io_pixelVal_in_0_5;
      end else if (10'h204 == _T_28[9:0]) begin
        image_0_516 <= io_pixelVal_in_0_4;
      end else if (10'h204 == _T_25[9:0]) begin
        image_0_516 <= io_pixelVal_in_0_3;
      end else if (10'h204 == _T_22[9:0]) begin
        image_0_516 <= io_pixelVal_in_0_2;
      end else if (10'h204 == _T_19[9:0]) begin
        image_0_516 <= io_pixelVal_in_0_1;
      end else if (10'h204 == _T_15[9:0]) begin
        image_0_516 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_517 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h205 == _T_37[9:0]) begin
        image_0_517 <= io_pixelVal_in_0_7;
      end else if (10'h205 == _T_34[9:0]) begin
        image_0_517 <= io_pixelVal_in_0_6;
      end else if (10'h205 == _T_31[9:0]) begin
        image_0_517 <= io_pixelVal_in_0_5;
      end else if (10'h205 == _T_28[9:0]) begin
        image_0_517 <= io_pixelVal_in_0_4;
      end else if (10'h205 == _T_25[9:0]) begin
        image_0_517 <= io_pixelVal_in_0_3;
      end else if (10'h205 == _T_22[9:0]) begin
        image_0_517 <= io_pixelVal_in_0_2;
      end else if (10'h205 == _T_19[9:0]) begin
        image_0_517 <= io_pixelVal_in_0_1;
      end else if (10'h205 == _T_15[9:0]) begin
        image_0_517 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_518 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h206 == _T_37[9:0]) begin
        image_0_518 <= io_pixelVal_in_0_7;
      end else if (10'h206 == _T_34[9:0]) begin
        image_0_518 <= io_pixelVal_in_0_6;
      end else if (10'h206 == _T_31[9:0]) begin
        image_0_518 <= io_pixelVal_in_0_5;
      end else if (10'h206 == _T_28[9:0]) begin
        image_0_518 <= io_pixelVal_in_0_4;
      end else if (10'h206 == _T_25[9:0]) begin
        image_0_518 <= io_pixelVal_in_0_3;
      end else if (10'h206 == _T_22[9:0]) begin
        image_0_518 <= io_pixelVal_in_0_2;
      end else if (10'h206 == _T_19[9:0]) begin
        image_0_518 <= io_pixelVal_in_0_1;
      end else if (10'h206 == _T_15[9:0]) begin
        image_0_518 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_519 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h207 == _T_37[9:0]) begin
        image_0_519 <= io_pixelVal_in_0_7;
      end else if (10'h207 == _T_34[9:0]) begin
        image_0_519 <= io_pixelVal_in_0_6;
      end else if (10'h207 == _T_31[9:0]) begin
        image_0_519 <= io_pixelVal_in_0_5;
      end else if (10'h207 == _T_28[9:0]) begin
        image_0_519 <= io_pixelVal_in_0_4;
      end else if (10'h207 == _T_25[9:0]) begin
        image_0_519 <= io_pixelVal_in_0_3;
      end else if (10'h207 == _T_22[9:0]) begin
        image_0_519 <= io_pixelVal_in_0_2;
      end else if (10'h207 == _T_19[9:0]) begin
        image_0_519 <= io_pixelVal_in_0_1;
      end else if (10'h207 == _T_15[9:0]) begin
        image_0_519 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_520 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h208 == _T_37[9:0]) begin
        image_0_520 <= io_pixelVal_in_0_7;
      end else if (10'h208 == _T_34[9:0]) begin
        image_0_520 <= io_pixelVal_in_0_6;
      end else if (10'h208 == _T_31[9:0]) begin
        image_0_520 <= io_pixelVal_in_0_5;
      end else if (10'h208 == _T_28[9:0]) begin
        image_0_520 <= io_pixelVal_in_0_4;
      end else if (10'h208 == _T_25[9:0]) begin
        image_0_520 <= io_pixelVal_in_0_3;
      end else if (10'h208 == _T_22[9:0]) begin
        image_0_520 <= io_pixelVal_in_0_2;
      end else if (10'h208 == _T_19[9:0]) begin
        image_0_520 <= io_pixelVal_in_0_1;
      end else if (10'h208 == _T_15[9:0]) begin
        image_0_520 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_521 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h209 == _T_37[9:0]) begin
        image_0_521 <= io_pixelVal_in_0_7;
      end else if (10'h209 == _T_34[9:0]) begin
        image_0_521 <= io_pixelVal_in_0_6;
      end else if (10'h209 == _T_31[9:0]) begin
        image_0_521 <= io_pixelVal_in_0_5;
      end else if (10'h209 == _T_28[9:0]) begin
        image_0_521 <= io_pixelVal_in_0_4;
      end else if (10'h209 == _T_25[9:0]) begin
        image_0_521 <= io_pixelVal_in_0_3;
      end else if (10'h209 == _T_22[9:0]) begin
        image_0_521 <= io_pixelVal_in_0_2;
      end else if (10'h209 == _T_19[9:0]) begin
        image_0_521 <= io_pixelVal_in_0_1;
      end else if (10'h209 == _T_15[9:0]) begin
        image_0_521 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_522 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h20a == _T_37[9:0]) begin
        image_0_522 <= io_pixelVal_in_0_7;
      end else if (10'h20a == _T_34[9:0]) begin
        image_0_522 <= io_pixelVal_in_0_6;
      end else if (10'h20a == _T_31[9:0]) begin
        image_0_522 <= io_pixelVal_in_0_5;
      end else if (10'h20a == _T_28[9:0]) begin
        image_0_522 <= io_pixelVal_in_0_4;
      end else if (10'h20a == _T_25[9:0]) begin
        image_0_522 <= io_pixelVal_in_0_3;
      end else if (10'h20a == _T_22[9:0]) begin
        image_0_522 <= io_pixelVal_in_0_2;
      end else if (10'h20a == _T_19[9:0]) begin
        image_0_522 <= io_pixelVal_in_0_1;
      end else if (10'h20a == _T_15[9:0]) begin
        image_0_522 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_523 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h20b == _T_37[9:0]) begin
        image_0_523 <= io_pixelVal_in_0_7;
      end else if (10'h20b == _T_34[9:0]) begin
        image_0_523 <= io_pixelVal_in_0_6;
      end else if (10'h20b == _T_31[9:0]) begin
        image_0_523 <= io_pixelVal_in_0_5;
      end else if (10'h20b == _T_28[9:0]) begin
        image_0_523 <= io_pixelVal_in_0_4;
      end else if (10'h20b == _T_25[9:0]) begin
        image_0_523 <= io_pixelVal_in_0_3;
      end else if (10'h20b == _T_22[9:0]) begin
        image_0_523 <= io_pixelVal_in_0_2;
      end else if (10'h20b == _T_19[9:0]) begin
        image_0_523 <= io_pixelVal_in_0_1;
      end else if (10'h20b == _T_15[9:0]) begin
        image_0_523 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_524 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h20c == _T_37[9:0]) begin
        image_0_524 <= io_pixelVal_in_0_7;
      end else if (10'h20c == _T_34[9:0]) begin
        image_0_524 <= io_pixelVal_in_0_6;
      end else if (10'h20c == _T_31[9:0]) begin
        image_0_524 <= io_pixelVal_in_0_5;
      end else if (10'h20c == _T_28[9:0]) begin
        image_0_524 <= io_pixelVal_in_0_4;
      end else if (10'h20c == _T_25[9:0]) begin
        image_0_524 <= io_pixelVal_in_0_3;
      end else if (10'h20c == _T_22[9:0]) begin
        image_0_524 <= io_pixelVal_in_0_2;
      end else if (10'h20c == _T_19[9:0]) begin
        image_0_524 <= io_pixelVal_in_0_1;
      end else if (10'h20c == _T_15[9:0]) begin
        image_0_524 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_525 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h20d == _T_37[9:0]) begin
        image_0_525 <= io_pixelVal_in_0_7;
      end else if (10'h20d == _T_34[9:0]) begin
        image_0_525 <= io_pixelVal_in_0_6;
      end else if (10'h20d == _T_31[9:0]) begin
        image_0_525 <= io_pixelVal_in_0_5;
      end else if (10'h20d == _T_28[9:0]) begin
        image_0_525 <= io_pixelVal_in_0_4;
      end else if (10'h20d == _T_25[9:0]) begin
        image_0_525 <= io_pixelVal_in_0_3;
      end else if (10'h20d == _T_22[9:0]) begin
        image_0_525 <= io_pixelVal_in_0_2;
      end else if (10'h20d == _T_19[9:0]) begin
        image_0_525 <= io_pixelVal_in_0_1;
      end else if (10'h20d == _T_15[9:0]) begin
        image_0_525 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_526 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h20e == _T_37[9:0]) begin
        image_0_526 <= io_pixelVal_in_0_7;
      end else if (10'h20e == _T_34[9:0]) begin
        image_0_526 <= io_pixelVal_in_0_6;
      end else if (10'h20e == _T_31[9:0]) begin
        image_0_526 <= io_pixelVal_in_0_5;
      end else if (10'h20e == _T_28[9:0]) begin
        image_0_526 <= io_pixelVal_in_0_4;
      end else if (10'h20e == _T_25[9:0]) begin
        image_0_526 <= io_pixelVal_in_0_3;
      end else if (10'h20e == _T_22[9:0]) begin
        image_0_526 <= io_pixelVal_in_0_2;
      end else if (10'h20e == _T_19[9:0]) begin
        image_0_526 <= io_pixelVal_in_0_1;
      end else if (10'h20e == _T_15[9:0]) begin
        image_0_526 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_527 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h20f == _T_37[9:0]) begin
        image_0_527 <= io_pixelVal_in_0_7;
      end else if (10'h20f == _T_34[9:0]) begin
        image_0_527 <= io_pixelVal_in_0_6;
      end else if (10'h20f == _T_31[9:0]) begin
        image_0_527 <= io_pixelVal_in_0_5;
      end else if (10'h20f == _T_28[9:0]) begin
        image_0_527 <= io_pixelVal_in_0_4;
      end else if (10'h20f == _T_25[9:0]) begin
        image_0_527 <= io_pixelVal_in_0_3;
      end else if (10'h20f == _T_22[9:0]) begin
        image_0_527 <= io_pixelVal_in_0_2;
      end else if (10'h20f == _T_19[9:0]) begin
        image_0_527 <= io_pixelVal_in_0_1;
      end else if (10'h20f == _T_15[9:0]) begin
        image_0_527 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_528 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h210 == _T_37[9:0]) begin
        image_0_528 <= io_pixelVal_in_0_7;
      end else if (10'h210 == _T_34[9:0]) begin
        image_0_528 <= io_pixelVal_in_0_6;
      end else if (10'h210 == _T_31[9:0]) begin
        image_0_528 <= io_pixelVal_in_0_5;
      end else if (10'h210 == _T_28[9:0]) begin
        image_0_528 <= io_pixelVal_in_0_4;
      end else if (10'h210 == _T_25[9:0]) begin
        image_0_528 <= io_pixelVal_in_0_3;
      end else if (10'h210 == _T_22[9:0]) begin
        image_0_528 <= io_pixelVal_in_0_2;
      end else if (10'h210 == _T_19[9:0]) begin
        image_0_528 <= io_pixelVal_in_0_1;
      end else if (10'h210 == _T_15[9:0]) begin
        image_0_528 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_529 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h211 == _T_37[9:0]) begin
        image_0_529 <= io_pixelVal_in_0_7;
      end else if (10'h211 == _T_34[9:0]) begin
        image_0_529 <= io_pixelVal_in_0_6;
      end else if (10'h211 == _T_31[9:0]) begin
        image_0_529 <= io_pixelVal_in_0_5;
      end else if (10'h211 == _T_28[9:0]) begin
        image_0_529 <= io_pixelVal_in_0_4;
      end else if (10'h211 == _T_25[9:0]) begin
        image_0_529 <= io_pixelVal_in_0_3;
      end else if (10'h211 == _T_22[9:0]) begin
        image_0_529 <= io_pixelVal_in_0_2;
      end else if (10'h211 == _T_19[9:0]) begin
        image_0_529 <= io_pixelVal_in_0_1;
      end else if (10'h211 == _T_15[9:0]) begin
        image_0_529 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_530 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h212 == _T_37[9:0]) begin
        image_0_530 <= io_pixelVal_in_0_7;
      end else if (10'h212 == _T_34[9:0]) begin
        image_0_530 <= io_pixelVal_in_0_6;
      end else if (10'h212 == _T_31[9:0]) begin
        image_0_530 <= io_pixelVal_in_0_5;
      end else if (10'h212 == _T_28[9:0]) begin
        image_0_530 <= io_pixelVal_in_0_4;
      end else if (10'h212 == _T_25[9:0]) begin
        image_0_530 <= io_pixelVal_in_0_3;
      end else if (10'h212 == _T_22[9:0]) begin
        image_0_530 <= io_pixelVal_in_0_2;
      end else if (10'h212 == _T_19[9:0]) begin
        image_0_530 <= io_pixelVal_in_0_1;
      end else if (10'h212 == _T_15[9:0]) begin
        image_0_530 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_531 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h213 == _T_37[9:0]) begin
        image_0_531 <= io_pixelVal_in_0_7;
      end else if (10'h213 == _T_34[9:0]) begin
        image_0_531 <= io_pixelVal_in_0_6;
      end else if (10'h213 == _T_31[9:0]) begin
        image_0_531 <= io_pixelVal_in_0_5;
      end else if (10'h213 == _T_28[9:0]) begin
        image_0_531 <= io_pixelVal_in_0_4;
      end else if (10'h213 == _T_25[9:0]) begin
        image_0_531 <= io_pixelVal_in_0_3;
      end else if (10'h213 == _T_22[9:0]) begin
        image_0_531 <= io_pixelVal_in_0_2;
      end else if (10'h213 == _T_19[9:0]) begin
        image_0_531 <= io_pixelVal_in_0_1;
      end else if (10'h213 == _T_15[9:0]) begin
        image_0_531 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_532 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h214 == _T_37[9:0]) begin
        image_0_532 <= io_pixelVal_in_0_7;
      end else if (10'h214 == _T_34[9:0]) begin
        image_0_532 <= io_pixelVal_in_0_6;
      end else if (10'h214 == _T_31[9:0]) begin
        image_0_532 <= io_pixelVal_in_0_5;
      end else if (10'h214 == _T_28[9:0]) begin
        image_0_532 <= io_pixelVal_in_0_4;
      end else if (10'h214 == _T_25[9:0]) begin
        image_0_532 <= io_pixelVal_in_0_3;
      end else if (10'h214 == _T_22[9:0]) begin
        image_0_532 <= io_pixelVal_in_0_2;
      end else if (10'h214 == _T_19[9:0]) begin
        image_0_532 <= io_pixelVal_in_0_1;
      end else if (10'h214 == _T_15[9:0]) begin
        image_0_532 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_533 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h215 == _T_37[9:0]) begin
        image_0_533 <= io_pixelVal_in_0_7;
      end else if (10'h215 == _T_34[9:0]) begin
        image_0_533 <= io_pixelVal_in_0_6;
      end else if (10'h215 == _T_31[9:0]) begin
        image_0_533 <= io_pixelVal_in_0_5;
      end else if (10'h215 == _T_28[9:0]) begin
        image_0_533 <= io_pixelVal_in_0_4;
      end else if (10'h215 == _T_25[9:0]) begin
        image_0_533 <= io_pixelVal_in_0_3;
      end else if (10'h215 == _T_22[9:0]) begin
        image_0_533 <= io_pixelVal_in_0_2;
      end else if (10'h215 == _T_19[9:0]) begin
        image_0_533 <= io_pixelVal_in_0_1;
      end else if (10'h215 == _T_15[9:0]) begin
        image_0_533 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_534 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h216 == _T_37[9:0]) begin
        image_0_534 <= io_pixelVal_in_0_7;
      end else if (10'h216 == _T_34[9:0]) begin
        image_0_534 <= io_pixelVal_in_0_6;
      end else if (10'h216 == _T_31[9:0]) begin
        image_0_534 <= io_pixelVal_in_0_5;
      end else if (10'h216 == _T_28[9:0]) begin
        image_0_534 <= io_pixelVal_in_0_4;
      end else if (10'h216 == _T_25[9:0]) begin
        image_0_534 <= io_pixelVal_in_0_3;
      end else if (10'h216 == _T_22[9:0]) begin
        image_0_534 <= io_pixelVal_in_0_2;
      end else if (10'h216 == _T_19[9:0]) begin
        image_0_534 <= io_pixelVal_in_0_1;
      end else if (10'h216 == _T_15[9:0]) begin
        image_0_534 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_535 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h217 == _T_37[9:0]) begin
        image_0_535 <= io_pixelVal_in_0_7;
      end else if (10'h217 == _T_34[9:0]) begin
        image_0_535 <= io_pixelVal_in_0_6;
      end else if (10'h217 == _T_31[9:0]) begin
        image_0_535 <= io_pixelVal_in_0_5;
      end else if (10'h217 == _T_28[9:0]) begin
        image_0_535 <= io_pixelVal_in_0_4;
      end else if (10'h217 == _T_25[9:0]) begin
        image_0_535 <= io_pixelVal_in_0_3;
      end else if (10'h217 == _T_22[9:0]) begin
        image_0_535 <= io_pixelVal_in_0_2;
      end else if (10'h217 == _T_19[9:0]) begin
        image_0_535 <= io_pixelVal_in_0_1;
      end else if (10'h217 == _T_15[9:0]) begin
        image_0_535 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_536 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h218 == _T_37[9:0]) begin
        image_0_536 <= io_pixelVal_in_0_7;
      end else if (10'h218 == _T_34[9:0]) begin
        image_0_536 <= io_pixelVal_in_0_6;
      end else if (10'h218 == _T_31[9:0]) begin
        image_0_536 <= io_pixelVal_in_0_5;
      end else if (10'h218 == _T_28[9:0]) begin
        image_0_536 <= io_pixelVal_in_0_4;
      end else if (10'h218 == _T_25[9:0]) begin
        image_0_536 <= io_pixelVal_in_0_3;
      end else if (10'h218 == _T_22[9:0]) begin
        image_0_536 <= io_pixelVal_in_0_2;
      end else if (10'h218 == _T_19[9:0]) begin
        image_0_536 <= io_pixelVal_in_0_1;
      end else if (10'h218 == _T_15[9:0]) begin
        image_0_536 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_537 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h219 == _T_37[9:0]) begin
        image_0_537 <= io_pixelVal_in_0_7;
      end else if (10'h219 == _T_34[9:0]) begin
        image_0_537 <= io_pixelVal_in_0_6;
      end else if (10'h219 == _T_31[9:0]) begin
        image_0_537 <= io_pixelVal_in_0_5;
      end else if (10'h219 == _T_28[9:0]) begin
        image_0_537 <= io_pixelVal_in_0_4;
      end else if (10'h219 == _T_25[9:0]) begin
        image_0_537 <= io_pixelVal_in_0_3;
      end else if (10'h219 == _T_22[9:0]) begin
        image_0_537 <= io_pixelVal_in_0_2;
      end else if (10'h219 == _T_19[9:0]) begin
        image_0_537 <= io_pixelVal_in_0_1;
      end else if (10'h219 == _T_15[9:0]) begin
        image_0_537 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_538 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h21a == _T_37[9:0]) begin
        image_0_538 <= io_pixelVal_in_0_7;
      end else if (10'h21a == _T_34[9:0]) begin
        image_0_538 <= io_pixelVal_in_0_6;
      end else if (10'h21a == _T_31[9:0]) begin
        image_0_538 <= io_pixelVal_in_0_5;
      end else if (10'h21a == _T_28[9:0]) begin
        image_0_538 <= io_pixelVal_in_0_4;
      end else if (10'h21a == _T_25[9:0]) begin
        image_0_538 <= io_pixelVal_in_0_3;
      end else if (10'h21a == _T_22[9:0]) begin
        image_0_538 <= io_pixelVal_in_0_2;
      end else if (10'h21a == _T_19[9:0]) begin
        image_0_538 <= io_pixelVal_in_0_1;
      end else if (10'h21a == _T_15[9:0]) begin
        image_0_538 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_539 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h21b == _T_37[9:0]) begin
        image_0_539 <= io_pixelVal_in_0_7;
      end else if (10'h21b == _T_34[9:0]) begin
        image_0_539 <= io_pixelVal_in_0_6;
      end else if (10'h21b == _T_31[9:0]) begin
        image_0_539 <= io_pixelVal_in_0_5;
      end else if (10'h21b == _T_28[9:0]) begin
        image_0_539 <= io_pixelVal_in_0_4;
      end else if (10'h21b == _T_25[9:0]) begin
        image_0_539 <= io_pixelVal_in_0_3;
      end else if (10'h21b == _T_22[9:0]) begin
        image_0_539 <= io_pixelVal_in_0_2;
      end else if (10'h21b == _T_19[9:0]) begin
        image_0_539 <= io_pixelVal_in_0_1;
      end else if (10'h21b == _T_15[9:0]) begin
        image_0_539 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_540 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h21c == _T_37[9:0]) begin
        image_0_540 <= io_pixelVal_in_0_7;
      end else if (10'h21c == _T_34[9:0]) begin
        image_0_540 <= io_pixelVal_in_0_6;
      end else if (10'h21c == _T_31[9:0]) begin
        image_0_540 <= io_pixelVal_in_0_5;
      end else if (10'h21c == _T_28[9:0]) begin
        image_0_540 <= io_pixelVal_in_0_4;
      end else if (10'h21c == _T_25[9:0]) begin
        image_0_540 <= io_pixelVal_in_0_3;
      end else if (10'h21c == _T_22[9:0]) begin
        image_0_540 <= io_pixelVal_in_0_2;
      end else if (10'h21c == _T_19[9:0]) begin
        image_0_540 <= io_pixelVal_in_0_1;
      end else if (10'h21c == _T_15[9:0]) begin
        image_0_540 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_541 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h21d == _T_37[9:0]) begin
        image_0_541 <= io_pixelVal_in_0_7;
      end else if (10'h21d == _T_34[9:0]) begin
        image_0_541 <= io_pixelVal_in_0_6;
      end else if (10'h21d == _T_31[9:0]) begin
        image_0_541 <= io_pixelVal_in_0_5;
      end else if (10'h21d == _T_28[9:0]) begin
        image_0_541 <= io_pixelVal_in_0_4;
      end else if (10'h21d == _T_25[9:0]) begin
        image_0_541 <= io_pixelVal_in_0_3;
      end else if (10'h21d == _T_22[9:0]) begin
        image_0_541 <= io_pixelVal_in_0_2;
      end else if (10'h21d == _T_19[9:0]) begin
        image_0_541 <= io_pixelVal_in_0_1;
      end else if (10'h21d == _T_15[9:0]) begin
        image_0_541 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_542 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h21e == _T_37[9:0]) begin
        image_0_542 <= io_pixelVal_in_0_7;
      end else if (10'h21e == _T_34[9:0]) begin
        image_0_542 <= io_pixelVal_in_0_6;
      end else if (10'h21e == _T_31[9:0]) begin
        image_0_542 <= io_pixelVal_in_0_5;
      end else if (10'h21e == _T_28[9:0]) begin
        image_0_542 <= io_pixelVal_in_0_4;
      end else if (10'h21e == _T_25[9:0]) begin
        image_0_542 <= io_pixelVal_in_0_3;
      end else if (10'h21e == _T_22[9:0]) begin
        image_0_542 <= io_pixelVal_in_0_2;
      end else if (10'h21e == _T_19[9:0]) begin
        image_0_542 <= io_pixelVal_in_0_1;
      end else if (10'h21e == _T_15[9:0]) begin
        image_0_542 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_543 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h21f == _T_37[9:0]) begin
        image_0_543 <= io_pixelVal_in_0_7;
      end else if (10'h21f == _T_34[9:0]) begin
        image_0_543 <= io_pixelVal_in_0_6;
      end else if (10'h21f == _T_31[9:0]) begin
        image_0_543 <= io_pixelVal_in_0_5;
      end else if (10'h21f == _T_28[9:0]) begin
        image_0_543 <= io_pixelVal_in_0_4;
      end else if (10'h21f == _T_25[9:0]) begin
        image_0_543 <= io_pixelVal_in_0_3;
      end else if (10'h21f == _T_22[9:0]) begin
        image_0_543 <= io_pixelVal_in_0_2;
      end else if (10'h21f == _T_19[9:0]) begin
        image_0_543 <= io_pixelVal_in_0_1;
      end else if (10'h21f == _T_15[9:0]) begin
        image_0_543 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_544 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h220 == _T_37[9:0]) begin
        image_0_544 <= io_pixelVal_in_0_7;
      end else if (10'h220 == _T_34[9:0]) begin
        image_0_544 <= io_pixelVal_in_0_6;
      end else if (10'h220 == _T_31[9:0]) begin
        image_0_544 <= io_pixelVal_in_0_5;
      end else if (10'h220 == _T_28[9:0]) begin
        image_0_544 <= io_pixelVal_in_0_4;
      end else if (10'h220 == _T_25[9:0]) begin
        image_0_544 <= io_pixelVal_in_0_3;
      end else if (10'h220 == _T_22[9:0]) begin
        image_0_544 <= io_pixelVal_in_0_2;
      end else if (10'h220 == _T_19[9:0]) begin
        image_0_544 <= io_pixelVal_in_0_1;
      end else if (10'h220 == _T_15[9:0]) begin
        image_0_544 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_545 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h221 == _T_37[9:0]) begin
        image_0_545 <= io_pixelVal_in_0_7;
      end else if (10'h221 == _T_34[9:0]) begin
        image_0_545 <= io_pixelVal_in_0_6;
      end else if (10'h221 == _T_31[9:0]) begin
        image_0_545 <= io_pixelVal_in_0_5;
      end else if (10'h221 == _T_28[9:0]) begin
        image_0_545 <= io_pixelVal_in_0_4;
      end else if (10'h221 == _T_25[9:0]) begin
        image_0_545 <= io_pixelVal_in_0_3;
      end else if (10'h221 == _T_22[9:0]) begin
        image_0_545 <= io_pixelVal_in_0_2;
      end else if (10'h221 == _T_19[9:0]) begin
        image_0_545 <= io_pixelVal_in_0_1;
      end else if (10'h221 == _T_15[9:0]) begin
        image_0_545 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_546 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h222 == _T_37[9:0]) begin
        image_0_546 <= io_pixelVal_in_0_7;
      end else if (10'h222 == _T_34[9:0]) begin
        image_0_546 <= io_pixelVal_in_0_6;
      end else if (10'h222 == _T_31[9:0]) begin
        image_0_546 <= io_pixelVal_in_0_5;
      end else if (10'h222 == _T_28[9:0]) begin
        image_0_546 <= io_pixelVal_in_0_4;
      end else if (10'h222 == _T_25[9:0]) begin
        image_0_546 <= io_pixelVal_in_0_3;
      end else if (10'h222 == _T_22[9:0]) begin
        image_0_546 <= io_pixelVal_in_0_2;
      end else if (10'h222 == _T_19[9:0]) begin
        image_0_546 <= io_pixelVal_in_0_1;
      end else if (10'h222 == _T_15[9:0]) begin
        image_0_546 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_547 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h223 == _T_37[9:0]) begin
        image_0_547 <= io_pixelVal_in_0_7;
      end else if (10'h223 == _T_34[9:0]) begin
        image_0_547 <= io_pixelVal_in_0_6;
      end else if (10'h223 == _T_31[9:0]) begin
        image_0_547 <= io_pixelVal_in_0_5;
      end else if (10'h223 == _T_28[9:0]) begin
        image_0_547 <= io_pixelVal_in_0_4;
      end else if (10'h223 == _T_25[9:0]) begin
        image_0_547 <= io_pixelVal_in_0_3;
      end else if (10'h223 == _T_22[9:0]) begin
        image_0_547 <= io_pixelVal_in_0_2;
      end else if (10'h223 == _T_19[9:0]) begin
        image_0_547 <= io_pixelVal_in_0_1;
      end else if (10'h223 == _T_15[9:0]) begin
        image_0_547 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_548 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h224 == _T_37[9:0]) begin
        image_0_548 <= io_pixelVal_in_0_7;
      end else if (10'h224 == _T_34[9:0]) begin
        image_0_548 <= io_pixelVal_in_0_6;
      end else if (10'h224 == _T_31[9:0]) begin
        image_0_548 <= io_pixelVal_in_0_5;
      end else if (10'h224 == _T_28[9:0]) begin
        image_0_548 <= io_pixelVal_in_0_4;
      end else if (10'h224 == _T_25[9:0]) begin
        image_0_548 <= io_pixelVal_in_0_3;
      end else if (10'h224 == _T_22[9:0]) begin
        image_0_548 <= io_pixelVal_in_0_2;
      end else if (10'h224 == _T_19[9:0]) begin
        image_0_548 <= io_pixelVal_in_0_1;
      end else if (10'h224 == _T_15[9:0]) begin
        image_0_548 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_549 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h225 == _T_37[9:0]) begin
        image_0_549 <= io_pixelVal_in_0_7;
      end else if (10'h225 == _T_34[9:0]) begin
        image_0_549 <= io_pixelVal_in_0_6;
      end else if (10'h225 == _T_31[9:0]) begin
        image_0_549 <= io_pixelVal_in_0_5;
      end else if (10'h225 == _T_28[9:0]) begin
        image_0_549 <= io_pixelVal_in_0_4;
      end else if (10'h225 == _T_25[9:0]) begin
        image_0_549 <= io_pixelVal_in_0_3;
      end else if (10'h225 == _T_22[9:0]) begin
        image_0_549 <= io_pixelVal_in_0_2;
      end else if (10'h225 == _T_19[9:0]) begin
        image_0_549 <= io_pixelVal_in_0_1;
      end else if (10'h225 == _T_15[9:0]) begin
        image_0_549 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_550 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h226 == _T_37[9:0]) begin
        image_0_550 <= io_pixelVal_in_0_7;
      end else if (10'h226 == _T_34[9:0]) begin
        image_0_550 <= io_pixelVal_in_0_6;
      end else if (10'h226 == _T_31[9:0]) begin
        image_0_550 <= io_pixelVal_in_0_5;
      end else if (10'h226 == _T_28[9:0]) begin
        image_0_550 <= io_pixelVal_in_0_4;
      end else if (10'h226 == _T_25[9:0]) begin
        image_0_550 <= io_pixelVal_in_0_3;
      end else if (10'h226 == _T_22[9:0]) begin
        image_0_550 <= io_pixelVal_in_0_2;
      end else if (10'h226 == _T_19[9:0]) begin
        image_0_550 <= io_pixelVal_in_0_1;
      end else if (10'h226 == _T_15[9:0]) begin
        image_0_550 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_551 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h227 == _T_37[9:0]) begin
        image_0_551 <= io_pixelVal_in_0_7;
      end else if (10'h227 == _T_34[9:0]) begin
        image_0_551 <= io_pixelVal_in_0_6;
      end else if (10'h227 == _T_31[9:0]) begin
        image_0_551 <= io_pixelVal_in_0_5;
      end else if (10'h227 == _T_28[9:0]) begin
        image_0_551 <= io_pixelVal_in_0_4;
      end else if (10'h227 == _T_25[9:0]) begin
        image_0_551 <= io_pixelVal_in_0_3;
      end else if (10'h227 == _T_22[9:0]) begin
        image_0_551 <= io_pixelVal_in_0_2;
      end else if (10'h227 == _T_19[9:0]) begin
        image_0_551 <= io_pixelVal_in_0_1;
      end else if (10'h227 == _T_15[9:0]) begin
        image_0_551 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_552 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h228 == _T_37[9:0]) begin
        image_0_552 <= io_pixelVal_in_0_7;
      end else if (10'h228 == _T_34[9:0]) begin
        image_0_552 <= io_pixelVal_in_0_6;
      end else if (10'h228 == _T_31[9:0]) begin
        image_0_552 <= io_pixelVal_in_0_5;
      end else if (10'h228 == _T_28[9:0]) begin
        image_0_552 <= io_pixelVal_in_0_4;
      end else if (10'h228 == _T_25[9:0]) begin
        image_0_552 <= io_pixelVal_in_0_3;
      end else if (10'h228 == _T_22[9:0]) begin
        image_0_552 <= io_pixelVal_in_0_2;
      end else if (10'h228 == _T_19[9:0]) begin
        image_0_552 <= io_pixelVal_in_0_1;
      end else if (10'h228 == _T_15[9:0]) begin
        image_0_552 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_553 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h229 == _T_37[9:0]) begin
        image_0_553 <= io_pixelVal_in_0_7;
      end else if (10'h229 == _T_34[9:0]) begin
        image_0_553 <= io_pixelVal_in_0_6;
      end else if (10'h229 == _T_31[9:0]) begin
        image_0_553 <= io_pixelVal_in_0_5;
      end else if (10'h229 == _T_28[9:0]) begin
        image_0_553 <= io_pixelVal_in_0_4;
      end else if (10'h229 == _T_25[9:0]) begin
        image_0_553 <= io_pixelVal_in_0_3;
      end else if (10'h229 == _T_22[9:0]) begin
        image_0_553 <= io_pixelVal_in_0_2;
      end else if (10'h229 == _T_19[9:0]) begin
        image_0_553 <= io_pixelVal_in_0_1;
      end else if (10'h229 == _T_15[9:0]) begin
        image_0_553 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_554 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h22a == _T_37[9:0]) begin
        image_0_554 <= io_pixelVal_in_0_7;
      end else if (10'h22a == _T_34[9:0]) begin
        image_0_554 <= io_pixelVal_in_0_6;
      end else if (10'h22a == _T_31[9:0]) begin
        image_0_554 <= io_pixelVal_in_0_5;
      end else if (10'h22a == _T_28[9:0]) begin
        image_0_554 <= io_pixelVal_in_0_4;
      end else if (10'h22a == _T_25[9:0]) begin
        image_0_554 <= io_pixelVal_in_0_3;
      end else if (10'h22a == _T_22[9:0]) begin
        image_0_554 <= io_pixelVal_in_0_2;
      end else if (10'h22a == _T_19[9:0]) begin
        image_0_554 <= io_pixelVal_in_0_1;
      end else if (10'h22a == _T_15[9:0]) begin
        image_0_554 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_555 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h22b == _T_37[9:0]) begin
        image_0_555 <= io_pixelVal_in_0_7;
      end else if (10'h22b == _T_34[9:0]) begin
        image_0_555 <= io_pixelVal_in_0_6;
      end else if (10'h22b == _T_31[9:0]) begin
        image_0_555 <= io_pixelVal_in_0_5;
      end else if (10'h22b == _T_28[9:0]) begin
        image_0_555 <= io_pixelVal_in_0_4;
      end else if (10'h22b == _T_25[9:0]) begin
        image_0_555 <= io_pixelVal_in_0_3;
      end else if (10'h22b == _T_22[9:0]) begin
        image_0_555 <= io_pixelVal_in_0_2;
      end else if (10'h22b == _T_19[9:0]) begin
        image_0_555 <= io_pixelVal_in_0_1;
      end else if (10'h22b == _T_15[9:0]) begin
        image_0_555 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_556 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h22c == _T_37[9:0]) begin
        image_0_556 <= io_pixelVal_in_0_7;
      end else if (10'h22c == _T_34[9:0]) begin
        image_0_556 <= io_pixelVal_in_0_6;
      end else if (10'h22c == _T_31[9:0]) begin
        image_0_556 <= io_pixelVal_in_0_5;
      end else if (10'h22c == _T_28[9:0]) begin
        image_0_556 <= io_pixelVal_in_0_4;
      end else if (10'h22c == _T_25[9:0]) begin
        image_0_556 <= io_pixelVal_in_0_3;
      end else if (10'h22c == _T_22[9:0]) begin
        image_0_556 <= io_pixelVal_in_0_2;
      end else if (10'h22c == _T_19[9:0]) begin
        image_0_556 <= io_pixelVal_in_0_1;
      end else if (10'h22c == _T_15[9:0]) begin
        image_0_556 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_557 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h22d == _T_37[9:0]) begin
        image_0_557 <= io_pixelVal_in_0_7;
      end else if (10'h22d == _T_34[9:0]) begin
        image_0_557 <= io_pixelVal_in_0_6;
      end else if (10'h22d == _T_31[9:0]) begin
        image_0_557 <= io_pixelVal_in_0_5;
      end else if (10'h22d == _T_28[9:0]) begin
        image_0_557 <= io_pixelVal_in_0_4;
      end else if (10'h22d == _T_25[9:0]) begin
        image_0_557 <= io_pixelVal_in_0_3;
      end else if (10'h22d == _T_22[9:0]) begin
        image_0_557 <= io_pixelVal_in_0_2;
      end else if (10'h22d == _T_19[9:0]) begin
        image_0_557 <= io_pixelVal_in_0_1;
      end else if (10'h22d == _T_15[9:0]) begin
        image_0_557 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_558 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h22e == _T_37[9:0]) begin
        image_0_558 <= io_pixelVal_in_0_7;
      end else if (10'h22e == _T_34[9:0]) begin
        image_0_558 <= io_pixelVal_in_0_6;
      end else if (10'h22e == _T_31[9:0]) begin
        image_0_558 <= io_pixelVal_in_0_5;
      end else if (10'h22e == _T_28[9:0]) begin
        image_0_558 <= io_pixelVal_in_0_4;
      end else if (10'h22e == _T_25[9:0]) begin
        image_0_558 <= io_pixelVal_in_0_3;
      end else if (10'h22e == _T_22[9:0]) begin
        image_0_558 <= io_pixelVal_in_0_2;
      end else if (10'h22e == _T_19[9:0]) begin
        image_0_558 <= io_pixelVal_in_0_1;
      end else if (10'h22e == _T_15[9:0]) begin
        image_0_558 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_559 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h22f == _T_37[9:0]) begin
        image_0_559 <= io_pixelVal_in_0_7;
      end else if (10'h22f == _T_34[9:0]) begin
        image_0_559 <= io_pixelVal_in_0_6;
      end else if (10'h22f == _T_31[9:0]) begin
        image_0_559 <= io_pixelVal_in_0_5;
      end else if (10'h22f == _T_28[9:0]) begin
        image_0_559 <= io_pixelVal_in_0_4;
      end else if (10'h22f == _T_25[9:0]) begin
        image_0_559 <= io_pixelVal_in_0_3;
      end else if (10'h22f == _T_22[9:0]) begin
        image_0_559 <= io_pixelVal_in_0_2;
      end else if (10'h22f == _T_19[9:0]) begin
        image_0_559 <= io_pixelVal_in_0_1;
      end else if (10'h22f == _T_15[9:0]) begin
        image_0_559 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_560 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h230 == _T_37[9:0]) begin
        image_0_560 <= io_pixelVal_in_0_7;
      end else if (10'h230 == _T_34[9:0]) begin
        image_0_560 <= io_pixelVal_in_0_6;
      end else if (10'h230 == _T_31[9:0]) begin
        image_0_560 <= io_pixelVal_in_0_5;
      end else if (10'h230 == _T_28[9:0]) begin
        image_0_560 <= io_pixelVal_in_0_4;
      end else if (10'h230 == _T_25[9:0]) begin
        image_0_560 <= io_pixelVal_in_0_3;
      end else if (10'h230 == _T_22[9:0]) begin
        image_0_560 <= io_pixelVal_in_0_2;
      end else if (10'h230 == _T_19[9:0]) begin
        image_0_560 <= io_pixelVal_in_0_1;
      end else if (10'h230 == _T_15[9:0]) begin
        image_0_560 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_561 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h231 == _T_37[9:0]) begin
        image_0_561 <= io_pixelVal_in_0_7;
      end else if (10'h231 == _T_34[9:0]) begin
        image_0_561 <= io_pixelVal_in_0_6;
      end else if (10'h231 == _T_31[9:0]) begin
        image_0_561 <= io_pixelVal_in_0_5;
      end else if (10'h231 == _T_28[9:0]) begin
        image_0_561 <= io_pixelVal_in_0_4;
      end else if (10'h231 == _T_25[9:0]) begin
        image_0_561 <= io_pixelVal_in_0_3;
      end else if (10'h231 == _T_22[9:0]) begin
        image_0_561 <= io_pixelVal_in_0_2;
      end else if (10'h231 == _T_19[9:0]) begin
        image_0_561 <= io_pixelVal_in_0_1;
      end else if (10'h231 == _T_15[9:0]) begin
        image_0_561 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_562 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h232 == _T_37[9:0]) begin
        image_0_562 <= io_pixelVal_in_0_7;
      end else if (10'h232 == _T_34[9:0]) begin
        image_0_562 <= io_pixelVal_in_0_6;
      end else if (10'h232 == _T_31[9:0]) begin
        image_0_562 <= io_pixelVal_in_0_5;
      end else if (10'h232 == _T_28[9:0]) begin
        image_0_562 <= io_pixelVal_in_0_4;
      end else if (10'h232 == _T_25[9:0]) begin
        image_0_562 <= io_pixelVal_in_0_3;
      end else if (10'h232 == _T_22[9:0]) begin
        image_0_562 <= io_pixelVal_in_0_2;
      end else if (10'h232 == _T_19[9:0]) begin
        image_0_562 <= io_pixelVal_in_0_1;
      end else if (10'h232 == _T_15[9:0]) begin
        image_0_562 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_563 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h233 == _T_37[9:0]) begin
        image_0_563 <= io_pixelVal_in_0_7;
      end else if (10'h233 == _T_34[9:0]) begin
        image_0_563 <= io_pixelVal_in_0_6;
      end else if (10'h233 == _T_31[9:0]) begin
        image_0_563 <= io_pixelVal_in_0_5;
      end else if (10'h233 == _T_28[9:0]) begin
        image_0_563 <= io_pixelVal_in_0_4;
      end else if (10'h233 == _T_25[9:0]) begin
        image_0_563 <= io_pixelVal_in_0_3;
      end else if (10'h233 == _T_22[9:0]) begin
        image_0_563 <= io_pixelVal_in_0_2;
      end else if (10'h233 == _T_19[9:0]) begin
        image_0_563 <= io_pixelVal_in_0_1;
      end else if (10'h233 == _T_15[9:0]) begin
        image_0_563 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_564 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h234 == _T_37[9:0]) begin
        image_0_564 <= io_pixelVal_in_0_7;
      end else if (10'h234 == _T_34[9:0]) begin
        image_0_564 <= io_pixelVal_in_0_6;
      end else if (10'h234 == _T_31[9:0]) begin
        image_0_564 <= io_pixelVal_in_0_5;
      end else if (10'h234 == _T_28[9:0]) begin
        image_0_564 <= io_pixelVal_in_0_4;
      end else if (10'h234 == _T_25[9:0]) begin
        image_0_564 <= io_pixelVal_in_0_3;
      end else if (10'h234 == _T_22[9:0]) begin
        image_0_564 <= io_pixelVal_in_0_2;
      end else if (10'h234 == _T_19[9:0]) begin
        image_0_564 <= io_pixelVal_in_0_1;
      end else if (10'h234 == _T_15[9:0]) begin
        image_0_564 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_565 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h235 == _T_37[9:0]) begin
        image_0_565 <= io_pixelVal_in_0_7;
      end else if (10'h235 == _T_34[9:0]) begin
        image_0_565 <= io_pixelVal_in_0_6;
      end else if (10'h235 == _T_31[9:0]) begin
        image_0_565 <= io_pixelVal_in_0_5;
      end else if (10'h235 == _T_28[9:0]) begin
        image_0_565 <= io_pixelVal_in_0_4;
      end else if (10'h235 == _T_25[9:0]) begin
        image_0_565 <= io_pixelVal_in_0_3;
      end else if (10'h235 == _T_22[9:0]) begin
        image_0_565 <= io_pixelVal_in_0_2;
      end else if (10'h235 == _T_19[9:0]) begin
        image_0_565 <= io_pixelVal_in_0_1;
      end else if (10'h235 == _T_15[9:0]) begin
        image_0_565 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_566 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h236 == _T_37[9:0]) begin
        image_0_566 <= io_pixelVal_in_0_7;
      end else if (10'h236 == _T_34[9:0]) begin
        image_0_566 <= io_pixelVal_in_0_6;
      end else if (10'h236 == _T_31[9:0]) begin
        image_0_566 <= io_pixelVal_in_0_5;
      end else if (10'h236 == _T_28[9:0]) begin
        image_0_566 <= io_pixelVal_in_0_4;
      end else if (10'h236 == _T_25[9:0]) begin
        image_0_566 <= io_pixelVal_in_0_3;
      end else if (10'h236 == _T_22[9:0]) begin
        image_0_566 <= io_pixelVal_in_0_2;
      end else if (10'h236 == _T_19[9:0]) begin
        image_0_566 <= io_pixelVal_in_0_1;
      end else if (10'h236 == _T_15[9:0]) begin
        image_0_566 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_567 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h237 == _T_37[9:0]) begin
        image_0_567 <= io_pixelVal_in_0_7;
      end else if (10'h237 == _T_34[9:0]) begin
        image_0_567 <= io_pixelVal_in_0_6;
      end else if (10'h237 == _T_31[9:0]) begin
        image_0_567 <= io_pixelVal_in_0_5;
      end else if (10'h237 == _T_28[9:0]) begin
        image_0_567 <= io_pixelVal_in_0_4;
      end else if (10'h237 == _T_25[9:0]) begin
        image_0_567 <= io_pixelVal_in_0_3;
      end else if (10'h237 == _T_22[9:0]) begin
        image_0_567 <= io_pixelVal_in_0_2;
      end else if (10'h237 == _T_19[9:0]) begin
        image_0_567 <= io_pixelVal_in_0_1;
      end else if (10'h237 == _T_15[9:0]) begin
        image_0_567 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_568 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h238 == _T_37[9:0]) begin
        image_0_568 <= io_pixelVal_in_0_7;
      end else if (10'h238 == _T_34[9:0]) begin
        image_0_568 <= io_pixelVal_in_0_6;
      end else if (10'h238 == _T_31[9:0]) begin
        image_0_568 <= io_pixelVal_in_0_5;
      end else if (10'h238 == _T_28[9:0]) begin
        image_0_568 <= io_pixelVal_in_0_4;
      end else if (10'h238 == _T_25[9:0]) begin
        image_0_568 <= io_pixelVal_in_0_3;
      end else if (10'h238 == _T_22[9:0]) begin
        image_0_568 <= io_pixelVal_in_0_2;
      end else if (10'h238 == _T_19[9:0]) begin
        image_0_568 <= io_pixelVal_in_0_1;
      end else if (10'h238 == _T_15[9:0]) begin
        image_0_568 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_569 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h239 == _T_37[9:0]) begin
        image_0_569 <= io_pixelVal_in_0_7;
      end else if (10'h239 == _T_34[9:0]) begin
        image_0_569 <= io_pixelVal_in_0_6;
      end else if (10'h239 == _T_31[9:0]) begin
        image_0_569 <= io_pixelVal_in_0_5;
      end else if (10'h239 == _T_28[9:0]) begin
        image_0_569 <= io_pixelVal_in_0_4;
      end else if (10'h239 == _T_25[9:0]) begin
        image_0_569 <= io_pixelVal_in_0_3;
      end else if (10'h239 == _T_22[9:0]) begin
        image_0_569 <= io_pixelVal_in_0_2;
      end else if (10'h239 == _T_19[9:0]) begin
        image_0_569 <= io_pixelVal_in_0_1;
      end else if (10'h239 == _T_15[9:0]) begin
        image_0_569 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_570 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h23a == _T_37[9:0]) begin
        image_0_570 <= io_pixelVal_in_0_7;
      end else if (10'h23a == _T_34[9:0]) begin
        image_0_570 <= io_pixelVal_in_0_6;
      end else if (10'h23a == _T_31[9:0]) begin
        image_0_570 <= io_pixelVal_in_0_5;
      end else if (10'h23a == _T_28[9:0]) begin
        image_0_570 <= io_pixelVal_in_0_4;
      end else if (10'h23a == _T_25[9:0]) begin
        image_0_570 <= io_pixelVal_in_0_3;
      end else if (10'h23a == _T_22[9:0]) begin
        image_0_570 <= io_pixelVal_in_0_2;
      end else if (10'h23a == _T_19[9:0]) begin
        image_0_570 <= io_pixelVal_in_0_1;
      end else if (10'h23a == _T_15[9:0]) begin
        image_0_570 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_571 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h23b == _T_37[9:0]) begin
        image_0_571 <= io_pixelVal_in_0_7;
      end else if (10'h23b == _T_34[9:0]) begin
        image_0_571 <= io_pixelVal_in_0_6;
      end else if (10'h23b == _T_31[9:0]) begin
        image_0_571 <= io_pixelVal_in_0_5;
      end else if (10'h23b == _T_28[9:0]) begin
        image_0_571 <= io_pixelVal_in_0_4;
      end else if (10'h23b == _T_25[9:0]) begin
        image_0_571 <= io_pixelVal_in_0_3;
      end else if (10'h23b == _T_22[9:0]) begin
        image_0_571 <= io_pixelVal_in_0_2;
      end else if (10'h23b == _T_19[9:0]) begin
        image_0_571 <= io_pixelVal_in_0_1;
      end else if (10'h23b == _T_15[9:0]) begin
        image_0_571 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_572 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h23c == _T_37[9:0]) begin
        image_0_572 <= io_pixelVal_in_0_7;
      end else if (10'h23c == _T_34[9:0]) begin
        image_0_572 <= io_pixelVal_in_0_6;
      end else if (10'h23c == _T_31[9:0]) begin
        image_0_572 <= io_pixelVal_in_0_5;
      end else if (10'h23c == _T_28[9:0]) begin
        image_0_572 <= io_pixelVal_in_0_4;
      end else if (10'h23c == _T_25[9:0]) begin
        image_0_572 <= io_pixelVal_in_0_3;
      end else if (10'h23c == _T_22[9:0]) begin
        image_0_572 <= io_pixelVal_in_0_2;
      end else if (10'h23c == _T_19[9:0]) begin
        image_0_572 <= io_pixelVal_in_0_1;
      end else if (10'h23c == _T_15[9:0]) begin
        image_0_572 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_573 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h23d == _T_37[9:0]) begin
        image_0_573 <= io_pixelVal_in_0_7;
      end else if (10'h23d == _T_34[9:0]) begin
        image_0_573 <= io_pixelVal_in_0_6;
      end else if (10'h23d == _T_31[9:0]) begin
        image_0_573 <= io_pixelVal_in_0_5;
      end else if (10'h23d == _T_28[9:0]) begin
        image_0_573 <= io_pixelVal_in_0_4;
      end else if (10'h23d == _T_25[9:0]) begin
        image_0_573 <= io_pixelVal_in_0_3;
      end else if (10'h23d == _T_22[9:0]) begin
        image_0_573 <= io_pixelVal_in_0_2;
      end else if (10'h23d == _T_19[9:0]) begin
        image_0_573 <= io_pixelVal_in_0_1;
      end else if (10'h23d == _T_15[9:0]) begin
        image_0_573 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_574 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h23e == _T_37[9:0]) begin
        image_0_574 <= io_pixelVal_in_0_7;
      end else if (10'h23e == _T_34[9:0]) begin
        image_0_574 <= io_pixelVal_in_0_6;
      end else if (10'h23e == _T_31[9:0]) begin
        image_0_574 <= io_pixelVal_in_0_5;
      end else if (10'h23e == _T_28[9:0]) begin
        image_0_574 <= io_pixelVal_in_0_4;
      end else if (10'h23e == _T_25[9:0]) begin
        image_0_574 <= io_pixelVal_in_0_3;
      end else if (10'h23e == _T_22[9:0]) begin
        image_0_574 <= io_pixelVal_in_0_2;
      end else if (10'h23e == _T_19[9:0]) begin
        image_0_574 <= io_pixelVal_in_0_1;
      end else if (10'h23e == _T_15[9:0]) begin
        image_0_574 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_575 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h23f == _T_37[9:0]) begin
        image_0_575 <= io_pixelVal_in_0_7;
      end else if (10'h23f == _T_34[9:0]) begin
        image_0_575 <= io_pixelVal_in_0_6;
      end else if (10'h23f == _T_31[9:0]) begin
        image_0_575 <= io_pixelVal_in_0_5;
      end else if (10'h23f == _T_28[9:0]) begin
        image_0_575 <= io_pixelVal_in_0_4;
      end else if (10'h23f == _T_25[9:0]) begin
        image_0_575 <= io_pixelVal_in_0_3;
      end else if (10'h23f == _T_22[9:0]) begin
        image_0_575 <= io_pixelVal_in_0_2;
      end else if (10'h23f == _T_19[9:0]) begin
        image_0_575 <= io_pixelVal_in_0_1;
      end else if (10'h23f == _T_15[9:0]) begin
        image_0_575 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_1_0 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h0 == _T_37[9:0]) begin
        image_1_0 <= io_pixelVal_in_1_7;
      end else if (10'h0 == _T_34[9:0]) begin
        image_1_0 <= io_pixelVal_in_1_6;
      end else if (10'h0 == _T_31[9:0]) begin
        image_1_0 <= io_pixelVal_in_1_5;
      end else if (10'h0 == _T_28[9:0]) begin
        image_1_0 <= io_pixelVal_in_1_4;
      end else if (10'h0 == _T_25[9:0]) begin
        image_1_0 <= io_pixelVal_in_1_3;
      end else if (10'h0 == _T_22[9:0]) begin
        image_1_0 <= io_pixelVal_in_1_2;
      end else if (10'h0 == _T_19[9:0]) begin
        image_1_0 <= io_pixelVal_in_1_1;
      end else if (10'h0 == _T_15[9:0]) begin
        image_1_0 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_1 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1 == _T_37[9:0]) begin
        image_1_1 <= io_pixelVal_in_1_7;
      end else if (10'h1 == _T_34[9:0]) begin
        image_1_1 <= io_pixelVal_in_1_6;
      end else if (10'h1 == _T_31[9:0]) begin
        image_1_1 <= io_pixelVal_in_1_5;
      end else if (10'h1 == _T_28[9:0]) begin
        image_1_1 <= io_pixelVal_in_1_4;
      end else if (10'h1 == _T_25[9:0]) begin
        image_1_1 <= io_pixelVal_in_1_3;
      end else if (10'h1 == _T_22[9:0]) begin
        image_1_1 <= io_pixelVal_in_1_2;
      end else if (10'h1 == _T_19[9:0]) begin
        image_1_1 <= io_pixelVal_in_1_1;
      end else if (10'h1 == _T_15[9:0]) begin
        image_1_1 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_2 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2 == _T_37[9:0]) begin
        image_1_2 <= io_pixelVal_in_1_7;
      end else if (10'h2 == _T_34[9:0]) begin
        image_1_2 <= io_pixelVal_in_1_6;
      end else if (10'h2 == _T_31[9:0]) begin
        image_1_2 <= io_pixelVal_in_1_5;
      end else if (10'h2 == _T_28[9:0]) begin
        image_1_2 <= io_pixelVal_in_1_4;
      end else if (10'h2 == _T_25[9:0]) begin
        image_1_2 <= io_pixelVal_in_1_3;
      end else if (10'h2 == _T_22[9:0]) begin
        image_1_2 <= io_pixelVal_in_1_2;
      end else if (10'h2 == _T_19[9:0]) begin
        image_1_2 <= io_pixelVal_in_1_1;
      end else if (10'h2 == _T_15[9:0]) begin
        image_1_2 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_3 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3 == _T_37[9:0]) begin
        image_1_3 <= io_pixelVal_in_1_7;
      end else if (10'h3 == _T_34[9:0]) begin
        image_1_3 <= io_pixelVal_in_1_6;
      end else if (10'h3 == _T_31[9:0]) begin
        image_1_3 <= io_pixelVal_in_1_5;
      end else if (10'h3 == _T_28[9:0]) begin
        image_1_3 <= io_pixelVal_in_1_4;
      end else if (10'h3 == _T_25[9:0]) begin
        image_1_3 <= io_pixelVal_in_1_3;
      end else if (10'h3 == _T_22[9:0]) begin
        image_1_3 <= io_pixelVal_in_1_2;
      end else if (10'h3 == _T_19[9:0]) begin
        image_1_3 <= io_pixelVal_in_1_1;
      end else if (10'h3 == _T_15[9:0]) begin
        image_1_3 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_4 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4 == _T_37[9:0]) begin
        image_1_4 <= io_pixelVal_in_1_7;
      end else if (10'h4 == _T_34[9:0]) begin
        image_1_4 <= io_pixelVal_in_1_6;
      end else if (10'h4 == _T_31[9:0]) begin
        image_1_4 <= io_pixelVal_in_1_5;
      end else if (10'h4 == _T_28[9:0]) begin
        image_1_4 <= io_pixelVal_in_1_4;
      end else if (10'h4 == _T_25[9:0]) begin
        image_1_4 <= io_pixelVal_in_1_3;
      end else if (10'h4 == _T_22[9:0]) begin
        image_1_4 <= io_pixelVal_in_1_2;
      end else if (10'h4 == _T_19[9:0]) begin
        image_1_4 <= io_pixelVal_in_1_1;
      end else if (10'h4 == _T_15[9:0]) begin
        image_1_4 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_5 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5 == _T_37[9:0]) begin
        image_1_5 <= io_pixelVal_in_1_7;
      end else if (10'h5 == _T_34[9:0]) begin
        image_1_5 <= io_pixelVal_in_1_6;
      end else if (10'h5 == _T_31[9:0]) begin
        image_1_5 <= io_pixelVal_in_1_5;
      end else if (10'h5 == _T_28[9:0]) begin
        image_1_5 <= io_pixelVal_in_1_4;
      end else if (10'h5 == _T_25[9:0]) begin
        image_1_5 <= io_pixelVal_in_1_3;
      end else if (10'h5 == _T_22[9:0]) begin
        image_1_5 <= io_pixelVal_in_1_2;
      end else if (10'h5 == _T_19[9:0]) begin
        image_1_5 <= io_pixelVal_in_1_1;
      end else if (10'h5 == _T_15[9:0]) begin
        image_1_5 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_6 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6 == _T_37[9:0]) begin
        image_1_6 <= io_pixelVal_in_1_7;
      end else if (10'h6 == _T_34[9:0]) begin
        image_1_6 <= io_pixelVal_in_1_6;
      end else if (10'h6 == _T_31[9:0]) begin
        image_1_6 <= io_pixelVal_in_1_5;
      end else if (10'h6 == _T_28[9:0]) begin
        image_1_6 <= io_pixelVal_in_1_4;
      end else if (10'h6 == _T_25[9:0]) begin
        image_1_6 <= io_pixelVal_in_1_3;
      end else if (10'h6 == _T_22[9:0]) begin
        image_1_6 <= io_pixelVal_in_1_2;
      end else if (10'h6 == _T_19[9:0]) begin
        image_1_6 <= io_pixelVal_in_1_1;
      end else if (10'h6 == _T_15[9:0]) begin
        image_1_6 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_7 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7 == _T_37[9:0]) begin
        image_1_7 <= io_pixelVal_in_1_7;
      end else if (10'h7 == _T_34[9:0]) begin
        image_1_7 <= io_pixelVal_in_1_6;
      end else if (10'h7 == _T_31[9:0]) begin
        image_1_7 <= io_pixelVal_in_1_5;
      end else if (10'h7 == _T_28[9:0]) begin
        image_1_7 <= io_pixelVal_in_1_4;
      end else if (10'h7 == _T_25[9:0]) begin
        image_1_7 <= io_pixelVal_in_1_3;
      end else if (10'h7 == _T_22[9:0]) begin
        image_1_7 <= io_pixelVal_in_1_2;
      end else if (10'h7 == _T_19[9:0]) begin
        image_1_7 <= io_pixelVal_in_1_1;
      end else if (10'h7 == _T_15[9:0]) begin
        image_1_7 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_8 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8 == _T_37[9:0]) begin
        image_1_8 <= io_pixelVal_in_1_7;
      end else if (10'h8 == _T_34[9:0]) begin
        image_1_8 <= io_pixelVal_in_1_6;
      end else if (10'h8 == _T_31[9:0]) begin
        image_1_8 <= io_pixelVal_in_1_5;
      end else if (10'h8 == _T_28[9:0]) begin
        image_1_8 <= io_pixelVal_in_1_4;
      end else if (10'h8 == _T_25[9:0]) begin
        image_1_8 <= io_pixelVal_in_1_3;
      end else if (10'h8 == _T_22[9:0]) begin
        image_1_8 <= io_pixelVal_in_1_2;
      end else if (10'h8 == _T_19[9:0]) begin
        image_1_8 <= io_pixelVal_in_1_1;
      end else if (10'h8 == _T_15[9:0]) begin
        image_1_8 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_9 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9 == _T_37[9:0]) begin
        image_1_9 <= io_pixelVal_in_1_7;
      end else if (10'h9 == _T_34[9:0]) begin
        image_1_9 <= io_pixelVal_in_1_6;
      end else if (10'h9 == _T_31[9:0]) begin
        image_1_9 <= io_pixelVal_in_1_5;
      end else if (10'h9 == _T_28[9:0]) begin
        image_1_9 <= io_pixelVal_in_1_4;
      end else if (10'h9 == _T_25[9:0]) begin
        image_1_9 <= io_pixelVal_in_1_3;
      end else if (10'h9 == _T_22[9:0]) begin
        image_1_9 <= io_pixelVal_in_1_2;
      end else if (10'h9 == _T_19[9:0]) begin
        image_1_9 <= io_pixelVal_in_1_1;
      end else if (10'h9 == _T_15[9:0]) begin
        image_1_9 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_10 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha == _T_37[9:0]) begin
        image_1_10 <= io_pixelVal_in_1_7;
      end else if (10'ha == _T_34[9:0]) begin
        image_1_10 <= io_pixelVal_in_1_6;
      end else if (10'ha == _T_31[9:0]) begin
        image_1_10 <= io_pixelVal_in_1_5;
      end else if (10'ha == _T_28[9:0]) begin
        image_1_10 <= io_pixelVal_in_1_4;
      end else if (10'ha == _T_25[9:0]) begin
        image_1_10 <= io_pixelVal_in_1_3;
      end else if (10'ha == _T_22[9:0]) begin
        image_1_10 <= io_pixelVal_in_1_2;
      end else if (10'ha == _T_19[9:0]) begin
        image_1_10 <= io_pixelVal_in_1_1;
      end else if (10'ha == _T_15[9:0]) begin
        image_1_10 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_11 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb == _T_37[9:0]) begin
        image_1_11 <= io_pixelVal_in_1_7;
      end else if (10'hb == _T_34[9:0]) begin
        image_1_11 <= io_pixelVal_in_1_6;
      end else if (10'hb == _T_31[9:0]) begin
        image_1_11 <= io_pixelVal_in_1_5;
      end else if (10'hb == _T_28[9:0]) begin
        image_1_11 <= io_pixelVal_in_1_4;
      end else if (10'hb == _T_25[9:0]) begin
        image_1_11 <= io_pixelVal_in_1_3;
      end else if (10'hb == _T_22[9:0]) begin
        image_1_11 <= io_pixelVal_in_1_2;
      end else if (10'hb == _T_19[9:0]) begin
        image_1_11 <= io_pixelVal_in_1_1;
      end else if (10'hb == _T_15[9:0]) begin
        image_1_11 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_12 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc == _T_37[9:0]) begin
        image_1_12 <= io_pixelVal_in_1_7;
      end else if (10'hc == _T_34[9:0]) begin
        image_1_12 <= io_pixelVal_in_1_6;
      end else if (10'hc == _T_31[9:0]) begin
        image_1_12 <= io_pixelVal_in_1_5;
      end else if (10'hc == _T_28[9:0]) begin
        image_1_12 <= io_pixelVal_in_1_4;
      end else if (10'hc == _T_25[9:0]) begin
        image_1_12 <= io_pixelVal_in_1_3;
      end else if (10'hc == _T_22[9:0]) begin
        image_1_12 <= io_pixelVal_in_1_2;
      end else if (10'hc == _T_19[9:0]) begin
        image_1_12 <= io_pixelVal_in_1_1;
      end else if (10'hc == _T_15[9:0]) begin
        image_1_12 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_13 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd == _T_37[9:0]) begin
        image_1_13 <= io_pixelVal_in_1_7;
      end else if (10'hd == _T_34[9:0]) begin
        image_1_13 <= io_pixelVal_in_1_6;
      end else if (10'hd == _T_31[9:0]) begin
        image_1_13 <= io_pixelVal_in_1_5;
      end else if (10'hd == _T_28[9:0]) begin
        image_1_13 <= io_pixelVal_in_1_4;
      end else if (10'hd == _T_25[9:0]) begin
        image_1_13 <= io_pixelVal_in_1_3;
      end else if (10'hd == _T_22[9:0]) begin
        image_1_13 <= io_pixelVal_in_1_2;
      end else if (10'hd == _T_19[9:0]) begin
        image_1_13 <= io_pixelVal_in_1_1;
      end else if (10'hd == _T_15[9:0]) begin
        image_1_13 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_14 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he == _T_37[9:0]) begin
        image_1_14 <= io_pixelVal_in_1_7;
      end else if (10'he == _T_34[9:0]) begin
        image_1_14 <= io_pixelVal_in_1_6;
      end else if (10'he == _T_31[9:0]) begin
        image_1_14 <= io_pixelVal_in_1_5;
      end else if (10'he == _T_28[9:0]) begin
        image_1_14 <= io_pixelVal_in_1_4;
      end else if (10'he == _T_25[9:0]) begin
        image_1_14 <= io_pixelVal_in_1_3;
      end else if (10'he == _T_22[9:0]) begin
        image_1_14 <= io_pixelVal_in_1_2;
      end else if (10'he == _T_19[9:0]) begin
        image_1_14 <= io_pixelVal_in_1_1;
      end else if (10'he == _T_15[9:0]) begin
        image_1_14 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_15 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf == _T_37[9:0]) begin
        image_1_15 <= io_pixelVal_in_1_7;
      end else if (10'hf == _T_34[9:0]) begin
        image_1_15 <= io_pixelVal_in_1_6;
      end else if (10'hf == _T_31[9:0]) begin
        image_1_15 <= io_pixelVal_in_1_5;
      end else if (10'hf == _T_28[9:0]) begin
        image_1_15 <= io_pixelVal_in_1_4;
      end else if (10'hf == _T_25[9:0]) begin
        image_1_15 <= io_pixelVal_in_1_3;
      end else if (10'hf == _T_22[9:0]) begin
        image_1_15 <= io_pixelVal_in_1_2;
      end else if (10'hf == _T_19[9:0]) begin
        image_1_15 <= io_pixelVal_in_1_1;
      end else if (10'hf == _T_15[9:0]) begin
        image_1_15 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_16 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10 == _T_37[9:0]) begin
        image_1_16 <= io_pixelVal_in_1_7;
      end else if (10'h10 == _T_34[9:0]) begin
        image_1_16 <= io_pixelVal_in_1_6;
      end else if (10'h10 == _T_31[9:0]) begin
        image_1_16 <= io_pixelVal_in_1_5;
      end else if (10'h10 == _T_28[9:0]) begin
        image_1_16 <= io_pixelVal_in_1_4;
      end else if (10'h10 == _T_25[9:0]) begin
        image_1_16 <= io_pixelVal_in_1_3;
      end else if (10'h10 == _T_22[9:0]) begin
        image_1_16 <= io_pixelVal_in_1_2;
      end else if (10'h10 == _T_19[9:0]) begin
        image_1_16 <= io_pixelVal_in_1_1;
      end else if (10'h10 == _T_15[9:0]) begin
        image_1_16 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_17 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11 == _T_37[9:0]) begin
        image_1_17 <= io_pixelVal_in_1_7;
      end else if (10'h11 == _T_34[9:0]) begin
        image_1_17 <= io_pixelVal_in_1_6;
      end else if (10'h11 == _T_31[9:0]) begin
        image_1_17 <= io_pixelVal_in_1_5;
      end else if (10'h11 == _T_28[9:0]) begin
        image_1_17 <= io_pixelVal_in_1_4;
      end else if (10'h11 == _T_25[9:0]) begin
        image_1_17 <= io_pixelVal_in_1_3;
      end else if (10'h11 == _T_22[9:0]) begin
        image_1_17 <= io_pixelVal_in_1_2;
      end else if (10'h11 == _T_19[9:0]) begin
        image_1_17 <= io_pixelVal_in_1_1;
      end else if (10'h11 == _T_15[9:0]) begin
        image_1_17 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_18 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12 == _T_37[9:0]) begin
        image_1_18 <= io_pixelVal_in_1_7;
      end else if (10'h12 == _T_34[9:0]) begin
        image_1_18 <= io_pixelVal_in_1_6;
      end else if (10'h12 == _T_31[9:0]) begin
        image_1_18 <= io_pixelVal_in_1_5;
      end else if (10'h12 == _T_28[9:0]) begin
        image_1_18 <= io_pixelVal_in_1_4;
      end else if (10'h12 == _T_25[9:0]) begin
        image_1_18 <= io_pixelVal_in_1_3;
      end else if (10'h12 == _T_22[9:0]) begin
        image_1_18 <= io_pixelVal_in_1_2;
      end else if (10'h12 == _T_19[9:0]) begin
        image_1_18 <= io_pixelVal_in_1_1;
      end else if (10'h12 == _T_15[9:0]) begin
        image_1_18 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_19 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13 == _T_37[9:0]) begin
        image_1_19 <= io_pixelVal_in_1_7;
      end else if (10'h13 == _T_34[9:0]) begin
        image_1_19 <= io_pixelVal_in_1_6;
      end else if (10'h13 == _T_31[9:0]) begin
        image_1_19 <= io_pixelVal_in_1_5;
      end else if (10'h13 == _T_28[9:0]) begin
        image_1_19 <= io_pixelVal_in_1_4;
      end else if (10'h13 == _T_25[9:0]) begin
        image_1_19 <= io_pixelVal_in_1_3;
      end else if (10'h13 == _T_22[9:0]) begin
        image_1_19 <= io_pixelVal_in_1_2;
      end else if (10'h13 == _T_19[9:0]) begin
        image_1_19 <= io_pixelVal_in_1_1;
      end else if (10'h13 == _T_15[9:0]) begin
        image_1_19 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_20 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14 == _T_37[9:0]) begin
        image_1_20 <= io_pixelVal_in_1_7;
      end else if (10'h14 == _T_34[9:0]) begin
        image_1_20 <= io_pixelVal_in_1_6;
      end else if (10'h14 == _T_31[9:0]) begin
        image_1_20 <= io_pixelVal_in_1_5;
      end else if (10'h14 == _T_28[9:0]) begin
        image_1_20 <= io_pixelVal_in_1_4;
      end else if (10'h14 == _T_25[9:0]) begin
        image_1_20 <= io_pixelVal_in_1_3;
      end else if (10'h14 == _T_22[9:0]) begin
        image_1_20 <= io_pixelVal_in_1_2;
      end else if (10'h14 == _T_19[9:0]) begin
        image_1_20 <= io_pixelVal_in_1_1;
      end else if (10'h14 == _T_15[9:0]) begin
        image_1_20 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_21 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15 == _T_37[9:0]) begin
        image_1_21 <= io_pixelVal_in_1_7;
      end else if (10'h15 == _T_34[9:0]) begin
        image_1_21 <= io_pixelVal_in_1_6;
      end else if (10'h15 == _T_31[9:0]) begin
        image_1_21 <= io_pixelVal_in_1_5;
      end else if (10'h15 == _T_28[9:0]) begin
        image_1_21 <= io_pixelVal_in_1_4;
      end else if (10'h15 == _T_25[9:0]) begin
        image_1_21 <= io_pixelVal_in_1_3;
      end else if (10'h15 == _T_22[9:0]) begin
        image_1_21 <= io_pixelVal_in_1_2;
      end else if (10'h15 == _T_19[9:0]) begin
        image_1_21 <= io_pixelVal_in_1_1;
      end else if (10'h15 == _T_15[9:0]) begin
        image_1_21 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_22 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16 == _T_37[9:0]) begin
        image_1_22 <= io_pixelVal_in_1_7;
      end else if (10'h16 == _T_34[9:0]) begin
        image_1_22 <= io_pixelVal_in_1_6;
      end else if (10'h16 == _T_31[9:0]) begin
        image_1_22 <= io_pixelVal_in_1_5;
      end else if (10'h16 == _T_28[9:0]) begin
        image_1_22 <= io_pixelVal_in_1_4;
      end else if (10'h16 == _T_25[9:0]) begin
        image_1_22 <= io_pixelVal_in_1_3;
      end else if (10'h16 == _T_22[9:0]) begin
        image_1_22 <= io_pixelVal_in_1_2;
      end else if (10'h16 == _T_19[9:0]) begin
        image_1_22 <= io_pixelVal_in_1_1;
      end else if (10'h16 == _T_15[9:0]) begin
        image_1_22 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_23 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17 == _T_37[9:0]) begin
        image_1_23 <= io_pixelVal_in_1_7;
      end else if (10'h17 == _T_34[9:0]) begin
        image_1_23 <= io_pixelVal_in_1_6;
      end else if (10'h17 == _T_31[9:0]) begin
        image_1_23 <= io_pixelVal_in_1_5;
      end else if (10'h17 == _T_28[9:0]) begin
        image_1_23 <= io_pixelVal_in_1_4;
      end else if (10'h17 == _T_25[9:0]) begin
        image_1_23 <= io_pixelVal_in_1_3;
      end else if (10'h17 == _T_22[9:0]) begin
        image_1_23 <= io_pixelVal_in_1_2;
      end else if (10'h17 == _T_19[9:0]) begin
        image_1_23 <= io_pixelVal_in_1_1;
      end else if (10'h17 == _T_15[9:0]) begin
        image_1_23 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_24 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18 == _T_37[9:0]) begin
        image_1_24 <= io_pixelVal_in_1_7;
      end else if (10'h18 == _T_34[9:0]) begin
        image_1_24 <= io_pixelVal_in_1_6;
      end else if (10'h18 == _T_31[9:0]) begin
        image_1_24 <= io_pixelVal_in_1_5;
      end else if (10'h18 == _T_28[9:0]) begin
        image_1_24 <= io_pixelVal_in_1_4;
      end else if (10'h18 == _T_25[9:0]) begin
        image_1_24 <= io_pixelVal_in_1_3;
      end else if (10'h18 == _T_22[9:0]) begin
        image_1_24 <= io_pixelVal_in_1_2;
      end else if (10'h18 == _T_19[9:0]) begin
        image_1_24 <= io_pixelVal_in_1_1;
      end else if (10'h18 == _T_15[9:0]) begin
        image_1_24 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_25 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19 == _T_37[9:0]) begin
        image_1_25 <= io_pixelVal_in_1_7;
      end else if (10'h19 == _T_34[9:0]) begin
        image_1_25 <= io_pixelVal_in_1_6;
      end else if (10'h19 == _T_31[9:0]) begin
        image_1_25 <= io_pixelVal_in_1_5;
      end else if (10'h19 == _T_28[9:0]) begin
        image_1_25 <= io_pixelVal_in_1_4;
      end else if (10'h19 == _T_25[9:0]) begin
        image_1_25 <= io_pixelVal_in_1_3;
      end else if (10'h19 == _T_22[9:0]) begin
        image_1_25 <= io_pixelVal_in_1_2;
      end else if (10'h19 == _T_19[9:0]) begin
        image_1_25 <= io_pixelVal_in_1_1;
      end else if (10'h19 == _T_15[9:0]) begin
        image_1_25 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_26 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a == _T_37[9:0]) begin
        image_1_26 <= io_pixelVal_in_1_7;
      end else if (10'h1a == _T_34[9:0]) begin
        image_1_26 <= io_pixelVal_in_1_6;
      end else if (10'h1a == _T_31[9:0]) begin
        image_1_26 <= io_pixelVal_in_1_5;
      end else if (10'h1a == _T_28[9:0]) begin
        image_1_26 <= io_pixelVal_in_1_4;
      end else if (10'h1a == _T_25[9:0]) begin
        image_1_26 <= io_pixelVal_in_1_3;
      end else if (10'h1a == _T_22[9:0]) begin
        image_1_26 <= io_pixelVal_in_1_2;
      end else if (10'h1a == _T_19[9:0]) begin
        image_1_26 <= io_pixelVal_in_1_1;
      end else if (10'h1a == _T_15[9:0]) begin
        image_1_26 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_27 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b == _T_37[9:0]) begin
        image_1_27 <= io_pixelVal_in_1_7;
      end else if (10'h1b == _T_34[9:0]) begin
        image_1_27 <= io_pixelVal_in_1_6;
      end else if (10'h1b == _T_31[9:0]) begin
        image_1_27 <= io_pixelVal_in_1_5;
      end else if (10'h1b == _T_28[9:0]) begin
        image_1_27 <= io_pixelVal_in_1_4;
      end else if (10'h1b == _T_25[9:0]) begin
        image_1_27 <= io_pixelVal_in_1_3;
      end else if (10'h1b == _T_22[9:0]) begin
        image_1_27 <= io_pixelVal_in_1_2;
      end else if (10'h1b == _T_19[9:0]) begin
        image_1_27 <= io_pixelVal_in_1_1;
      end else if (10'h1b == _T_15[9:0]) begin
        image_1_27 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_28 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c == _T_37[9:0]) begin
        image_1_28 <= io_pixelVal_in_1_7;
      end else if (10'h1c == _T_34[9:0]) begin
        image_1_28 <= io_pixelVal_in_1_6;
      end else if (10'h1c == _T_31[9:0]) begin
        image_1_28 <= io_pixelVal_in_1_5;
      end else if (10'h1c == _T_28[9:0]) begin
        image_1_28 <= io_pixelVal_in_1_4;
      end else if (10'h1c == _T_25[9:0]) begin
        image_1_28 <= io_pixelVal_in_1_3;
      end else if (10'h1c == _T_22[9:0]) begin
        image_1_28 <= io_pixelVal_in_1_2;
      end else if (10'h1c == _T_19[9:0]) begin
        image_1_28 <= io_pixelVal_in_1_1;
      end else if (10'h1c == _T_15[9:0]) begin
        image_1_28 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_29 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d == _T_37[9:0]) begin
        image_1_29 <= io_pixelVal_in_1_7;
      end else if (10'h1d == _T_34[9:0]) begin
        image_1_29 <= io_pixelVal_in_1_6;
      end else if (10'h1d == _T_31[9:0]) begin
        image_1_29 <= io_pixelVal_in_1_5;
      end else if (10'h1d == _T_28[9:0]) begin
        image_1_29 <= io_pixelVal_in_1_4;
      end else if (10'h1d == _T_25[9:0]) begin
        image_1_29 <= io_pixelVal_in_1_3;
      end else if (10'h1d == _T_22[9:0]) begin
        image_1_29 <= io_pixelVal_in_1_2;
      end else if (10'h1d == _T_19[9:0]) begin
        image_1_29 <= io_pixelVal_in_1_1;
      end else if (10'h1d == _T_15[9:0]) begin
        image_1_29 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_30 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e == _T_37[9:0]) begin
        image_1_30 <= io_pixelVal_in_1_7;
      end else if (10'h1e == _T_34[9:0]) begin
        image_1_30 <= io_pixelVal_in_1_6;
      end else if (10'h1e == _T_31[9:0]) begin
        image_1_30 <= io_pixelVal_in_1_5;
      end else if (10'h1e == _T_28[9:0]) begin
        image_1_30 <= io_pixelVal_in_1_4;
      end else if (10'h1e == _T_25[9:0]) begin
        image_1_30 <= io_pixelVal_in_1_3;
      end else if (10'h1e == _T_22[9:0]) begin
        image_1_30 <= io_pixelVal_in_1_2;
      end else if (10'h1e == _T_19[9:0]) begin
        image_1_30 <= io_pixelVal_in_1_1;
      end else if (10'h1e == _T_15[9:0]) begin
        image_1_30 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_31 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f == _T_37[9:0]) begin
        image_1_31 <= io_pixelVal_in_1_7;
      end else if (10'h1f == _T_34[9:0]) begin
        image_1_31 <= io_pixelVal_in_1_6;
      end else if (10'h1f == _T_31[9:0]) begin
        image_1_31 <= io_pixelVal_in_1_5;
      end else if (10'h1f == _T_28[9:0]) begin
        image_1_31 <= io_pixelVal_in_1_4;
      end else if (10'h1f == _T_25[9:0]) begin
        image_1_31 <= io_pixelVal_in_1_3;
      end else if (10'h1f == _T_22[9:0]) begin
        image_1_31 <= io_pixelVal_in_1_2;
      end else if (10'h1f == _T_19[9:0]) begin
        image_1_31 <= io_pixelVal_in_1_1;
      end else if (10'h1f == _T_15[9:0]) begin
        image_1_31 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_32 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20 == _T_37[9:0]) begin
        image_1_32 <= io_pixelVal_in_1_7;
      end else if (10'h20 == _T_34[9:0]) begin
        image_1_32 <= io_pixelVal_in_1_6;
      end else if (10'h20 == _T_31[9:0]) begin
        image_1_32 <= io_pixelVal_in_1_5;
      end else if (10'h20 == _T_28[9:0]) begin
        image_1_32 <= io_pixelVal_in_1_4;
      end else if (10'h20 == _T_25[9:0]) begin
        image_1_32 <= io_pixelVal_in_1_3;
      end else if (10'h20 == _T_22[9:0]) begin
        image_1_32 <= io_pixelVal_in_1_2;
      end else if (10'h20 == _T_19[9:0]) begin
        image_1_32 <= io_pixelVal_in_1_1;
      end else if (10'h20 == _T_15[9:0]) begin
        image_1_32 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_33 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21 == _T_37[9:0]) begin
        image_1_33 <= io_pixelVal_in_1_7;
      end else if (10'h21 == _T_34[9:0]) begin
        image_1_33 <= io_pixelVal_in_1_6;
      end else if (10'h21 == _T_31[9:0]) begin
        image_1_33 <= io_pixelVal_in_1_5;
      end else if (10'h21 == _T_28[9:0]) begin
        image_1_33 <= io_pixelVal_in_1_4;
      end else if (10'h21 == _T_25[9:0]) begin
        image_1_33 <= io_pixelVal_in_1_3;
      end else if (10'h21 == _T_22[9:0]) begin
        image_1_33 <= io_pixelVal_in_1_2;
      end else if (10'h21 == _T_19[9:0]) begin
        image_1_33 <= io_pixelVal_in_1_1;
      end else if (10'h21 == _T_15[9:0]) begin
        image_1_33 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_34 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22 == _T_37[9:0]) begin
        image_1_34 <= io_pixelVal_in_1_7;
      end else if (10'h22 == _T_34[9:0]) begin
        image_1_34 <= io_pixelVal_in_1_6;
      end else if (10'h22 == _T_31[9:0]) begin
        image_1_34 <= io_pixelVal_in_1_5;
      end else if (10'h22 == _T_28[9:0]) begin
        image_1_34 <= io_pixelVal_in_1_4;
      end else if (10'h22 == _T_25[9:0]) begin
        image_1_34 <= io_pixelVal_in_1_3;
      end else if (10'h22 == _T_22[9:0]) begin
        image_1_34 <= io_pixelVal_in_1_2;
      end else if (10'h22 == _T_19[9:0]) begin
        image_1_34 <= io_pixelVal_in_1_1;
      end else if (10'h22 == _T_15[9:0]) begin
        image_1_34 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_35 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23 == _T_37[9:0]) begin
        image_1_35 <= io_pixelVal_in_1_7;
      end else if (10'h23 == _T_34[9:0]) begin
        image_1_35 <= io_pixelVal_in_1_6;
      end else if (10'h23 == _T_31[9:0]) begin
        image_1_35 <= io_pixelVal_in_1_5;
      end else if (10'h23 == _T_28[9:0]) begin
        image_1_35 <= io_pixelVal_in_1_4;
      end else if (10'h23 == _T_25[9:0]) begin
        image_1_35 <= io_pixelVal_in_1_3;
      end else if (10'h23 == _T_22[9:0]) begin
        image_1_35 <= io_pixelVal_in_1_2;
      end else if (10'h23 == _T_19[9:0]) begin
        image_1_35 <= io_pixelVal_in_1_1;
      end else if (10'h23 == _T_15[9:0]) begin
        image_1_35 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_36 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h24 == _T_37[9:0]) begin
        image_1_36 <= io_pixelVal_in_1_7;
      end else if (10'h24 == _T_34[9:0]) begin
        image_1_36 <= io_pixelVal_in_1_6;
      end else if (10'h24 == _T_31[9:0]) begin
        image_1_36 <= io_pixelVal_in_1_5;
      end else if (10'h24 == _T_28[9:0]) begin
        image_1_36 <= io_pixelVal_in_1_4;
      end else if (10'h24 == _T_25[9:0]) begin
        image_1_36 <= io_pixelVal_in_1_3;
      end else if (10'h24 == _T_22[9:0]) begin
        image_1_36 <= io_pixelVal_in_1_2;
      end else if (10'h24 == _T_19[9:0]) begin
        image_1_36 <= io_pixelVal_in_1_1;
      end else if (10'h24 == _T_15[9:0]) begin
        image_1_36 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_37 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h25 == _T_37[9:0]) begin
        image_1_37 <= io_pixelVal_in_1_7;
      end else if (10'h25 == _T_34[9:0]) begin
        image_1_37 <= io_pixelVal_in_1_6;
      end else if (10'h25 == _T_31[9:0]) begin
        image_1_37 <= io_pixelVal_in_1_5;
      end else if (10'h25 == _T_28[9:0]) begin
        image_1_37 <= io_pixelVal_in_1_4;
      end else if (10'h25 == _T_25[9:0]) begin
        image_1_37 <= io_pixelVal_in_1_3;
      end else if (10'h25 == _T_22[9:0]) begin
        image_1_37 <= io_pixelVal_in_1_2;
      end else if (10'h25 == _T_19[9:0]) begin
        image_1_37 <= io_pixelVal_in_1_1;
      end else if (10'h25 == _T_15[9:0]) begin
        image_1_37 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_38 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h26 == _T_37[9:0]) begin
        image_1_38 <= io_pixelVal_in_1_7;
      end else if (10'h26 == _T_34[9:0]) begin
        image_1_38 <= io_pixelVal_in_1_6;
      end else if (10'h26 == _T_31[9:0]) begin
        image_1_38 <= io_pixelVal_in_1_5;
      end else if (10'h26 == _T_28[9:0]) begin
        image_1_38 <= io_pixelVal_in_1_4;
      end else if (10'h26 == _T_25[9:0]) begin
        image_1_38 <= io_pixelVal_in_1_3;
      end else if (10'h26 == _T_22[9:0]) begin
        image_1_38 <= io_pixelVal_in_1_2;
      end else if (10'h26 == _T_19[9:0]) begin
        image_1_38 <= io_pixelVal_in_1_1;
      end else if (10'h26 == _T_15[9:0]) begin
        image_1_38 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_39 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h27 == _T_37[9:0]) begin
        image_1_39 <= io_pixelVal_in_1_7;
      end else if (10'h27 == _T_34[9:0]) begin
        image_1_39 <= io_pixelVal_in_1_6;
      end else if (10'h27 == _T_31[9:0]) begin
        image_1_39 <= io_pixelVal_in_1_5;
      end else if (10'h27 == _T_28[9:0]) begin
        image_1_39 <= io_pixelVal_in_1_4;
      end else if (10'h27 == _T_25[9:0]) begin
        image_1_39 <= io_pixelVal_in_1_3;
      end else if (10'h27 == _T_22[9:0]) begin
        image_1_39 <= io_pixelVal_in_1_2;
      end else if (10'h27 == _T_19[9:0]) begin
        image_1_39 <= io_pixelVal_in_1_1;
      end else if (10'h27 == _T_15[9:0]) begin
        image_1_39 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_40 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h28 == _T_37[9:0]) begin
        image_1_40 <= io_pixelVal_in_1_7;
      end else if (10'h28 == _T_34[9:0]) begin
        image_1_40 <= io_pixelVal_in_1_6;
      end else if (10'h28 == _T_31[9:0]) begin
        image_1_40 <= io_pixelVal_in_1_5;
      end else if (10'h28 == _T_28[9:0]) begin
        image_1_40 <= io_pixelVal_in_1_4;
      end else if (10'h28 == _T_25[9:0]) begin
        image_1_40 <= io_pixelVal_in_1_3;
      end else if (10'h28 == _T_22[9:0]) begin
        image_1_40 <= io_pixelVal_in_1_2;
      end else if (10'h28 == _T_19[9:0]) begin
        image_1_40 <= io_pixelVal_in_1_1;
      end else if (10'h28 == _T_15[9:0]) begin
        image_1_40 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_41 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h29 == _T_37[9:0]) begin
        image_1_41 <= io_pixelVal_in_1_7;
      end else if (10'h29 == _T_34[9:0]) begin
        image_1_41 <= io_pixelVal_in_1_6;
      end else if (10'h29 == _T_31[9:0]) begin
        image_1_41 <= io_pixelVal_in_1_5;
      end else if (10'h29 == _T_28[9:0]) begin
        image_1_41 <= io_pixelVal_in_1_4;
      end else if (10'h29 == _T_25[9:0]) begin
        image_1_41 <= io_pixelVal_in_1_3;
      end else if (10'h29 == _T_22[9:0]) begin
        image_1_41 <= io_pixelVal_in_1_2;
      end else if (10'h29 == _T_19[9:0]) begin
        image_1_41 <= io_pixelVal_in_1_1;
      end else if (10'h29 == _T_15[9:0]) begin
        image_1_41 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_42 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2a == _T_37[9:0]) begin
        image_1_42 <= io_pixelVal_in_1_7;
      end else if (10'h2a == _T_34[9:0]) begin
        image_1_42 <= io_pixelVal_in_1_6;
      end else if (10'h2a == _T_31[9:0]) begin
        image_1_42 <= io_pixelVal_in_1_5;
      end else if (10'h2a == _T_28[9:0]) begin
        image_1_42 <= io_pixelVal_in_1_4;
      end else if (10'h2a == _T_25[9:0]) begin
        image_1_42 <= io_pixelVal_in_1_3;
      end else if (10'h2a == _T_22[9:0]) begin
        image_1_42 <= io_pixelVal_in_1_2;
      end else if (10'h2a == _T_19[9:0]) begin
        image_1_42 <= io_pixelVal_in_1_1;
      end else if (10'h2a == _T_15[9:0]) begin
        image_1_42 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_43 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2b == _T_37[9:0]) begin
        image_1_43 <= io_pixelVal_in_1_7;
      end else if (10'h2b == _T_34[9:0]) begin
        image_1_43 <= io_pixelVal_in_1_6;
      end else if (10'h2b == _T_31[9:0]) begin
        image_1_43 <= io_pixelVal_in_1_5;
      end else if (10'h2b == _T_28[9:0]) begin
        image_1_43 <= io_pixelVal_in_1_4;
      end else if (10'h2b == _T_25[9:0]) begin
        image_1_43 <= io_pixelVal_in_1_3;
      end else if (10'h2b == _T_22[9:0]) begin
        image_1_43 <= io_pixelVal_in_1_2;
      end else if (10'h2b == _T_19[9:0]) begin
        image_1_43 <= io_pixelVal_in_1_1;
      end else if (10'h2b == _T_15[9:0]) begin
        image_1_43 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_44 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2c == _T_37[9:0]) begin
        image_1_44 <= io_pixelVal_in_1_7;
      end else if (10'h2c == _T_34[9:0]) begin
        image_1_44 <= io_pixelVal_in_1_6;
      end else if (10'h2c == _T_31[9:0]) begin
        image_1_44 <= io_pixelVal_in_1_5;
      end else if (10'h2c == _T_28[9:0]) begin
        image_1_44 <= io_pixelVal_in_1_4;
      end else if (10'h2c == _T_25[9:0]) begin
        image_1_44 <= io_pixelVal_in_1_3;
      end else if (10'h2c == _T_22[9:0]) begin
        image_1_44 <= io_pixelVal_in_1_2;
      end else if (10'h2c == _T_19[9:0]) begin
        image_1_44 <= io_pixelVal_in_1_1;
      end else if (10'h2c == _T_15[9:0]) begin
        image_1_44 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_45 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2d == _T_37[9:0]) begin
        image_1_45 <= io_pixelVal_in_1_7;
      end else if (10'h2d == _T_34[9:0]) begin
        image_1_45 <= io_pixelVal_in_1_6;
      end else if (10'h2d == _T_31[9:0]) begin
        image_1_45 <= io_pixelVal_in_1_5;
      end else if (10'h2d == _T_28[9:0]) begin
        image_1_45 <= io_pixelVal_in_1_4;
      end else if (10'h2d == _T_25[9:0]) begin
        image_1_45 <= io_pixelVal_in_1_3;
      end else if (10'h2d == _T_22[9:0]) begin
        image_1_45 <= io_pixelVal_in_1_2;
      end else if (10'h2d == _T_19[9:0]) begin
        image_1_45 <= io_pixelVal_in_1_1;
      end else if (10'h2d == _T_15[9:0]) begin
        image_1_45 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_46 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2e == _T_37[9:0]) begin
        image_1_46 <= io_pixelVal_in_1_7;
      end else if (10'h2e == _T_34[9:0]) begin
        image_1_46 <= io_pixelVal_in_1_6;
      end else if (10'h2e == _T_31[9:0]) begin
        image_1_46 <= io_pixelVal_in_1_5;
      end else if (10'h2e == _T_28[9:0]) begin
        image_1_46 <= io_pixelVal_in_1_4;
      end else if (10'h2e == _T_25[9:0]) begin
        image_1_46 <= io_pixelVal_in_1_3;
      end else if (10'h2e == _T_22[9:0]) begin
        image_1_46 <= io_pixelVal_in_1_2;
      end else if (10'h2e == _T_19[9:0]) begin
        image_1_46 <= io_pixelVal_in_1_1;
      end else if (10'h2e == _T_15[9:0]) begin
        image_1_46 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_47 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2f == _T_37[9:0]) begin
        image_1_47 <= io_pixelVal_in_1_7;
      end else if (10'h2f == _T_34[9:0]) begin
        image_1_47 <= io_pixelVal_in_1_6;
      end else if (10'h2f == _T_31[9:0]) begin
        image_1_47 <= io_pixelVal_in_1_5;
      end else if (10'h2f == _T_28[9:0]) begin
        image_1_47 <= io_pixelVal_in_1_4;
      end else if (10'h2f == _T_25[9:0]) begin
        image_1_47 <= io_pixelVal_in_1_3;
      end else if (10'h2f == _T_22[9:0]) begin
        image_1_47 <= io_pixelVal_in_1_2;
      end else if (10'h2f == _T_19[9:0]) begin
        image_1_47 <= io_pixelVal_in_1_1;
      end else if (10'h2f == _T_15[9:0]) begin
        image_1_47 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_48 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h30 == _T_37[9:0]) begin
        image_1_48 <= io_pixelVal_in_1_7;
      end else if (10'h30 == _T_34[9:0]) begin
        image_1_48 <= io_pixelVal_in_1_6;
      end else if (10'h30 == _T_31[9:0]) begin
        image_1_48 <= io_pixelVal_in_1_5;
      end else if (10'h30 == _T_28[9:0]) begin
        image_1_48 <= io_pixelVal_in_1_4;
      end else if (10'h30 == _T_25[9:0]) begin
        image_1_48 <= io_pixelVal_in_1_3;
      end else if (10'h30 == _T_22[9:0]) begin
        image_1_48 <= io_pixelVal_in_1_2;
      end else if (10'h30 == _T_19[9:0]) begin
        image_1_48 <= io_pixelVal_in_1_1;
      end else if (10'h30 == _T_15[9:0]) begin
        image_1_48 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_49 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h31 == _T_37[9:0]) begin
        image_1_49 <= io_pixelVal_in_1_7;
      end else if (10'h31 == _T_34[9:0]) begin
        image_1_49 <= io_pixelVal_in_1_6;
      end else if (10'h31 == _T_31[9:0]) begin
        image_1_49 <= io_pixelVal_in_1_5;
      end else if (10'h31 == _T_28[9:0]) begin
        image_1_49 <= io_pixelVal_in_1_4;
      end else if (10'h31 == _T_25[9:0]) begin
        image_1_49 <= io_pixelVal_in_1_3;
      end else if (10'h31 == _T_22[9:0]) begin
        image_1_49 <= io_pixelVal_in_1_2;
      end else if (10'h31 == _T_19[9:0]) begin
        image_1_49 <= io_pixelVal_in_1_1;
      end else if (10'h31 == _T_15[9:0]) begin
        image_1_49 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_50 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h32 == _T_37[9:0]) begin
        image_1_50 <= io_pixelVal_in_1_7;
      end else if (10'h32 == _T_34[9:0]) begin
        image_1_50 <= io_pixelVal_in_1_6;
      end else if (10'h32 == _T_31[9:0]) begin
        image_1_50 <= io_pixelVal_in_1_5;
      end else if (10'h32 == _T_28[9:0]) begin
        image_1_50 <= io_pixelVal_in_1_4;
      end else if (10'h32 == _T_25[9:0]) begin
        image_1_50 <= io_pixelVal_in_1_3;
      end else if (10'h32 == _T_22[9:0]) begin
        image_1_50 <= io_pixelVal_in_1_2;
      end else if (10'h32 == _T_19[9:0]) begin
        image_1_50 <= io_pixelVal_in_1_1;
      end else if (10'h32 == _T_15[9:0]) begin
        image_1_50 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_51 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h33 == _T_37[9:0]) begin
        image_1_51 <= io_pixelVal_in_1_7;
      end else if (10'h33 == _T_34[9:0]) begin
        image_1_51 <= io_pixelVal_in_1_6;
      end else if (10'h33 == _T_31[9:0]) begin
        image_1_51 <= io_pixelVal_in_1_5;
      end else if (10'h33 == _T_28[9:0]) begin
        image_1_51 <= io_pixelVal_in_1_4;
      end else if (10'h33 == _T_25[9:0]) begin
        image_1_51 <= io_pixelVal_in_1_3;
      end else if (10'h33 == _T_22[9:0]) begin
        image_1_51 <= io_pixelVal_in_1_2;
      end else if (10'h33 == _T_19[9:0]) begin
        image_1_51 <= io_pixelVal_in_1_1;
      end else if (10'h33 == _T_15[9:0]) begin
        image_1_51 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_52 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h34 == _T_37[9:0]) begin
        image_1_52 <= io_pixelVal_in_1_7;
      end else if (10'h34 == _T_34[9:0]) begin
        image_1_52 <= io_pixelVal_in_1_6;
      end else if (10'h34 == _T_31[9:0]) begin
        image_1_52 <= io_pixelVal_in_1_5;
      end else if (10'h34 == _T_28[9:0]) begin
        image_1_52 <= io_pixelVal_in_1_4;
      end else if (10'h34 == _T_25[9:0]) begin
        image_1_52 <= io_pixelVal_in_1_3;
      end else if (10'h34 == _T_22[9:0]) begin
        image_1_52 <= io_pixelVal_in_1_2;
      end else if (10'h34 == _T_19[9:0]) begin
        image_1_52 <= io_pixelVal_in_1_1;
      end else if (10'h34 == _T_15[9:0]) begin
        image_1_52 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_53 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h35 == _T_37[9:0]) begin
        image_1_53 <= io_pixelVal_in_1_7;
      end else if (10'h35 == _T_34[9:0]) begin
        image_1_53 <= io_pixelVal_in_1_6;
      end else if (10'h35 == _T_31[9:0]) begin
        image_1_53 <= io_pixelVal_in_1_5;
      end else if (10'h35 == _T_28[9:0]) begin
        image_1_53 <= io_pixelVal_in_1_4;
      end else if (10'h35 == _T_25[9:0]) begin
        image_1_53 <= io_pixelVal_in_1_3;
      end else if (10'h35 == _T_22[9:0]) begin
        image_1_53 <= io_pixelVal_in_1_2;
      end else if (10'h35 == _T_19[9:0]) begin
        image_1_53 <= io_pixelVal_in_1_1;
      end else if (10'h35 == _T_15[9:0]) begin
        image_1_53 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_54 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h36 == _T_37[9:0]) begin
        image_1_54 <= io_pixelVal_in_1_7;
      end else if (10'h36 == _T_34[9:0]) begin
        image_1_54 <= io_pixelVal_in_1_6;
      end else if (10'h36 == _T_31[9:0]) begin
        image_1_54 <= io_pixelVal_in_1_5;
      end else if (10'h36 == _T_28[9:0]) begin
        image_1_54 <= io_pixelVal_in_1_4;
      end else if (10'h36 == _T_25[9:0]) begin
        image_1_54 <= io_pixelVal_in_1_3;
      end else if (10'h36 == _T_22[9:0]) begin
        image_1_54 <= io_pixelVal_in_1_2;
      end else if (10'h36 == _T_19[9:0]) begin
        image_1_54 <= io_pixelVal_in_1_1;
      end else if (10'h36 == _T_15[9:0]) begin
        image_1_54 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_55 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h37 == _T_37[9:0]) begin
        image_1_55 <= io_pixelVal_in_1_7;
      end else if (10'h37 == _T_34[9:0]) begin
        image_1_55 <= io_pixelVal_in_1_6;
      end else if (10'h37 == _T_31[9:0]) begin
        image_1_55 <= io_pixelVal_in_1_5;
      end else if (10'h37 == _T_28[9:0]) begin
        image_1_55 <= io_pixelVal_in_1_4;
      end else if (10'h37 == _T_25[9:0]) begin
        image_1_55 <= io_pixelVal_in_1_3;
      end else if (10'h37 == _T_22[9:0]) begin
        image_1_55 <= io_pixelVal_in_1_2;
      end else if (10'h37 == _T_19[9:0]) begin
        image_1_55 <= io_pixelVal_in_1_1;
      end else if (10'h37 == _T_15[9:0]) begin
        image_1_55 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_56 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h38 == _T_37[9:0]) begin
        image_1_56 <= io_pixelVal_in_1_7;
      end else if (10'h38 == _T_34[9:0]) begin
        image_1_56 <= io_pixelVal_in_1_6;
      end else if (10'h38 == _T_31[9:0]) begin
        image_1_56 <= io_pixelVal_in_1_5;
      end else if (10'h38 == _T_28[9:0]) begin
        image_1_56 <= io_pixelVal_in_1_4;
      end else if (10'h38 == _T_25[9:0]) begin
        image_1_56 <= io_pixelVal_in_1_3;
      end else if (10'h38 == _T_22[9:0]) begin
        image_1_56 <= io_pixelVal_in_1_2;
      end else if (10'h38 == _T_19[9:0]) begin
        image_1_56 <= io_pixelVal_in_1_1;
      end else if (10'h38 == _T_15[9:0]) begin
        image_1_56 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_57 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h39 == _T_37[9:0]) begin
        image_1_57 <= io_pixelVal_in_1_7;
      end else if (10'h39 == _T_34[9:0]) begin
        image_1_57 <= io_pixelVal_in_1_6;
      end else if (10'h39 == _T_31[9:0]) begin
        image_1_57 <= io_pixelVal_in_1_5;
      end else if (10'h39 == _T_28[9:0]) begin
        image_1_57 <= io_pixelVal_in_1_4;
      end else if (10'h39 == _T_25[9:0]) begin
        image_1_57 <= io_pixelVal_in_1_3;
      end else if (10'h39 == _T_22[9:0]) begin
        image_1_57 <= io_pixelVal_in_1_2;
      end else if (10'h39 == _T_19[9:0]) begin
        image_1_57 <= io_pixelVal_in_1_1;
      end else if (10'h39 == _T_15[9:0]) begin
        image_1_57 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_58 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3a == _T_37[9:0]) begin
        image_1_58 <= io_pixelVal_in_1_7;
      end else if (10'h3a == _T_34[9:0]) begin
        image_1_58 <= io_pixelVal_in_1_6;
      end else if (10'h3a == _T_31[9:0]) begin
        image_1_58 <= io_pixelVal_in_1_5;
      end else if (10'h3a == _T_28[9:0]) begin
        image_1_58 <= io_pixelVal_in_1_4;
      end else if (10'h3a == _T_25[9:0]) begin
        image_1_58 <= io_pixelVal_in_1_3;
      end else if (10'h3a == _T_22[9:0]) begin
        image_1_58 <= io_pixelVal_in_1_2;
      end else if (10'h3a == _T_19[9:0]) begin
        image_1_58 <= io_pixelVal_in_1_1;
      end else if (10'h3a == _T_15[9:0]) begin
        image_1_58 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_59 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3b == _T_37[9:0]) begin
        image_1_59 <= io_pixelVal_in_1_7;
      end else if (10'h3b == _T_34[9:0]) begin
        image_1_59 <= io_pixelVal_in_1_6;
      end else if (10'h3b == _T_31[9:0]) begin
        image_1_59 <= io_pixelVal_in_1_5;
      end else if (10'h3b == _T_28[9:0]) begin
        image_1_59 <= io_pixelVal_in_1_4;
      end else if (10'h3b == _T_25[9:0]) begin
        image_1_59 <= io_pixelVal_in_1_3;
      end else if (10'h3b == _T_22[9:0]) begin
        image_1_59 <= io_pixelVal_in_1_2;
      end else if (10'h3b == _T_19[9:0]) begin
        image_1_59 <= io_pixelVal_in_1_1;
      end else if (10'h3b == _T_15[9:0]) begin
        image_1_59 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_60 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3c == _T_37[9:0]) begin
        image_1_60 <= io_pixelVal_in_1_7;
      end else if (10'h3c == _T_34[9:0]) begin
        image_1_60 <= io_pixelVal_in_1_6;
      end else if (10'h3c == _T_31[9:0]) begin
        image_1_60 <= io_pixelVal_in_1_5;
      end else if (10'h3c == _T_28[9:0]) begin
        image_1_60 <= io_pixelVal_in_1_4;
      end else if (10'h3c == _T_25[9:0]) begin
        image_1_60 <= io_pixelVal_in_1_3;
      end else if (10'h3c == _T_22[9:0]) begin
        image_1_60 <= io_pixelVal_in_1_2;
      end else if (10'h3c == _T_19[9:0]) begin
        image_1_60 <= io_pixelVal_in_1_1;
      end else if (10'h3c == _T_15[9:0]) begin
        image_1_60 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_61 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3d == _T_37[9:0]) begin
        image_1_61 <= io_pixelVal_in_1_7;
      end else if (10'h3d == _T_34[9:0]) begin
        image_1_61 <= io_pixelVal_in_1_6;
      end else if (10'h3d == _T_31[9:0]) begin
        image_1_61 <= io_pixelVal_in_1_5;
      end else if (10'h3d == _T_28[9:0]) begin
        image_1_61 <= io_pixelVal_in_1_4;
      end else if (10'h3d == _T_25[9:0]) begin
        image_1_61 <= io_pixelVal_in_1_3;
      end else if (10'h3d == _T_22[9:0]) begin
        image_1_61 <= io_pixelVal_in_1_2;
      end else if (10'h3d == _T_19[9:0]) begin
        image_1_61 <= io_pixelVal_in_1_1;
      end else if (10'h3d == _T_15[9:0]) begin
        image_1_61 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_62 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3e == _T_37[9:0]) begin
        image_1_62 <= io_pixelVal_in_1_7;
      end else if (10'h3e == _T_34[9:0]) begin
        image_1_62 <= io_pixelVal_in_1_6;
      end else if (10'h3e == _T_31[9:0]) begin
        image_1_62 <= io_pixelVal_in_1_5;
      end else if (10'h3e == _T_28[9:0]) begin
        image_1_62 <= io_pixelVal_in_1_4;
      end else if (10'h3e == _T_25[9:0]) begin
        image_1_62 <= io_pixelVal_in_1_3;
      end else if (10'h3e == _T_22[9:0]) begin
        image_1_62 <= io_pixelVal_in_1_2;
      end else if (10'h3e == _T_19[9:0]) begin
        image_1_62 <= io_pixelVal_in_1_1;
      end else if (10'h3e == _T_15[9:0]) begin
        image_1_62 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_63 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3f == _T_37[9:0]) begin
        image_1_63 <= io_pixelVal_in_1_7;
      end else if (10'h3f == _T_34[9:0]) begin
        image_1_63 <= io_pixelVal_in_1_6;
      end else if (10'h3f == _T_31[9:0]) begin
        image_1_63 <= io_pixelVal_in_1_5;
      end else if (10'h3f == _T_28[9:0]) begin
        image_1_63 <= io_pixelVal_in_1_4;
      end else if (10'h3f == _T_25[9:0]) begin
        image_1_63 <= io_pixelVal_in_1_3;
      end else if (10'h3f == _T_22[9:0]) begin
        image_1_63 <= io_pixelVal_in_1_2;
      end else if (10'h3f == _T_19[9:0]) begin
        image_1_63 <= io_pixelVal_in_1_1;
      end else if (10'h3f == _T_15[9:0]) begin
        image_1_63 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_64 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h40 == _T_37[9:0]) begin
        image_1_64 <= io_pixelVal_in_1_7;
      end else if (10'h40 == _T_34[9:0]) begin
        image_1_64 <= io_pixelVal_in_1_6;
      end else if (10'h40 == _T_31[9:0]) begin
        image_1_64 <= io_pixelVal_in_1_5;
      end else if (10'h40 == _T_28[9:0]) begin
        image_1_64 <= io_pixelVal_in_1_4;
      end else if (10'h40 == _T_25[9:0]) begin
        image_1_64 <= io_pixelVal_in_1_3;
      end else if (10'h40 == _T_22[9:0]) begin
        image_1_64 <= io_pixelVal_in_1_2;
      end else if (10'h40 == _T_19[9:0]) begin
        image_1_64 <= io_pixelVal_in_1_1;
      end else if (10'h40 == _T_15[9:0]) begin
        image_1_64 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_65 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h41 == _T_37[9:0]) begin
        image_1_65 <= io_pixelVal_in_1_7;
      end else if (10'h41 == _T_34[9:0]) begin
        image_1_65 <= io_pixelVal_in_1_6;
      end else if (10'h41 == _T_31[9:0]) begin
        image_1_65 <= io_pixelVal_in_1_5;
      end else if (10'h41 == _T_28[9:0]) begin
        image_1_65 <= io_pixelVal_in_1_4;
      end else if (10'h41 == _T_25[9:0]) begin
        image_1_65 <= io_pixelVal_in_1_3;
      end else if (10'h41 == _T_22[9:0]) begin
        image_1_65 <= io_pixelVal_in_1_2;
      end else if (10'h41 == _T_19[9:0]) begin
        image_1_65 <= io_pixelVal_in_1_1;
      end else if (10'h41 == _T_15[9:0]) begin
        image_1_65 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_66 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h42 == _T_37[9:0]) begin
        image_1_66 <= io_pixelVal_in_1_7;
      end else if (10'h42 == _T_34[9:0]) begin
        image_1_66 <= io_pixelVal_in_1_6;
      end else if (10'h42 == _T_31[9:0]) begin
        image_1_66 <= io_pixelVal_in_1_5;
      end else if (10'h42 == _T_28[9:0]) begin
        image_1_66 <= io_pixelVal_in_1_4;
      end else if (10'h42 == _T_25[9:0]) begin
        image_1_66 <= io_pixelVal_in_1_3;
      end else if (10'h42 == _T_22[9:0]) begin
        image_1_66 <= io_pixelVal_in_1_2;
      end else if (10'h42 == _T_19[9:0]) begin
        image_1_66 <= io_pixelVal_in_1_1;
      end else if (10'h42 == _T_15[9:0]) begin
        image_1_66 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_67 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h43 == _T_37[9:0]) begin
        image_1_67 <= io_pixelVal_in_1_7;
      end else if (10'h43 == _T_34[9:0]) begin
        image_1_67 <= io_pixelVal_in_1_6;
      end else if (10'h43 == _T_31[9:0]) begin
        image_1_67 <= io_pixelVal_in_1_5;
      end else if (10'h43 == _T_28[9:0]) begin
        image_1_67 <= io_pixelVal_in_1_4;
      end else if (10'h43 == _T_25[9:0]) begin
        image_1_67 <= io_pixelVal_in_1_3;
      end else if (10'h43 == _T_22[9:0]) begin
        image_1_67 <= io_pixelVal_in_1_2;
      end else if (10'h43 == _T_19[9:0]) begin
        image_1_67 <= io_pixelVal_in_1_1;
      end else if (10'h43 == _T_15[9:0]) begin
        image_1_67 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_68 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h44 == _T_37[9:0]) begin
        image_1_68 <= io_pixelVal_in_1_7;
      end else if (10'h44 == _T_34[9:0]) begin
        image_1_68 <= io_pixelVal_in_1_6;
      end else if (10'h44 == _T_31[9:0]) begin
        image_1_68 <= io_pixelVal_in_1_5;
      end else if (10'h44 == _T_28[9:0]) begin
        image_1_68 <= io_pixelVal_in_1_4;
      end else if (10'h44 == _T_25[9:0]) begin
        image_1_68 <= io_pixelVal_in_1_3;
      end else if (10'h44 == _T_22[9:0]) begin
        image_1_68 <= io_pixelVal_in_1_2;
      end else if (10'h44 == _T_19[9:0]) begin
        image_1_68 <= io_pixelVal_in_1_1;
      end else if (10'h44 == _T_15[9:0]) begin
        image_1_68 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_69 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h45 == _T_37[9:0]) begin
        image_1_69 <= io_pixelVal_in_1_7;
      end else if (10'h45 == _T_34[9:0]) begin
        image_1_69 <= io_pixelVal_in_1_6;
      end else if (10'h45 == _T_31[9:0]) begin
        image_1_69 <= io_pixelVal_in_1_5;
      end else if (10'h45 == _T_28[9:0]) begin
        image_1_69 <= io_pixelVal_in_1_4;
      end else if (10'h45 == _T_25[9:0]) begin
        image_1_69 <= io_pixelVal_in_1_3;
      end else if (10'h45 == _T_22[9:0]) begin
        image_1_69 <= io_pixelVal_in_1_2;
      end else if (10'h45 == _T_19[9:0]) begin
        image_1_69 <= io_pixelVal_in_1_1;
      end else if (10'h45 == _T_15[9:0]) begin
        image_1_69 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_70 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h46 == _T_37[9:0]) begin
        image_1_70 <= io_pixelVal_in_1_7;
      end else if (10'h46 == _T_34[9:0]) begin
        image_1_70 <= io_pixelVal_in_1_6;
      end else if (10'h46 == _T_31[9:0]) begin
        image_1_70 <= io_pixelVal_in_1_5;
      end else if (10'h46 == _T_28[9:0]) begin
        image_1_70 <= io_pixelVal_in_1_4;
      end else if (10'h46 == _T_25[9:0]) begin
        image_1_70 <= io_pixelVal_in_1_3;
      end else if (10'h46 == _T_22[9:0]) begin
        image_1_70 <= io_pixelVal_in_1_2;
      end else if (10'h46 == _T_19[9:0]) begin
        image_1_70 <= io_pixelVal_in_1_1;
      end else if (10'h46 == _T_15[9:0]) begin
        image_1_70 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_71 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h47 == _T_37[9:0]) begin
        image_1_71 <= io_pixelVal_in_1_7;
      end else if (10'h47 == _T_34[9:0]) begin
        image_1_71 <= io_pixelVal_in_1_6;
      end else if (10'h47 == _T_31[9:0]) begin
        image_1_71 <= io_pixelVal_in_1_5;
      end else if (10'h47 == _T_28[9:0]) begin
        image_1_71 <= io_pixelVal_in_1_4;
      end else if (10'h47 == _T_25[9:0]) begin
        image_1_71 <= io_pixelVal_in_1_3;
      end else if (10'h47 == _T_22[9:0]) begin
        image_1_71 <= io_pixelVal_in_1_2;
      end else if (10'h47 == _T_19[9:0]) begin
        image_1_71 <= io_pixelVal_in_1_1;
      end else if (10'h47 == _T_15[9:0]) begin
        image_1_71 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_72 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h48 == _T_37[9:0]) begin
        image_1_72 <= io_pixelVal_in_1_7;
      end else if (10'h48 == _T_34[9:0]) begin
        image_1_72 <= io_pixelVal_in_1_6;
      end else if (10'h48 == _T_31[9:0]) begin
        image_1_72 <= io_pixelVal_in_1_5;
      end else if (10'h48 == _T_28[9:0]) begin
        image_1_72 <= io_pixelVal_in_1_4;
      end else if (10'h48 == _T_25[9:0]) begin
        image_1_72 <= io_pixelVal_in_1_3;
      end else if (10'h48 == _T_22[9:0]) begin
        image_1_72 <= io_pixelVal_in_1_2;
      end else if (10'h48 == _T_19[9:0]) begin
        image_1_72 <= io_pixelVal_in_1_1;
      end else if (10'h48 == _T_15[9:0]) begin
        image_1_72 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_73 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h49 == _T_37[9:0]) begin
        image_1_73 <= io_pixelVal_in_1_7;
      end else if (10'h49 == _T_34[9:0]) begin
        image_1_73 <= io_pixelVal_in_1_6;
      end else if (10'h49 == _T_31[9:0]) begin
        image_1_73 <= io_pixelVal_in_1_5;
      end else if (10'h49 == _T_28[9:0]) begin
        image_1_73 <= io_pixelVal_in_1_4;
      end else if (10'h49 == _T_25[9:0]) begin
        image_1_73 <= io_pixelVal_in_1_3;
      end else if (10'h49 == _T_22[9:0]) begin
        image_1_73 <= io_pixelVal_in_1_2;
      end else if (10'h49 == _T_19[9:0]) begin
        image_1_73 <= io_pixelVal_in_1_1;
      end else if (10'h49 == _T_15[9:0]) begin
        image_1_73 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_74 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4a == _T_37[9:0]) begin
        image_1_74 <= io_pixelVal_in_1_7;
      end else if (10'h4a == _T_34[9:0]) begin
        image_1_74 <= io_pixelVal_in_1_6;
      end else if (10'h4a == _T_31[9:0]) begin
        image_1_74 <= io_pixelVal_in_1_5;
      end else if (10'h4a == _T_28[9:0]) begin
        image_1_74 <= io_pixelVal_in_1_4;
      end else if (10'h4a == _T_25[9:0]) begin
        image_1_74 <= io_pixelVal_in_1_3;
      end else if (10'h4a == _T_22[9:0]) begin
        image_1_74 <= io_pixelVal_in_1_2;
      end else if (10'h4a == _T_19[9:0]) begin
        image_1_74 <= io_pixelVal_in_1_1;
      end else if (10'h4a == _T_15[9:0]) begin
        image_1_74 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_75 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4b == _T_37[9:0]) begin
        image_1_75 <= io_pixelVal_in_1_7;
      end else if (10'h4b == _T_34[9:0]) begin
        image_1_75 <= io_pixelVal_in_1_6;
      end else if (10'h4b == _T_31[9:0]) begin
        image_1_75 <= io_pixelVal_in_1_5;
      end else if (10'h4b == _T_28[9:0]) begin
        image_1_75 <= io_pixelVal_in_1_4;
      end else if (10'h4b == _T_25[9:0]) begin
        image_1_75 <= io_pixelVal_in_1_3;
      end else if (10'h4b == _T_22[9:0]) begin
        image_1_75 <= io_pixelVal_in_1_2;
      end else if (10'h4b == _T_19[9:0]) begin
        image_1_75 <= io_pixelVal_in_1_1;
      end else if (10'h4b == _T_15[9:0]) begin
        image_1_75 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_76 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4c == _T_37[9:0]) begin
        image_1_76 <= io_pixelVal_in_1_7;
      end else if (10'h4c == _T_34[9:0]) begin
        image_1_76 <= io_pixelVal_in_1_6;
      end else if (10'h4c == _T_31[9:0]) begin
        image_1_76 <= io_pixelVal_in_1_5;
      end else if (10'h4c == _T_28[9:0]) begin
        image_1_76 <= io_pixelVal_in_1_4;
      end else if (10'h4c == _T_25[9:0]) begin
        image_1_76 <= io_pixelVal_in_1_3;
      end else if (10'h4c == _T_22[9:0]) begin
        image_1_76 <= io_pixelVal_in_1_2;
      end else if (10'h4c == _T_19[9:0]) begin
        image_1_76 <= io_pixelVal_in_1_1;
      end else if (10'h4c == _T_15[9:0]) begin
        image_1_76 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_77 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4d == _T_37[9:0]) begin
        image_1_77 <= io_pixelVal_in_1_7;
      end else if (10'h4d == _T_34[9:0]) begin
        image_1_77 <= io_pixelVal_in_1_6;
      end else if (10'h4d == _T_31[9:0]) begin
        image_1_77 <= io_pixelVal_in_1_5;
      end else if (10'h4d == _T_28[9:0]) begin
        image_1_77 <= io_pixelVal_in_1_4;
      end else if (10'h4d == _T_25[9:0]) begin
        image_1_77 <= io_pixelVal_in_1_3;
      end else if (10'h4d == _T_22[9:0]) begin
        image_1_77 <= io_pixelVal_in_1_2;
      end else if (10'h4d == _T_19[9:0]) begin
        image_1_77 <= io_pixelVal_in_1_1;
      end else if (10'h4d == _T_15[9:0]) begin
        image_1_77 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_78 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4e == _T_37[9:0]) begin
        image_1_78 <= io_pixelVal_in_1_7;
      end else if (10'h4e == _T_34[9:0]) begin
        image_1_78 <= io_pixelVal_in_1_6;
      end else if (10'h4e == _T_31[9:0]) begin
        image_1_78 <= io_pixelVal_in_1_5;
      end else if (10'h4e == _T_28[9:0]) begin
        image_1_78 <= io_pixelVal_in_1_4;
      end else if (10'h4e == _T_25[9:0]) begin
        image_1_78 <= io_pixelVal_in_1_3;
      end else if (10'h4e == _T_22[9:0]) begin
        image_1_78 <= io_pixelVal_in_1_2;
      end else if (10'h4e == _T_19[9:0]) begin
        image_1_78 <= io_pixelVal_in_1_1;
      end else if (10'h4e == _T_15[9:0]) begin
        image_1_78 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_79 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4f == _T_37[9:0]) begin
        image_1_79 <= io_pixelVal_in_1_7;
      end else if (10'h4f == _T_34[9:0]) begin
        image_1_79 <= io_pixelVal_in_1_6;
      end else if (10'h4f == _T_31[9:0]) begin
        image_1_79 <= io_pixelVal_in_1_5;
      end else if (10'h4f == _T_28[9:0]) begin
        image_1_79 <= io_pixelVal_in_1_4;
      end else if (10'h4f == _T_25[9:0]) begin
        image_1_79 <= io_pixelVal_in_1_3;
      end else if (10'h4f == _T_22[9:0]) begin
        image_1_79 <= io_pixelVal_in_1_2;
      end else if (10'h4f == _T_19[9:0]) begin
        image_1_79 <= io_pixelVal_in_1_1;
      end else if (10'h4f == _T_15[9:0]) begin
        image_1_79 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_80 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h50 == _T_37[9:0]) begin
        image_1_80 <= io_pixelVal_in_1_7;
      end else if (10'h50 == _T_34[9:0]) begin
        image_1_80 <= io_pixelVal_in_1_6;
      end else if (10'h50 == _T_31[9:0]) begin
        image_1_80 <= io_pixelVal_in_1_5;
      end else if (10'h50 == _T_28[9:0]) begin
        image_1_80 <= io_pixelVal_in_1_4;
      end else if (10'h50 == _T_25[9:0]) begin
        image_1_80 <= io_pixelVal_in_1_3;
      end else if (10'h50 == _T_22[9:0]) begin
        image_1_80 <= io_pixelVal_in_1_2;
      end else if (10'h50 == _T_19[9:0]) begin
        image_1_80 <= io_pixelVal_in_1_1;
      end else if (10'h50 == _T_15[9:0]) begin
        image_1_80 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_81 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h51 == _T_37[9:0]) begin
        image_1_81 <= io_pixelVal_in_1_7;
      end else if (10'h51 == _T_34[9:0]) begin
        image_1_81 <= io_pixelVal_in_1_6;
      end else if (10'h51 == _T_31[9:0]) begin
        image_1_81 <= io_pixelVal_in_1_5;
      end else if (10'h51 == _T_28[9:0]) begin
        image_1_81 <= io_pixelVal_in_1_4;
      end else if (10'h51 == _T_25[9:0]) begin
        image_1_81 <= io_pixelVal_in_1_3;
      end else if (10'h51 == _T_22[9:0]) begin
        image_1_81 <= io_pixelVal_in_1_2;
      end else if (10'h51 == _T_19[9:0]) begin
        image_1_81 <= io_pixelVal_in_1_1;
      end else if (10'h51 == _T_15[9:0]) begin
        image_1_81 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_82 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h52 == _T_37[9:0]) begin
        image_1_82 <= io_pixelVal_in_1_7;
      end else if (10'h52 == _T_34[9:0]) begin
        image_1_82 <= io_pixelVal_in_1_6;
      end else if (10'h52 == _T_31[9:0]) begin
        image_1_82 <= io_pixelVal_in_1_5;
      end else if (10'h52 == _T_28[9:0]) begin
        image_1_82 <= io_pixelVal_in_1_4;
      end else if (10'h52 == _T_25[9:0]) begin
        image_1_82 <= io_pixelVal_in_1_3;
      end else if (10'h52 == _T_22[9:0]) begin
        image_1_82 <= io_pixelVal_in_1_2;
      end else if (10'h52 == _T_19[9:0]) begin
        image_1_82 <= io_pixelVal_in_1_1;
      end else if (10'h52 == _T_15[9:0]) begin
        image_1_82 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_83 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h53 == _T_37[9:0]) begin
        image_1_83 <= io_pixelVal_in_1_7;
      end else if (10'h53 == _T_34[9:0]) begin
        image_1_83 <= io_pixelVal_in_1_6;
      end else if (10'h53 == _T_31[9:0]) begin
        image_1_83 <= io_pixelVal_in_1_5;
      end else if (10'h53 == _T_28[9:0]) begin
        image_1_83 <= io_pixelVal_in_1_4;
      end else if (10'h53 == _T_25[9:0]) begin
        image_1_83 <= io_pixelVal_in_1_3;
      end else if (10'h53 == _T_22[9:0]) begin
        image_1_83 <= io_pixelVal_in_1_2;
      end else if (10'h53 == _T_19[9:0]) begin
        image_1_83 <= io_pixelVal_in_1_1;
      end else if (10'h53 == _T_15[9:0]) begin
        image_1_83 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_84 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h54 == _T_37[9:0]) begin
        image_1_84 <= io_pixelVal_in_1_7;
      end else if (10'h54 == _T_34[9:0]) begin
        image_1_84 <= io_pixelVal_in_1_6;
      end else if (10'h54 == _T_31[9:0]) begin
        image_1_84 <= io_pixelVal_in_1_5;
      end else if (10'h54 == _T_28[9:0]) begin
        image_1_84 <= io_pixelVal_in_1_4;
      end else if (10'h54 == _T_25[9:0]) begin
        image_1_84 <= io_pixelVal_in_1_3;
      end else if (10'h54 == _T_22[9:0]) begin
        image_1_84 <= io_pixelVal_in_1_2;
      end else if (10'h54 == _T_19[9:0]) begin
        image_1_84 <= io_pixelVal_in_1_1;
      end else if (10'h54 == _T_15[9:0]) begin
        image_1_84 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_85 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h55 == _T_37[9:0]) begin
        image_1_85 <= io_pixelVal_in_1_7;
      end else if (10'h55 == _T_34[9:0]) begin
        image_1_85 <= io_pixelVal_in_1_6;
      end else if (10'h55 == _T_31[9:0]) begin
        image_1_85 <= io_pixelVal_in_1_5;
      end else if (10'h55 == _T_28[9:0]) begin
        image_1_85 <= io_pixelVal_in_1_4;
      end else if (10'h55 == _T_25[9:0]) begin
        image_1_85 <= io_pixelVal_in_1_3;
      end else if (10'h55 == _T_22[9:0]) begin
        image_1_85 <= io_pixelVal_in_1_2;
      end else if (10'h55 == _T_19[9:0]) begin
        image_1_85 <= io_pixelVal_in_1_1;
      end else if (10'h55 == _T_15[9:0]) begin
        image_1_85 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_86 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h56 == _T_37[9:0]) begin
        image_1_86 <= io_pixelVal_in_1_7;
      end else if (10'h56 == _T_34[9:0]) begin
        image_1_86 <= io_pixelVal_in_1_6;
      end else if (10'h56 == _T_31[9:0]) begin
        image_1_86 <= io_pixelVal_in_1_5;
      end else if (10'h56 == _T_28[9:0]) begin
        image_1_86 <= io_pixelVal_in_1_4;
      end else if (10'h56 == _T_25[9:0]) begin
        image_1_86 <= io_pixelVal_in_1_3;
      end else if (10'h56 == _T_22[9:0]) begin
        image_1_86 <= io_pixelVal_in_1_2;
      end else if (10'h56 == _T_19[9:0]) begin
        image_1_86 <= io_pixelVal_in_1_1;
      end else if (10'h56 == _T_15[9:0]) begin
        image_1_86 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_87 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h57 == _T_37[9:0]) begin
        image_1_87 <= io_pixelVal_in_1_7;
      end else if (10'h57 == _T_34[9:0]) begin
        image_1_87 <= io_pixelVal_in_1_6;
      end else if (10'h57 == _T_31[9:0]) begin
        image_1_87 <= io_pixelVal_in_1_5;
      end else if (10'h57 == _T_28[9:0]) begin
        image_1_87 <= io_pixelVal_in_1_4;
      end else if (10'h57 == _T_25[9:0]) begin
        image_1_87 <= io_pixelVal_in_1_3;
      end else if (10'h57 == _T_22[9:0]) begin
        image_1_87 <= io_pixelVal_in_1_2;
      end else if (10'h57 == _T_19[9:0]) begin
        image_1_87 <= io_pixelVal_in_1_1;
      end else if (10'h57 == _T_15[9:0]) begin
        image_1_87 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_88 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h58 == _T_37[9:0]) begin
        image_1_88 <= io_pixelVal_in_1_7;
      end else if (10'h58 == _T_34[9:0]) begin
        image_1_88 <= io_pixelVal_in_1_6;
      end else if (10'h58 == _T_31[9:0]) begin
        image_1_88 <= io_pixelVal_in_1_5;
      end else if (10'h58 == _T_28[9:0]) begin
        image_1_88 <= io_pixelVal_in_1_4;
      end else if (10'h58 == _T_25[9:0]) begin
        image_1_88 <= io_pixelVal_in_1_3;
      end else if (10'h58 == _T_22[9:0]) begin
        image_1_88 <= io_pixelVal_in_1_2;
      end else if (10'h58 == _T_19[9:0]) begin
        image_1_88 <= io_pixelVal_in_1_1;
      end else if (10'h58 == _T_15[9:0]) begin
        image_1_88 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_89 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h59 == _T_37[9:0]) begin
        image_1_89 <= io_pixelVal_in_1_7;
      end else if (10'h59 == _T_34[9:0]) begin
        image_1_89 <= io_pixelVal_in_1_6;
      end else if (10'h59 == _T_31[9:0]) begin
        image_1_89 <= io_pixelVal_in_1_5;
      end else if (10'h59 == _T_28[9:0]) begin
        image_1_89 <= io_pixelVal_in_1_4;
      end else if (10'h59 == _T_25[9:0]) begin
        image_1_89 <= io_pixelVal_in_1_3;
      end else if (10'h59 == _T_22[9:0]) begin
        image_1_89 <= io_pixelVal_in_1_2;
      end else if (10'h59 == _T_19[9:0]) begin
        image_1_89 <= io_pixelVal_in_1_1;
      end else if (10'h59 == _T_15[9:0]) begin
        image_1_89 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_90 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5a == _T_37[9:0]) begin
        image_1_90 <= io_pixelVal_in_1_7;
      end else if (10'h5a == _T_34[9:0]) begin
        image_1_90 <= io_pixelVal_in_1_6;
      end else if (10'h5a == _T_31[9:0]) begin
        image_1_90 <= io_pixelVal_in_1_5;
      end else if (10'h5a == _T_28[9:0]) begin
        image_1_90 <= io_pixelVal_in_1_4;
      end else if (10'h5a == _T_25[9:0]) begin
        image_1_90 <= io_pixelVal_in_1_3;
      end else if (10'h5a == _T_22[9:0]) begin
        image_1_90 <= io_pixelVal_in_1_2;
      end else if (10'h5a == _T_19[9:0]) begin
        image_1_90 <= io_pixelVal_in_1_1;
      end else if (10'h5a == _T_15[9:0]) begin
        image_1_90 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_91 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5b == _T_37[9:0]) begin
        image_1_91 <= io_pixelVal_in_1_7;
      end else if (10'h5b == _T_34[9:0]) begin
        image_1_91 <= io_pixelVal_in_1_6;
      end else if (10'h5b == _T_31[9:0]) begin
        image_1_91 <= io_pixelVal_in_1_5;
      end else if (10'h5b == _T_28[9:0]) begin
        image_1_91 <= io_pixelVal_in_1_4;
      end else if (10'h5b == _T_25[9:0]) begin
        image_1_91 <= io_pixelVal_in_1_3;
      end else if (10'h5b == _T_22[9:0]) begin
        image_1_91 <= io_pixelVal_in_1_2;
      end else if (10'h5b == _T_19[9:0]) begin
        image_1_91 <= io_pixelVal_in_1_1;
      end else if (10'h5b == _T_15[9:0]) begin
        image_1_91 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_92 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5c == _T_37[9:0]) begin
        image_1_92 <= io_pixelVal_in_1_7;
      end else if (10'h5c == _T_34[9:0]) begin
        image_1_92 <= io_pixelVal_in_1_6;
      end else if (10'h5c == _T_31[9:0]) begin
        image_1_92 <= io_pixelVal_in_1_5;
      end else if (10'h5c == _T_28[9:0]) begin
        image_1_92 <= io_pixelVal_in_1_4;
      end else if (10'h5c == _T_25[9:0]) begin
        image_1_92 <= io_pixelVal_in_1_3;
      end else if (10'h5c == _T_22[9:0]) begin
        image_1_92 <= io_pixelVal_in_1_2;
      end else if (10'h5c == _T_19[9:0]) begin
        image_1_92 <= io_pixelVal_in_1_1;
      end else if (10'h5c == _T_15[9:0]) begin
        image_1_92 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_93 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5d == _T_37[9:0]) begin
        image_1_93 <= io_pixelVal_in_1_7;
      end else if (10'h5d == _T_34[9:0]) begin
        image_1_93 <= io_pixelVal_in_1_6;
      end else if (10'h5d == _T_31[9:0]) begin
        image_1_93 <= io_pixelVal_in_1_5;
      end else if (10'h5d == _T_28[9:0]) begin
        image_1_93 <= io_pixelVal_in_1_4;
      end else if (10'h5d == _T_25[9:0]) begin
        image_1_93 <= io_pixelVal_in_1_3;
      end else if (10'h5d == _T_22[9:0]) begin
        image_1_93 <= io_pixelVal_in_1_2;
      end else if (10'h5d == _T_19[9:0]) begin
        image_1_93 <= io_pixelVal_in_1_1;
      end else if (10'h5d == _T_15[9:0]) begin
        image_1_93 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_94 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5e == _T_37[9:0]) begin
        image_1_94 <= io_pixelVal_in_1_7;
      end else if (10'h5e == _T_34[9:0]) begin
        image_1_94 <= io_pixelVal_in_1_6;
      end else if (10'h5e == _T_31[9:0]) begin
        image_1_94 <= io_pixelVal_in_1_5;
      end else if (10'h5e == _T_28[9:0]) begin
        image_1_94 <= io_pixelVal_in_1_4;
      end else if (10'h5e == _T_25[9:0]) begin
        image_1_94 <= io_pixelVal_in_1_3;
      end else if (10'h5e == _T_22[9:0]) begin
        image_1_94 <= io_pixelVal_in_1_2;
      end else if (10'h5e == _T_19[9:0]) begin
        image_1_94 <= io_pixelVal_in_1_1;
      end else if (10'h5e == _T_15[9:0]) begin
        image_1_94 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_95 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5f == _T_37[9:0]) begin
        image_1_95 <= io_pixelVal_in_1_7;
      end else if (10'h5f == _T_34[9:0]) begin
        image_1_95 <= io_pixelVal_in_1_6;
      end else if (10'h5f == _T_31[9:0]) begin
        image_1_95 <= io_pixelVal_in_1_5;
      end else if (10'h5f == _T_28[9:0]) begin
        image_1_95 <= io_pixelVal_in_1_4;
      end else if (10'h5f == _T_25[9:0]) begin
        image_1_95 <= io_pixelVal_in_1_3;
      end else if (10'h5f == _T_22[9:0]) begin
        image_1_95 <= io_pixelVal_in_1_2;
      end else if (10'h5f == _T_19[9:0]) begin
        image_1_95 <= io_pixelVal_in_1_1;
      end else if (10'h5f == _T_15[9:0]) begin
        image_1_95 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_96 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h60 == _T_37[9:0]) begin
        image_1_96 <= io_pixelVal_in_1_7;
      end else if (10'h60 == _T_34[9:0]) begin
        image_1_96 <= io_pixelVal_in_1_6;
      end else if (10'h60 == _T_31[9:0]) begin
        image_1_96 <= io_pixelVal_in_1_5;
      end else if (10'h60 == _T_28[9:0]) begin
        image_1_96 <= io_pixelVal_in_1_4;
      end else if (10'h60 == _T_25[9:0]) begin
        image_1_96 <= io_pixelVal_in_1_3;
      end else if (10'h60 == _T_22[9:0]) begin
        image_1_96 <= io_pixelVal_in_1_2;
      end else if (10'h60 == _T_19[9:0]) begin
        image_1_96 <= io_pixelVal_in_1_1;
      end else if (10'h60 == _T_15[9:0]) begin
        image_1_96 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_97 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h61 == _T_37[9:0]) begin
        image_1_97 <= io_pixelVal_in_1_7;
      end else if (10'h61 == _T_34[9:0]) begin
        image_1_97 <= io_pixelVal_in_1_6;
      end else if (10'h61 == _T_31[9:0]) begin
        image_1_97 <= io_pixelVal_in_1_5;
      end else if (10'h61 == _T_28[9:0]) begin
        image_1_97 <= io_pixelVal_in_1_4;
      end else if (10'h61 == _T_25[9:0]) begin
        image_1_97 <= io_pixelVal_in_1_3;
      end else if (10'h61 == _T_22[9:0]) begin
        image_1_97 <= io_pixelVal_in_1_2;
      end else if (10'h61 == _T_19[9:0]) begin
        image_1_97 <= io_pixelVal_in_1_1;
      end else if (10'h61 == _T_15[9:0]) begin
        image_1_97 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_98 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h62 == _T_37[9:0]) begin
        image_1_98 <= io_pixelVal_in_1_7;
      end else if (10'h62 == _T_34[9:0]) begin
        image_1_98 <= io_pixelVal_in_1_6;
      end else if (10'h62 == _T_31[9:0]) begin
        image_1_98 <= io_pixelVal_in_1_5;
      end else if (10'h62 == _T_28[9:0]) begin
        image_1_98 <= io_pixelVal_in_1_4;
      end else if (10'h62 == _T_25[9:0]) begin
        image_1_98 <= io_pixelVal_in_1_3;
      end else if (10'h62 == _T_22[9:0]) begin
        image_1_98 <= io_pixelVal_in_1_2;
      end else if (10'h62 == _T_19[9:0]) begin
        image_1_98 <= io_pixelVal_in_1_1;
      end else if (10'h62 == _T_15[9:0]) begin
        image_1_98 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_99 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h63 == _T_37[9:0]) begin
        image_1_99 <= io_pixelVal_in_1_7;
      end else if (10'h63 == _T_34[9:0]) begin
        image_1_99 <= io_pixelVal_in_1_6;
      end else if (10'h63 == _T_31[9:0]) begin
        image_1_99 <= io_pixelVal_in_1_5;
      end else if (10'h63 == _T_28[9:0]) begin
        image_1_99 <= io_pixelVal_in_1_4;
      end else if (10'h63 == _T_25[9:0]) begin
        image_1_99 <= io_pixelVal_in_1_3;
      end else if (10'h63 == _T_22[9:0]) begin
        image_1_99 <= io_pixelVal_in_1_2;
      end else if (10'h63 == _T_19[9:0]) begin
        image_1_99 <= io_pixelVal_in_1_1;
      end else if (10'h63 == _T_15[9:0]) begin
        image_1_99 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_100 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h64 == _T_37[9:0]) begin
        image_1_100 <= io_pixelVal_in_1_7;
      end else if (10'h64 == _T_34[9:0]) begin
        image_1_100 <= io_pixelVal_in_1_6;
      end else if (10'h64 == _T_31[9:0]) begin
        image_1_100 <= io_pixelVal_in_1_5;
      end else if (10'h64 == _T_28[9:0]) begin
        image_1_100 <= io_pixelVal_in_1_4;
      end else if (10'h64 == _T_25[9:0]) begin
        image_1_100 <= io_pixelVal_in_1_3;
      end else if (10'h64 == _T_22[9:0]) begin
        image_1_100 <= io_pixelVal_in_1_2;
      end else if (10'h64 == _T_19[9:0]) begin
        image_1_100 <= io_pixelVal_in_1_1;
      end else if (10'h64 == _T_15[9:0]) begin
        image_1_100 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_101 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h65 == _T_37[9:0]) begin
        image_1_101 <= io_pixelVal_in_1_7;
      end else if (10'h65 == _T_34[9:0]) begin
        image_1_101 <= io_pixelVal_in_1_6;
      end else if (10'h65 == _T_31[9:0]) begin
        image_1_101 <= io_pixelVal_in_1_5;
      end else if (10'h65 == _T_28[9:0]) begin
        image_1_101 <= io_pixelVal_in_1_4;
      end else if (10'h65 == _T_25[9:0]) begin
        image_1_101 <= io_pixelVal_in_1_3;
      end else if (10'h65 == _T_22[9:0]) begin
        image_1_101 <= io_pixelVal_in_1_2;
      end else if (10'h65 == _T_19[9:0]) begin
        image_1_101 <= io_pixelVal_in_1_1;
      end else if (10'h65 == _T_15[9:0]) begin
        image_1_101 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_102 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h66 == _T_37[9:0]) begin
        image_1_102 <= io_pixelVal_in_1_7;
      end else if (10'h66 == _T_34[9:0]) begin
        image_1_102 <= io_pixelVal_in_1_6;
      end else if (10'h66 == _T_31[9:0]) begin
        image_1_102 <= io_pixelVal_in_1_5;
      end else if (10'h66 == _T_28[9:0]) begin
        image_1_102 <= io_pixelVal_in_1_4;
      end else if (10'h66 == _T_25[9:0]) begin
        image_1_102 <= io_pixelVal_in_1_3;
      end else if (10'h66 == _T_22[9:0]) begin
        image_1_102 <= io_pixelVal_in_1_2;
      end else if (10'h66 == _T_19[9:0]) begin
        image_1_102 <= io_pixelVal_in_1_1;
      end else if (10'h66 == _T_15[9:0]) begin
        image_1_102 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_103 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h67 == _T_37[9:0]) begin
        image_1_103 <= io_pixelVal_in_1_7;
      end else if (10'h67 == _T_34[9:0]) begin
        image_1_103 <= io_pixelVal_in_1_6;
      end else if (10'h67 == _T_31[9:0]) begin
        image_1_103 <= io_pixelVal_in_1_5;
      end else if (10'h67 == _T_28[9:0]) begin
        image_1_103 <= io_pixelVal_in_1_4;
      end else if (10'h67 == _T_25[9:0]) begin
        image_1_103 <= io_pixelVal_in_1_3;
      end else if (10'h67 == _T_22[9:0]) begin
        image_1_103 <= io_pixelVal_in_1_2;
      end else if (10'h67 == _T_19[9:0]) begin
        image_1_103 <= io_pixelVal_in_1_1;
      end else if (10'h67 == _T_15[9:0]) begin
        image_1_103 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_104 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h68 == _T_37[9:0]) begin
        image_1_104 <= io_pixelVal_in_1_7;
      end else if (10'h68 == _T_34[9:0]) begin
        image_1_104 <= io_pixelVal_in_1_6;
      end else if (10'h68 == _T_31[9:0]) begin
        image_1_104 <= io_pixelVal_in_1_5;
      end else if (10'h68 == _T_28[9:0]) begin
        image_1_104 <= io_pixelVal_in_1_4;
      end else if (10'h68 == _T_25[9:0]) begin
        image_1_104 <= io_pixelVal_in_1_3;
      end else if (10'h68 == _T_22[9:0]) begin
        image_1_104 <= io_pixelVal_in_1_2;
      end else if (10'h68 == _T_19[9:0]) begin
        image_1_104 <= io_pixelVal_in_1_1;
      end else if (10'h68 == _T_15[9:0]) begin
        image_1_104 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_105 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h69 == _T_37[9:0]) begin
        image_1_105 <= io_pixelVal_in_1_7;
      end else if (10'h69 == _T_34[9:0]) begin
        image_1_105 <= io_pixelVal_in_1_6;
      end else if (10'h69 == _T_31[9:0]) begin
        image_1_105 <= io_pixelVal_in_1_5;
      end else if (10'h69 == _T_28[9:0]) begin
        image_1_105 <= io_pixelVal_in_1_4;
      end else if (10'h69 == _T_25[9:0]) begin
        image_1_105 <= io_pixelVal_in_1_3;
      end else if (10'h69 == _T_22[9:0]) begin
        image_1_105 <= io_pixelVal_in_1_2;
      end else if (10'h69 == _T_19[9:0]) begin
        image_1_105 <= io_pixelVal_in_1_1;
      end else if (10'h69 == _T_15[9:0]) begin
        image_1_105 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_106 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6a == _T_37[9:0]) begin
        image_1_106 <= io_pixelVal_in_1_7;
      end else if (10'h6a == _T_34[9:0]) begin
        image_1_106 <= io_pixelVal_in_1_6;
      end else if (10'h6a == _T_31[9:0]) begin
        image_1_106 <= io_pixelVal_in_1_5;
      end else if (10'h6a == _T_28[9:0]) begin
        image_1_106 <= io_pixelVal_in_1_4;
      end else if (10'h6a == _T_25[9:0]) begin
        image_1_106 <= io_pixelVal_in_1_3;
      end else if (10'h6a == _T_22[9:0]) begin
        image_1_106 <= io_pixelVal_in_1_2;
      end else if (10'h6a == _T_19[9:0]) begin
        image_1_106 <= io_pixelVal_in_1_1;
      end else if (10'h6a == _T_15[9:0]) begin
        image_1_106 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_107 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6b == _T_37[9:0]) begin
        image_1_107 <= io_pixelVal_in_1_7;
      end else if (10'h6b == _T_34[9:0]) begin
        image_1_107 <= io_pixelVal_in_1_6;
      end else if (10'h6b == _T_31[9:0]) begin
        image_1_107 <= io_pixelVal_in_1_5;
      end else if (10'h6b == _T_28[9:0]) begin
        image_1_107 <= io_pixelVal_in_1_4;
      end else if (10'h6b == _T_25[9:0]) begin
        image_1_107 <= io_pixelVal_in_1_3;
      end else if (10'h6b == _T_22[9:0]) begin
        image_1_107 <= io_pixelVal_in_1_2;
      end else if (10'h6b == _T_19[9:0]) begin
        image_1_107 <= io_pixelVal_in_1_1;
      end else if (10'h6b == _T_15[9:0]) begin
        image_1_107 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_108 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6c == _T_37[9:0]) begin
        image_1_108 <= io_pixelVal_in_1_7;
      end else if (10'h6c == _T_34[9:0]) begin
        image_1_108 <= io_pixelVal_in_1_6;
      end else if (10'h6c == _T_31[9:0]) begin
        image_1_108 <= io_pixelVal_in_1_5;
      end else if (10'h6c == _T_28[9:0]) begin
        image_1_108 <= io_pixelVal_in_1_4;
      end else if (10'h6c == _T_25[9:0]) begin
        image_1_108 <= io_pixelVal_in_1_3;
      end else if (10'h6c == _T_22[9:0]) begin
        image_1_108 <= io_pixelVal_in_1_2;
      end else if (10'h6c == _T_19[9:0]) begin
        image_1_108 <= io_pixelVal_in_1_1;
      end else if (10'h6c == _T_15[9:0]) begin
        image_1_108 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_109 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6d == _T_37[9:0]) begin
        image_1_109 <= io_pixelVal_in_1_7;
      end else if (10'h6d == _T_34[9:0]) begin
        image_1_109 <= io_pixelVal_in_1_6;
      end else if (10'h6d == _T_31[9:0]) begin
        image_1_109 <= io_pixelVal_in_1_5;
      end else if (10'h6d == _T_28[9:0]) begin
        image_1_109 <= io_pixelVal_in_1_4;
      end else if (10'h6d == _T_25[9:0]) begin
        image_1_109 <= io_pixelVal_in_1_3;
      end else if (10'h6d == _T_22[9:0]) begin
        image_1_109 <= io_pixelVal_in_1_2;
      end else if (10'h6d == _T_19[9:0]) begin
        image_1_109 <= io_pixelVal_in_1_1;
      end else if (10'h6d == _T_15[9:0]) begin
        image_1_109 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_110 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6e == _T_37[9:0]) begin
        image_1_110 <= io_pixelVal_in_1_7;
      end else if (10'h6e == _T_34[9:0]) begin
        image_1_110 <= io_pixelVal_in_1_6;
      end else if (10'h6e == _T_31[9:0]) begin
        image_1_110 <= io_pixelVal_in_1_5;
      end else if (10'h6e == _T_28[9:0]) begin
        image_1_110 <= io_pixelVal_in_1_4;
      end else if (10'h6e == _T_25[9:0]) begin
        image_1_110 <= io_pixelVal_in_1_3;
      end else if (10'h6e == _T_22[9:0]) begin
        image_1_110 <= io_pixelVal_in_1_2;
      end else if (10'h6e == _T_19[9:0]) begin
        image_1_110 <= io_pixelVal_in_1_1;
      end else if (10'h6e == _T_15[9:0]) begin
        image_1_110 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_111 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6f == _T_37[9:0]) begin
        image_1_111 <= io_pixelVal_in_1_7;
      end else if (10'h6f == _T_34[9:0]) begin
        image_1_111 <= io_pixelVal_in_1_6;
      end else if (10'h6f == _T_31[9:0]) begin
        image_1_111 <= io_pixelVal_in_1_5;
      end else if (10'h6f == _T_28[9:0]) begin
        image_1_111 <= io_pixelVal_in_1_4;
      end else if (10'h6f == _T_25[9:0]) begin
        image_1_111 <= io_pixelVal_in_1_3;
      end else if (10'h6f == _T_22[9:0]) begin
        image_1_111 <= io_pixelVal_in_1_2;
      end else if (10'h6f == _T_19[9:0]) begin
        image_1_111 <= io_pixelVal_in_1_1;
      end else if (10'h6f == _T_15[9:0]) begin
        image_1_111 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_112 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h70 == _T_37[9:0]) begin
        image_1_112 <= io_pixelVal_in_1_7;
      end else if (10'h70 == _T_34[9:0]) begin
        image_1_112 <= io_pixelVal_in_1_6;
      end else if (10'h70 == _T_31[9:0]) begin
        image_1_112 <= io_pixelVal_in_1_5;
      end else if (10'h70 == _T_28[9:0]) begin
        image_1_112 <= io_pixelVal_in_1_4;
      end else if (10'h70 == _T_25[9:0]) begin
        image_1_112 <= io_pixelVal_in_1_3;
      end else if (10'h70 == _T_22[9:0]) begin
        image_1_112 <= io_pixelVal_in_1_2;
      end else if (10'h70 == _T_19[9:0]) begin
        image_1_112 <= io_pixelVal_in_1_1;
      end else if (10'h70 == _T_15[9:0]) begin
        image_1_112 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_113 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h71 == _T_37[9:0]) begin
        image_1_113 <= io_pixelVal_in_1_7;
      end else if (10'h71 == _T_34[9:0]) begin
        image_1_113 <= io_pixelVal_in_1_6;
      end else if (10'h71 == _T_31[9:0]) begin
        image_1_113 <= io_pixelVal_in_1_5;
      end else if (10'h71 == _T_28[9:0]) begin
        image_1_113 <= io_pixelVal_in_1_4;
      end else if (10'h71 == _T_25[9:0]) begin
        image_1_113 <= io_pixelVal_in_1_3;
      end else if (10'h71 == _T_22[9:0]) begin
        image_1_113 <= io_pixelVal_in_1_2;
      end else if (10'h71 == _T_19[9:0]) begin
        image_1_113 <= io_pixelVal_in_1_1;
      end else if (10'h71 == _T_15[9:0]) begin
        image_1_113 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_114 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h72 == _T_37[9:0]) begin
        image_1_114 <= io_pixelVal_in_1_7;
      end else if (10'h72 == _T_34[9:0]) begin
        image_1_114 <= io_pixelVal_in_1_6;
      end else if (10'h72 == _T_31[9:0]) begin
        image_1_114 <= io_pixelVal_in_1_5;
      end else if (10'h72 == _T_28[9:0]) begin
        image_1_114 <= io_pixelVal_in_1_4;
      end else if (10'h72 == _T_25[9:0]) begin
        image_1_114 <= io_pixelVal_in_1_3;
      end else if (10'h72 == _T_22[9:0]) begin
        image_1_114 <= io_pixelVal_in_1_2;
      end else if (10'h72 == _T_19[9:0]) begin
        image_1_114 <= io_pixelVal_in_1_1;
      end else if (10'h72 == _T_15[9:0]) begin
        image_1_114 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_115 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h73 == _T_37[9:0]) begin
        image_1_115 <= io_pixelVal_in_1_7;
      end else if (10'h73 == _T_34[9:0]) begin
        image_1_115 <= io_pixelVal_in_1_6;
      end else if (10'h73 == _T_31[9:0]) begin
        image_1_115 <= io_pixelVal_in_1_5;
      end else if (10'h73 == _T_28[9:0]) begin
        image_1_115 <= io_pixelVal_in_1_4;
      end else if (10'h73 == _T_25[9:0]) begin
        image_1_115 <= io_pixelVal_in_1_3;
      end else if (10'h73 == _T_22[9:0]) begin
        image_1_115 <= io_pixelVal_in_1_2;
      end else if (10'h73 == _T_19[9:0]) begin
        image_1_115 <= io_pixelVal_in_1_1;
      end else if (10'h73 == _T_15[9:0]) begin
        image_1_115 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_116 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h74 == _T_37[9:0]) begin
        image_1_116 <= io_pixelVal_in_1_7;
      end else if (10'h74 == _T_34[9:0]) begin
        image_1_116 <= io_pixelVal_in_1_6;
      end else if (10'h74 == _T_31[9:0]) begin
        image_1_116 <= io_pixelVal_in_1_5;
      end else if (10'h74 == _T_28[9:0]) begin
        image_1_116 <= io_pixelVal_in_1_4;
      end else if (10'h74 == _T_25[9:0]) begin
        image_1_116 <= io_pixelVal_in_1_3;
      end else if (10'h74 == _T_22[9:0]) begin
        image_1_116 <= io_pixelVal_in_1_2;
      end else if (10'h74 == _T_19[9:0]) begin
        image_1_116 <= io_pixelVal_in_1_1;
      end else if (10'h74 == _T_15[9:0]) begin
        image_1_116 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_117 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h75 == _T_37[9:0]) begin
        image_1_117 <= io_pixelVal_in_1_7;
      end else if (10'h75 == _T_34[9:0]) begin
        image_1_117 <= io_pixelVal_in_1_6;
      end else if (10'h75 == _T_31[9:0]) begin
        image_1_117 <= io_pixelVal_in_1_5;
      end else if (10'h75 == _T_28[9:0]) begin
        image_1_117 <= io_pixelVal_in_1_4;
      end else if (10'h75 == _T_25[9:0]) begin
        image_1_117 <= io_pixelVal_in_1_3;
      end else if (10'h75 == _T_22[9:0]) begin
        image_1_117 <= io_pixelVal_in_1_2;
      end else if (10'h75 == _T_19[9:0]) begin
        image_1_117 <= io_pixelVal_in_1_1;
      end else if (10'h75 == _T_15[9:0]) begin
        image_1_117 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_118 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h76 == _T_37[9:0]) begin
        image_1_118 <= io_pixelVal_in_1_7;
      end else if (10'h76 == _T_34[9:0]) begin
        image_1_118 <= io_pixelVal_in_1_6;
      end else if (10'h76 == _T_31[9:0]) begin
        image_1_118 <= io_pixelVal_in_1_5;
      end else if (10'h76 == _T_28[9:0]) begin
        image_1_118 <= io_pixelVal_in_1_4;
      end else if (10'h76 == _T_25[9:0]) begin
        image_1_118 <= io_pixelVal_in_1_3;
      end else if (10'h76 == _T_22[9:0]) begin
        image_1_118 <= io_pixelVal_in_1_2;
      end else if (10'h76 == _T_19[9:0]) begin
        image_1_118 <= io_pixelVal_in_1_1;
      end else if (10'h76 == _T_15[9:0]) begin
        image_1_118 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_119 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h77 == _T_37[9:0]) begin
        image_1_119 <= io_pixelVal_in_1_7;
      end else if (10'h77 == _T_34[9:0]) begin
        image_1_119 <= io_pixelVal_in_1_6;
      end else if (10'h77 == _T_31[9:0]) begin
        image_1_119 <= io_pixelVal_in_1_5;
      end else if (10'h77 == _T_28[9:0]) begin
        image_1_119 <= io_pixelVal_in_1_4;
      end else if (10'h77 == _T_25[9:0]) begin
        image_1_119 <= io_pixelVal_in_1_3;
      end else if (10'h77 == _T_22[9:0]) begin
        image_1_119 <= io_pixelVal_in_1_2;
      end else if (10'h77 == _T_19[9:0]) begin
        image_1_119 <= io_pixelVal_in_1_1;
      end else if (10'h77 == _T_15[9:0]) begin
        image_1_119 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_120 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h78 == _T_37[9:0]) begin
        image_1_120 <= io_pixelVal_in_1_7;
      end else if (10'h78 == _T_34[9:0]) begin
        image_1_120 <= io_pixelVal_in_1_6;
      end else if (10'h78 == _T_31[9:0]) begin
        image_1_120 <= io_pixelVal_in_1_5;
      end else if (10'h78 == _T_28[9:0]) begin
        image_1_120 <= io_pixelVal_in_1_4;
      end else if (10'h78 == _T_25[9:0]) begin
        image_1_120 <= io_pixelVal_in_1_3;
      end else if (10'h78 == _T_22[9:0]) begin
        image_1_120 <= io_pixelVal_in_1_2;
      end else if (10'h78 == _T_19[9:0]) begin
        image_1_120 <= io_pixelVal_in_1_1;
      end else if (10'h78 == _T_15[9:0]) begin
        image_1_120 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_121 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h79 == _T_37[9:0]) begin
        image_1_121 <= io_pixelVal_in_1_7;
      end else if (10'h79 == _T_34[9:0]) begin
        image_1_121 <= io_pixelVal_in_1_6;
      end else if (10'h79 == _T_31[9:0]) begin
        image_1_121 <= io_pixelVal_in_1_5;
      end else if (10'h79 == _T_28[9:0]) begin
        image_1_121 <= io_pixelVal_in_1_4;
      end else if (10'h79 == _T_25[9:0]) begin
        image_1_121 <= io_pixelVal_in_1_3;
      end else if (10'h79 == _T_22[9:0]) begin
        image_1_121 <= io_pixelVal_in_1_2;
      end else if (10'h79 == _T_19[9:0]) begin
        image_1_121 <= io_pixelVal_in_1_1;
      end else if (10'h79 == _T_15[9:0]) begin
        image_1_121 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_122 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7a == _T_37[9:0]) begin
        image_1_122 <= io_pixelVal_in_1_7;
      end else if (10'h7a == _T_34[9:0]) begin
        image_1_122 <= io_pixelVal_in_1_6;
      end else if (10'h7a == _T_31[9:0]) begin
        image_1_122 <= io_pixelVal_in_1_5;
      end else if (10'h7a == _T_28[9:0]) begin
        image_1_122 <= io_pixelVal_in_1_4;
      end else if (10'h7a == _T_25[9:0]) begin
        image_1_122 <= io_pixelVal_in_1_3;
      end else if (10'h7a == _T_22[9:0]) begin
        image_1_122 <= io_pixelVal_in_1_2;
      end else if (10'h7a == _T_19[9:0]) begin
        image_1_122 <= io_pixelVal_in_1_1;
      end else if (10'h7a == _T_15[9:0]) begin
        image_1_122 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_123 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7b == _T_37[9:0]) begin
        image_1_123 <= io_pixelVal_in_1_7;
      end else if (10'h7b == _T_34[9:0]) begin
        image_1_123 <= io_pixelVal_in_1_6;
      end else if (10'h7b == _T_31[9:0]) begin
        image_1_123 <= io_pixelVal_in_1_5;
      end else if (10'h7b == _T_28[9:0]) begin
        image_1_123 <= io_pixelVal_in_1_4;
      end else if (10'h7b == _T_25[9:0]) begin
        image_1_123 <= io_pixelVal_in_1_3;
      end else if (10'h7b == _T_22[9:0]) begin
        image_1_123 <= io_pixelVal_in_1_2;
      end else if (10'h7b == _T_19[9:0]) begin
        image_1_123 <= io_pixelVal_in_1_1;
      end else if (10'h7b == _T_15[9:0]) begin
        image_1_123 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_124 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7c == _T_37[9:0]) begin
        image_1_124 <= io_pixelVal_in_1_7;
      end else if (10'h7c == _T_34[9:0]) begin
        image_1_124 <= io_pixelVal_in_1_6;
      end else if (10'h7c == _T_31[9:0]) begin
        image_1_124 <= io_pixelVal_in_1_5;
      end else if (10'h7c == _T_28[9:0]) begin
        image_1_124 <= io_pixelVal_in_1_4;
      end else if (10'h7c == _T_25[9:0]) begin
        image_1_124 <= io_pixelVal_in_1_3;
      end else if (10'h7c == _T_22[9:0]) begin
        image_1_124 <= io_pixelVal_in_1_2;
      end else if (10'h7c == _T_19[9:0]) begin
        image_1_124 <= io_pixelVal_in_1_1;
      end else if (10'h7c == _T_15[9:0]) begin
        image_1_124 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_125 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7d == _T_37[9:0]) begin
        image_1_125 <= io_pixelVal_in_1_7;
      end else if (10'h7d == _T_34[9:0]) begin
        image_1_125 <= io_pixelVal_in_1_6;
      end else if (10'h7d == _T_31[9:0]) begin
        image_1_125 <= io_pixelVal_in_1_5;
      end else if (10'h7d == _T_28[9:0]) begin
        image_1_125 <= io_pixelVal_in_1_4;
      end else if (10'h7d == _T_25[9:0]) begin
        image_1_125 <= io_pixelVal_in_1_3;
      end else if (10'h7d == _T_22[9:0]) begin
        image_1_125 <= io_pixelVal_in_1_2;
      end else if (10'h7d == _T_19[9:0]) begin
        image_1_125 <= io_pixelVal_in_1_1;
      end else if (10'h7d == _T_15[9:0]) begin
        image_1_125 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_126 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7e == _T_37[9:0]) begin
        image_1_126 <= io_pixelVal_in_1_7;
      end else if (10'h7e == _T_34[9:0]) begin
        image_1_126 <= io_pixelVal_in_1_6;
      end else if (10'h7e == _T_31[9:0]) begin
        image_1_126 <= io_pixelVal_in_1_5;
      end else if (10'h7e == _T_28[9:0]) begin
        image_1_126 <= io_pixelVal_in_1_4;
      end else if (10'h7e == _T_25[9:0]) begin
        image_1_126 <= io_pixelVal_in_1_3;
      end else if (10'h7e == _T_22[9:0]) begin
        image_1_126 <= io_pixelVal_in_1_2;
      end else if (10'h7e == _T_19[9:0]) begin
        image_1_126 <= io_pixelVal_in_1_1;
      end else if (10'h7e == _T_15[9:0]) begin
        image_1_126 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_127 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7f == _T_37[9:0]) begin
        image_1_127 <= io_pixelVal_in_1_7;
      end else if (10'h7f == _T_34[9:0]) begin
        image_1_127 <= io_pixelVal_in_1_6;
      end else if (10'h7f == _T_31[9:0]) begin
        image_1_127 <= io_pixelVal_in_1_5;
      end else if (10'h7f == _T_28[9:0]) begin
        image_1_127 <= io_pixelVal_in_1_4;
      end else if (10'h7f == _T_25[9:0]) begin
        image_1_127 <= io_pixelVal_in_1_3;
      end else if (10'h7f == _T_22[9:0]) begin
        image_1_127 <= io_pixelVal_in_1_2;
      end else if (10'h7f == _T_19[9:0]) begin
        image_1_127 <= io_pixelVal_in_1_1;
      end else if (10'h7f == _T_15[9:0]) begin
        image_1_127 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_128 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h80 == _T_37[9:0]) begin
        image_1_128 <= io_pixelVal_in_1_7;
      end else if (10'h80 == _T_34[9:0]) begin
        image_1_128 <= io_pixelVal_in_1_6;
      end else if (10'h80 == _T_31[9:0]) begin
        image_1_128 <= io_pixelVal_in_1_5;
      end else if (10'h80 == _T_28[9:0]) begin
        image_1_128 <= io_pixelVal_in_1_4;
      end else if (10'h80 == _T_25[9:0]) begin
        image_1_128 <= io_pixelVal_in_1_3;
      end else if (10'h80 == _T_22[9:0]) begin
        image_1_128 <= io_pixelVal_in_1_2;
      end else if (10'h80 == _T_19[9:0]) begin
        image_1_128 <= io_pixelVal_in_1_1;
      end else if (10'h80 == _T_15[9:0]) begin
        image_1_128 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_129 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h81 == _T_37[9:0]) begin
        image_1_129 <= io_pixelVal_in_1_7;
      end else if (10'h81 == _T_34[9:0]) begin
        image_1_129 <= io_pixelVal_in_1_6;
      end else if (10'h81 == _T_31[9:0]) begin
        image_1_129 <= io_pixelVal_in_1_5;
      end else if (10'h81 == _T_28[9:0]) begin
        image_1_129 <= io_pixelVal_in_1_4;
      end else if (10'h81 == _T_25[9:0]) begin
        image_1_129 <= io_pixelVal_in_1_3;
      end else if (10'h81 == _T_22[9:0]) begin
        image_1_129 <= io_pixelVal_in_1_2;
      end else if (10'h81 == _T_19[9:0]) begin
        image_1_129 <= io_pixelVal_in_1_1;
      end else if (10'h81 == _T_15[9:0]) begin
        image_1_129 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_130 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h82 == _T_37[9:0]) begin
        image_1_130 <= io_pixelVal_in_1_7;
      end else if (10'h82 == _T_34[9:0]) begin
        image_1_130 <= io_pixelVal_in_1_6;
      end else if (10'h82 == _T_31[9:0]) begin
        image_1_130 <= io_pixelVal_in_1_5;
      end else if (10'h82 == _T_28[9:0]) begin
        image_1_130 <= io_pixelVal_in_1_4;
      end else if (10'h82 == _T_25[9:0]) begin
        image_1_130 <= io_pixelVal_in_1_3;
      end else if (10'h82 == _T_22[9:0]) begin
        image_1_130 <= io_pixelVal_in_1_2;
      end else if (10'h82 == _T_19[9:0]) begin
        image_1_130 <= io_pixelVal_in_1_1;
      end else if (10'h82 == _T_15[9:0]) begin
        image_1_130 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_131 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h83 == _T_37[9:0]) begin
        image_1_131 <= io_pixelVal_in_1_7;
      end else if (10'h83 == _T_34[9:0]) begin
        image_1_131 <= io_pixelVal_in_1_6;
      end else if (10'h83 == _T_31[9:0]) begin
        image_1_131 <= io_pixelVal_in_1_5;
      end else if (10'h83 == _T_28[9:0]) begin
        image_1_131 <= io_pixelVal_in_1_4;
      end else if (10'h83 == _T_25[9:0]) begin
        image_1_131 <= io_pixelVal_in_1_3;
      end else if (10'h83 == _T_22[9:0]) begin
        image_1_131 <= io_pixelVal_in_1_2;
      end else if (10'h83 == _T_19[9:0]) begin
        image_1_131 <= io_pixelVal_in_1_1;
      end else if (10'h83 == _T_15[9:0]) begin
        image_1_131 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_132 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h84 == _T_37[9:0]) begin
        image_1_132 <= io_pixelVal_in_1_7;
      end else if (10'h84 == _T_34[9:0]) begin
        image_1_132 <= io_pixelVal_in_1_6;
      end else if (10'h84 == _T_31[9:0]) begin
        image_1_132 <= io_pixelVal_in_1_5;
      end else if (10'h84 == _T_28[9:0]) begin
        image_1_132 <= io_pixelVal_in_1_4;
      end else if (10'h84 == _T_25[9:0]) begin
        image_1_132 <= io_pixelVal_in_1_3;
      end else if (10'h84 == _T_22[9:0]) begin
        image_1_132 <= io_pixelVal_in_1_2;
      end else if (10'h84 == _T_19[9:0]) begin
        image_1_132 <= io_pixelVal_in_1_1;
      end else if (10'h84 == _T_15[9:0]) begin
        image_1_132 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_133 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h85 == _T_37[9:0]) begin
        image_1_133 <= io_pixelVal_in_1_7;
      end else if (10'h85 == _T_34[9:0]) begin
        image_1_133 <= io_pixelVal_in_1_6;
      end else if (10'h85 == _T_31[9:0]) begin
        image_1_133 <= io_pixelVal_in_1_5;
      end else if (10'h85 == _T_28[9:0]) begin
        image_1_133 <= io_pixelVal_in_1_4;
      end else if (10'h85 == _T_25[9:0]) begin
        image_1_133 <= io_pixelVal_in_1_3;
      end else if (10'h85 == _T_22[9:0]) begin
        image_1_133 <= io_pixelVal_in_1_2;
      end else if (10'h85 == _T_19[9:0]) begin
        image_1_133 <= io_pixelVal_in_1_1;
      end else if (10'h85 == _T_15[9:0]) begin
        image_1_133 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_134 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h86 == _T_37[9:0]) begin
        image_1_134 <= io_pixelVal_in_1_7;
      end else if (10'h86 == _T_34[9:0]) begin
        image_1_134 <= io_pixelVal_in_1_6;
      end else if (10'h86 == _T_31[9:0]) begin
        image_1_134 <= io_pixelVal_in_1_5;
      end else if (10'h86 == _T_28[9:0]) begin
        image_1_134 <= io_pixelVal_in_1_4;
      end else if (10'h86 == _T_25[9:0]) begin
        image_1_134 <= io_pixelVal_in_1_3;
      end else if (10'h86 == _T_22[9:0]) begin
        image_1_134 <= io_pixelVal_in_1_2;
      end else if (10'h86 == _T_19[9:0]) begin
        image_1_134 <= io_pixelVal_in_1_1;
      end else if (10'h86 == _T_15[9:0]) begin
        image_1_134 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_135 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h87 == _T_37[9:0]) begin
        image_1_135 <= io_pixelVal_in_1_7;
      end else if (10'h87 == _T_34[9:0]) begin
        image_1_135 <= io_pixelVal_in_1_6;
      end else if (10'h87 == _T_31[9:0]) begin
        image_1_135 <= io_pixelVal_in_1_5;
      end else if (10'h87 == _T_28[9:0]) begin
        image_1_135 <= io_pixelVal_in_1_4;
      end else if (10'h87 == _T_25[9:0]) begin
        image_1_135 <= io_pixelVal_in_1_3;
      end else if (10'h87 == _T_22[9:0]) begin
        image_1_135 <= io_pixelVal_in_1_2;
      end else if (10'h87 == _T_19[9:0]) begin
        image_1_135 <= io_pixelVal_in_1_1;
      end else if (10'h87 == _T_15[9:0]) begin
        image_1_135 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_136 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h88 == _T_37[9:0]) begin
        image_1_136 <= io_pixelVal_in_1_7;
      end else if (10'h88 == _T_34[9:0]) begin
        image_1_136 <= io_pixelVal_in_1_6;
      end else if (10'h88 == _T_31[9:0]) begin
        image_1_136 <= io_pixelVal_in_1_5;
      end else if (10'h88 == _T_28[9:0]) begin
        image_1_136 <= io_pixelVal_in_1_4;
      end else if (10'h88 == _T_25[9:0]) begin
        image_1_136 <= io_pixelVal_in_1_3;
      end else if (10'h88 == _T_22[9:0]) begin
        image_1_136 <= io_pixelVal_in_1_2;
      end else if (10'h88 == _T_19[9:0]) begin
        image_1_136 <= io_pixelVal_in_1_1;
      end else if (10'h88 == _T_15[9:0]) begin
        image_1_136 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_137 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h89 == _T_37[9:0]) begin
        image_1_137 <= io_pixelVal_in_1_7;
      end else if (10'h89 == _T_34[9:0]) begin
        image_1_137 <= io_pixelVal_in_1_6;
      end else if (10'h89 == _T_31[9:0]) begin
        image_1_137 <= io_pixelVal_in_1_5;
      end else if (10'h89 == _T_28[9:0]) begin
        image_1_137 <= io_pixelVal_in_1_4;
      end else if (10'h89 == _T_25[9:0]) begin
        image_1_137 <= io_pixelVal_in_1_3;
      end else if (10'h89 == _T_22[9:0]) begin
        image_1_137 <= io_pixelVal_in_1_2;
      end else if (10'h89 == _T_19[9:0]) begin
        image_1_137 <= io_pixelVal_in_1_1;
      end else if (10'h89 == _T_15[9:0]) begin
        image_1_137 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_138 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8a == _T_37[9:0]) begin
        image_1_138 <= io_pixelVal_in_1_7;
      end else if (10'h8a == _T_34[9:0]) begin
        image_1_138 <= io_pixelVal_in_1_6;
      end else if (10'h8a == _T_31[9:0]) begin
        image_1_138 <= io_pixelVal_in_1_5;
      end else if (10'h8a == _T_28[9:0]) begin
        image_1_138 <= io_pixelVal_in_1_4;
      end else if (10'h8a == _T_25[9:0]) begin
        image_1_138 <= io_pixelVal_in_1_3;
      end else if (10'h8a == _T_22[9:0]) begin
        image_1_138 <= io_pixelVal_in_1_2;
      end else if (10'h8a == _T_19[9:0]) begin
        image_1_138 <= io_pixelVal_in_1_1;
      end else if (10'h8a == _T_15[9:0]) begin
        image_1_138 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_139 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8b == _T_37[9:0]) begin
        image_1_139 <= io_pixelVal_in_1_7;
      end else if (10'h8b == _T_34[9:0]) begin
        image_1_139 <= io_pixelVal_in_1_6;
      end else if (10'h8b == _T_31[9:0]) begin
        image_1_139 <= io_pixelVal_in_1_5;
      end else if (10'h8b == _T_28[9:0]) begin
        image_1_139 <= io_pixelVal_in_1_4;
      end else if (10'h8b == _T_25[9:0]) begin
        image_1_139 <= io_pixelVal_in_1_3;
      end else if (10'h8b == _T_22[9:0]) begin
        image_1_139 <= io_pixelVal_in_1_2;
      end else if (10'h8b == _T_19[9:0]) begin
        image_1_139 <= io_pixelVal_in_1_1;
      end else if (10'h8b == _T_15[9:0]) begin
        image_1_139 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_140 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8c == _T_37[9:0]) begin
        image_1_140 <= io_pixelVal_in_1_7;
      end else if (10'h8c == _T_34[9:0]) begin
        image_1_140 <= io_pixelVal_in_1_6;
      end else if (10'h8c == _T_31[9:0]) begin
        image_1_140 <= io_pixelVal_in_1_5;
      end else if (10'h8c == _T_28[9:0]) begin
        image_1_140 <= io_pixelVal_in_1_4;
      end else if (10'h8c == _T_25[9:0]) begin
        image_1_140 <= io_pixelVal_in_1_3;
      end else if (10'h8c == _T_22[9:0]) begin
        image_1_140 <= io_pixelVal_in_1_2;
      end else if (10'h8c == _T_19[9:0]) begin
        image_1_140 <= io_pixelVal_in_1_1;
      end else if (10'h8c == _T_15[9:0]) begin
        image_1_140 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_141 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8d == _T_37[9:0]) begin
        image_1_141 <= io_pixelVal_in_1_7;
      end else if (10'h8d == _T_34[9:0]) begin
        image_1_141 <= io_pixelVal_in_1_6;
      end else if (10'h8d == _T_31[9:0]) begin
        image_1_141 <= io_pixelVal_in_1_5;
      end else if (10'h8d == _T_28[9:0]) begin
        image_1_141 <= io_pixelVal_in_1_4;
      end else if (10'h8d == _T_25[9:0]) begin
        image_1_141 <= io_pixelVal_in_1_3;
      end else if (10'h8d == _T_22[9:0]) begin
        image_1_141 <= io_pixelVal_in_1_2;
      end else if (10'h8d == _T_19[9:0]) begin
        image_1_141 <= io_pixelVal_in_1_1;
      end else if (10'h8d == _T_15[9:0]) begin
        image_1_141 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_142 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8e == _T_37[9:0]) begin
        image_1_142 <= io_pixelVal_in_1_7;
      end else if (10'h8e == _T_34[9:0]) begin
        image_1_142 <= io_pixelVal_in_1_6;
      end else if (10'h8e == _T_31[9:0]) begin
        image_1_142 <= io_pixelVal_in_1_5;
      end else if (10'h8e == _T_28[9:0]) begin
        image_1_142 <= io_pixelVal_in_1_4;
      end else if (10'h8e == _T_25[9:0]) begin
        image_1_142 <= io_pixelVal_in_1_3;
      end else if (10'h8e == _T_22[9:0]) begin
        image_1_142 <= io_pixelVal_in_1_2;
      end else if (10'h8e == _T_19[9:0]) begin
        image_1_142 <= io_pixelVal_in_1_1;
      end else if (10'h8e == _T_15[9:0]) begin
        image_1_142 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_143 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8f == _T_37[9:0]) begin
        image_1_143 <= io_pixelVal_in_1_7;
      end else if (10'h8f == _T_34[9:0]) begin
        image_1_143 <= io_pixelVal_in_1_6;
      end else if (10'h8f == _T_31[9:0]) begin
        image_1_143 <= io_pixelVal_in_1_5;
      end else if (10'h8f == _T_28[9:0]) begin
        image_1_143 <= io_pixelVal_in_1_4;
      end else if (10'h8f == _T_25[9:0]) begin
        image_1_143 <= io_pixelVal_in_1_3;
      end else if (10'h8f == _T_22[9:0]) begin
        image_1_143 <= io_pixelVal_in_1_2;
      end else if (10'h8f == _T_19[9:0]) begin
        image_1_143 <= io_pixelVal_in_1_1;
      end else if (10'h8f == _T_15[9:0]) begin
        image_1_143 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_144 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h90 == _T_37[9:0]) begin
        image_1_144 <= io_pixelVal_in_1_7;
      end else if (10'h90 == _T_34[9:0]) begin
        image_1_144 <= io_pixelVal_in_1_6;
      end else if (10'h90 == _T_31[9:0]) begin
        image_1_144 <= io_pixelVal_in_1_5;
      end else if (10'h90 == _T_28[9:0]) begin
        image_1_144 <= io_pixelVal_in_1_4;
      end else if (10'h90 == _T_25[9:0]) begin
        image_1_144 <= io_pixelVal_in_1_3;
      end else if (10'h90 == _T_22[9:0]) begin
        image_1_144 <= io_pixelVal_in_1_2;
      end else if (10'h90 == _T_19[9:0]) begin
        image_1_144 <= io_pixelVal_in_1_1;
      end else if (10'h90 == _T_15[9:0]) begin
        image_1_144 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_145 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h91 == _T_37[9:0]) begin
        image_1_145 <= io_pixelVal_in_1_7;
      end else if (10'h91 == _T_34[9:0]) begin
        image_1_145 <= io_pixelVal_in_1_6;
      end else if (10'h91 == _T_31[9:0]) begin
        image_1_145 <= io_pixelVal_in_1_5;
      end else if (10'h91 == _T_28[9:0]) begin
        image_1_145 <= io_pixelVal_in_1_4;
      end else if (10'h91 == _T_25[9:0]) begin
        image_1_145 <= io_pixelVal_in_1_3;
      end else if (10'h91 == _T_22[9:0]) begin
        image_1_145 <= io_pixelVal_in_1_2;
      end else if (10'h91 == _T_19[9:0]) begin
        image_1_145 <= io_pixelVal_in_1_1;
      end else if (10'h91 == _T_15[9:0]) begin
        image_1_145 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_146 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h92 == _T_37[9:0]) begin
        image_1_146 <= io_pixelVal_in_1_7;
      end else if (10'h92 == _T_34[9:0]) begin
        image_1_146 <= io_pixelVal_in_1_6;
      end else if (10'h92 == _T_31[9:0]) begin
        image_1_146 <= io_pixelVal_in_1_5;
      end else if (10'h92 == _T_28[9:0]) begin
        image_1_146 <= io_pixelVal_in_1_4;
      end else if (10'h92 == _T_25[9:0]) begin
        image_1_146 <= io_pixelVal_in_1_3;
      end else if (10'h92 == _T_22[9:0]) begin
        image_1_146 <= io_pixelVal_in_1_2;
      end else if (10'h92 == _T_19[9:0]) begin
        image_1_146 <= io_pixelVal_in_1_1;
      end else if (10'h92 == _T_15[9:0]) begin
        image_1_146 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_147 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h93 == _T_37[9:0]) begin
        image_1_147 <= io_pixelVal_in_1_7;
      end else if (10'h93 == _T_34[9:0]) begin
        image_1_147 <= io_pixelVal_in_1_6;
      end else if (10'h93 == _T_31[9:0]) begin
        image_1_147 <= io_pixelVal_in_1_5;
      end else if (10'h93 == _T_28[9:0]) begin
        image_1_147 <= io_pixelVal_in_1_4;
      end else if (10'h93 == _T_25[9:0]) begin
        image_1_147 <= io_pixelVal_in_1_3;
      end else if (10'h93 == _T_22[9:0]) begin
        image_1_147 <= io_pixelVal_in_1_2;
      end else if (10'h93 == _T_19[9:0]) begin
        image_1_147 <= io_pixelVal_in_1_1;
      end else if (10'h93 == _T_15[9:0]) begin
        image_1_147 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_148 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h94 == _T_37[9:0]) begin
        image_1_148 <= io_pixelVal_in_1_7;
      end else if (10'h94 == _T_34[9:0]) begin
        image_1_148 <= io_pixelVal_in_1_6;
      end else if (10'h94 == _T_31[9:0]) begin
        image_1_148 <= io_pixelVal_in_1_5;
      end else if (10'h94 == _T_28[9:0]) begin
        image_1_148 <= io_pixelVal_in_1_4;
      end else if (10'h94 == _T_25[9:0]) begin
        image_1_148 <= io_pixelVal_in_1_3;
      end else if (10'h94 == _T_22[9:0]) begin
        image_1_148 <= io_pixelVal_in_1_2;
      end else if (10'h94 == _T_19[9:0]) begin
        image_1_148 <= io_pixelVal_in_1_1;
      end else if (10'h94 == _T_15[9:0]) begin
        image_1_148 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_149 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h95 == _T_37[9:0]) begin
        image_1_149 <= io_pixelVal_in_1_7;
      end else if (10'h95 == _T_34[9:0]) begin
        image_1_149 <= io_pixelVal_in_1_6;
      end else if (10'h95 == _T_31[9:0]) begin
        image_1_149 <= io_pixelVal_in_1_5;
      end else if (10'h95 == _T_28[9:0]) begin
        image_1_149 <= io_pixelVal_in_1_4;
      end else if (10'h95 == _T_25[9:0]) begin
        image_1_149 <= io_pixelVal_in_1_3;
      end else if (10'h95 == _T_22[9:0]) begin
        image_1_149 <= io_pixelVal_in_1_2;
      end else if (10'h95 == _T_19[9:0]) begin
        image_1_149 <= io_pixelVal_in_1_1;
      end else if (10'h95 == _T_15[9:0]) begin
        image_1_149 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_150 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h96 == _T_37[9:0]) begin
        image_1_150 <= io_pixelVal_in_1_7;
      end else if (10'h96 == _T_34[9:0]) begin
        image_1_150 <= io_pixelVal_in_1_6;
      end else if (10'h96 == _T_31[9:0]) begin
        image_1_150 <= io_pixelVal_in_1_5;
      end else if (10'h96 == _T_28[9:0]) begin
        image_1_150 <= io_pixelVal_in_1_4;
      end else if (10'h96 == _T_25[9:0]) begin
        image_1_150 <= io_pixelVal_in_1_3;
      end else if (10'h96 == _T_22[9:0]) begin
        image_1_150 <= io_pixelVal_in_1_2;
      end else if (10'h96 == _T_19[9:0]) begin
        image_1_150 <= io_pixelVal_in_1_1;
      end else if (10'h96 == _T_15[9:0]) begin
        image_1_150 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_151 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h97 == _T_37[9:0]) begin
        image_1_151 <= io_pixelVal_in_1_7;
      end else if (10'h97 == _T_34[9:0]) begin
        image_1_151 <= io_pixelVal_in_1_6;
      end else if (10'h97 == _T_31[9:0]) begin
        image_1_151 <= io_pixelVal_in_1_5;
      end else if (10'h97 == _T_28[9:0]) begin
        image_1_151 <= io_pixelVal_in_1_4;
      end else if (10'h97 == _T_25[9:0]) begin
        image_1_151 <= io_pixelVal_in_1_3;
      end else if (10'h97 == _T_22[9:0]) begin
        image_1_151 <= io_pixelVal_in_1_2;
      end else if (10'h97 == _T_19[9:0]) begin
        image_1_151 <= io_pixelVal_in_1_1;
      end else if (10'h97 == _T_15[9:0]) begin
        image_1_151 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_152 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h98 == _T_37[9:0]) begin
        image_1_152 <= io_pixelVal_in_1_7;
      end else if (10'h98 == _T_34[9:0]) begin
        image_1_152 <= io_pixelVal_in_1_6;
      end else if (10'h98 == _T_31[9:0]) begin
        image_1_152 <= io_pixelVal_in_1_5;
      end else if (10'h98 == _T_28[9:0]) begin
        image_1_152 <= io_pixelVal_in_1_4;
      end else if (10'h98 == _T_25[9:0]) begin
        image_1_152 <= io_pixelVal_in_1_3;
      end else if (10'h98 == _T_22[9:0]) begin
        image_1_152 <= io_pixelVal_in_1_2;
      end else if (10'h98 == _T_19[9:0]) begin
        image_1_152 <= io_pixelVal_in_1_1;
      end else if (10'h98 == _T_15[9:0]) begin
        image_1_152 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_153 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h99 == _T_37[9:0]) begin
        image_1_153 <= io_pixelVal_in_1_7;
      end else if (10'h99 == _T_34[9:0]) begin
        image_1_153 <= io_pixelVal_in_1_6;
      end else if (10'h99 == _T_31[9:0]) begin
        image_1_153 <= io_pixelVal_in_1_5;
      end else if (10'h99 == _T_28[9:0]) begin
        image_1_153 <= io_pixelVal_in_1_4;
      end else if (10'h99 == _T_25[9:0]) begin
        image_1_153 <= io_pixelVal_in_1_3;
      end else if (10'h99 == _T_22[9:0]) begin
        image_1_153 <= io_pixelVal_in_1_2;
      end else if (10'h99 == _T_19[9:0]) begin
        image_1_153 <= io_pixelVal_in_1_1;
      end else if (10'h99 == _T_15[9:0]) begin
        image_1_153 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_154 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9a == _T_37[9:0]) begin
        image_1_154 <= io_pixelVal_in_1_7;
      end else if (10'h9a == _T_34[9:0]) begin
        image_1_154 <= io_pixelVal_in_1_6;
      end else if (10'h9a == _T_31[9:0]) begin
        image_1_154 <= io_pixelVal_in_1_5;
      end else if (10'h9a == _T_28[9:0]) begin
        image_1_154 <= io_pixelVal_in_1_4;
      end else if (10'h9a == _T_25[9:0]) begin
        image_1_154 <= io_pixelVal_in_1_3;
      end else if (10'h9a == _T_22[9:0]) begin
        image_1_154 <= io_pixelVal_in_1_2;
      end else if (10'h9a == _T_19[9:0]) begin
        image_1_154 <= io_pixelVal_in_1_1;
      end else if (10'h9a == _T_15[9:0]) begin
        image_1_154 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_155 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9b == _T_37[9:0]) begin
        image_1_155 <= io_pixelVal_in_1_7;
      end else if (10'h9b == _T_34[9:0]) begin
        image_1_155 <= io_pixelVal_in_1_6;
      end else if (10'h9b == _T_31[9:0]) begin
        image_1_155 <= io_pixelVal_in_1_5;
      end else if (10'h9b == _T_28[9:0]) begin
        image_1_155 <= io_pixelVal_in_1_4;
      end else if (10'h9b == _T_25[9:0]) begin
        image_1_155 <= io_pixelVal_in_1_3;
      end else if (10'h9b == _T_22[9:0]) begin
        image_1_155 <= io_pixelVal_in_1_2;
      end else if (10'h9b == _T_19[9:0]) begin
        image_1_155 <= io_pixelVal_in_1_1;
      end else if (10'h9b == _T_15[9:0]) begin
        image_1_155 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_156 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9c == _T_37[9:0]) begin
        image_1_156 <= io_pixelVal_in_1_7;
      end else if (10'h9c == _T_34[9:0]) begin
        image_1_156 <= io_pixelVal_in_1_6;
      end else if (10'h9c == _T_31[9:0]) begin
        image_1_156 <= io_pixelVal_in_1_5;
      end else if (10'h9c == _T_28[9:0]) begin
        image_1_156 <= io_pixelVal_in_1_4;
      end else if (10'h9c == _T_25[9:0]) begin
        image_1_156 <= io_pixelVal_in_1_3;
      end else if (10'h9c == _T_22[9:0]) begin
        image_1_156 <= io_pixelVal_in_1_2;
      end else if (10'h9c == _T_19[9:0]) begin
        image_1_156 <= io_pixelVal_in_1_1;
      end else if (10'h9c == _T_15[9:0]) begin
        image_1_156 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_157 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9d == _T_37[9:0]) begin
        image_1_157 <= io_pixelVal_in_1_7;
      end else if (10'h9d == _T_34[9:0]) begin
        image_1_157 <= io_pixelVal_in_1_6;
      end else if (10'h9d == _T_31[9:0]) begin
        image_1_157 <= io_pixelVal_in_1_5;
      end else if (10'h9d == _T_28[9:0]) begin
        image_1_157 <= io_pixelVal_in_1_4;
      end else if (10'h9d == _T_25[9:0]) begin
        image_1_157 <= io_pixelVal_in_1_3;
      end else if (10'h9d == _T_22[9:0]) begin
        image_1_157 <= io_pixelVal_in_1_2;
      end else if (10'h9d == _T_19[9:0]) begin
        image_1_157 <= io_pixelVal_in_1_1;
      end else if (10'h9d == _T_15[9:0]) begin
        image_1_157 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_158 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9e == _T_37[9:0]) begin
        image_1_158 <= io_pixelVal_in_1_7;
      end else if (10'h9e == _T_34[9:0]) begin
        image_1_158 <= io_pixelVal_in_1_6;
      end else if (10'h9e == _T_31[9:0]) begin
        image_1_158 <= io_pixelVal_in_1_5;
      end else if (10'h9e == _T_28[9:0]) begin
        image_1_158 <= io_pixelVal_in_1_4;
      end else if (10'h9e == _T_25[9:0]) begin
        image_1_158 <= io_pixelVal_in_1_3;
      end else if (10'h9e == _T_22[9:0]) begin
        image_1_158 <= io_pixelVal_in_1_2;
      end else if (10'h9e == _T_19[9:0]) begin
        image_1_158 <= io_pixelVal_in_1_1;
      end else if (10'h9e == _T_15[9:0]) begin
        image_1_158 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_159 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9f == _T_37[9:0]) begin
        image_1_159 <= io_pixelVal_in_1_7;
      end else if (10'h9f == _T_34[9:0]) begin
        image_1_159 <= io_pixelVal_in_1_6;
      end else if (10'h9f == _T_31[9:0]) begin
        image_1_159 <= io_pixelVal_in_1_5;
      end else if (10'h9f == _T_28[9:0]) begin
        image_1_159 <= io_pixelVal_in_1_4;
      end else if (10'h9f == _T_25[9:0]) begin
        image_1_159 <= io_pixelVal_in_1_3;
      end else if (10'h9f == _T_22[9:0]) begin
        image_1_159 <= io_pixelVal_in_1_2;
      end else if (10'h9f == _T_19[9:0]) begin
        image_1_159 <= io_pixelVal_in_1_1;
      end else if (10'h9f == _T_15[9:0]) begin
        image_1_159 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_160 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha0 == _T_37[9:0]) begin
        image_1_160 <= io_pixelVal_in_1_7;
      end else if (10'ha0 == _T_34[9:0]) begin
        image_1_160 <= io_pixelVal_in_1_6;
      end else if (10'ha0 == _T_31[9:0]) begin
        image_1_160 <= io_pixelVal_in_1_5;
      end else if (10'ha0 == _T_28[9:0]) begin
        image_1_160 <= io_pixelVal_in_1_4;
      end else if (10'ha0 == _T_25[9:0]) begin
        image_1_160 <= io_pixelVal_in_1_3;
      end else if (10'ha0 == _T_22[9:0]) begin
        image_1_160 <= io_pixelVal_in_1_2;
      end else if (10'ha0 == _T_19[9:0]) begin
        image_1_160 <= io_pixelVal_in_1_1;
      end else if (10'ha0 == _T_15[9:0]) begin
        image_1_160 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_161 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha1 == _T_37[9:0]) begin
        image_1_161 <= io_pixelVal_in_1_7;
      end else if (10'ha1 == _T_34[9:0]) begin
        image_1_161 <= io_pixelVal_in_1_6;
      end else if (10'ha1 == _T_31[9:0]) begin
        image_1_161 <= io_pixelVal_in_1_5;
      end else if (10'ha1 == _T_28[9:0]) begin
        image_1_161 <= io_pixelVal_in_1_4;
      end else if (10'ha1 == _T_25[9:0]) begin
        image_1_161 <= io_pixelVal_in_1_3;
      end else if (10'ha1 == _T_22[9:0]) begin
        image_1_161 <= io_pixelVal_in_1_2;
      end else if (10'ha1 == _T_19[9:0]) begin
        image_1_161 <= io_pixelVal_in_1_1;
      end else if (10'ha1 == _T_15[9:0]) begin
        image_1_161 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_162 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha2 == _T_37[9:0]) begin
        image_1_162 <= io_pixelVal_in_1_7;
      end else if (10'ha2 == _T_34[9:0]) begin
        image_1_162 <= io_pixelVal_in_1_6;
      end else if (10'ha2 == _T_31[9:0]) begin
        image_1_162 <= io_pixelVal_in_1_5;
      end else if (10'ha2 == _T_28[9:0]) begin
        image_1_162 <= io_pixelVal_in_1_4;
      end else if (10'ha2 == _T_25[9:0]) begin
        image_1_162 <= io_pixelVal_in_1_3;
      end else if (10'ha2 == _T_22[9:0]) begin
        image_1_162 <= io_pixelVal_in_1_2;
      end else if (10'ha2 == _T_19[9:0]) begin
        image_1_162 <= io_pixelVal_in_1_1;
      end else if (10'ha2 == _T_15[9:0]) begin
        image_1_162 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_163 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha3 == _T_37[9:0]) begin
        image_1_163 <= io_pixelVal_in_1_7;
      end else if (10'ha3 == _T_34[9:0]) begin
        image_1_163 <= io_pixelVal_in_1_6;
      end else if (10'ha3 == _T_31[9:0]) begin
        image_1_163 <= io_pixelVal_in_1_5;
      end else if (10'ha3 == _T_28[9:0]) begin
        image_1_163 <= io_pixelVal_in_1_4;
      end else if (10'ha3 == _T_25[9:0]) begin
        image_1_163 <= io_pixelVal_in_1_3;
      end else if (10'ha3 == _T_22[9:0]) begin
        image_1_163 <= io_pixelVal_in_1_2;
      end else if (10'ha3 == _T_19[9:0]) begin
        image_1_163 <= io_pixelVal_in_1_1;
      end else if (10'ha3 == _T_15[9:0]) begin
        image_1_163 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_164 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha4 == _T_37[9:0]) begin
        image_1_164 <= io_pixelVal_in_1_7;
      end else if (10'ha4 == _T_34[9:0]) begin
        image_1_164 <= io_pixelVal_in_1_6;
      end else if (10'ha4 == _T_31[9:0]) begin
        image_1_164 <= io_pixelVal_in_1_5;
      end else if (10'ha4 == _T_28[9:0]) begin
        image_1_164 <= io_pixelVal_in_1_4;
      end else if (10'ha4 == _T_25[9:0]) begin
        image_1_164 <= io_pixelVal_in_1_3;
      end else if (10'ha4 == _T_22[9:0]) begin
        image_1_164 <= io_pixelVal_in_1_2;
      end else if (10'ha4 == _T_19[9:0]) begin
        image_1_164 <= io_pixelVal_in_1_1;
      end else if (10'ha4 == _T_15[9:0]) begin
        image_1_164 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_165 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha5 == _T_37[9:0]) begin
        image_1_165 <= io_pixelVal_in_1_7;
      end else if (10'ha5 == _T_34[9:0]) begin
        image_1_165 <= io_pixelVal_in_1_6;
      end else if (10'ha5 == _T_31[9:0]) begin
        image_1_165 <= io_pixelVal_in_1_5;
      end else if (10'ha5 == _T_28[9:0]) begin
        image_1_165 <= io_pixelVal_in_1_4;
      end else if (10'ha5 == _T_25[9:0]) begin
        image_1_165 <= io_pixelVal_in_1_3;
      end else if (10'ha5 == _T_22[9:0]) begin
        image_1_165 <= io_pixelVal_in_1_2;
      end else if (10'ha5 == _T_19[9:0]) begin
        image_1_165 <= io_pixelVal_in_1_1;
      end else if (10'ha5 == _T_15[9:0]) begin
        image_1_165 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_166 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha6 == _T_37[9:0]) begin
        image_1_166 <= io_pixelVal_in_1_7;
      end else if (10'ha6 == _T_34[9:0]) begin
        image_1_166 <= io_pixelVal_in_1_6;
      end else if (10'ha6 == _T_31[9:0]) begin
        image_1_166 <= io_pixelVal_in_1_5;
      end else if (10'ha6 == _T_28[9:0]) begin
        image_1_166 <= io_pixelVal_in_1_4;
      end else if (10'ha6 == _T_25[9:0]) begin
        image_1_166 <= io_pixelVal_in_1_3;
      end else if (10'ha6 == _T_22[9:0]) begin
        image_1_166 <= io_pixelVal_in_1_2;
      end else if (10'ha6 == _T_19[9:0]) begin
        image_1_166 <= io_pixelVal_in_1_1;
      end else if (10'ha6 == _T_15[9:0]) begin
        image_1_166 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_167 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha7 == _T_37[9:0]) begin
        image_1_167 <= io_pixelVal_in_1_7;
      end else if (10'ha7 == _T_34[9:0]) begin
        image_1_167 <= io_pixelVal_in_1_6;
      end else if (10'ha7 == _T_31[9:0]) begin
        image_1_167 <= io_pixelVal_in_1_5;
      end else if (10'ha7 == _T_28[9:0]) begin
        image_1_167 <= io_pixelVal_in_1_4;
      end else if (10'ha7 == _T_25[9:0]) begin
        image_1_167 <= io_pixelVal_in_1_3;
      end else if (10'ha7 == _T_22[9:0]) begin
        image_1_167 <= io_pixelVal_in_1_2;
      end else if (10'ha7 == _T_19[9:0]) begin
        image_1_167 <= io_pixelVal_in_1_1;
      end else if (10'ha7 == _T_15[9:0]) begin
        image_1_167 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_168 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha8 == _T_37[9:0]) begin
        image_1_168 <= io_pixelVal_in_1_7;
      end else if (10'ha8 == _T_34[9:0]) begin
        image_1_168 <= io_pixelVal_in_1_6;
      end else if (10'ha8 == _T_31[9:0]) begin
        image_1_168 <= io_pixelVal_in_1_5;
      end else if (10'ha8 == _T_28[9:0]) begin
        image_1_168 <= io_pixelVal_in_1_4;
      end else if (10'ha8 == _T_25[9:0]) begin
        image_1_168 <= io_pixelVal_in_1_3;
      end else if (10'ha8 == _T_22[9:0]) begin
        image_1_168 <= io_pixelVal_in_1_2;
      end else if (10'ha8 == _T_19[9:0]) begin
        image_1_168 <= io_pixelVal_in_1_1;
      end else if (10'ha8 == _T_15[9:0]) begin
        image_1_168 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_169 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha9 == _T_37[9:0]) begin
        image_1_169 <= io_pixelVal_in_1_7;
      end else if (10'ha9 == _T_34[9:0]) begin
        image_1_169 <= io_pixelVal_in_1_6;
      end else if (10'ha9 == _T_31[9:0]) begin
        image_1_169 <= io_pixelVal_in_1_5;
      end else if (10'ha9 == _T_28[9:0]) begin
        image_1_169 <= io_pixelVal_in_1_4;
      end else if (10'ha9 == _T_25[9:0]) begin
        image_1_169 <= io_pixelVal_in_1_3;
      end else if (10'ha9 == _T_22[9:0]) begin
        image_1_169 <= io_pixelVal_in_1_2;
      end else if (10'ha9 == _T_19[9:0]) begin
        image_1_169 <= io_pixelVal_in_1_1;
      end else if (10'ha9 == _T_15[9:0]) begin
        image_1_169 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_170 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'haa == _T_37[9:0]) begin
        image_1_170 <= io_pixelVal_in_1_7;
      end else if (10'haa == _T_34[9:0]) begin
        image_1_170 <= io_pixelVal_in_1_6;
      end else if (10'haa == _T_31[9:0]) begin
        image_1_170 <= io_pixelVal_in_1_5;
      end else if (10'haa == _T_28[9:0]) begin
        image_1_170 <= io_pixelVal_in_1_4;
      end else if (10'haa == _T_25[9:0]) begin
        image_1_170 <= io_pixelVal_in_1_3;
      end else if (10'haa == _T_22[9:0]) begin
        image_1_170 <= io_pixelVal_in_1_2;
      end else if (10'haa == _T_19[9:0]) begin
        image_1_170 <= io_pixelVal_in_1_1;
      end else if (10'haa == _T_15[9:0]) begin
        image_1_170 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_171 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hab == _T_37[9:0]) begin
        image_1_171 <= io_pixelVal_in_1_7;
      end else if (10'hab == _T_34[9:0]) begin
        image_1_171 <= io_pixelVal_in_1_6;
      end else if (10'hab == _T_31[9:0]) begin
        image_1_171 <= io_pixelVal_in_1_5;
      end else if (10'hab == _T_28[9:0]) begin
        image_1_171 <= io_pixelVal_in_1_4;
      end else if (10'hab == _T_25[9:0]) begin
        image_1_171 <= io_pixelVal_in_1_3;
      end else if (10'hab == _T_22[9:0]) begin
        image_1_171 <= io_pixelVal_in_1_2;
      end else if (10'hab == _T_19[9:0]) begin
        image_1_171 <= io_pixelVal_in_1_1;
      end else if (10'hab == _T_15[9:0]) begin
        image_1_171 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_172 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hac == _T_37[9:0]) begin
        image_1_172 <= io_pixelVal_in_1_7;
      end else if (10'hac == _T_34[9:0]) begin
        image_1_172 <= io_pixelVal_in_1_6;
      end else if (10'hac == _T_31[9:0]) begin
        image_1_172 <= io_pixelVal_in_1_5;
      end else if (10'hac == _T_28[9:0]) begin
        image_1_172 <= io_pixelVal_in_1_4;
      end else if (10'hac == _T_25[9:0]) begin
        image_1_172 <= io_pixelVal_in_1_3;
      end else if (10'hac == _T_22[9:0]) begin
        image_1_172 <= io_pixelVal_in_1_2;
      end else if (10'hac == _T_19[9:0]) begin
        image_1_172 <= io_pixelVal_in_1_1;
      end else if (10'hac == _T_15[9:0]) begin
        image_1_172 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_173 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'had == _T_37[9:0]) begin
        image_1_173 <= io_pixelVal_in_1_7;
      end else if (10'had == _T_34[9:0]) begin
        image_1_173 <= io_pixelVal_in_1_6;
      end else if (10'had == _T_31[9:0]) begin
        image_1_173 <= io_pixelVal_in_1_5;
      end else if (10'had == _T_28[9:0]) begin
        image_1_173 <= io_pixelVal_in_1_4;
      end else if (10'had == _T_25[9:0]) begin
        image_1_173 <= io_pixelVal_in_1_3;
      end else if (10'had == _T_22[9:0]) begin
        image_1_173 <= io_pixelVal_in_1_2;
      end else if (10'had == _T_19[9:0]) begin
        image_1_173 <= io_pixelVal_in_1_1;
      end else if (10'had == _T_15[9:0]) begin
        image_1_173 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_174 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hae == _T_37[9:0]) begin
        image_1_174 <= io_pixelVal_in_1_7;
      end else if (10'hae == _T_34[9:0]) begin
        image_1_174 <= io_pixelVal_in_1_6;
      end else if (10'hae == _T_31[9:0]) begin
        image_1_174 <= io_pixelVal_in_1_5;
      end else if (10'hae == _T_28[9:0]) begin
        image_1_174 <= io_pixelVal_in_1_4;
      end else if (10'hae == _T_25[9:0]) begin
        image_1_174 <= io_pixelVal_in_1_3;
      end else if (10'hae == _T_22[9:0]) begin
        image_1_174 <= io_pixelVal_in_1_2;
      end else if (10'hae == _T_19[9:0]) begin
        image_1_174 <= io_pixelVal_in_1_1;
      end else if (10'hae == _T_15[9:0]) begin
        image_1_174 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_175 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'haf == _T_37[9:0]) begin
        image_1_175 <= io_pixelVal_in_1_7;
      end else if (10'haf == _T_34[9:0]) begin
        image_1_175 <= io_pixelVal_in_1_6;
      end else if (10'haf == _T_31[9:0]) begin
        image_1_175 <= io_pixelVal_in_1_5;
      end else if (10'haf == _T_28[9:0]) begin
        image_1_175 <= io_pixelVal_in_1_4;
      end else if (10'haf == _T_25[9:0]) begin
        image_1_175 <= io_pixelVal_in_1_3;
      end else if (10'haf == _T_22[9:0]) begin
        image_1_175 <= io_pixelVal_in_1_2;
      end else if (10'haf == _T_19[9:0]) begin
        image_1_175 <= io_pixelVal_in_1_1;
      end else if (10'haf == _T_15[9:0]) begin
        image_1_175 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_176 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb0 == _T_37[9:0]) begin
        image_1_176 <= io_pixelVal_in_1_7;
      end else if (10'hb0 == _T_34[9:0]) begin
        image_1_176 <= io_pixelVal_in_1_6;
      end else if (10'hb0 == _T_31[9:0]) begin
        image_1_176 <= io_pixelVal_in_1_5;
      end else if (10'hb0 == _T_28[9:0]) begin
        image_1_176 <= io_pixelVal_in_1_4;
      end else if (10'hb0 == _T_25[9:0]) begin
        image_1_176 <= io_pixelVal_in_1_3;
      end else if (10'hb0 == _T_22[9:0]) begin
        image_1_176 <= io_pixelVal_in_1_2;
      end else if (10'hb0 == _T_19[9:0]) begin
        image_1_176 <= io_pixelVal_in_1_1;
      end else if (10'hb0 == _T_15[9:0]) begin
        image_1_176 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_177 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb1 == _T_37[9:0]) begin
        image_1_177 <= io_pixelVal_in_1_7;
      end else if (10'hb1 == _T_34[9:0]) begin
        image_1_177 <= io_pixelVal_in_1_6;
      end else if (10'hb1 == _T_31[9:0]) begin
        image_1_177 <= io_pixelVal_in_1_5;
      end else if (10'hb1 == _T_28[9:0]) begin
        image_1_177 <= io_pixelVal_in_1_4;
      end else if (10'hb1 == _T_25[9:0]) begin
        image_1_177 <= io_pixelVal_in_1_3;
      end else if (10'hb1 == _T_22[9:0]) begin
        image_1_177 <= io_pixelVal_in_1_2;
      end else if (10'hb1 == _T_19[9:0]) begin
        image_1_177 <= io_pixelVal_in_1_1;
      end else if (10'hb1 == _T_15[9:0]) begin
        image_1_177 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_178 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb2 == _T_37[9:0]) begin
        image_1_178 <= io_pixelVal_in_1_7;
      end else if (10'hb2 == _T_34[9:0]) begin
        image_1_178 <= io_pixelVal_in_1_6;
      end else if (10'hb2 == _T_31[9:0]) begin
        image_1_178 <= io_pixelVal_in_1_5;
      end else if (10'hb2 == _T_28[9:0]) begin
        image_1_178 <= io_pixelVal_in_1_4;
      end else if (10'hb2 == _T_25[9:0]) begin
        image_1_178 <= io_pixelVal_in_1_3;
      end else if (10'hb2 == _T_22[9:0]) begin
        image_1_178 <= io_pixelVal_in_1_2;
      end else if (10'hb2 == _T_19[9:0]) begin
        image_1_178 <= io_pixelVal_in_1_1;
      end else if (10'hb2 == _T_15[9:0]) begin
        image_1_178 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_179 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb3 == _T_37[9:0]) begin
        image_1_179 <= io_pixelVal_in_1_7;
      end else if (10'hb3 == _T_34[9:0]) begin
        image_1_179 <= io_pixelVal_in_1_6;
      end else if (10'hb3 == _T_31[9:0]) begin
        image_1_179 <= io_pixelVal_in_1_5;
      end else if (10'hb3 == _T_28[9:0]) begin
        image_1_179 <= io_pixelVal_in_1_4;
      end else if (10'hb3 == _T_25[9:0]) begin
        image_1_179 <= io_pixelVal_in_1_3;
      end else if (10'hb3 == _T_22[9:0]) begin
        image_1_179 <= io_pixelVal_in_1_2;
      end else if (10'hb3 == _T_19[9:0]) begin
        image_1_179 <= io_pixelVal_in_1_1;
      end else if (10'hb3 == _T_15[9:0]) begin
        image_1_179 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_180 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb4 == _T_37[9:0]) begin
        image_1_180 <= io_pixelVal_in_1_7;
      end else if (10'hb4 == _T_34[9:0]) begin
        image_1_180 <= io_pixelVal_in_1_6;
      end else if (10'hb4 == _T_31[9:0]) begin
        image_1_180 <= io_pixelVal_in_1_5;
      end else if (10'hb4 == _T_28[9:0]) begin
        image_1_180 <= io_pixelVal_in_1_4;
      end else if (10'hb4 == _T_25[9:0]) begin
        image_1_180 <= io_pixelVal_in_1_3;
      end else if (10'hb4 == _T_22[9:0]) begin
        image_1_180 <= io_pixelVal_in_1_2;
      end else if (10'hb4 == _T_19[9:0]) begin
        image_1_180 <= io_pixelVal_in_1_1;
      end else if (10'hb4 == _T_15[9:0]) begin
        image_1_180 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_181 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb5 == _T_37[9:0]) begin
        image_1_181 <= io_pixelVal_in_1_7;
      end else if (10'hb5 == _T_34[9:0]) begin
        image_1_181 <= io_pixelVal_in_1_6;
      end else if (10'hb5 == _T_31[9:0]) begin
        image_1_181 <= io_pixelVal_in_1_5;
      end else if (10'hb5 == _T_28[9:0]) begin
        image_1_181 <= io_pixelVal_in_1_4;
      end else if (10'hb5 == _T_25[9:0]) begin
        image_1_181 <= io_pixelVal_in_1_3;
      end else if (10'hb5 == _T_22[9:0]) begin
        image_1_181 <= io_pixelVal_in_1_2;
      end else if (10'hb5 == _T_19[9:0]) begin
        image_1_181 <= io_pixelVal_in_1_1;
      end else if (10'hb5 == _T_15[9:0]) begin
        image_1_181 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_182 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb6 == _T_37[9:0]) begin
        image_1_182 <= io_pixelVal_in_1_7;
      end else if (10'hb6 == _T_34[9:0]) begin
        image_1_182 <= io_pixelVal_in_1_6;
      end else if (10'hb6 == _T_31[9:0]) begin
        image_1_182 <= io_pixelVal_in_1_5;
      end else if (10'hb6 == _T_28[9:0]) begin
        image_1_182 <= io_pixelVal_in_1_4;
      end else if (10'hb6 == _T_25[9:0]) begin
        image_1_182 <= io_pixelVal_in_1_3;
      end else if (10'hb6 == _T_22[9:0]) begin
        image_1_182 <= io_pixelVal_in_1_2;
      end else if (10'hb6 == _T_19[9:0]) begin
        image_1_182 <= io_pixelVal_in_1_1;
      end else if (10'hb6 == _T_15[9:0]) begin
        image_1_182 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_183 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb7 == _T_37[9:0]) begin
        image_1_183 <= io_pixelVal_in_1_7;
      end else if (10'hb7 == _T_34[9:0]) begin
        image_1_183 <= io_pixelVal_in_1_6;
      end else if (10'hb7 == _T_31[9:0]) begin
        image_1_183 <= io_pixelVal_in_1_5;
      end else if (10'hb7 == _T_28[9:0]) begin
        image_1_183 <= io_pixelVal_in_1_4;
      end else if (10'hb7 == _T_25[9:0]) begin
        image_1_183 <= io_pixelVal_in_1_3;
      end else if (10'hb7 == _T_22[9:0]) begin
        image_1_183 <= io_pixelVal_in_1_2;
      end else if (10'hb7 == _T_19[9:0]) begin
        image_1_183 <= io_pixelVal_in_1_1;
      end else if (10'hb7 == _T_15[9:0]) begin
        image_1_183 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_184 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb8 == _T_37[9:0]) begin
        image_1_184 <= io_pixelVal_in_1_7;
      end else if (10'hb8 == _T_34[9:0]) begin
        image_1_184 <= io_pixelVal_in_1_6;
      end else if (10'hb8 == _T_31[9:0]) begin
        image_1_184 <= io_pixelVal_in_1_5;
      end else if (10'hb8 == _T_28[9:0]) begin
        image_1_184 <= io_pixelVal_in_1_4;
      end else if (10'hb8 == _T_25[9:0]) begin
        image_1_184 <= io_pixelVal_in_1_3;
      end else if (10'hb8 == _T_22[9:0]) begin
        image_1_184 <= io_pixelVal_in_1_2;
      end else if (10'hb8 == _T_19[9:0]) begin
        image_1_184 <= io_pixelVal_in_1_1;
      end else if (10'hb8 == _T_15[9:0]) begin
        image_1_184 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_185 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb9 == _T_37[9:0]) begin
        image_1_185 <= io_pixelVal_in_1_7;
      end else if (10'hb9 == _T_34[9:0]) begin
        image_1_185 <= io_pixelVal_in_1_6;
      end else if (10'hb9 == _T_31[9:0]) begin
        image_1_185 <= io_pixelVal_in_1_5;
      end else if (10'hb9 == _T_28[9:0]) begin
        image_1_185 <= io_pixelVal_in_1_4;
      end else if (10'hb9 == _T_25[9:0]) begin
        image_1_185 <= io_pixelVal_in_1_3;
      end else if (10'hb9 == _T_22[9:0]) begin
        image_1_185 <= io_pixelVal_in_1_2;
      end else if (10'hb9 == _T_19[9:0]) begin
        image_1_185 <= io_pixelVal_in_1_1;
      end else if (10'hb9 == _T_15[9:0]) begin
        image_1_185 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_186 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hba == _T_37[9:0]) begin
        image_1_186 <= io_pixelVal_in_1_7;
      end else if (10'hba == _T_34[9:0]) begin
        image_1_186 <= io_pixelVal_in_1_6;
      end else if (10'hba == _T_31[9:0]) begin
        image_1_186 <= io_pixelVal_in_1_5;
      end else if (10'hba == _T_28[9:0]) begin
        image_1_186 <= io_pixelVal_in_1_4;
      end else if (10'hba == _T_25[9:0]) begin
        image_1_186 <= io_pixelVal_in_1_3;
      end else if (10'hba == _T_22[9:0]) begin
        image_1_186 <= io_pixelVal_in_1_2;
      end else if (10'hba == _T_19[9:0]) begin
        image_1_186 <= io_pixelVal_in_1_1;
      end else if (10'hba == _T_15[9:0]) begin
        image_1_186 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_187 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hbb == _T_37[9:0]) begin
        image_1_187 <= io_pixelVal_in_1_7;
      end else if (10'hbb == _T_34[9:0]) begin
        image_1_187 <= io_pixelVal_in_1_6;
      end else if (10'hbb == _T_31[9:0]) begin
        image_1_187 <= io_pixelVal_in_1_5;
      end else if (10'hbb == _T_28[9:0]) begin
        image_1_187 <= io_pixelVal_in_1_4;
      end else if (10'hbb == _T_25[9:0]) begin
        image_1_187 <= io_pixelVal_in_1_3;
      end else if (10'hbb == _T_22[9:0]) begin
        image_1_187 <= io_pixelVal_in_1_2;
      end else if (10'hbb == _T_19[9:0]) begin
        image_1_187 <= io_pixelVal_in_1_1;
      end else if (10'hbb == _T_15[9:0]) begin
        image_1_187 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_188 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hbc == _T_37[9:0]) begin
        image_1_188 <= io_pixelVal_in_1_7;
      end else if (10'hbc == _T_34[9:0]) begin
        image_1_188 <= io_pixelVal_in_1_6;
      end else if (10'hbc == _T_31[9:0]) begin
        image_1_188 <= io_pixelVal_in_1_5;
      end else if (10'hbc == _T_28[9:0]) begin
        image_1_188 <= io_pixelVal_in_1_4;
      end else if (10'hbc == _T_25[9:0]) begin
        image_1_188 <= io_pixelVal_in_1_3;
      end else if (10'hbc == _T_22[9:0]) begin
        image_1_188 <= io_pixelVal_in_1_2;
      end else if (10'hbc == _T_19[9:0]) begin
        image_1_188 <= io_pixelVal_in_1_1;
      end else if (10'hbc == _T_15[9:0]) begin
        image_1_188 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_189 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hbd == _T_37[9:0]) begin
        image_1_189 <= io_pixelVal_in_1_7;
      end else if (10'hbd == _T_34[9:0]) begin
        image_1_189 <= io_pixelVal_in_1_6;
      end else if (10'hbd == _T_31[9:0]) begin
        image_1_189 <= io_pixelVal_in_1_5;
      end else if (10'hbd == _T_28[9:0]) begin
        image_1_189 <= io_pixelVal_in_1_4;
      end else if (10'hbd == _T_25[9:0]) begin
        image_1_189 <= io_pixelVal_in_1_3;
      end else if (10'hbd == _T_22[9:0]) begin
        image_1_189 <= io_pixelVal_in_1_2;
      end else if (10'hbd == _T_19[9:0]) begin
        image_1_189 <= io_pixelVal_in_1_1;
      end else if (10'hbd == _T_15[9:0]) begin
        image_1_189 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_190 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hbe == _T_37[9:0]) begin
        image_1_190 <= io_pixelVal_in_1_7;
      end else if (10'hbe == _T_34[9:0]) begin
        image_1_190 <= io_pixelVal_in_1_6;
      end else if (10'hbe == _T_31[9:0]) begin
        image_1_190 <= io_pixelVal_in_1_5;
      end else if (10'hbe == _T_28[9:0]) begin
        image_1_190 <= io_pixelVal_in_1_4;
      end else if (10'hbe == _T_25[9:0]) begin
        image_1_190 <= io_pixelVal_in_1_3;
      end else if (10'hbe == _T_22[9:0]) begin
        image_1_190 <= io_pixelVal_in_1_2;
      end else if (10'hbe == _T_19[9:0]) begin
        image_1_190 <= io_pixelVal_in_1_1;
      end else if (10'hbe == _T_15[9:0]) begin
        image_1_190 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_191 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hbf == _T_37[9:0]) begin
        image_1_191 <= io_pixelVal_in_1_7;
      end else if (10'hbf == _T_34[9:0]) begin
        image_1_191 <= io_pixelVal_in_1_6;
      end else if (10'hbf == _T_31[9:0]) begin
        image_1_191 <= io_pixelVal_in_1_5;
      end else if (10'hbf == _T_28[9:0]) begin
        image_1_191 <= io_pixelVal_in_1_4;
      end else if (10'hbf == _T_25[9:0]) begin
        image_1_191 <= io_pixelVal_in_1_3;
      end else if (10'hbf == _T_22[9:0]) begin
        image_1_191 <= io_pixelVal_in_1_2;
      end else if (10'hbf == _T_19[9:0]) begin
        image_1_191 <= io_pixelVal_in_1_1;
      end else if (10'hbf == _T_15[9:0]) begin
        image_1_191 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_192 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc0 == _T_37[9:0]) begin
        image_1_192 <= io_pixelVal_in_1_7;
      end else if (10'hc0 == _T_34[9:0]) begin
        image_1_192 <= io_pixelVal_in_1_6;
      end else if (10'hc0 == _T_31[9:0]) begin
        image_1_192 <= io_pixelVal_in_1_5;
      end else if (10'hc0 == _T_28[9:0]) begin
        image_1_192 <= io_pixelVal_in_1_4;
      end else if (10'hc0 == _T_25[9:0]) begin
        image_1_192 <= io_pixelVal_in_1_3;
      end else if (10'hc0 == _T_22[9:0]) begin
        image_1_192 <= io_pixelVal_in_1_2;
      end else if (10'hc0 == _T_19[9:0]) begin
        image_1_192 <= io_pixelVal_in_1_1;
      end else if (10'hc0 == _T_15[9:0]) begin
        image_1_192 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_193 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc1 == _T_37[9:0]) begin
        image_1_193 <= io_pixelVal_in_1_7;
      end else if (10'hc1 == _T_34[9:0]) begin
        image_1_193 <= io_pixelVal_in_1_6;
      end else if (10'hc1 == _T_31[9:0]) begin
        image_1_193 <= io_pixelVal_in_1_5;
      end else if (10'hc1 == _T_28[9:0]) begin
        image_1_193 <= io_pixelVal_in_1_4;
      end else if (10'hc1 == _T_25[9:0]) begin
        image_1_193 <= io_pixelVal_in_1_3;
      end else if (10'hc1 == _T_22[9:0]) begin
        image_1_193 <= io_pixelVal_in_1_2;
      end else if (10'hc1 == _T_19[9:0]) begin
        image_1_193 <= io_pixelVal_in_1_1;
      end else if (10'hc1 == _T_15[9:0]) begin
        image_1_193 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_194 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc2 == _T_37[9:0]) begin
        image_1_194 <= io_pixelVal_in_1_7;
      end else if (10'hc2 == _T_34[9:0]) begin
        image_1_194 <= io_pixelVal_in_1_6;
      end else if (10'hc2 == _T_31[9:0]) begin
        image_1_194 <= io_pixelVal_in_1_5;
      end else if (10'hc2 == _T_28[9:0]) begin
        image_1_194 <= io_pixelVal_in_1_4;
      end else if (10'hc2 == _T_25[9:0]) begin
        image_1_194 <= io_pixelVal_in_1_3;
      end else if (10'hc2 == _T_22[9:0]) begin
        image_1_194 <= io_pixelVal_in_1_2;
      end else if (10'hc2 == _T_19[9:0]) begin
        image_1_194 <= io_pixelVal_in_1_1;
      end else if (10'hc2 == _T_15[9:0]) begin
        image_1_194 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_195 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc3 == _T_37[9:0]) begin
        image_1_195 <= io_pixelVal_in_1_7;
      end else if (10'hc3 == _T_34[9:0]) begin
        image_1_195 <= io_pixelVal_in_1_6;
      end else if (10'hc3 == _T_31[9:0]) begin
        image_1_195 <= io_pixelVal_in_1_5;
      end else if (10'hc3 == _T_28[9:0]) begin
        image_1_195 <= io_pixelVal_in_1_4;
      end else if (10'hc3 == _T_25[9:0]) begin
        image_1_195 <= io_pixelVal_in_1_3;
      end else if (10'hc3 == _T_22[9:0]) begin
        image_1_195 <= io_pixelVal_in_1_2;
      end else if (10'hc3 == _T_19[9:0]) begin
        image_1_195 <= io_pixelVal_in_1_1;
      end else if (10'hc3 == _T_15[9:0]) begin
        image_1_195 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_196 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc4 == _T_37[9:0]) begin
        image_1_196 <= io_pixelVal_in_1_7;
      end else if (10'hc4 == _T_34[9:0]) begin
        image_1_196 <= io_pixelVal_in_1_6;
      end else if (10'hc4 == _T_31[9:0]) begin
        image_1_196 <= io_pixelVal_in_1_5;
      end else if (10'hc4 == _T_28[9:0]) begin
        image_1_196 <= io_pixelVal_in_1_4;
      end else if (10'hc4 == _T_25[9:0]) begin
        image_1_196 <= io_pixelVal_in_1_3;
      end else if (10'hc4 == _T_22[9:0]) begin
        image_1_196 <= io_pixelVal_in_1_2;
      end else if (10'hc4 == _T_19[9:0]) begin
        image_1_196 <= io_pixelVal_in_1_1;
      end else if (10'hc4 == _T_15[9:0]) begin
        image_1_196 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_197 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc5 == _T_37[9:0]) begin
        image_1_197 <= io_pixelVal_in_1_7;
      end else if (10'hc5 == _T_34[9:0]) begin
        image_1_197 <= io_pixelVal_in_1_6;
      end else if (10'hc5 == _T_31[9:0]) begin
        image_1_197 <= io_pixelVal_in_1_5;
      end else if (10'hc5 == _T_28[9:0]) begin
        image_1_197 <= io_pixelVal_in_1_4;
      end else if (10'hc5 == _T_25[9:0]) begin
        image_1_197 <= io_pixelVal_in_1_3;
      end else if (10'hc5 == _T_22[9:0]) begin
        image_1_197 <= io_pixelVal_in_1_2;
      end else if (10'hc5 == _T_19[9:0]) begin
        image_1_197 <= io_pixelVal_in_1_1;
      end else if (10'hc5 == _T_15[9:0]) begin
        image_1_197 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_198 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc6 == _T_37[9:0]) begin
        image_1_198 <= io_pixelVal_in_1_7;
      end else if (10'hc6 == _T_34[9:0]) begin
        image_1_198 <= io_pixelVal_in_1_6;
      end else if (10'hc6 == _T_31[9:0]) begin
        image_1_198 <= io_pixelVal_in_1_5;
      end else if (10'hc6 == _T_28[9:0]) begin
        image_1_198 <= io_pixelVal_in_1_4;
      end else if (10'hc6 == _T_25[9:0]) begin
        image_1_198 <= io_pixelVal_in_1_3;
      end else if (10'hc6 == _T_22[9:0]) begin
        image_1_198 <= io_pixelVal_in_1_2;
      end else if (10'hc6 == _T_19[9:0]) begin
        image_1_198 <= io_pixelVal_in_1_1;
      end else if (10'hc6 == _T_15[9:0]) begin
        image_1_198 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_199 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc7 == _T_37[9:0]) begin
        image_1_199 <= io_pixelVal_in_1_7;
      end else if (10'hc7 == _T_34[9:0]) begin
        image_1_199 <= io_pixelVal_in_1_6;
      end else if (10'hc7 == _T_31[9:0]) begin
        image_1_199 <= io_pixelVal_in_1_5;
      end else if (10'hc7 == _T_28[9:0]) begin
        image_1_199 <= io_pixelVal_in_1_4;
      end else if (10'hc7 == _T_25[9:0]) begin
        image_1_199 <= io_pixelVal_in_1_3;
      end else if (10'hc7 == _T_22[9:0]) begin
        image_1_199 <= io_pixelVal_in_1_2;
      end else if (10'hc7 == _T_19[9:0]) begin
        image_1_199 <= io_pixelVal_in_1_1;
      end else if (10'hc7 == _T_15[9:0]) begin
        image_1_199 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_200 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc8 == _T_37[9:0]) begin
        image_1_200 <= io_pixelVal_in_1_7;
      end else if (10'hc8 == _T_34[9:0]) begin
        image_1_200 <= io_pixelVal_in_1_6;
      end else if (10'hc8 == _T_31[9:0]) begin
        image_1_200 <= io_pixelVal_in_1_5;
      end else if (10'hc8 == _T_28[9:0]) begin
        image_1_200 <= io_pixelVal_in_1_4;
      end else if (10'hc8 == _T_25[9:0]) begin
        image_1_200 <= io_pixelVal_in_1_3;
      end else if (10'hc8 == _T_22[9:0]) begin
        image_1_200 <= io_pixelVal_in_1_2;
      end else if (10'hc8 == _T_19[9:0]) begin
        image_1_200 <= io_pixelVal_in_1_1;
      end else if (10'hc8 == _T_15[9:0]) begin
        image_1_200 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_201 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc9 == _T_37[9:0]) begin
        image_1_201 <= io_pixelVal_in_1_7;
      end else if (10'hc9 == _T_34[9:0]) begin
        image_1_201 <= io_pixelVal_in_1_6;
      end else if (10'hc9 == _T_31[9:0]) begin
        image_1_201 <= io_pixelVal_in_1_5;
      end else if (10'hc9 == _T_28[9:0]) begin
        image_1_201 <= io_pixelVal_in_1_4;
      end else if (10'hc9 == _T_25[9:0]) begin
        image_1_201 <= io_pixelVal_in_1_3;
      end else if (10'hc9 == _T_22[9:0]) begin
        image_1_201 <= io_pixelVal_in_1_2;
      end else if (10'hc9 == _T_19[9:0]) begin
        image_1_201 <= io_pixelVal_in_1_1;
      end else if (10'hc9 == _T_15[9:0]) begin
        image_1_201 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_202 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hca == _T_37[9:0]) begin
        image_1_202 <= io_pixelVal_in_1_7;
      end else if (10'hca == _T_34[9:0]) begin
        image_1_202 <= io_pixelVal_in_1_6;
      end else if (10'hca == _T_31[9:0]) begin
        image_1_202 <= io_pixelVal_in_1_5;
      end else if (10'hca == _T_28[9:0]) begin
        image_1_202 <= io_pixelVal_in_1_4;
      end else if (10'hca == _T_25[9:0]) begin
        image_1_202 <= io_pixelVal_in_1_3;
      end else if (10'hca == _T_22[9:0]) begin
        image_1_202 <= io_pixelVal_in_1_2;
      end else if (10'hca == _T_19[9:0]) begin
        image_1_202 <= io_pixelVal_in_1_1;
      end else if (10'hca == _T_15[9:0]) begin
        image_1_202 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_203 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hcb == _T_37[9:0]) begin
        image_1_203 <= io_pixelVal_in_1_7;
      end else if (10'hcb == _T_34[9:0]) begin
        image_1_203 <= io_pixelVal_in_1_6;
      end else if (10'hcb == _T_31[9:0]) begin
        image_1_203 <= io_pixelVal_in_1_5;
      end else if (10'hcb == _T_28[9:0]) begin
        image_1_203 <= io_pixelVal_in_1_4;
      end else if (10'hcb == _T_25[9:0]) begin
        image_1_203 <= io_pixelVal_in_1_3;
      end else if (10'hcb == _T_22[9:0]) begin
        image_1_203 <= io_pixelVal_in_1_2;
      end else if (10'hcb == _T_19[9:0]) begin
        image_1_203 <= io_pixelVal_in_1_1;
      end else if (10'hcb == _T_15[9:0]) begin
        image_1_203 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_204 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hcc == _T_37[9:0]) begin
        image_1_204 <= io_pixelVal_in_1_7;
      end else if (10'hcc == _T_34[9:0]) begin
        image_1_204 <= io_pixelVal_in_1_6;
      end else if (10'hcc == _T_31[9:0]) begin
        image_1_204 <= io_pixelVal_in_1_5;
      end else if (10'hcc == _T_28[9:0]) begin
        image_1_204 <= io_pixelVal_in_1_4;
      end else if (10'hcc == _T_25[9:0]) begin
        image_1_204 <= io_pixelVal_in_1_3;
      end else if (10'hcc == _T_22[9:0]) begin
        image_1_204 <= io_pixelVal_in_1_2;
      end else if (10'hcc == _T_19[9:0]) begin
        image_1_204 <= io_pixelVal_in_1_1;
      end else if (10'hcc == _T_15[9:0]) begin
        image_1_204 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_205 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hcd == _T_37[9:0]) begin
        image_1_205 <= io_pixelVal_in_1_7;
      end else if (10'hcd == _T_34[9:0]) begin
        image_1_205 <= io_pixelVal_in_1_6;
      end else if (10'hcd == _T_31[9:0]) begin
        image_1_205 <= io_pixelVal_in_1_5;
      end else if (10'hcd == _T_28[9:0]) begin
        image_1_205 <= io_pixelVal_in_1_4;
      end else if (10'hcd == _T_25[9:0]) begin
        image_1_205 <= io_pixelVal_in_1_3;
      end else if (10'hcd == _T_22[9:0]) begin
        image_1_205 <= io_pixelVal_in_1_2;
      end else if (10'hcd == _T_19[9:0]) begin
        image_1_205 <= io_pixelVal_in_1_1;
      end else if (10'hcd == _T_15[9:0]) begin
        image_1_205 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_206 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hce == _T_37[9:0]) begin
        image_1_206 <= io_pixelVal_in_1_7;
      end else if (10'hce == _T_34[9:0]) begin
        image_1_206 <= io_pixelVal_in_1_6;
      end else if (10'hce == _T_31[9:0]) begin
        image_1_206 <= io_pixelVal_in_1_5;
      end else if (10'hce == _T_28[9:0]) begin
        image_1_206 <= io_pixelVal_in_1_4;
      end else if (10'hce == _T_25[9:0]) begin
        image_1_206 <= io_pixelVal_in_1_3;
      end else if (10'hce == _T_22[9:0]) begin
        image_1_206 <= io_pixelVal_in_1_2;
      end else if (10'hce == _T_19[9:0]) begin
        image_1_206 <= io_pixelVal_in_1_1;
      end else if (10'hce == _T_15[9:0]) begin
        image_1_206 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_207 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hcf == _T_37[9:0]) begin
        image_1_207 <= io_pixelVal_in_1_7;
      end else if (10'hcf == _T_34[9:0]) begin
        image_1_207 <= io_pixelVal_in_1_6;
      end else if (10'hcf == _T_31[9:0]) begin
        image_1_207 <= io_pixelVal_in_1_5;
      end else if (10'hcf == _T_28[9:0]) begin
        image_1_207 <= io_pixelVal_in_1_4;
      end else if (10'hcf == _T_25[9:0]) begin
        image_1_207 <= io_pixelVal_in_1_3;
      end else if (10'hcf == _T_22[9:0]) begin
        image_1_207 <= io_pixelVal_in_1_2;
      end else if (10'hcf == _T_19[9:0]) begin
        image_1_207 <= io_pixelVal_in_1_1;
      end else if (10'hcf == _T_15[9:0]) begin
        image_1_207 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_208 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd0 == _T_37[9:0]) begin
        image_1_208 <= io_pixelVal_in_1_7;
      end else if (10'hd0 == _T_34[9:0]) begin
        image_1_208 <= io_pixelVal_in_1_6;
      end else if (10'hd0 == _T_31[9:0]) begin
        image_1_208 <= io_pixelVal_in_1_5;
      end else if (10'hd0 == _T_28[9:0]) begin
        image_1_208 <= io_pixelVal_in_1_4;
      end else if (10'hd0 == _T_25[9:0]) begin
        image_1_208 <= io_pixelVal_in_1_3;
      end else if (10'hd0 == _T_22[9:0]) begin
        image_1_208 <= io_pixelVal_in_1_2;
      end else if (10'hd0 == _T_19[9:0]) begin
        image_1_208 <= io_pixelVal_in_1_1;
      end else if (10'hd0 == _T_15[9:0]) begin
        image_1_208 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_209 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd1 == _T_37[9:0]) begin
        image_1_209 <= io_pixelVal_in_1_7;
      end else if (10'hd1 == _T_34[9:0]) begin
        image_1_209 <= io_pixelVal_in_1_6;
      end else if (10'hd1 == _T_31[9:0]) begin
        image_1_209 <= io_pixelVal_in_1_5;
      end else if (10'hd1 == _T_28[9:0]) begin
        image_1_209 <= io_pixelVal_in_1_4;
      end else if (10'hd1 == _T_25[9:0]) begin
        image_1_209 <= io_pixelVal_in_1_3;
      end else if (10'hd1 == _T_22[9:0]) begin
        image_1_209 <= io_pixelVal_in_1_2;
      end else if (10'hd1 == _T_19[9:0]) begin
        image_1_209 <= io_pixelVal_in_1_1;
      end else if (10'hd1 == _T_15[9:0]) begin
        image_1_209 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_210 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd2 == _T_37[9:0]) begin
        image_1_210 <= io_pixelVal_in_1_7;
      end else if (10'hd2 == _T_34[9:0]) begin
        image_1_210 <= io_pixelVal_in_1_6;
      end else if (10'hd2 == _T_31[9:0]) begin
        image_1_210 <= io_pixelVal_in_1_5;
      end else if (10'hd2 == _T_28[9:0]) begin
        image_1_210 <= io_pixelVal_in_1_4;
      end else if (10'hd2 == _T_25[9:0]) begin
        image_1_210 <= io_pixelVal_in_1_3;
      end else if (10'hd2 == _T_22[9:0]) begin
        image_1_210 <= io_pixelVal_in_1_2;
      end else if (10'hd2 == _T_19[9:0]) begin
        image_1_210 <= io_pixelVal_in_1_1;
      end else if (10'hd2 == _T_15[9:0]) begin
        image_1_210 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_211 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd3 == _T_37[9:0]) begin
        image_1_211 <= io_pixelVal_in_1_7;
      end else if (10'hd3 == _T_34[9:0]) begin
        image_1_211 <= io_pixelVal_in_1_6;
      end else if (10'hd3 == _T_31[9:0]) begin
        image_1_211 <= io_pixelVal_in_1_5;
      end else if (10'hd3 == _T_28[9:0]) begin
        image_1_211 <= io_pixelVal_in_1_4;
      end else if (10'hd3 == _T_25[9:0]) begin
        image_1_211 <= io_pixelVal_in_1_3;
      end else if (10'hd3 == _T_22[9:0]) begin
        image_1_211 <= io_pixelVal_in_1_2;
      end else if (10'hd3 == _T_19[9:0]) begin
        image_1_211 <= io_pixelVal_in_1_1;
      end else if (10'hd3 == _T_15[9:0]) begin
        image_1_211 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_212 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd4 == _T_37[9:0]) begin
        image_1_212 <= io_pixelVal_in_1_7;
      end else if (10'hd4 == _T_34[9:0]) begin
        image_1_212 <= io_pixelVal_in_1_6;
      end else if (10'hd4 == _T_31[9:0]) begin
        image_1_212 <= io_pixelVal_in_1_5;
      end else if (10'hd4 == _T_28[9:0]) begin
        image_1_212 <= io_pixelVal_in_1_4;
      end else if (10'hd4 == _T_25[9:0]) begin
        image_1_212 <= io_pixelVal_in_1_3;
      end else if (10'hd4 == _T_22[9:0]) begin
        image_1_212 <= io_pixelVal_in_1_2;
      end else if (10'hd4 == _T_19[9:0]) begin
        image_1_212 <= io_pixelVal_in_1_1;
      end else if (10'hd4 == _T_15[9:0]) begin
        image_1_212 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_213 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd5 == _T_37[9:0]) begin
        image_1_213 <= io_pixelVal_in_1_7;
      end else if (10'hd5 == _T_34[9:0]) begin
        image_1_213 <= io_pixelVal_in_1_6;
      end else if (10'hd5 == _T_31[9:0]) begin
        image_1_213 <= io_pixelVal_in_1_5;
      end else if (10'hd5 == _T_28[9:0]) begin
        image_1_213 <= io_pixelVal_in_1_4;
      end else if (10'hd5 == _T_25[9:0]) begin
        image_1_213 <= io_pixelVal_in_1_3;
      end else if (10'hd5 == _T_22[9:0]) begin
        image_1_213 <= io_pixelVal_in_1_2;
      end else if (10'hd5 == _T_19[9:0]) begin
        image_1_213 <= io_pixelVal_in_1_1;
      end else if (10'hd5 == _T_15[9:0]) begin
        image_1_213 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_214 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd6 == _T_37[9:0]) begin
        image_1_214 <= io_pixelVal_in_1_7;
      end else if (10'hd6 == _T_34[9:0]) begin
        image_1_214 <= io_pixelVal_in_1_6;
      end else if (10'hd6 == _T_31[9:0]) begin
        image_1_214 <= io_pixelVal_in_1_5;
      end else if (10'hd6 == _T_28[9:0]) begin
        image_1_214 <= io_pixelVal_in_1_4;
      end else if (10'hd6 == _T_25[9:0]) begin
        image_1_214 <= io_pixelVal_in_1_3;
      end else if (10'hd6 == _T_22[9:0]) begin
        image_1_214 <= io_pixelVal_in_1_2;
      end else if (10'hd6 == _T_19[9:0]) begin
        image_1_214 <= io_pixelVal_in_1_1;
      end else if (10'hd6 == _T_15[9:0]) begin
        image_1_214 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_215 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd7 == _T_37[9:0]) begin
        image_1_215 <= io_pixelVal_in_1_7;
      end else if (10'hd7 == _T_34[9:0]) begin
        image_1_215 <= io_pixelVal_in_1_6;
      end else if (10'hd7 == _T_31[9:0]) begin
        image_1_215 <= io_pixelVal_in_1_5;
      end else if (10'hd7 == _T_28[9:0]) begin
        image_1_215 <= io_pixelVal_in_1_4;
      end else if (10'hd7 == _T_25[9:0]) begin
        image_1_215 <= io_pixelVal_in_1_3;
      end else if (10'hd7 == _T_22[9:0]) begin
        image_1_215 <= io_pixelVal_in_1_2;
      end else if (10'hd7 == _T_19[9:0]) begin
        image_1_215 <= io_pixelVal_in_1_1;
      end else if (10'hd7 == _T_15[9:0]) begin
        image_1_215 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_216 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd8 == _T_37[9:0]) begin
        image_1_216 <= io_pixelVal_in_1_7;
      end else if (10'hd8 == _T_34[9:0]) begin
        image_1_216 <= io_pixelVal_in_1_6;
      end else if (10'hd8 == _T_31[9:0]) begin
        image_1_216 <= io_pixelVal_in_1_5;
      end else if (10'hd8 == _T_28[9:0]) begin
        image_1_216 <= io_pixelVal_in_1_4;
      end else if (10'hd8 == _T_25[9:0]) begin
        image_1_216 <= io_pixelVal_in_1_3;
      end else if (10'hd8 == _T_22[9:0]) begin
        image_1_216 <= io_pixelVal_in_1_2;
      end else if (10'hd8 == _T_19[9:0]) begin
        image_1_216 <= io_pixelVal_in_1_1;
      end else if (10'hd8 == _T_15[9:0]) begin
        image_1_216 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_217 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd9 == _T_37[9:0]) begin
        image_1_217 <= io_pixelVal_in_1_7;
      end else if (10'hd9 == _T_34[9:0]) begin
        image_1_217 <= io_pixelVal_in_1_6;
      end else if (10'hd9 == _T_31[9:0]) begin
        image_1_217 <= io_pixelVal_in_1_5;
      end else if (10'hd9 == _T_28[9:0]) begin
        image_1_217 <= io_pixelVal_in_1_4;
      end else if (10'hd9 == _T_25[9:0]) begin
        image_1_217 <= io_pixelVal_in_1_3;
      end else if (10'hd9 == _T_22[9:0]) begin
        image_1_217 <= io_pixelVal_in_1_2;
      end else if (10'hd9 == _T_19[9:0]) begin
        image_1_217 <= io_pixelVal_in_1_1;
      end else if (10'hd9 == _T_15[9:0]) begin
        image_1_217 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_218 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hda == _T_37[9:0]) begin
        image_1_218 <= io_pixelVal_in_1_7;
      end else if (10'hda == _T_34[9:0]) begin
        image_1_218 <= io_pixelVal_in_1_6;
      end else if (10'hda == _T_31[9:0]) begin
        image_1_218 <= io_pixelVal_in_1_5;
      end else if (10'hda == _T_28[9:0]) begin
        image_1_218 <= io_pixelVal_in_1_4;
      end else if (10'hda == _T_25[9:0]) begin
        image_1_218 <= io_pixelVal_in_1_3;
      end else if (10'hda == _T_22[9:0]) begin
        image_1_218 <= io_pixelVal_in_1_2;
      end else if (10'hda == _T_19[9:0]) begin
        image_1_218 <= io_pixelVal_in_1_1;
      end else if (10'hda == _T_15[9:0]) begin
        image_1_218 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_219 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hdb == _T_37[9:0]) begin
        image_1_219 <= io_pixelVal_in_1_7;
      end else if (10'hdb == _T_34[9:0]) begin
        image_1_219 <= io_pixelVal_in_1_6;
      end else if (10'hdb == _T_31[9:0]) begin
        image_1_219 <= io_pixelVal_in_1_5;
      end else if (10'hdb == _T_28[9:0]) begin
        image_1_219 <= io_pixelVal_in_1_4;
      end else if (10'hdb == _T_25[9:0]) begin
        image_1_219 <= io_pixelVal_in_1_3;
      end else if (10'hdb == _T_22[9:0]) begin
        image_1_219 <= io_pixelVal_in_1_2;
      end else if (10'hdb == _T_19[9:0]) begin
        image_1_219 <= io_pixelVal_in_1_1;
      end else if (10'hdb == _T_15[9:0]) begin
        image_1_219 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_220 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hdc == _T_37[9:0]) begin
        image_1_220 <= io_pixelVal_in_1_7;
      end else if (10'hdc == _T_34[9:0]) begin
        image_1_220 <= io_pixelVal_in_1_6;
      end else if (10'hdc == _T_31[9:0]) begin
        image_1_220 <= io_pixelVal_in_1_5;
      end else if (10'hdc == _T_28[9:0]) begin
        image_1_220 <= io_pixelVal_in_1_4;
      end else if (10'hdc == _T_25[9:0]) begin
        image_1_220 <= io_pixelVal_in_1_3;
      end else if (10'hdc == _T_22[9:0]) begin
        image_1_220 <= io_pixelVal_in_1_2;
      end else if (10'hdc == _T_19[9:0]) begin
        image_1_220 <= io_pixelVal_in_1_1;
      end else if (10'hdc == _T_15[9:0]) begin
        image_1_220 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_221 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hdd == _T_37[9:0]) begin
        image_1_221 <= io_pixelVal_in_1_7;
      end else if (10'hdd == _T_34[9:0]) begin
        image_1_221 <= io_pixelVal_in_1_6;
      end else if (10'hdd == _T_31[9:0]) begin
        image_1_221 <= io_pixelVal_in_1_5;
      end else if (10'hdd == _T_28[9:0]) begin
        image_1_221 <= io_pixelVal_in_1_4;
      end else if (10'hdd == _T_25[9:0]) begin
        image_1_221 <= io_pixelVal_in_1_3;
      end else if (10'hdd == _T_22[9:0]) begin
        image_1_221 <= io_pixelVal_in_1_2;
      end else if (10'hdd == _T_19[9:0]) begin
        image_1_221 <= io_pixelVal_in_1_1;
      end else if (10'hdd == _T_15[9:0]) begin
        image_1_221 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_222 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hde == _T_37[9:0]) begin
        image_1_222 <= io_pixelVal_in_1_7;
      end else if (10'hde == _T_34[9:0]) begin
        image_1_222 <= io_pixelVal_in_1_6;
      end else if (10'hde == _T_31[9:0]) begin
        image_1_222 <= io_pixelVal_in_1_5;
      end else if (10'hde == _T_28[9:0]) begin
        image_1_222 <= io_pixelVal_in_1_4;
      end else if (10'hde == _T_25[9:0]) begin
        image_1_222 <= io_pixelVal_in_1_3;
      end else if (10'hde == _T_22[9:0]) begin
        image_1_222 <= io_pixelVal_in_1_2;
      end else if (10'hde == _T_19[9:0]) begin
        image_1_222 <= io_pixelVal_in_1_1;
      end else if (10'hde == _T_15[9:0]) begin
        image_1_222 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_223 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hdf == _T_37[9:0]) begin
        image_1_223 <= io_pixelVal_in_1_7;
      end else if (10'hdf == _T_34[9:0]) begin
        image_1_223 <= io_pixelVal_in_1_6;
      end else if (10'hdf == _T_31[9:0]) begin
        image_1_223 <= io_pixelVal_in_1_5;
      end else if (10'hdf == _T_28[9:0]) begin
        image_1_223 <= io_pixelVal_in_1_4;
      end else if (10'hdf == _T_25[9:0]) begin
        image_1_223 <= io_pixelVal_in_1_3;
      end else if (10'hdf == _T_22[9:0]) begin
        image_1_223 <= io_pixelVal_in_1_2;
      end else if (10'hdf == _T_19[9:0]) begin
        image_1_223 <= io_pixelVal_in_1_1;
      end else if (10'hdf == _T_15[9:0]) begin
        image_1_223 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_224 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he0 == _T_37[9:0]) begin
        image_1_224 <= io_pixelVal_in_1_7;
      end else if (10'he0 == _T_34[9:0]) begin
        image_1_224 <= io_pixelVal_in_1_6;
      end else if (10'he0 == _T_31[9:0]) begin
        image_1_224 <= io_pixelVal_in_1_5;
      end else if (10'he0 == _T_28[9:0]) begin
        image_1_224 <= io_pixelVal_in_1_4;
      end else if (10'he0 == _T_25[9:0]) begin
        image_1_224 <= io_pixelVal_in_1_3;
      end else if (10'he0 == _T_22[9:0]) begin
        image_1_224 <= io_pixelVal_in_1_2;
      end else if (10'he0 == _T_19[9:0]) begin
        image_1_224 <= io_pixelVal_in_1_1;
      end else if (10'he0 == _T_15[9:0]) begin
        image_1_224 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_225 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he1 == _T_37[9:0]) begin
        image_1_225 <= io_pixelVal_in_1_7;
      end else if (10'he1 == _T_34[9:0]) begin
        image_1_225 <= io_pixelVal_in_1_6;
      end else if (10'he1 == _T_31[9:0]) begin
        image_1_225 <= io_pixelVal_in_1_5;
      end else if (10'he1 == _T_28[9:0]) begin
        image_1_225 <= io_pixelVal_in_1_4;
      end else if (10'he1 == _T_25[9:0]) begin
        image_1_225 <= io_pixelVal_in_1_3;
      end else if (10'he1 == _T_22[9:0]) begin
        image_1_225 <= io_pixelVal_in_1_2;
      end else if (10'he1 == _T_19[9:0]) begin
        image_1_225 <= io_pixelVal_in_1_1;
      end else if (10'he1 == _T_15[9:0]) begin
        image_1_225 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_226 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he2 == _T_37[9:0]) begin
        image_1_226 <= io_pixelVal_in_1_7;
      end else if (10'he2 == _T_34[9:0]) begin
        image_1_226 <= io_pixelVal_in_1_6;
      end else if (10'he2 == _T_31[9:0]) begin
        image_1_226 <= io_pixelVal_in_1_5;
      end else if (10'he2 == _T_28[9:0]) begin
        image_1_226 <= io_pixelVal_in_1_4;
      end else if (10'he2 == _T_25[9:0]) begin
        image_1_226 <= io_pixelVal_in_1_3;
      end else if (10'he2 == _T_22[9:0]) begin
        image_1_226 <= io_pixelVal_in_1_2;
      end else if (10'he2 == _T_19[9:0]) begin
        image_1_226 <= io_pixelVal_in_1_1;
      end else if (10'he2 == _T_15[9:0]) begin
        image_1_226 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_227 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he3 == _T_37[9:0]) begin
        image_1_227 <= io_pixelVal_in_1_7;
      end else if (10'he3 == _T_34[9:0]) begin
        image_1_227 <= io_pixelVal_in_1_6;
      end else if (10'he3 == _T_31[9:0]) begin
        image_1_227 <= io_pixelVal_in_1_5;
      end else if (10'he3 == _T_28[9:0]) begin
        image_1_227 <= io_pixelVal_in_1_4;
      end else if (10'he3 == _T_25[9:0]) begin
        image_1_227 <= io_pixelVal_in_1_3;
      end else if (10'he3 == _T_22[9:0]) begin
        image_1_227 <= io_pixelVal_in_1_2;
      end else if (10'he3 == _T_19[9:0]) begin
        image_1_227 <= io_pixelVal_in_1_1;
      end else if (10'he3 == _T_15[9:0]) begin
        image_1_227 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_228 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he4 == _T_37[9:0]) begin
        image_1_228 <= io_pixelVal_in_1_7;
      end else if (10'he4 == _T_34[9:0]) begin
        image_1_228 <= io_pixelVal_in_1_6;
      end else if (10'he4 == _T_31[9:0]) begin
        image_1_228 <= io_pixelVal_in_1_5;
      end else if (10'he4 == _T_28[9:0]) begin
        image_1_228 <= io_pixelVal_in_1_4;
      end else if (10'he4 == _T_25[9:0]) begin
        image_1_228 <= io_pixelVal_in_1_3;
      end else if (10'he4 == _T_22[9:0]) begin
        image_1_228 <= io_pixelVal_in_1_2;
      end else if (10'he4 == _T_19[9:0]) begin
        image_1_228 <= io_pixelVal_in_1_1;
      end else if (10'he4 == _T_15[9:0]) begin
        image_1_228 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_229 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he5 == _T_37[9:0]) begin
        image_1_229 <= io_pixelVal_in_1_7;
      end else if (10'he5 == _T_34[9:0]) begin
        image_1_229 <= io_pixelVal_in_1_6;
      end else if (10'he5 == _T_31[9:0]) begin
        image_1_229 <= io_pixelVal_in_1_5;
      end else if (10'he5 == _T_28[9:0]) begin
        image_1_229 <= io_pixelVal_in_1_4;
      end else if (10'he5 == _T_25[9:0]) begin
        image_1_229 <= io_pixelVal_in_1_3;
      end else if (10'he5 == _T_22[9:0]) begin
        image_1_229 <= io_pixelVal_in_1_2;
      end else if (10'he5 == _T_19[9:0]) begin
        image_1_229 <= io_pixelVal_in_1_1;
      end else if (10'he5 == _T_15[9:0]) begin
        image_1_229 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_230 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he6 == _T_37[9:0]) begin
        image_1_230 <= io_pixelVal_in_1_7;
      end else if (10'he6 == _T_34[9:0]) begin
        image_1_230 <= io_pixelVal_in_1_6;
      end else if (10'he6 == _T_31[9:0]) begin
        image_1_230 <= io_pixelVal_in_1_5;
      end else if (10'he6 == _T_28[9:0]) begin
        image_1_230 <= io_pixelVal_in_1_4;
      end else if (10'he6 == _T_25[9:0]) begin
        image_1_230 <= io_pixelVal_in_1_3;
      end else if (10'he6 == _T_22[9:0]) begin
        image_1_230 <= io_pixelVal_in_1_2;
      end else if (10'he6 == _T_19[9:0]) begin
        image_1_230 <= io_pixelVal_in_1_1;
      end else if (10'he6 == _T_15[9:0]) begin
        image_1_230 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_231 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he7 == _T_37[9:0]) begin
        image_1_231 <= io_pixelVal_in_1_7;
      end else if (10'he7 == _T_34[9:0]) begin
        image_1_231 <= io_pixelVal_in_1_6;
      end else if (10'he7 == _T_31[9:0]) begin
        image_1_231 <= io_pixelVal_in_1_5;
      end else if (10'he7 == _T_28[9:0]) begin
        image_1_231 <= io_pixelVal_in_1_4;
      end else if (10'he7 == _T_25[9:0]) begin
        image_1_231 <= io_pixelVal_in_1_3;
      end else if (10'he7 == _T_22[9:0]) begin
        image_1_231 <= io_pixelVal_in_1_2;
      end else if (10'he7 == _T_19[9:0]) begin
        image_1_231 <= io_pixelVal_in_1_1;
      end else if (10'he7 == _T_15[9:0]) begin
        image_1_231 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_232 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he8 == _T_37[9:0]) begin
        image_1_232 <= io_pixelVal_in_1_7;
      end else if (10'he8 == _T_34[9:0]) begin
        image_1_232 <= io_pixelVal_in_1_6;
      end else if (10'he8 == _T_31[9:0]) begin
        image_1_232 <= io_pixelVal_in_1_5;
      end else if (10'he8 == _T_28[9:0]) begin
        image_1_232 <= io_pixelVal_in_1_4;
      end else if (10'he8 == _T_25[9:0]) begin
        image_1_232 <= io_pixelVal_in_1_3;
      end else if (10'he8 == _T_22[9:0]) begin
        image_1_232 <= io_pixelVal_in_1_2;
      end else if (10'he8 == _T_19[9:0]) begin
        image_1_232 <= io_pixelVal_in_1_1;
      end else if (10'he8 == _T_15[9:0]) begin
        image_1_232 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_233 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he9 == _T_37[9:0]) begin
        image_1_233 <= io_pixelVal_in_1_7;
      end else if (10'he9 == _T_34[9:0]) begin
        image_1_233 <= io_pixelVal_in_1_6;
      end else if (10'he9 == _T_31[9:0]) begin
        image_1_233 <= io_pixelVal_in_1_5;
      end else if (10'he9 == _T_28[9:0]) begin
        image_1_233 <= io_pixelVal_in_1_4;
      end else if (10'he9 == _T_25[9:0]) begin
        image_1_233 <= io_pixelVal_in_1_3;
      end else if (10'he9 == _T_22[9:0]) begin
        image_1_233 <= io_pixelVal_in_1_2;
      end else if (10'he9 == _T_19[9:0]) begin
        image_1_233 <= io_pixelVal_in_1_1;
      end else if (10'he9 == _T_15[9:0]) begin
        image_1_233 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_234 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hea == _T_37[9:0]) begin
        image_1_234 <= io_pixelVal_in_1_7;
      end else if (10'hea == _T_34[9:0]) begin
        image_1_234 <= io_pixelVal_in_1_6;
      end else if (10'hea == _T_31[9:0]) begin
        image_1_234 <= io_pixelVal_in_1_5;
      end else if (10'hea == _T_28[9:0]) begin
        image_1_234 <= io_pixelVal_in_1_4;
      end else if (10'hea == _T_25[9:0]) begin
        image_1_234 <= io_pixelVal_in_1_3;
      end else if (10'hea == _T_22[9:0]) begin
        image_1_234 <= io_pixelVal_in_1_2;
      end else if (10'hea == _T_19[9:0]) begin
        image_1_234 <= io_pixelVal_in_1_1;
      end else if (10'hea == _T_15[9:0]) begin
        image_1_234 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_235 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'heb == _T_37[9:0]) begin
        image_1_235 <= io_pixelVal_in_1_7;
      end else if (10'heb == _T_34[9:0]) begin
        image_1_235 <= io_pixelVal_in_1_6;
      end else if (10'heb == _T_31[9:0]) begin
        image_1_235 <= io_pixelVal_in_1_5;
      end else if (10'heb == _T_28[9:0]) begin
        image_1_235 <= io_pixelVal_in_1_4;
      end else if (10'heb == _T_25[9:0]) begin
        image_1_235 <= io_pixelVal_in_1_3;
      end else if (10'heb == _T_22[9:0]) begin
        image_1_235 <= io_pixelVal_in_1_2;
      end else if (10'heb == _T_19[9:0]) begin
        image_1_235 <= io_pixelVal_in_1_1;
      end else if (10'heb == _T_15[9:0]) begin
        image_1_235 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_236 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hec == _T_37[9:0]) begin
        image_1_236 <= io_pixelVal_in_1_7;
      end else if (10'hec == _T_34[9:0]) begin
        image_1_236 <= io_pixelVal_in_1_6;
      end else if (10'hec == _T_31[9:0]) begin
        image_1_236 <= io_pixelVal_in_1_5;
      end else if (10'hec == _T_28[9:0]) begin
        image_1_236 <= io_pixelVal_in_1_4;
      end else if (10'hec == _T_25[9:0]) begin
        image_1_236 <= io_pixelVal_in_1_3;
      end else if (10'hec == _T_22[9:0]) begin
        image_1_236 <= io_pixelVal_in_1_2;
      end else if (10'hec == _T_19[9:0]) begin
        image_1_236 <= io_pixelVal_in_1_1;
      end else if (10'hec == _T_15[9:0]) begin
        image_1_236 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_237 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hed == _T_37[9:0]) begin
        image_1_237 <= io_pixelVal_in_1_7;
      end else if (10'hed == _T_34[9:0]) begin
        image_1_237 <= io_pixelVal_in_1_6;
      end else if (10'hed == _T_31[9:0]) begin
        image_1_237 <= io_pixelVal_in_1_5;
      end else if (10'hed == _T_28[9:0]) begin
        image_1_237 <= io_pixelVal_in_1_4;
      end else if (10'hed == _T_25[9:0]) begin
        image_1_237 <= io_pixelVal_in_1_3;
      end else if (10'hed == _T_22[9:0]) begin
        image_1_237 <= io_pixelVal_in_1_2;
      end else if (10'hed == _T_19[9:0]) begin
        image_1_237 <= io_pixelVal_in_1_1;
      end else if (10'hed == _T_15[9:0]) begin
        image_1_237 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_238 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hee == _T_37[9:0]) begin
        image_1_238 <= io_pixelVal_in_1_7;
      end else if (10'hee == _T_34[9:0]) begin
        image_1_238 <= io_pixelVal_in_1_6;
      end else if (10'hee == _T_31[9:0]) begin
        image_1_238 <= io_pixelVal_in_1_5;
      end else if (10'hee == _T_28[9:0]) begin
        image_1_238 <= io_pixelVal_in_1_4;
      end else if (10'hee == _T_25[9:0]) begin
        image_1_238 <= io_pixelVal_in_1_3;
      end else if (10'hee == _T_22[9:0]) begin
        image_1_238 <= io_pixelVal_in_1_2;
      end else if (10'hee == _T_19[9:0]) begin
        image_1_238 <= io_pixelVal_in_1_1;
      end else if (10'hee == _T_15[9:0]) begin
        image_1_238 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_239 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hef == _T_37[9:0]) begin
        image_1_239 <= io_pixelVal_in_1_7;
      end else if (10'hef == _T_34[9:0]) begin
        image_1_239 <= io_pixelVal_in_1_6;
      end else if (10'hef == _T_31[9:0]) begin
        image_1_239 <= io_pixelVal_in_1_5;
      end else if (10'hef == _T_28[9:0]) begin
        image_1_239 <= io_pixelVal_in_1_4;
      end else if (10'hef == _T_25[9:0]) begin
        image_1_239 <= io_pixelVal_in_1_3;
      end else if (10'hef == _T_22[9:0]) begin
        image_1_239 <= io_pixelVal_in_1_2;
      end else if (10'hef == _T_19[9:0]) begin
        image_1_239 <= io_pixelVal_in_1_1;
      end else if (10'hef == _T_15[9:0]) begin
        image_1_239 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_240 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf0 == _T_37[9:0]) begin
        image_1_240 <= io_pixelVal_in_1_7;
      end else if (10'hf0 == _T_34[9:0]) begin
        image_1_240 <= io_pixelVal_in_1_6;
      end else if (10'hf0 == _T_31[9:0]) begin
        image_1_240 <= io_pixelVal_in_1_5;
      end else if (10'hf0 == _T_28[9:0]) begin
        image_1_240 <= io_pixelVal_in_1_4;
      end else if (10'hf0 == _T_25[9:0]) begin
        image_1_240 <= io_pixelVal_in_1_3;
      end else if (10'hf0 == _T_22[9:0]) begin
        image_1_240 <= io_pixelVal_in_1_2;
      end else if (10'hf0 == _T_19[9:0]) begin
        image_1_240 <= io_pixelVal_in_1_1;
      end else if (10'hf0 == _T_15[9:0]) begin
        image_1_240 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_241 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf1 == _T_37[9:0]) begin
        image_1_241 <= io_pixelVal_in_1_7;
      end else if (10'hf1 == _T_34[9:0]) begin
        image_1_241 <= io_pixelVal_in_1_6;
      end else if (10'hf1 == _T_31[9:0]) begin
        image_1_241 <= io_pixelVal_in_1_5;
      end else if (10'hf1 == _T_28[9:0]) begin
        image_1_241 <= io_pixelVal_in_1_4;
      end else if (10'hf1 == _T_25[9:0]) begin
        image_1_241 <= io_pixelVal_in_1_3;
      end else if (10'hf1 == _T_22[9:0]) begin
        image_1_241 <= io_pixelVal_in_1_2;
      end else if (10'hf1 == _T_19[9:0]) begin
        image_1_241 <= io_pixelVal_in_1_1;
      end else if (10'hf1 == _T_15[9:0]) begin
        image_1_241 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_242 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf2 == _T_37[9:0]) begin
        image_1_242 <= io_pixelVal_in_1_7;
      end else if (10'hf2 == _T_34[9:0]) begin
        image_1_242 <= io_pixelVal_in_1_6;
      end else if (10'hf2 == _T_31[9:0]) begin
        image_1_242 <= io_pixelVal_in_1_5;
      end else if (10'hf2 == _T_28[9:0]) begin
        image_1_242 <= io_pixelVal_in_1_4;
      end else if (10'hf2 == _T_25[9:0]) begin
        image_1_242 <= io_pixelVal_in_1_3;
      end else if (10'hf2 == _T_22[9:0]) begin
        image_1_242 <= io_pixelVal_in_1_2;
      end else if (10'hf2 == _T_19[9:0]) begin
        image_1_242 <= io_pixelVal_in_1_1;
      end else if (10'hf2 == _T_15[9:0]) begin
        image_1_242 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_243 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf3 == _T_37[9:0]) begin
        image_1_243 <= io_pixelVal_in_1_7;
      end else if (10'hf3 == _T_34[9:0]) begin
        image_1_243 <= io_pixelVal_in_1_6;
      end else if (10'hf3 == _T_31[9:0]) begin
        image_1_243 <= io_pixelVal_in_1_5;
      end else if (10'hf3 == _T_28[9:0]) begin
        image_1_243 <= io_pixelVal_in_1_4;
      end else if (10'hf3 == _T_25[9:0]) begin
        image_1_243 <= io_pixelVal_in_1_3;
      end else if (10'hf3 == _T_22[9:0]) begin
        image_1_243 <= io_pixelVal_in_1_2;
      end else if (10'hf3 == _T_19[9:0]) begin
        image_1_243 <= io_pixelVal_in_1_1;
      end else if (10'hf3 == _T_15[9:0]) begin
        image_1_243 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_244 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf4 == _T_37[9:0]) begin
        image_1_244 <= io_pixelVal_in_1_7;
      end else if (10'hf4 == _T_34[9:0]) begin
        image_1_244 <= io_pixelVal_in_1_6;
      end else if (10'hf4 == _T_31[9:0]) begin
        image_1_244 <= io_pixelVal_in_1_5;
      end else if (10'hf4 == _T_28[9:0]) begin
        image_1_244 <= io_pixelVal_in_1_4;
      end else if (10'hf4 == _T_25[9:0]) begin
        image_1_244 <= io_pixelVal_in_1_3;
      end else if (10'hf4 == _T_22[9:0]) begin
        image_1_244 <= io_pixelVal_in_1_2;
      end else if (10'hf4 == _T_19[9:0]) begin
        image_1_244 <= io_pixelVal_in_1_1;
      end else if (10'hf4 == _T_15[9:0]) begin
        image_1_244 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_245 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf5 == _T_37[9:0]) begin
        image_1_245 <= io_pixelVal_in_1_7;
      end else if (10'hf5 == _T_34[9:0]) begin
        image_1_245 <= io_pixelVal_in_1_6;
      end else if (10'hf5 == _T_31[9:0]) begin
        image_1_245 <= io_pixelVal_in_1_5;
      end else if (10'hf5 == _T_28[9:0]) begin
        image_1_245 <= io_pixelVal_in_1_4;
      end else if (10'hf5 == _T_25[9:0]) begin
        image_1_245 <= io_pixelVal_in_1_3;
      end else if (10'hf5 == _T_22[9:0]) begin
        image_1_245 <= io_pixelVal_in_1_2;
      end else if (10'hf5 == _T_19[9:0]) begin
        image_1_245 <= io_pixelVal_in_1_1;
      end else if (10'hf5 == _T_15[9:0]) begin
        image_1_245 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_246 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf6 == _T_37[9:0]) begin
        image_1_246 <= io_pixelVal_in_1_7;
      end else if (10'hf6 == _T_34[9:0]) begin
        image_1_246 <= io_pixelVal_in_1_6;
      end else if (10'hf6 == _T_31[9:0]) begin
        image_1_246 <= io_pixelVal_in_1_5;
      end else if (10'hf6 == _T_28[9:0]) begin
        image_1_246 <= io_pixelVal_in_1_4;
      end else if (10'hf6 == _T_25[9:0]) begin
        image_1_246 <= io_pixelVal_in_1_3;
      end else if (10'hf6 == _T_22[9:0]) begin
        image_1_246 <= io_pixelVal_in_1_2;
      end else if (10'hf6 == _T_19[9:0]) begin
        image_1_246 <= io_pixelVal_in_1_1;
      end else if (10'hf6 == _T_15[9:0]) begin
        image_1_246 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_247 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf7 == _T_37[9:0]) begin
        image_1_247 <= io_pixelVal_in_1_7;
      end else if (10'hf7 == _T_34[9:0]) begin
        image_1_247 <= io_pixelVal_in_1_6;
      end else if (10'hf7 == _T_31[9:0]) begin
        image_1_247 <= io_pixelVal_in_1_5;
      end else if (10'hf7 == _T_28[9:0]) begin
        image_1_247 <= io_pixelVal_in_1_4;
      end else if (10'hf7 == _T_25[9:0]) begin
        image_1_247 <= io_pixelVal_in_1_3;
      end else if (10'hf7 == _T_22[9:0]) begin
        image_1_247 <= io_pixelVal_in_1_2;
      end else if (10'hf7 == _T_19[9:0]) begin
        image_1_247 <= io_pixelVal_in_1_1;
      end else if (10'hf7 == _T_15[9:0]) begin
        image_1_247 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_248 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf8 == _T_37[9:0]) begin
        image_1_248 <= io_pixelVal_in_1_7;
      end else if (10'hf8 == _T_34[9:0]) begin
        image_1_248 <= io_pixelVal_in_1_6;
      end else if (10'hf8 == _T_31[9:0]) begin
        image_1_248 <= io_pixelVal_in_1_5;
      end else if (10'hf8 == _T_28[9:0]) begin
        image_1_248 <= io_pixelVal_in_1_4;
      end else if (10'hf8 == _T_25[9:0]) begin
        image_1_248 <= io_pixelVal_in_1_3;
      end else if (10'hf8 == _T_22[9:0]) begin
        image_1_248 <= io_pixelVal_in_1_2;
      end else if (10'hf8 == _T_19[9:0]) begin
        image_1_248 <= io_pixelVal_in_1_1;
      end else if (10'hf8 == _T_15[9:0]) begin
        image_1_248 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_249 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf9 == _T_37[9:0]) begin
        image_1_249 <= io_pixelVal_in_1_7;
      end else if (10'hf9 == _T_34[9:0]) begin
        image_1_249 <= io_pixelVal_in_1_6;
      end else if (10'hf9 == _T_31[9:0]) begin
        image_1_249 <= io_pixelVal_in_1_5;
      end else if (10'hf9 == _T_28[9:0]) begin
        image_1_249 <= io_pixelVal_in_1_4;
      end else if (10'hf9 == _T_25[9:0]) begin
        image_1_249 <= io_pixelVal_in_1_3;
      end else if (10'hf9 == _T_22[9:0]) begin
        image_1_249 <= io_pixelVal_in_1_2;
      end else if (10'hf9 == _T_19[9:0]) begin
        image_1_249 <= io_pixelVal_in_1_1;
      end else if (10'hf9 == _T_15[9:0]) begin
        image_1_249 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_250 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hfa == _T_37[9:0]) begin
        image_1_250 <= io_pixelVal_in_1_7;
      end else if (10'hfa == _T_34[9:0]) begin
        image_1_250 <= io_pixelVal_in_1_6;
      end else if (10'hfa == _T_31[9:0]) begin
        image_1_250 <= io_pixelVal_in_1_5;
      end else if (10'hfa == _T_28[9:0]) begin
        image_1_250 <= io_pixelVal_in_1_4;
      end else if (10'hfa == _T_25[9:0]) begin
        image_1_250 <= io_pixelVal_in_1_3;
      end else if (10'hfa == _T_22[9:0]) begin
        image_1_250 <= io_pixelVal_in_1_2;
      end else if (10'hfa == _T_19[9:0]) begin
        image_1_250 <= io_pixelVal_in_1_1;
      end else if (10'hfa == _T_15[9:0]) begin
        image_1_250 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_251 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hfb == _T_37[9:0]) begin
        image_1_251 <= io_pixelVal_in_1_7;
      end else if (10'hfb == _T_34[9:0]) begin
        image_1_251 <= io_pixelVal_in_1_6;
      end else if (10'hfb == _T_31[9:0]) begin
        image_1_251 <= io_pixelVal_in_1_5;
      end else if (10'hfb == _T_28[9:0]) begin
        image_1_251 <= io_pixelVal_in_1_4;
      end else if (10'hfb == _T_25[9:0]) begin
        image_1_251 <= io_pixelVal_in_1_3;
      end else if (10'hfb == _T_22[9:0]) begin
        image_1_251 <= io_pixelVal_in_1_2;
      end else if (10'hfb == _T_19[9:0]) begin
        image_1_251 <= io_pixelVal_in_1_1;
      end else if (10'hfb == _T_15[9:0]) begin
        image_1_251 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_252 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hfc == _T_37[9:0]) begin
        image_1_252 <= io_pixelVal_in_1_7;
      end else if (10'hfc == _T_34[9:0]) begin
        image_1_252 <= io_pixelVal_in_1_6;
      end else if (10'hfc == _T_31[9:0]) begin
        image_1_252 <= io_pixelVal_in_1_5;
      end else if (10'hfc == _T_28[9:0]) begin
        image_1_252 <= io_pixelVal_in_1_4;
      end else if (10'hfc == _T_25[9:0]) begin
        image_1_252 <= io_pixelVal_in_1_3;
      end else if (10'hfc == _T_22[9:0]) begin
        image_1_252 <= io_pixelVal_in_1_2;
      end else if (10'hfc == _T_19[9:0]) begin
        image_1_252 <= io_pixelVal_in_1_1;
      end else if (10'hfc == _T_15[9:0]) begin
        image_1_252 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_253 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hfd == _T_37[9:0]) begin
        image_1_253 <= io_pixelVal_in_1_7;
      end else if (10'hfd == _T_34[9:0]) begin
        image_1_253 <= io_pixelVal_in_1_6;
      end else if (10'hfd == _T_31[9:0]) begin
        image_1_253 <= io_pixelVal_in_1_5;
      end else if (10'hfd == _T_28[9:0]) begin
        image_1_253 <= io_pixelVal_in_1_4;
      end else if (10'hfd == _T_25[9:0]) begin
        image_1_253 <= io_pixelVal_in_1_3;
      end else if (10'hfd == _T_22[9:0]) begin
        image_1_253 <= io_pixelVal_in_1_2;
      end else if (10'hfd == _T_19[9:0]) begin
        image_1_253 <= io_pixelVal_in_1_1;
      end else if (10'hfd == _T_15[9:0]) begin
        image_1_253 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_254 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hfe == _T_37[9:0]) begin
        image_1_254 <= io_pixelVal_in_1_7;
      end else if (10'hfe == _T_34[9:0]) begin
        image_1_254 <= io_pixelVal_in_1_6;
      end else if (10'hfe == _T_31[9:0]) begin
        image_1_254 <= io_pixelVal_in_1_5;
      end else if (10'hfe == _T_28[9:0]) begin
        image_1_254 <= io_pixelVal_in_1_4;
      end else if (10'hfe == _T_25[9:0]) begin
        image_1_254 <= io_pixelVal_in_1_3;
      end else if (10'hfe == _T_22[9:0]) begin
        image_1_254 <= io_pixelVal_in_1_2;
      end else if (10'hfe == _T_19[9:0]) begin
        image_1_254 <= io_pixelVal_in_1_1;
      end else if (10'hfe == _T_15[9:0]) begin
        image_1_254 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_255 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hff == _T_37[9:0]) begin
        image_1_255 <= io_pixelVal_in_1_7;
      end else if (10'hff == _T_34[9:0]) begin
        image_1_255 <= io_pixelVal_in_1_6;
      end else if (10'hff == _T_31[9:0]) begin
        image_1_255 <= io_pixelVal_in_1_5;
      end else if (10'hff == _T_28[9:0]) begin
        image_1_255 <= io_pixelVal_in_1_4;
      end else if (10'hff == _T_25[9:0]) begin
        image_1_255 <= io_pixelVal_in_1_3;
      end else if (10'hff == _T_22[9:0]) begin
        image_1_255 <= io_pixelVal_in_1_2;
      end else if (10'hff == _T_19[9:0]) begin
        image_1_255 <= io_pixelVal_in_1_1;
      end else if (10'hff == _T_15[9:0]) begin
        image_1_255 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_256 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h100 == _T_37[9:0]) begin
        image_1_256 <= io_pixelVal_in_1_7;
      end else if (10'h100 == _T_34[9:0]) begin
        image_1_256 <= io_pixelVal_in_1_6;
      end else if (10'h100 == _T_31[9:0]) begin
        image_1_256 <= io_pixelVal_in_1_5;
      end else if (10'h100 == _T_28[9:0]) begin
        image_1_256 <= io_pixelVal_in_1_4;
      end else if (10'h100 == _T_25[9:0]) begin
        image_1_256 <= io_pixelVal_in_1_3;
      end else if (10'h100 == _T_22[9:0]) begin
        image_1_256 <= io_pixelVal_in_1_2;
      end else if (10'h100 == _T_19[9:0]) begin
        image_1_256 <= io_pixelVal_in_1_1;
      end else if (10'h100 == _T_15[9:0]) begin
        image_1_256 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_257 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h101 == _T_37[9:0]) begin
        image_1_257 <= io_pixelVal_in_1_7;
      end else if (10'h101 == _T_34[9:0]) begin
        image_1_257 <= io_pixelVal_in_1_6;
      end else if (10'h101 == _T_31[9:0]) begin
        image_1_257 <= io_pixelVal_in_1_5;
      end else if (10'h101 == _T_28[9:0]) begin
        image_1_257 <= io_pixelVal_in_1_4;
      end else if (10'h101 == _T_25[9:0]) begin
        image_1_257 <= io_pixelVal_in_1_3;
      end else if (10'h101 == _T_22[9:0]) begin
        image_1_257 <= io_pixelVal_in_1_2;
      end else if (10'h101 == _T_19[9:0]) begin
        image_1_257 <= io_pixelVal_in_1_1;
      end else if (10'h101 == _T_15[9:0]) begin
        image_1_257 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_258 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h102 == _T_37[9:0]) begin
        image_1_258 <= io_pixelVal_in_1_7;
      end else if (10'h102 == _T_34[9:0]) begin
        image_1_258 <= io_pixelVal_in_1_6;
      end else if (10'h102 == _T_31[9:0]) begin
        image_1_258 <= io_pixelVal_in_1_5;
      end else if (10'h102 == _T_28[9:0]) begin
        image_1_258 <= io_pixelVal_in_1_4;
      end else if (10'h102 == _T_25[9:0]) begin
        image_1_258 <= io_pixelVal_in_1_3;
      end else if (10'h102 == _T_22[9:0]) begin
        image_1_258 <= io_pixelVal_in_1_2;
      end else if (10'h102 == _T_19[9:0]) begin
        image_1_258 <= io_pixelVal_in_1_1;
      end else if (10'h102 == _T_15[9:0]) begin
        image_1_258 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_259 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h103 == _T_37[9:0]) begin
        image_1_259 <= io_pixelVal_in_1_7;
      end else if (10'h103 == _T_34[9:0]) begin
        image_1_259 <= io_pixelVal_in_1_6;
      end else if (10'h103 == _T_31[9:0]) begin
        image_1_259 <= io_pixelVal_in_1_5;
      end else if (10'h103 == _T_28[9:0]) begin
        image_1_259 <= io_pixelVal_in_1_4;
      end else if (10'h103 == _T_25[9:0]) begin
        image_1_259 <= io_pixelVal_in_1_3;
      end else if (10'h103 == _T_22[9:0]) begin
        image_1_259 <= io_pixelVal_in_1_2;
      end else if (10'h103 == _T_19[9:0]) begin
        image_1_259 <= io_pixelVal_in_1_1;
      end else if (10'h103 == _T_15[9:0]) begin
        image_1_259 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_260 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h104 == _T_37[9:0]) begin
        image_1_260 <= io_pixelVal_in_1_7;
      end else if (10'h104 == _T_34[9:0]) begin
        image_1_260 <= io_pixelVal_in_1_6;
      end else if (10'h104 == _T_31[9:0]) begin
        image_1_260 <= io_pixelVal_in_1_5;
      end else if (10'h104 == _T_28[9:0]) begin
        image_1_260 <= io_pixelVal_in_1_4;
      end else if (10'h104 == _T_25[9:0]) begin
        image_1_260 <= io_pixelVal_in_1_3;
      end else if (10'h104 == _T_22[9:0]) begin
        image_1_260 <= io_pixelVal_in_1_2;
      end else if (10'h104 == _T_19[9:0]) begin
        image_1_260 <= io_pixelVal_in_1_1;
      end else if (10'h104 == _T_15[9:0]) begin
        image_1_260 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_261 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h105 == _T_37[9:0]) begin
        image_1_261 <= io_pixelVal_in_1_7;
      end else if (10'h105 == _T_34[9:0]) begin
        image_1_261 <= io_pixelVal_in_1_6;
      end else if (10'h105 == _T_31[9:0]) begin
        image_1_261 <= io_pixelVal_in_1_5;
      end else if (10'h105 == _T_28[9:0]) begin
        image_1_261 <= io_pixelVal_in_1_4;
      end else if (10'h105 == _T_25[9:0]) begin
        image_1_261 <= io_pixelVal_in_1_3;
      end else if (10'h105 == _T_22[9:0]) begin
        image_1_261 <= io_pixelVal_in_1_2;
      end else if (10'h105 == _T_19[9:0]) begin
        image_1_261 <= io_pixelVal_in_1_1;
      end else if (10'h105 == _T_15[9:0]) begin
        image_1_261 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_262 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h106 == _T_37[9:0]) begin
        image_1_262 <= io_pixelVal_in_1_7;
      end else if (10'h106 == _T_34[9:0]) begin
        image_1_262 <= io_pixelVal_in_1_6;
      end else if (10'h106 == _T_31[9:0]) begin
        image_1_262 <= io_pixelVal_in_1_5;
      end else if (10'h106 == _T_28[9:0]) begin
        image_1_262 <= io_pixelVal_in_1_4;
      end else if (10'h106 == _T_25[9:0]) begin
        image_1_262 <= io_pixelVal_in_1_3;
      end else if (10'h106 == _T_22[9:0]) begin
        image_1_262 <= io_pixelVal_in_1_2;
      end else if (10'h106 == _T_19[9:0]) begin
        image_1_262 <= io_pixelVal_in_1_1;
      end else if (10'h106 == _T_15[9:0]) begin
        image_1_262 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_263 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h107 == _T_37[9:0]) begin
        image_1_263 <= io_pixelVal_in_1_7;
      end else if (10'h107 == _T_34[9:0]) begin
        image_1_263 <= io_pixelVal_in_1_6;
      end else if (10'h107 == _T_31[9:0]) begin
        image_1_263 <= io_pixelVal_in_1_5;
      end else if (10'h107 == _T_28[9:0]) begin
        image_1_263 <= io_pixelVal_in_1_4;
      end else if (10'h107 == _T_25[9:0]) begin
        image_1_263 <= io_pixelVal_in_1_3;
      end else if (10'h107 == _T_22[9:0]) begin
        image_1_263 <= io_pixelVal_in_1_2;
      end else if (10'h107 == _T_19[9:0]) begin
        image_1_263 <= io_pixelVal_in_1_1;
      end else if (10'h107 == _T_15[9:0]) begin
        image_1_263 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_264 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h108 == _T_37[9:0]) begin
        image_1_264 <= io_pixelVal_in_1_7;
      end else if (10'h108 == _T_34[9:0]) begin
        image_1_264 <= io_pixelVal_in_1_6;
      end else if (10'h108 == _T_31[9:0]) begin
        image_1_264 <= io_pixelVal_in_1_5;
      end else if (10'h108 == _T_28[9:0]) begin
        image_1_264 <= io_pixelVal_in_1_4;
      end else if (10'h108 == _T_25[9:0]) begin
        image_1_264 <= io_pixelVal_in_1_3;
      end else if (10'h108 == _T_22[9:0]) begin
        image_1_264 <= io_pixelVal_in_1_2;
      end else if (10'h108 == _T_19[9:0]) begin
        image_1_264 <= io_pixelVal_in_1_1;
      end else if (10'h108 == _T_15[9:0]) begin
        image_1_264 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_265 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h109 == _T_37[9:0]) begin
        image_1_265 <= io_pixelVal_in_1_7;
      end else if (10'h109 == _T_34[9:0]) begin
        image_1_265 <= io_pixelVal_in_1_6;
      end else if (10'h109 == _T_31[9:0]) begin
        image_1_265 <= io_pixelVal_in_1_5;
      end else if (10'h109 == _T_28[9:0]) begin
        image_1_265 <= io_pixelVal_in_1_4;
      end else if (10'h109 == _T_25[9:0]) begin
        image_1_265 <= io_pixelVal_in_1_3;
      end else if (10'h109 == _T_22[9:0]) begin
        image_1_265 <= io_pixelVal_in_1_2;
      end else if (10'h109 == _T_19[9:0]) begin
        image_1_265 <= io_pixelVal_in_1_1;
      end else if (10'h109 == _T_15[9:0]) begin
        image_1_265 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_266 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10a == _T_37[9:0]) begin
        image_1_266 <= io_pixelVal_in_1_7;
      end else if (10'h10a == _T_34[9:0]) begin
        image_1_266 <= io_pixelVal_in_1_6;
      end else if (10'h10a == _T_31[9:0]) begin
        image_1_266 <= io_pixelVal_in_1_5;
      end else if (10'h10a == _T_28[9:0]) begin
        image_1_266 <= io_pixelVal_in_1_4;
      end else if (10'h10a == _T_25[9:0]) begin
        image_1_266 <= io_pixelVal_in_1_3;
      end else if (10'h10a == _T_22[9:0]) begin
        image_1_266 <= io_pixelVal_in_1_2;
      end else if (10'h10a == _T_19[9:0]) begin
        image_1_266 <= io_pixelVal_in_1_1;
      end else if (10'h10a == _T_15[9:0]) begin
        image_1_266 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_267 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10b == _T_37[9:0]) begin
        image_1_267 <= io_pixelVal_in_1_7;
      end else if (10'h10b == _T_34[9:0]) begin
        image_1_267 <= io_pixelVal_in_1_6;
      end else if (10'h10b == _T_31[9:0]) begin
        image_1_267 <= io_pixelVal_in_1_5;
      end else if (10'h10b == _T_28[9:0]) begin
        image_1_267 <= io_pixelVal_in_1_4;
      end else if (10'h10b == _T_25[9:0]) begin
        image_1_267 <= io_pixelVal_in_1_3;
      end else if (10'h10b == _T_22[9:0]) begin
        image_1_267 <= io_pixelVal_in_1_2;
      end else if (10'h10b == _T_19[9:0]) begin
        image_1_267 <= io_pixelVal_in_1_1;
      end else if (10'h10b == _T_15[9:0]) begin
        image_1_267 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_268 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10c == _T_37[9:0]) begin
        image_1_268 <= io_pixelVal_in_1_7;
      end else if (10'h10c == _T_34[9:0]) begin
        image_1_268 <= io_pixelVal_in_1_6;
      end else if (10'h10c == _T_31[9:0]) begin
        image_1_268 <= io_pixelVal_in_1_5;
      end else if (10'h10c == _T_28[9:0]) begin
        image_1_268 <= io_pixelVal_in_1_4;
      end else if (10'h10c == _T_25[9:0]) begin
        image_1_268 <= io_pixelVal_in_1_3;
      end else if (10'h10c == _T_22[9:0]) begin
        image_1_268 <= io_pixelVal_in_1_2;
      end else if (10'h10c == _T_19[9:0]) begin
        image_1_268 <= io_pixelVal_in_1_1;
      end else if (10'h10c == _T_15[9:0]) begin
        image_1_268 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_269 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10d == _T_37[9:0]) begin
        image_1_269 <= io_pixelVal_in_1_7;
      end else if (10'h10d == _T_34[9:0]) begin
        image_1_269 <= io_pixelVal_in_1_6;
      end else if (10'h10d == _T_31[9:0]) begin
        image_1_269 <= io_pixelVal_in_1_5;
      end else if (10'h10d == _T_28[9:0]) begin
        image_1_269 <= io_pixelVal_in_1_4;
      end else if (10'h10d == _T_25[9:0]) begin
        image_1_269 <= io_pixelVal_in_1_3;
      end else if (10'h10d == _T_22[9:0]) begin
        image_1_269 <= io_pixelVal_in_1_2;
      end else if (10'h10d == _T_19[9:0]) begin
        image_1_269 <= io_pixelVal_in_1_1;
      end else if (10'h10d == _T_15[9:0]) begin
        image_1_269 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_270 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10e == _T_37[9:0]) begin
        image_1_270 <= io_pixelVal_in_1_7;
      end else if (10'h10e == _T_34[9:0]) begin
        image_1_270 <= io_pixelVal_in_1_6;
      end else if (10'h10e == _T_31[9:0]) begin
        image_1_270 <= io_pixelVal_in_1_5;
      end else if (10'h10e == _T_28[9:0]) begin
        image_1_270 <= io_pixelVal_in_1_4;
      end else if (10'h10e == _T_25[9:0]) begin
        image_1_270 <= io_pixelVal_in_1_3;
      end else if (10'h10e == _T_22[9:0]) begin
        image_1_270 <= io_pixelVal_in_1_2;
      end else if (10'h10e == _T_19[9:0]) begin
        image_1_270 <= io_pixelVal_in_1_1;
      end else if (10'h10e == _T_15[9:0]) begin
        image_1_270 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_271 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10f == _T_37[9:0]) begin
        image_1_271 <= io_pixelVal_in_1_7;
      end else if (10'h10f == _T_34[9:0]) begin
        image_1_271 <= io_pixelVal_in_1_6;
      end else if (10'h10f == _T_31[9:0]) begin
        image_1_271 <= io_pixelVal_in_1_5;
      end else if (10'h10f == _T_28[9:0]) begin
        image_1_271 <= io_pixelVal_in_1_4;
      end else if (10'h10f == _T_25[9:0]) begin
        image_1_271 <= io_pixelVal_in_1_3;
      end else if (10'h10f == _T_22[9:0]) begin
        image_1_271 <= io_pixelVal_in_1_2;
      end else if (10'h10f == _T_19[9:0]) begin
        image_1_271 <= io_pixelVal_in_1_1;
      end else if (10'h10f == _T_15[9:0]) begin
        image_1_271 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_272 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h110 == _T_37[9:0]) begin
        image_1_272 <= io_pixelVal_in_1_7;
      end else if (10'h110 == _T_34[9:0]) begin
        image_1_272 <= io_pixelVal_in_1_6;
      end else if (10'h110 == _T_31[9:0]) begin
        image_1_272 <= io_pixelVal_in_1_5;
      end else if (10'h110 == _T_28[9:0]) begin
        image_1_272 <= io_pixelVal_in_1_4;
      end else if (10'h110 == _T_25[9:0]) begin
        image_1_272 <= io_pixelVal_in_1_3;
      end else if (10'h110 == _T_22[9:0]) begin
        image_1_272 <= io_pixelVal_in_1_2;
      end else if (10'h110 == _T_19[9:0]) begin
        image_1_272 <= io_pixelVal_in_1_1;
      end else if (10'h110 == _T_15[9:0]) begin
        image_1_272 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_273 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h111 == _T_37[9:0]) begin
        image_1_273 <= io_pixelVal_in_1_7;
      end else if (10'h111 == _T_34[9:0]) begin
        image_1_273 <= io_pixelVal_in_1_6;
      end else if (10'h111 == _T_31[9:0]) begin
        image_1_273 <= io_pixelVal_in_1_5;
      end else if (10'h111 == _T_28[9:0]) begin
        image_1_273 <= io_pixelVal_in_1_4;
      end else if (10'h111 == _T_25[9:0]) begin
        image_1_273 <= io_pixelVal_in_1_3;
      end else if (10'h111 == _T_22[9:0]) begin
        image_1_273 <= io_pixelVal_in_1_2;
      end else if (10'h111 == _T_19[9:0]) begin
        image_1_273 <= io_pixelVal_in_1_1;
      end else if (10'h111 == _T_15[9:0]) begin
        image_1_273 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_274 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h112 == _T_37[9:0]) begin
        image_1_274 <= io_pixelVal_in_1_7;
      end else if (10'h112 == _T_34[9:0]) begin
        image_1_274 <= io_pixelVal_in_1_6;
      end else if (10'h112 == _T_31[9:0]) begin
        image_1_274 <= io_pixelVal_in_1_5;
      end else if (10'h112 == _T_28[9:0]) begin
        image_1_274 <= io_pixelVal_in_1_4;
      end else if (10'h112 == _T_25[9:0]) begin
        image_1_274 <= io_pixelVal_in_1_3;
      end else if (10'h112 == _T_22[9:0]) begin
        image_1_274 <= io_pixelVal_in_1_2;
      end else if (10'h112 == _T_19[9:0]) begin
        image_1_274 <= io_pixelVal_in_1_1;
      end else if (10'h112 == _T_15[9:0]) begin
        image_1_274 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_275 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h113 == _T_37[9:0]) begin
        image_1_275 <= io_pixelVal_in_1_7;
      end else if (10'h113 == _T_34[9:0]) begin
        image_1_275 <= io_pixelVal_in_1_6;
      end else if (10'h113 == _T_31[9:0]) begin
        image_1_275 <= io_pixelVal_in_1_5;
      end else if (10'h113 == _T_28[9:0]) begin
        image_1_275 <= io_pixelVal_in_1_4;
      end else if (10'h113 == _T_25[9:0]) begin
        image_1_275 <= io_pixelVal_in_1_3;
      end else if (10'h113 == _T_22[9:0]) begin
        image_1_275 <= io_pixelVal_in_1_2;
      end else if (10'h113 == _T_19[9:0]) begin
        image_1_275 <= io_pixelVal_in_1_1;
      end else if (10'h113 == _T_15[9:0]) begin
        image_1_275 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_276 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h114 == _T_37[9:0]) begin
        image_1_276 <= io_pixelVal_in_1_7;
      end else if (10'h114 == _T_34[9:0]) begin
        image_1_276 <= io_pixelVal_in_1_6;
      end else if (10'h114 == _T_31[9:0]) begin
        image_1_276 <= io_pixelVal_in_1_5;
      end else if (10'h114 == _T_28[9:0]) begin
        image_1_276 <= io_pixelVal_in_1_4;
      end else if (10'h114 == _T_25[9:0]) begin
        image_1_276 <= io_pixelVal_in_1_3;
      end else if (10'h114 == _T_22[9:0]) begin
        image_1_276 <= io_pixelVal_in_1_2;
      end else if (10'h114 == _T_19[9:0]) begin
        image_1_276 <= io_pixelVal_in_1_1;
      end else if (10'h114 == _T_15[9:0]) begin
        image_1_276 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_277 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h115 == _T_37[9:0]) begin
        image_1_277 <= io_pixelVal_in_1_7;
      end else if (10'h115 == _T_34[9:0]) begin
        image_1_277 <= io_pixelVal_in_1_6;
      end else if (10'h115 == _T_31[9:0]) begin
        image_1_277 <= io_pixelVal_in_1_5;
      end else if (10'h115 == _T_28[9:0]) begin
        image_1_277 <= io_pixelVal_in_1_4;
      end else if (10'h115 == _T_25[9:0]) begin
        image_1_277 <= io_pixelVal_in_1_3;
      end else if (10'h115 == _T_22[9:0]) begin
        image_1_277 <= io_pixelVal_in_1_2;
      end else if (10'h115 == _T_19[9:0]) begin
        image_1_277 <= io_pixelVal_in_1_1;
      end else if (10'h115 == _T_15[9:0]) begin
        image_1_277 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_278 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h116 == _T_37[9:0]) begin
        image_1_278 <= io_pixelVal_in_1_7;
      end else if (10'h116 == _T_34[9:0]) begin
        image_1_278 <= io_pixelVal_in_1_6;
      end else if (10'h116 == _T_31[9:0]) begin
        image_1_278 <= io_pixelVal_in_1_5;
      end else if (10'h116 == _T_28[9:0]) begin
        image_1_278 <= io_pixelVal_in_1_4;
      end else if (10'h116 == _T_25[9:0]) begin
        image_1_278 <= io_pixelVal_in_1_3;
      end else if (10'h116 == _T_22[9:0]) begin
        image_1_278 <= io_pixelVal_in_1_2;
      end else if (10'h116 == _T_19[9:0]) begin
        image_1_278 <= io_pixelVal_in_1_1;
      end else if (10'h116 == _T_15[9:0]) begin
        image_1_278 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_279 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h117 == _T_37[9:0]) begin
        image_1_279 <= io_pixelVal_in_1_7;
      end else if (10'h117 == _T_34[9:0]) begin
        image_1_279 <= io_pixelVal_in_1_6;
      end else if (10'h117 == _T_31[9:0]) begin
        image_1_279 <= io_pixelVal_in_1_5;
      end else if (10'h117 == _T_28[9:0]) begin
        image_1_279 <= io_pixelVal_in_1_4;
      end else if (10'h117 == _T_25[9:0]) begin
        image_1_279 <= io_pixelVal_in_1_3;
      end else if (10'h117 == _T_22[9:0]) begin
        image_1_279 <= io_pixelVal_in_1_2;
      end else if (10'h117 == _T_19[9:0]) begin
        image_1_279 <= io_pixelVal_in_1_1;
      end else if (10'h117 == _T_15[9:0]) begin
        image_1_279 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_280 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h118 == _T_37[9:0]) begin
        image_1_280 <= io_pixelVal_in_1_7;
      end else if (10'h118 == _T_34[9:0]) begin
        image_1_280 <= io_pixelVal_in_1_6;
      end else if (10'h118 == _T_31[9:0]) begin
        image_1_280 <= io_pixelVal_in_1_5;
      end else if (10'h118 == _T_28[9:0]) begin
        image_1_280 <= io_pixelVal_in_1_4;
      end else if (10'h118 == _T_25[9:0]) begin
        image_1_280 <= io_pixelVal_in_1_3;
      end else if (10'h118 == _T_22[9:0]) begin
        image_1_280 <= io_pixelVal_in_1_2;
      end else if (10'h118 == _T_19[9:0]) begin
        image_1_280 <= io_pixelVal_in_1_1;
      end else if (10'h118 == _T_15[9:0]) begin
        image_1_280 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_281 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h119 == _T_37[9:0]) begin
        image_1_281 <= io_pixelVal_in_1_7;
      end else if (10'h119 == _T_34[9:0]) begin
        image_1_281 <= io_pixelVal_in_1_6;
      end else if (10'h119 == _T_31[9:0]) begin
        image_1_281 <= io_pixelVal_in_1_5;
      end else if (10'h119 == _T_28[9:0]) begin
        image_1_281 <= io_pixelVal_in_1_4;
      end else if (10'h119 == _T_25[9:0]) begin
        image_1_281 <= io_pixelVal_in_1_3;
      end else if (10'h119 == _T_22[9:0]) begin
        image_1_281 <= io_pixelVal_in_1_2;
      end else if (10'h119 == _T_19[9:0]) begin
        image_1_281 <= io_pixelVal_in_1_1;
      end else if (10'h119 == _T_15[9:0]) begin
        image_1_281 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_282 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11a == _T_37[9:0]) begin
        image_1_282 <= io_pixelVal_in_1_7;
      end else if (10'h11a == _T_34[9:0]) begin
        image_1_282 <= io_pixelVal_in_1_6;
      end else if (10'h11a == _T_31[9:0]) begin
        image_1_282 <= io_pixelVal_in_1_5;
      end else if (10'h11a == _T_28[9:0]) begin
        image_1_282 <= io_pixelVal_in_1_4;
      end else if (10'h11a == _T_25[9:0]) begin
        image_1_282 <= io_pixelVal_in_1_3;
      end else if (10'h11a == _T_22[9:0]) begin
        image_1_282 <= io_pixelVal_in_1_2;
      end else if (10'h11a == _T_19[9:0]) begin
        image_1_282 <= io_pixelVal_in_1_1;
      end else if (10'h11a == _T_15[9:0]) begin
        image_1_282 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_283 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11b == _T_37[9:0]) begin
        image_1_283 <= io_pixelVal_in_1_7;
      end else if (10'h11b == _T_34[9:0]) begin
        image_1_283 <= io_pixelVal_in_1_6;
      end else if (10'h11b == _T_31[9:0]) begin
        image_1_283 <= io_pixelVal_in_1_5;
      end else if (10'h11b == _T_28[9:0]) begin
        image_1_283 <= io_pixelVal_in_1_4;
      end else if (10'h11b == _T_25[9:0]) begin
        image_1_283 <= io_pixelVal_in_1_3;
      end else if (10'h11b == _T_22[9:0]) begin
        image_1_283 <= io_pixelVal_in_1_2;
      end else if (10'h11b == _T_19[9:0]) begin
        image_1_283 <= io_pixelVal_in_1_1;
      end else if (10'h11b == _T_15[9:0]) begin
        image_1_283 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_284 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11c == _T_37[9:0]) begin
        image_1_284 <= io_pixelVal_in_1_7;
      end else if (10'h11c == _T_34[9:0]) begin
        image_1_284 <= io_pixelVal_in_1_6;
      end else if (10'h11c == _T_31[9:0]) begin
        image_1_284 <= io_pixelVal_in_1_5;
      end else if (10'h11c == _T_28[9:0]) begin
        image_1_284 <= io_pixelVal_in_1_4;
      end else if (10'h11c == _T_25[9:0]) begin
        image_1_284 <= io_pixelVal_in_1_3;
      end else if (10'h11c == _T_22[9:0]) begin
        image_1_284 <= io_pixelVal_in_1_2;
      end else if (10'h11c == _T_19[9:0]) begin
        image_1_284 <= io_pixelVal_in_1_1;
      end else if (10'h11c == _T_15[9:0]) begin
        image_1_284 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_285 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11d == _T_37[9:0]) begin
        image_1_285 <= io_pixelVal_in_1_7;
      end else if (10'h11d == _T_34[9:0]) begin
        image_1_285 <= io_pixelVal_in_1_6;
      end else if (10'h11d == _T_31[9:0]) begin
        image_1_285 <= io_pixelVal_in_1_5;
      end else if (10'h11d == _T_28[9:0]) begin
        image_1_285 <= io_pixelVal_in_1_4;
      end else if (10'h11d == _T_25[9:0]) begin
        image_1_285 <= io_pixelVal_in_1_3;
      end else if (10'h11d == _T_22[9:0]) begin
        image_1_285 <= io_pixelVal_in_1_2;
      end else if (10'h11d == _T_19[9:0]) begin
        image_1_285 <= io_pixelVal_in_1_1;
      end else if (10'h11d == _T_15[9:0]) begin
        image_1_285 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_286 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11e == _T_37[9:0]) begin
        image_1_286 <= io_pixelVal_in_1_7;
      end else if (10'h11e == _T_34[9:0]) begin
        image_1_286 <= io_pixelVal_in_1_6;
      end else if (10'h11e == _T_31[9:0]) begin
        image_1_286 <= io_pixelVal_in_1_5;
      end else if (10'h11e == _T_28[9:0]) begin
        image_1_286 <= io_pixelVal_in_1_4;
      end else if (10'h11e == _T_25[9:0]) begin
        image_1_286 <= io_pixelVal_in_1_3;
      end else if (10'h11e == _T_22[9:0]) begin
        image_1_286 <= io_pixelVal_in_1_2;
      end else if (10'h11e == _T_19[9:0]) begin
        image_1_286 <= io_pixelVal_in_1_1;
      end else if (10'h11e == _T_15[9:0]) begin
        image_1_286 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_287 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11f == _T_37[9:0]) begin
        image_1_287 <= io_pixelVal_in_1_7;
      end else if (10'h11f == _T_34[9:0]) begin
        image_1_287 <= io_pixelVal_in_1_6;
      end else if (10'h11f == _T_31[9:0]) begin
        image_1_287 <= io_pixelVal_in_1_5;
      end else if (10'h11f == _T_28[9:0]) begin
        image_1_287 <= io_pixelVal_in_1_4;
      end else if (10'h11f == _T_25[9:0]) begin
        image_1_287 <= io_pixelVal_in_1_3;
      end else if (10'h11f == _T_22[9:0]) begin
        image_1_287 <= io_pixelVal_in_1_2;
      end else if (10'h11f == _T_19[9:0]) begin
        image_1_287 <= io_pixelVal_in_1_1;
      end else if (10'h11f == _T_15[9:0]) begin
        image_1_287 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_288 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h120 == _T_37[9:0]) begin
        image_1_288 <= io_pixelVal_in_1_7;
      end else if (10'h120 == _T_34[9:0]) begin
        image_1_288 <= io_pixelVal_in_1_6;
      end else if (10'h120 == _T_31[9:0]) begin
        image_1_288 <= io_pixelVal_in_1_5;
      end else if (10'h120 == _T_28[9:0]) begin
        image_1_288 <= io_pixelVal_in_1_4;
      end else if (10'h120 == _T_25[9:0]) begin
        image_1_288 <= io_pixelVal_in_1_3;
      end else if (10'h120 == _T_22[9:0]) begin
        image_1_288 <= io_pixelVal_in_1_2;
      end else if (10'h120 == _T_19[9:0]) begin
        image_1_288 <= io_pixelVal_in_1_1;
      end else if (10'h120 == _T_15[9:0]) begin
        image_1_288 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_289 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h121 == _T_37[9:0]) begin
        image_1_289 <= io_pixelVal_in_1_7;
      end else if (10'h121 == _T_34[9:0]) begin
        image_1_289 <= io_pixelVal_in_1_6;
      end else if (10'h121 == _T_31[9:0]) begin
        image_1_289 <= io_pixelVal_in_1_5;
      end else if (10'h121 == _T_28[9:0]) begin
        image_1_289 <= io_pixelVal_in_1_4;
      end else if (10'h121 == _T_25[9:0]) begin
        image_1_289 <= io_pixelVal_in_1_3;
      end else if (10'h121 == _T_22[9:0]) begin
        image_1_289 <= io_pixelVal_in_1_2;
      end else if (10'h121 == _T_19[9:0]) begin
        image_1_289 <= io_pixelVal_in_1_1;
      end else if (10'h121 == _T_15[9:0]) begin
        image_1_289 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_290 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h122 == _T_37[9:0]) begin
        image_1_290 <= io_pixelVal_in_1_7;
      end else if (10'h122 == _T_34[9:0]) begin
        image_1_290 <= io_pixelVal_in_1_6;
      end else if (10'h122 == _T_31[9:0]) begin
        image_1_290 <= io_pixelVal_in_1_5;
      end else if (10'h122 == _T_28[9:0]) begin
        image_1_290 <= io_pixelVal_in_1_4;
      end else if (10'h122 == _T_25[9:0]) begin
        image_1_290 <= io_pixelVal_in_1_3;
      end else if (10'h122 == _T_22[9:0]) begin
        image_1_290 <= io_pixelVal_in_1_2;
      end else if (10'h122 == _T_19[9:0]) begin
        image_1_290 <= io_pixelVal_in_1_1;
      end else if (10'h122 == _T_15[9:0]) begin
        image_1_290 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_291 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h123 == _T_37[9:0]) begin
        image_1_291 <= io_pixelVal_in_1_7;
      end else if (10'h123 == _T_34[9:0]) begin
        image_1_291 <= io_pixelVal_in_1_6;
      end else if (10'h123 == _T_31[9:0]) begin
        image_1_291 <= io_pixelVal_in_1_5;
      end else if (10'h123 == _T_28[9:0]) begin
        image_1_291 <= io_pixelVal_in_1_4;
      end else if (10'h123 == _T_25[9:0]) begin
        image_1_291 <= io_pixelVal_in_1_3;
      end else if (10'h123 == _T_22[9:0]) begin
        image_1_291 <= io_pixelVal_in_1_2;
      end else if (10'h123 == _T_19[9:0]) begin
        image_1_291 <= io_pixelVal_in_1_1;
      end else if (10'h123 == _T_15[9:0]) begin
        image_1_291 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_292 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h124 == _T_37[9:0]) begin
        image_1_292 <= io_pixelVal_in_1_7;
      end else if (10'h124 == _T_34[9:0]) begin
        image_1_292 <= io_pixelVal_in_1_6;
      end else if (10'h124 == _T_31[9:0]) begin
        image_1_292 <= io_pixelVal_in_1_5;
      end else if (10'h124 == _T_28[9:0]) begin
        image_1_292 <= io_pixelVal_in_1_4;
      end else if (10'h124 == _T_25[9:0]) begin
        image_1_292 <= io_pixelVal_in_1_3;
      end else if (10'h124 == _T_22[9:0]) begin
        image_1_292 <= io_pixelVal_in_1_2;
      end else if (10'h124 == _T_19[9:0]) begin
        image_1_292 <= io_pixelVal_in_1_1;
      end else if (10'h124 == _T_15[9:0]) begin
        image_1_292 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_293 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h125 == _T_37[9:0]) begin
        image_1_293 <= io_pixelVal_in_1_7;
      end else if (10'h125 == _T_34[9:0]) begin
        image_1_293 <= io_pixelVal_in_1_6;
      end else if (10'h125 == _T_31[9:0]) begin
        image_1_293 <= io_pixelVal_in_1_5;
      end else if (10'h125 == _T_28[9:0]) begin
        image_1_293 <= io_pixelVal_in_1_4;
      end else if (10'h125 == _T_25[9:0]) begin
        image_1_293 <= io_pixelVal_in_1_3;
      end else if (10'h125 == _T_22[9:0]) begin
        image_1_293 <= io_pixelVal_in_1_2;
      end else if (10'h125 == _T_19[9:0]) begin
        image_1_293 <= io_pixelVal_in_1_1;
      end else if (10'h125 == _T_15[9:0]) begin
        image_1_293 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_294 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h126 == _T_37[9:0]) begin
        image_1_294 <= io_pixelVal_in_1_7;
      end else if (10'h126 == _T_34[9:0]) begin
        image_1_294 <= io_pixelVal_in_1_6;
      end else if (10'h126 == _T_31[9:0]) begin
        image_1_294 <= io_pixelVal_in_1_5;
      end else if (10'h126 == _T_28[9:0]) begin
        image_1_294 <= io_pixelVal_in_1_4;
      end else if (10'h126 == _T_25[9:0]) begin
        image_1_294 <= io_pixelVal_in_1_3;
      end else if (10'h126 == _T_22[9:0]) begin
        image_1_294 <= io_pixelVal_in_1_2;
      end else if (10'h126 == _T_19[9:0]) begin
        image_1_294 <= io_pixelVal_in_1_1;
      end else if (10'h126 == _T_15[9:0]) begin
        image_1_294 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_295 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h127 == _T_37[9:0]) begin
        image_1_295 <= io_pixelVal_in_1_7;
      end else if (10'h127 == _T_34[9:0]) begin
        image_1_295 <= io_pixelVal_in_1_6;
      end else if (10'h127 == _T_31[9:0]) begin
        image_1_295 <= io_pixelVal_in_1_5;
      end else if (10'h127 == _T_28[9:0]) begin
        image_1_295 <= io_pixelVal_in_1_4;
      end else if (10'h127 == _T_25[9:0]) begin
        image_1_295 <= io_pixelVal_in_1_3;
      end else if (10'h127 == _T_22[9:0]) begin
        image_1_295 <= io_pixelVal_in_1_2;
      end else if (10'h127 == _T_19[9:0]) begin
        image_1_295 <= io_pixelVal_in_1_1;
      end else if (10'h127 == _T_15[9:0]) begin
        image_1_295 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_296 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h128 == _T_37[9:0]) begin
        image_1_296 <= io_pixelVal_in_1_7;
      end else if (10'h128 == _T_34[9:0]) begin
        image_1_296 <= io_pixelVal_in_1_6;
      end else if (10'h128 == _T_31[9:0]) begin
        image_1_296 <= io_pixelVal_in_1_5;
      end else if (10'h128 == _T_28[9:0]) begin
        image_1_296 <= io_pixelVal_in_1_4;
      end else if (10'h128 == _T_25[9:0]) begin
        image_1_296 <= io_pixelVal_in_1_3;
      end else if (10'h128 == _T_22[9:0]) begin
        image_1_296 <= io_pixelVal_in_1_2;
      end else if (10'h128 == _T_19[9:0]) begin
        image_1_296 <= io_pixelVal_in_1_1;
      end else if (10'h128 == _T_15[9:0]) begin
        image_1_296 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_297 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h129 == _T_37[9:0]) begin
        image_1_297 <= io_pixelVal_in_1_7;
      end else if (10'h129 == _T_34[9:0]) begin
        image_1_297 <= io_pixelVal_in_1_6;
      end else if (10'h129 == _T_31[9:0]) begin
        image_1_297 <= io_pixelVal_in_1_5;
      end else if (10'h129 == _T_28[9:0]) begin
        image_1_297 <= io_pixelVal_in_1_4;
      end else if (10'h129 == _T_25[9:0]) begin
        image_1_297 <= io_pixelVal_in_1_3;
      end else if (10'h129 == _T_22[9:0]) begin
        image_1_297 <= io_pixelVal_in_1_2;
      end else if (10'h129 == _T_19[9:0]) begin
        image_1_297 <= io_pixelVal_in_1_1;
      end else if (10'h129 == _T_15[9:0]) begin
        image_1_297 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_298 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12a == _T_37[9:0]) begin
        image_1_298 <= io_pixelVal_in_1_7;
      end else if (10'h12a == _T_34[9:0]) begin
        image_1_298 <= io_pixelVal_in_1_6;
      end else if (10'h12a == _T_31[9:0]) begin
        image_1_298 <= io_pixelVal_in_1_5;
      end else if (10'h12a == _T_28[9:0]) begin
        image_1_298 <= io_pixelVal_in_1_4;
      end else if (10'h12a == _T_25[9:0]) begin
        image_1_298 <= io_pixelVal_in_1_3;
      end else if (10'h12a == _T_22[9:0]) begin
        image_1_298 <= io_pixelVal_in_1_2;
      end else if (10'h12a == _T_19[9:0]) begin
        image_1_298 <= io_pixelVal_in_1_1;
      end else if (10'h12a == _T_15[9:0]) begin
        image_1_298 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_299 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12b == _T_37[9:0]) begin
        image_1_299 <= io_pixelVal_in_1_7;
      end else if (10'h12b == _T_34[9:0]) begin
        image_1_299 <= io_pixelVal_in_1_6;
      end else if (10'h12b == _T_31[9:0]) begin
        image_1_299 <= io_pixelVal_in_1_5;
      end else if (10'h12b == _T_28[9:0]) begin
        image_1_299 <= io_pixelVal_in_1_4;
      end else if (10'h12b == _T_25[9:0]) begin
        image_1_299 <= io_pixelVal_in_1_3;
      end else if (10'h12b == _T_22[9:0]) begin
        image_1_299 <= io_pixelVal_in_1_2;
      end else if (10'h12b == _T_19[9:0]) begin
        image_1_299 <= io_pixelVal_in_1_1;
      end else if (10'h12b == _T_15[9:0]) begin
        image_1_299 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_300 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12c == _T_37[9:0]) begin
        image_1_300 <= io_pixelVal_in_1_7;
      end else if (10'h12c == _T_34[9:0]) begin
        image_1_300 <= io_pixelVal_in_1_6;
      end else if (10'h12c == _T_31[9:0]) begin
        image_1_300 <= io_pixelVal_in_1_5;
      end else if (10'h12c == _T_28[9:0]) begin
        image_1_300 <= io_pixelVal_in_1_4;
      end else if (10'h12c == _T_25[9:0]) begin
        image_1_300 <= io_pixelVal_in_1_3;
      end else if (10'h12c == _T_22[9:0]) begin
        image_1_300 <= io_pixelVal_in_1_2;
      end else if (10'h12c == _T_19[9:0]) begin
        image_1_300 <= io_pixelVal_in_1_1;
      end else if (10'h12c == _T_15[9:0]) begin
        image_1_300 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_301 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12d == _T_37[9:0]) begin
        image_1_301 <= io_pixelVal_in_1_7;
      end else if (10'h12d == _T_34[9:0]) begin
        image_1_301 <= io_pixelVal_in_1_6;
      end else if (10'h12d == _T_31[9:0]) begin
        image_1_301 <= io_pixelVal_in_1_5;
      end else if (10'h12d == _T_28[9:0]) begin
        image_1_301 <= io_pixelVal_in_1_4;
      end else if (10'h12d == _T_25[9:0]) begin
        image_1_301 <= io_pixelVal_in_1_3;
      end else if (10'h12d == _T_22[9:0]) begin
        image_1_301 <= io_pixelVal_in_1_2;
      end else if (10'h12d == _T_19[9:0]) begin
        image_1_301 <= io_pixelVal_in_1_1;
      end else if (10'h12d == _T_15[9:0]) begin
        image_1_301 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_302 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12e == _T_37[9:0]) begin
        image_1_302 <= io_pixelVal_in_1_7;
      end else if (10'h12e == _T_34[9:0]) begin
        image_1_302 <= io_pixelVal_in_1_6;
      end else if (10'h12e == _T_31[9:0]) begin
        image_1_302 <= io_pixelVal_in_1_5;
      end else if (10'h12e == _T_28[9:0]) begin
        image_1_302 <= io_pixelVal_in_1_4;
      end else if (10'h12e == _T_25[9:0]) begin
        image_1_302 <= io_pixelVal_in_1_3;
      end else if (10'h12e == _T_22[9:0]) begin
        image_1_302 <= io_pixelVal_in_1_2;
      end else if (10'h12e == _T_19[9:0]) begin
        image_1_302 <= io_pixelVal_in_1_1;
      end else if (10'h12e == _T_15[9:0]) begin
        image_1_302 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_303 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12f == _T_37[9:0]) begin
        image_1_303 <= io_pixelVal_in_1_7;
      end else if (10'h12f == _T_34[9:0]) begin
        image_1_303 <= io_pixelVal_in_1_6;
      end else if (10'h12f == _T_31[9:0]) begin
        image_1_303 <= io_pixelVal_in_1_5;
      end else if (10'h12f == _T_28[9:0]) begin
        image_1_303 <= io_pixelVal_in_1_4;
      end else if (10'h12f == _T_25[9:0]) begin
        image_1_303 <= io_pixelVal_in_1_3;
      end else if (10'h12f == _T_22[9:0]) begin
        image_1_303 <= io_pixelVal_in_1_2;
      end else if (10'h12f == _T_19[9:0]) begin
        image_1_303 <= io_pixelVal_in_1_1;
      end else if (10'h12f == _T_15[9:0]) begin
        image_1_303 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_304 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h130 == _T_37[9:0]) begin
        image_1_304 <= io_pixelVal_in_1_7;
      end else if (10'h130 == _T_34[9:0]) begin
        image_1_304 <= io_pixelVal_in_1_6;
      end else if (10'h130 == _T_31[9:0]) begin
        image_1_304 <= io_pixelVal_in_1_5;
      end else if (10'h130 == _T_28[9:0]) begin
        image_1_304 <= io_pixelVal_in_1_4;
      end else if (10'h130 == _T_25[9:0]) begin
        image_1_304 <= io_pixelVal_in_1_3;
      end else if (10'h130 == _T_22[9:0]) begin
        image_1_304 <= io_pixelVal_in_1_2;
      end else if (10'h130 == _T_19[9:0]) begin
        image_1_304 <= io_pixelVal_in_1_1;
      end else if (10'h130 == _T_15[9:0]) begin
        image_1_304 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_305 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h131 == _T_37[9:0]) begin
        image_1_305 <= io_pixelVal_in_1_7;
      end else if (10'h131 == _T_34[9:0]) begin
        image_1_305 <= io_pixelVal_in_1_6;
      end else if (10'h131 == _T_31[9:0]) begin
        image_1_305 <= io_pixelVal_in_1_5;
      end else if (10'h131 == _T_28[9:0]) begin
        image_1_305 <= io_pixelVal_in_1_4;
      end else if (10'h131 == _T_25[9:0]) begin
        image_1_305 <= io_pixelVal_in_1_3;
      end else if (10'h131 == _T_22[9:0]) begin
        image_1_305 <= io_pixelVal_in_1_2;
      end else if (10'h131 == _T_19[9:0]) begin
        image_1_305 <= io_pixelVal_in_1_1;
      end else if (10'h131 == _T_15[9:0]) begin
        image_1_305 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_306 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h132 == _T_37[9:0]) begin
        image_1_306 <= io_pixelVal_in_1_7;
      end else if (10'h132 == _T_34[9:0]) begin
        image_1_306 <= io_pixelVal_in_1_6;
      end else if (10'h132 == _T_31[9:0]) begin
        image_1_306 <= io_pixelVal_in_1_5;
      end else if (10'h132 == _T_28[9:0]) begin
        image_1_306 <= io_pixelVal_in_1_4;
      end else if (10'h132 == _T_25[9:0]) begin
        image_1_306 <= io_pixelVal_in_1_3;
      end else if (10'h132 == _T_22[9:0]) begin
        image_1_306 <= io_pixelVal_in_1_2;
      end else if (10'h132 == _T_19[9:0]) begin
        image_1_306 <= io_pixelVal_in_1_1;
      end else if (10'h132 == _T_15[9:0]) begin
        image_1_306 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_307 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h133 == _T_37[9:0]) begin
        image_1_307 <= io_pixelVal_in_1_7;
      end else if (10'h133 == _T_34[9:0]) begin
        image_1_307 <= io_pixelVal_in_1_6;
      end else if (10'h133 == _T_31[9:0]) begin
        image_1_307 <= io_pixelVal_in_1_5;
      end else if (10'h133 == _T_28[9:0]) begin
        image_1_307 <= io_pixelVal_in_1_4;
      end else if (10'h133 == _T_25[9:0]) begin
        image_1_307 <= io_pixelVal_in_1_3;
      end else if (10'h133 == _T_22[9:0]) begin
        image_1_307 <= io_pixelVal_in_1_2;
      end else if (10'h133 == _T_19[9:0]) begin
        image_1_307 <= io_pixelVal_in_1_1;
      end else if (10'h133 == _T_15[9:0]) begin
        image_1_307 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_308 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h134 == _T_37[9:0]) begin
        image_1_308 <= io_pixelVal_in_1_7;
      end else if (10'h134 == _T_34[9:0]) begin
        image_1_308 <= io_pixelVal_in_1_6;
      end else if (10'h134 == _T_31[9:0]) begin
        image_1_308 <= io_pixelVal_in_1_5;
      end else if (10'h134 == _T_28[9:0]) begin
        image_1_308 <= io_pixelVal_in_1_4;
      end else if (10'h134 == _T_25[9:0]) begin
        image_1_308 <= io_pixelVal_in_1_3;
      end else if (10'h134 == _T_22[9:0]) begin
        image_1_308 <= io_pixelVal_in_1_2;
      end else if (10'h134 == _T_19[9:0]) begin
        image_1_308 <= io_pixelVal_in_1_1;
      end else if (10'h134 == _T_15[9:0]) begin
        image_1_308 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_309 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h135 == _T_37[9:0]) begin
        image_1_309 <= io_pixelVal_in_1_7;
      end else if (10'h135 == _T_34[9:0]) begin
        image_1_309 <= io_pixelVal_in_1_6;
      end else if (10'h135 == _T_31[9:0]) begin
        image_1_309 <= io_pixelVal_in_1_5;
      end else if (10'h135 == _T_28[9:0]) begin
        image_1_309 <= io_pixelVal_in_1_4;
      end else if (10'h135 == _T_25[9:0]) begin
        image_1_309 <= io_pixelVal_in_1_3;
      end else if (10'h135 == _T_22[9:0]) begin
        image_1_309 <= io_pixelVal_in_1_2;
      end else if (10'h135 == _T_19[9:0]) begin
        image_1_309 <= io_pixelVal_in_1_1;
      end else if (10'h135 == _T_15[9:0]) begin
        image_1_309 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_310 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h136 == _T_37[9:0]) begin
        image_1_310 <= io_pixelVal_in_1_7;
      end else if (10'h136 == _T_34[9:0]) begin
        image_1_310 <= io_pixelVal_in_1_6;
      end else if (10'h136 == _T_31[9:0]) begin
        image_1_310 <= io_pixelVal_in_1_5;
      end else if (10'h136 == _T_28[9:0]) begin
        image_1_310 <= io_pixelVal_in_1_4;
      end else if (10'h136 == _T_25[9:0]) begin
        image_1_310 <= io_pixelVal_in_1_3;
      end else if (10'h136 == _T_22[9:0]) begin
        image_1_310 <= io_pixelVal_in_1_2;
      end else if (10'h136 == _T_19[9:0]) begin
        image_1_310 <= io_pixelVal_in_1_1;
      end else if (10'h136 == _T_15[9:0]) begin
        image_1_310 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_311 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h137 == _T_37[9:0]) begin
        image_1_311 <= io_pixelVal_in_1_7;
      end else if (10'h137 == _T_34[9:0]) begin
        image_1_311 <= io_pixelVal_in_1_6;
      end else if (10'h137 == _T_31[9:0]) begin
        image_1_311 <= io_pixelVal_in_1_5;
      end else if (10'h137 == _T_28[9:0]) begin
        image_1_311 <= io_pixelVal_in_1_4;
      end else if (10'h137 == _T_25[9:0]) begin
        image_1_311 <= io_pixelVal_in_1_3;
      end else if (10'h137 == _T_22[9:0]) begin
        image_1_311 <= io_pixelVal_in_1_2;
      end else if (10'h137 == _T_19[9:0]) begin
        image_1_311 <= io_pixelVal_in_1_1;
      end else if (10'h137 == _T_15[9:0]) begin
        image_1_311 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_312 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h138 == _T_37[9:0]) begin
        image_1_312 <= io_pixelVal_in_1_7;
      end else if (10'h138 == _T_34[9:0]) begin
        image_1_312 <= io_pixelVal_in_1_6;
      end else if (10'h138 == _T_31[9:0]) begin
        image_1_312 <= io_pixelVal_in_1_5;
      end else if (10'h138 == _T_28[9:0]) begin
        image_1_312 <= io_pixelVal_in_1_4;
      end else if (10'h138 == _T_25[9:0]) begin
        image_1_312 <= io_pixelVal_in_1_3;
      end else if (10'h138 == _T_22[9:0]) begin
        image_1_312 <= io_pixelVal_in_1_2;
      end else if (10'h138 == _T_19[9:0]) begin
        image_1_312 <= io_pixelVal_in_1_1;
      end else if (10'h138 == _T_15[9:0]) begin
        image_1_312 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_313 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h139 == _T_37[9:0]) begin
        image_1_313 <= io_pixelVal_in_1_7;
      end else if (10'h139 == _T_34[9:0]) begin
        image_1_313 <= io_pixelVal_in_1_6;
      end else if (10'h139 == _T_31[9:0]) begin
        image_1_313 <= io_pixelVal_in_1_5;
      end else if (10'h139 == _T_28[9:0]) begin
        image_1_313 <= io_pixelVal_in_1_4;
      end else if (10'h139 == _T_25[9:0]) begin
        image_1_313 <= io_pixelVal_in_1_3;
      end else if (10'h139 == _T_22[9:0]) begin
        image_1_313 <= io_pixelVal_in_1_2;
      end else if (10'h139 == _T_19[9:0]) begin
        image_1_313 <= io_pixelVal_in_1_1;
      end else if (10'h139 == _T_15[9:0]) begin
        image_1_313 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_314 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13a == _T_37[9:0]) begin
        image_1_314 <= io_pixelVal_in_1_7;
      end else if (10'h13a == _T_34[9:0]) begin
        image_1_314 <= io_pixelVal_in_1_6;
      end else if (10'h13a == _T_31[9:0]) begin
        image_1_314 <= io_pixelVal_in_1_5;
      end else if (10'h13a == _T_28[9:0]) begin
        image_1_314 <= io_pixelVal_in_1_4;
      end else if (10'h13a == _T_25[9:0]) begin
        image_1_314 <= io_pixelVal_in_1_3;
      end else if (10'h13a == _T_22[9:0]) begin
        image_1_314 <= io_pixelVal_in_1_2;
      end else if (10'h13a == _T_19[9:0]) begin
        image_1_314 <= io_pixelVal_in_1_1;
      end else if (10'h13a == _T_15[9:0]) begin
        image_1_314 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_315 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13b == _T_37[9:0]) begin
        image_1_315 <= io_pixelVal_in_1_7;
      end else if (10'h13b == _T_34[9:0]) begin
        image_1_315 <= io_pixelVal_in_1_6;
      end else if (10'h13b == _T_31[9:0]) begin
        image_1_315 <= io_pixelVal_in_1_5;
      end else if (10'h13b == _T_28[9:0]) begin
        image_1_315 <= io_pixelVal_in_1_4;
      end else if (10'h13b == _T_25[9:0]) begin
        image_1_315 <= io_pixelVal_in_1_3;
      end else if (10'h13b == _T_22[9:0]) begin
        image_1_315 <= io_pixelVal_in_1_2;
      end else if (10'h13b == _T_19[9:0]) begin
        image_1_315 <= io_pixelVal_in_1_1;
      end else if (10'h13b == _T_15[9:0]) begin
        image_1_315 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_316 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13c == _T_37[9:0]) begin
        image_1_316 <= io_pixelVal_in_1_7;
      end else if (10'h13c == _T_34[9:0]) begin
        image_1_316 <= io_pixelVal_in_1_6;
      end else if (10'h13c == _T_31[9:0]) begin
        image_1_316 <= io_pixelVal_in_1_5;
      end else if (10'h13c == _T_28[9:0]) begin
        image_1_316 <= io_pixelVal_in_1_4;
      end else if (10'h13c == _T_25[9:0]) begin
        image_1_316 <= io_pixelVal_in_1_3;
      end else if (10'h13c == _T_22[9:0]) begin
        image_1_316 <= io_pixelVal_in_1_2;
      end else if (10'h13c == _T_19[9:0]) begin
        image_1_316 <= io_pixelVal_in_1_1;
      end else if (10'h13c == _T_15[9:0]) begin
        image_1_316 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_317 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13d == _T_37[9:0]) begin
        image_1_317 <= io_pixelVal_in_1_7;
      end else if (10'h13d == _T_34[9:0]) begin
        image_1_317 <= io_pixelVal_in_1_6;
      end else if (10'h13d == _T_31[9:0]) begin
        image_1_317 <= io_pixelVal_in_1_5;
      end else if (10'h13d == _T_28[9:0]) begin
        image_1_317 <= io_pixelVal_in_1_4;
      end else if (10'h13d == _T_25[9:0]) begin
        image_1_317 <= io_pixelVal_in_1_3;
      end else if (10'h13d == _T_22[9:0]) begin
        image_1_317 <= io_pixelVal_in_1_2;
      end else if (10'h13d == _T_19[9:0]) begin
        image_1_317 <= io_pixelVal_in_1_1;
      end else if (10'h13d == _T_15[9:0]) begin
        image_1_317 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_318 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13e == _T_37[9:0]) begin
        image_1_318 <= io_pixelVal_in_1_7;
      end else if (10'h13e == _T_34[9:0]) begin
        image_1_318 <= io_pixelVal_in_1_6;
      end else if (10'h13e == _T_31[9:0]) begin
        image_1_318 <= io_pixelVal_in_1_5;
      end else if (10'h13e == _T_28[9:0]) begin
        image_1_318 <= io_pixelVal_in_1_4;
      end else if (10'h13e == _T_25[9:0]) begin
        image_1_318 <= io_pixelVal_in_1_3;
      end else if (10'h13e == _T_22[9:0]) begin
        image_1_318 <= io_pixelVal_in_1_2;
      end else if (10'h13e == _T_19[9:0]) begin
        image_1_318 <= io_pixelVal_in_1_1;
      end else if (10'h13e == _T_15[9:0]) begin
        image_1_318 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_319 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13f == _T_37[9:0]) begin
        image_1_319 <= io_pixelVal_in_1_7;
      end else if (10'h13f == _T_34[9:0]) begin
        image_1_319 <= io_pixelVal_in_1_6;
      end else if (10'h13f == _T_31[9:0]) begin
        image_1_319 <= io_pixelVal_in_1_5;
      end else if (10'h13f == _T_28[9:0]) begin
        image_1_319 <= io_pixelVal_in_1_4;
      end else if (10'h13f == _T_25[9:0]) begin
        image_1_319 <= io_pixelVal_in_1_3;
      end else if (10'h13f == _T_22[9:0]) begin
        image_1_319 <= io_pixelVal_in_1_2;
      end else if (10'h13f == _T_19[9:0]) begin
        image_1_319 <= io_pixelVal_in_1_1;
      end else if (10'h13f == _T_15[9:0]) begin
        image_1_319 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_320 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h140 == _T_37[9:0]) begin
        image_1_320 <= io_pixelVal_in_1_7;
      end else if (10'h140 == _T_34[9:0]) begin
        image_1_320 <= io_pixelVal_in_1_6;
      end else if (10'h140 == _T_31[9:0]) begin
        image_1_320 <= io_pixelVal_in_1_5;
      end else if (10'h140 == _T_28[9:0]) begin
        image_1_320 <= io_pixelVal_in_1_4;
      end else if (10'h140 == _T_25[9:0]) begin
        image_1_320 <= io_pixelVal_in_1_3;
      end else if (10'h140 == _T_22[9:0]) begin
        image_1_320 <= io_pixelVal_in_1_2;
      end else if (10'h140 == _T_19[9:0]) begin
        image_1_320 <= io_pixelVal_in_1_1;
      end else if (10'h140 == _T_15[9:0]) begin
        image_1_320 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_321 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h141 == _T_37[9:0]) begin
        image_1_321 <= io_pixelVal_in_1_7;
      end else if (10'h141 == _T_34[9:0]) begin
        image_1_321 <= io_pixelVal_in_1_6;
      end else if (10'h141 == _T_31[9:0]) begin
        image_1_321 <= io_pixelVal_in_1_5;
      end else if (10'h141 == _T_28[9:0]) begin
        image_1_321 <= io_pixelVal_in_1_4;
      end else if (10'h141 == _T_25[9:0]) begin
        image_1_321 <= io_pixelVal_in_1_3;
      end else if (10'h141 == _T_22[9:0]) begin
        image_1_321 <= io_pixelVal_in_1_2;
      end else if (10'h141 == _T_19[9:0]) begin
        image_1_321 <= io_pixelVal_in_1_1;
      end else if (10'h141 == _T_15[9:0]) begin
        image_1_321 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_322 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h142 == _T_37[9:0]) begin
        image_1_322 <= io_pixelVal_in_1_7;
      end else if (10'h142 == _T_34[9:0]) begin
        image_1_322 <= io_pixelVal_in_1_6;
      end else if (10'h142 == _T_31[9:0]) begin
        image_1_322 <= io_pixelVal_in_1_5;
      end else if (10'h142 == _T_28[9:0]) begin
        image_1_322 <= io_pixelVal_in_1_4;
      end else if (10'h142 == _T_25[9:0]) begin
        image_1_322 <= io_pixelVal_in_1_3;
      end else if (10'h142 == _T_22[9:0]) begin
        image_1_322 <= io_pixelVal_in_1_2;
      end else if (10'h142 == _T_19[9:0]) begin
        image_1_322 <= io_pixelVal_in_1_1;
      end else if (10'h142 == _T_15[9:0]) begin
        image_1_322 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_323 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h143 == _T_37[9:0]) begin
        image_1_323 <= io_pixelVal_in_1_7;
      end else if (10'h143 == _T_34[9:0]) begin
        image_1_323 <= io_pixelVal_in_1_6;
      end else if (10'h143 == _T_31[9:0]) begin
        image_1_323 <= io_pixelVal_in_1_5;
      end else if (10'h143 == _T_28[9:0]) begin
        image_1_323 <= io_pixelVal_in_1_4;
      end else if (10'h143 == _T_25[9:0]) begin
        image_1_323 <= io_pixelVal_in_1_3;
      end else if (10'h143 == _T_22[9:0]) begin
        image_1_323 <= io_pixelVal_in_1_2;
      end else if (10'h143 == _T_19[9:0]) begin
        image_1_323 <= io_pixelVal_in_1_1;
      end else if (10'h143 == _T_15[9:0]) begin
        image_1_323 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_324 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h144 == _T_37[9:0]) begin
        image_1_324 <= io_pixelVal_in_1_7;
      end else if (10'h144 == _T_34[9:0]) begin
        image_1_324 <= io_pixelVal_in_1_6;
      end else if (10'h144 == _T_31[9:0]) begin
        image_1_324 <= io_pixelVal_in_1_5;
      end else if (10'h144 == _T_28[9:0]) begin
        image_1_324 <= io_pixelVal_in_1_4;
      end else if (10'h144 == _T_25[9:0]) begin
        image_1_324 <= io_pixelVal_in_1_3;
      end else if (10'h144 == _T_22[9:0]) begin
        image_1_324 <= io_pixelVal_in_1_2;
      end else if (10'h144 == _T_19[9:0]) begin
        image_1_324 <= io_pixelVal_in_1_1;
      end else if (10'h144 == _T_15[9:0]) begin
        image_1_324 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_325 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h145 == _T_37[9:0]) begin
        image_1_325 <= io_pixelVal_in_1_7;
      end else if (10'h145 == _T_34[9:0]) begin
        image_1_325 <= io_pixelVal_in_1_6;
      end else if (10'h145 == _T_31[9:0]) begin
        image_1_325 <= io_pixelVal_in_1_5;
      end else if (10'h145 == _T_28[9:0]) begin
        image_1_325 <= io_pixelVal_in_1_4;
      end else if (10'h145 == _T_25[9:0]) begin
        image_1_325 <= io_pixelVal_in_1_3;
      end else if (10'h145 == _T_22[9:0]) begin
        image_1_325 <= io_pixelVal_in_1_2;
      end else if (10'h145 == _T_19[9:0]) begin
        image_1_325 <= io_pixelVal_in_1_1;
      end else if (10'h145 == _T_15[9:0]) begin
        image_1_325 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_326 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h146 == _T_37[9:0]) begin
        image_1_326 <= io_pixelVal_in_1_7;
      end else if (10'h146 == _T_34[9:0]) begin
        image_1_326 <= io_pixelVal_in_1_6;
      end else if (10'h146 == _T_31[9:0]) begin
        image_1_326 <= io_pixelVal_in_1_5;
      end else if (10'h146 == _T_28[9:0]) begin
        image_1_326 <= io_pixelVal_in_1_4;
      end else if (10'h146 == _T_25[9:0]) begin
        image_1_326 <= io_pixelVal_in_1_3;
      end else if (10'h146 == _T_22[9:0]) begin
        image_1_326 <= io_pixelVal_in_1_2;
      end else if (10'h146 == _T_19[9:0]) begin
        image_1_326 <= io_pixelVal_in_1_1;
      end else if (10'h146 == _T_15[9:0]) begin
        image_1_326 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_327 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h147 == _T_37[9:0]) begin
        image_1_327 <= io_pixelVal_in_1_7;
      end else if (10'h147 == _T_34[9:0]) begin
        image_1_327 <= io_pixelVal_in_1_6;
      end else if (10'h147 == _T_31[9:0]) begin
        image_1_327 <= io_pixelVal_in_1_5;
      end else if (10'h147 == _T_28[9:0]) begin
        image_1_327 <= io_pixelVal_in_1_4;
      end else if (10'h147 == _T_25[9:0]) begin
        image_1_327 <= io_pixelVal_in_1_3;
      end else if (10'h147 == _T_22[9:0]) begin
        image_1_327 <= io_pixelVal_in_1_2;
      end else if (10'h147 == _T_19[9:0]) begin
        image_1_327 <= io_pixelVal_in_1_1;
      end else if (10'h147 == _T_15[9:0]) begin
        image_1_327 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_328 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h148 == _T_37[9:0]) begin
        image_1_328 <= io_pixelVal_in_1_7;
      end else if (10'h148 == _T_34[9:0]) begin
        image_1_328 <= io_pixelVal_in_1_6;
      end else if (10'h148 == _T_31[9:0]) begin
        image_1_328 <= io_pixelVal_in_1_5;
      end else if (10'h148 == _T_28[9:0]) begin
        image_1_328 <= io_pixelVal_in_1_4;
      end else if (10'h148 == _T_25[9:0]) begin
        image_1_328 <= io_pixelVal_in_1_3;
      end else if (10'h148 == _T_22[9:0]) begin
        image_1_328 <= io_pixelVal_in_1_2;
      end else if (10'h148 == _T_19[9:0]) begin
        image_1_328 <= io_pixelVal_in_1_1;
      end else if (10'h148 == _T_15[9:0]) begin
        image_1_328 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_329 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h149 == _T_37[9:0]) begin
        image_1_329 <= io_pixelVal_in_1_7;
      end else if (10'h149 == _T_34[9:0]) begin
        image_1_329 <= io_pixelVal_in_1_6;
      end else if (10'h149 == _T_31[9:0]) begin
        image_1_329 <= io_pixelVal_in_1_5;
      end else if (10'h149 == _T_28[9:0]) begin
        image_1_329 <= io_pixelVal_in_1_4;
      end else if (10'h149 == _T_25[9:0]) begin
        image_1_329 <= io_pixelVal_in_1_3;
      end else if (10'h149 == _T_22[9:0]) begin
        image_1_329 <= io_pixelVal_in_1_2;
      end else if (10'h149 == _T_19[9:0]) begin
        image_1_329 <= io_pixelVal_in_1_1;
      end else if (10'h149 == _T_15[9:0]) begin
        image_1_329 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_330 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14a == _T_37[9:0]) begin
        image_1_330 <= io_pixelVal_in_1_7;
      end else if (10'h14a == _T_34[9:0]) begin
        image_1_330 <= io_pixelVal_in_1_6;
      end else if (10'h14a == _T_31[9:0]) begin
        image_1_330 <= io_pixelVal_in_1_5;
      end else if (10'h14a == _T_28[9:0]) begin
        image_1_330 <= io_pixelVal_in_1_4;
      end else if (10'h14a == _T_25[9:0]) begin
        image_1_330 <= io_pixelVal_in_1_3;
      end else if (10'h14a == _T_22[9:0]) begin
        image_1_330 <= io_pixelVal_in_1_2;
      end else if (10'h14a == _T_19[9:0]) begin
        image_1_330 <= io_pixelVal_in_1_1;
      end else if (10'h14a == _T_15[9:0]) begin
        image_1_330 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_331 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14b == _T_37[9:0]) begin
        image_1_331 <= io_pixelVal_in_1_7;
      end else if (10'h14b == _T_34[9:0]) begin
        image_1_331 <= io_pixelVal_in_1_6;
      end else if (10'h14b == _T_31[9:0]) begin
        image_1_331 <= io_pixelVal_in_1_5;
      end else if (10'h14b == _T_28[9:0]) begin
        image_1_331 <= io_pixelVal_in_1_4;
      end else if (10'h14b == _T_25[9:0]) begin
        image_1_331 <= io_pixelVal_in_1_3;
      end else if (10'h14b == _T_22[9:0]) begin
        image_1_331 <= io_pixelVal_in_1_2;
      end else if (10'h14b == _T_19[9:0]) begin
        image_1_331 <= io_pixelVal_in_1_1;
      end else if (10'h14b == _T_15[9:0]) begin
        image_1_331 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_332 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14c == _T_37[9:0]) begin
        image_1_332 <= io_pixelVal_in_1_7;
      end else if (10'h14c == _T_34[9:0]) begin
        image_1_332 <= io_pixelVal_in_1_6;
      end else if (10'h14c == _T_31[9:0]) begin
        image_1_332 <= io_pixelVal_in_1_5;
      end else if (10'h14c == _T_28[9:0]) begin
        image_1_332 <= io_pixelVal_in_1_4;
      end else if (10'h14c == _T_25[9:0]) begin
        image_1_332 <= io_pixelVal_in_1_3;
      end else if (10'h14c == _T_22[9:0]) begin
        image_1_332 <= io_pixelVal_in_1_2;
      end else if (10'h14c == _T_19[9:0]) begin
        image_1_332 <= io_pixelVal_in_1_1;
      end else if (10'h14c == _T_15[9:0]) begin
        image_1_332 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_333 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14d == _T_37[9:0]) begin
        image_1_333 <= io_pixelVal_in_1_7;
      end else if (10'h14d == _T_34[9:0]) begin
        image_1_333 <= io_pixelVal_in_1_6;
      end else if (10'h14d == _T_31[9:0]) begin
        image_1_333 <= io_pixelVal_in_1_5;
      end else if (10'h14d == _T_28[9:0]) begin
        image_1_333 <= io_pixelVal_in_1_4;
      end else if (10'h14d == _T_25[9:0]) begin
        image_1_333 <= io_pixelVal_in_1_3;
      end else if (10'h14d == _T_22[9:0]) begin
        image_1_333 <= io_pixelVal_in_1_2;
      end else if (10'h14d == _T_19[9:0]) begin
        image_1_333 <= io_pixelVal_in_1_1;
      end else if (10'h14d == _T_15[9:0]) begin
        image_1_333 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_334 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14e == _T_37[9:0]) begin
        image_1_334 <= io_pixelVal_in_1_7;
      end else if (10'h14e == _T_34[9:0]) begin
        image_1_334 <= io_pixelVal_in_1_6;
      end else if (10'h14e == _T_31[9:0]) begin
        image_1_334 <= io_pixelVal_in_1_5;
      end else if (10'h14e == _T_28[9:0]) begin
        image_1_334 <= io_pixelVal_in_1_4;
      end else if (10'h14e == _T_25[9:0]) begin
        image_1_334 <= io_pixelVal_in_1_3;
      end else if (10'h14e == _T_22[9:0]) begin
        image_1_334 <= io_pixelVal_in_1_2;
      end else if (10'h14e == _T_19[9:0]) begin
        image_1_334 <= io_pixelVal_in_1_1;
      end else if (10'h14e == _T_15[9:0]) begin
        image_1_334 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_335 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14f == _T_37[9:0]) begin
        image_1_335 <= io_pixelVal_in_1_7;
      end else if (10'h14f == _T_34[9:0]) begin
        image_1_335 <= io_pixelVal_in_1_6;
      end else if (10'h14f == _T_31[9:0]) begin
        image_1_335 <= io_pixelVal_in_1_5;
      end else if (10'h14f == _T_28[9:0]) begin
        image_1_335 <= io_pixelVal_in_1_4;
      end else if (10'h14f == _T_25[9:0]) begin
        image_1_335 <= io_pixelVal_in_1_3;
      end else if (10'h14f == _T_22[9:0]) begin
        image_1_335 <= io_pixelVal_in_1_2;
      end else if (10'h14f == _T_19[9:0]) begin
        image_1_335 <= io_pixelVal_in_1_1;
      end else if (10'h14f == _T_15[9:0]) begin
        image_1_335 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_336 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h150 == _T_37[9:0]) begin
        image_1_336 <= io_pixelVal_in_1_7;
      end else if (10'h150 == _T_34[9:0]) begin
        image_1_336 <= io_pixelVal_in_1_6;
      end else if (10'h150 == _T_31[9:0]) begin
        image_1_336 <= io_pixelVal_in_1_5;
      end else if (10'h150 == _T_28[9:0]) begin
        image_1_336 <= io_pixelVal_in_1_4;
      end else if (10'h150 == _T_25[9:0]) begin
        image_1_336 <= io_pixelVal_in_1_3;
      end else if (10'h150 == _T_22[9:0]) begin
        image_1_336 <= io_pixelVal_in_1_2;
      end else if (10'h150 == _T_19[9:0]) begin
        image_1_336 <= io_pixelVal_in_1_1;
      end else if (10'h150 == _T_15[9:0]) begin
        image_1_336 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_337 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h151 == _T_37[9:0]) begin
        image_1_337 <= io_pixelVal_in_1_7;
      end else if (10'h151 == _T_34[9:0]) begin
        image_1_337 <= io_pixelVal_in_1_6;
      end else if (10'h151 == _T_31[9:0]) begin
        image_1_337 <= io_pixelVal_in_1_5;
      end else if (10'h151 == _T_28[9:0]) begin
        image_1_337 <= io_pixelVal_in_1_4;
      end else if (10'h151 == _T_25[9:0]) begin
        image_1_337 <= io_pixelVal_in_1_3;
      end else if (10'h151 == _T_22[9:0]) begin
        image_1_337 <= io_pixelVal_in_1_2;
      end else if (10'h151 == _T_19[9:0]) begin
        image_1_337 <= io_pixelVal_in_1_1;
      end else if (10'h151 == _T_15[9:0]) begin
        image_1_337 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_338 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h152 == _T_37[9:0]) begin
        image_1_338 <= io_pixelVal_in_1_7;
      end else if (10'h152 == _T_34[9:0]) begin
        image_1_338 <= io_pixelVal_in_1_6;
      end else if (10'h152 == _T_31[9:0]) begin
        image_1_338 <= io_pixelVal_in_1_5;
      end else if (10'h152 == _T_28[9:0]) begin
        image_1_338 <= io_pixelVal_in_1_4;
      end else if (10'h152 == _T_25[9:0]) begin
        image_1_338 <= io_pixelVal_in_1_3;
      end else if (10'h152 == _T_22[9:0]) begin
        image_1_338 <= io_pixelVal_in_1_2;
      end else if (10'h152 == _T_19[9:0]) begin
        image_1_338 <= io_pixelVal_in_1_1;
      end else if (10'h152 == _T_15[9:0]) begin
        image_1_338 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_339 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h153 == _T_37[9:0]) begin
        image_1_339 <= io_pixelVal_in_1_7;
      end else if (10'h153 == _T_34[9:0]) begin
        image_1_339 <= io_pixelVal_in_1_6;
      end else if (10'h153 == _T_31[9:0]) begin
        image_1_339 <= io_pixelVal_in_1_5;
      end else if (10'h153 == _T_28[9:0]) begin
        image_1_339 <= io_pixelVal_in_1_4;
      end else if (10'h153 == _T_25[9:0]) begin
        image_1_339 <= io_pixelVal_in_1_3;
      end else if (10'h153 == _T_22[9:0]) begin
        image_1_339 <= io_pixelVal_in_1_2;
      end else if (10'h153 == _T_19[9:0]) begin
        image_1_339 <= io_pixelVal_in_1_1;
      end else if (10'h153 == _T_15[9:0]) begin
        image_1_339 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_340 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h154 == _T_37[9:0]) begin
        image_1_340 <= io_pixelVal_in_1_7;
      end else if (10'h154 == _T_34[9:0]) begin
        image_1_340 <= io_pixelVal_in_1_6;
      end else if (10'h154 == _T_31[9:0]) begin
        image_1_340 <= io_pixelVal_in_1_5;
      end else if (10'h154 == _T_28[9:0]) begin
        image_1_340 <= io_pixelVal_in_1_4;
      end else if (10'h154 == _T_25[9:0]) begin
        image_1_340 <= io_pixelVal_in_1_3;
      end else if (10'h154 == _T_22[9:0]) begin
        image_1_340 <= io_pixelVal_in_1_2;
      end else if (10'h154 == _T_19[9:0]) begin
        image_1_340 <= io_pixelVal_in_1_1;
      end else if (10'h154 == _T_15[9:0]) begin
        image_1_340 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_341 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h155 == _T_37[9:0]) begin
        image_1_341 <= io_pixelVal_in_1_7;
      end else if (10'h155 == _T_34[9:0]) begin
        image_1_341 <= io_pixelVal_in_1_6;
      end else if (10'h155 == _T_31[9:0]) begin
        image_1_341 <= io_pixelVal_in_1_5;
      end else if (10'h155 == _T_28[9:0]) begin
        image_1_341 <= io_pixelVal_in_1_4;
      end else if (10'h155 == _T_25[9:0]) begin
        image_1_341 <= io_pixelVal_in_1_3;
      end else if (10'h155 == _T_22[9:0]) begin
        image_1_341 <= io_pixelVal_in_1_2;
      end else if (10'h155 == _T_19[9:0]) begin
        image_1_341 <= io_pixelVal_in_1_1;
      end else if (10'h155 == _T_15[9:0]) begin
        image_1_341 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_342 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h156 == _T_37[9:0]) begin
        image_1_342 <= io_pixelVal_in_1_7;
      end else if (10'h156 == _T_34[9:0]) begin
        image_1_342 <= io_pixelVal_in_1_6;
      end else if (10'h156 == _T_31[9:0]) begin
        image_1_342 <= io_pixelVal_in_1_5;
      end else if (10'h156 == _T_28[9:0]) begin
        image_1_342 <= io_pixelVal_in_1_4;
      end else if (10'h156 == _T_25[9:0]) begin
        image_1_342 <= io_pixelVal_in_1_3;
      end else if (10'h156 == _T_22[9:0]) begin
        image_1_342 <= io_pixelVal_in_1_2;
      end else if (10'h156 == _T_19[9:0]) begin
        image_1_342 <= io_pixelVal_in_1_1;
      end else if (10'h156 == _T_15[9:0]) begin
        image_1_342 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_343 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h157 == _T_37[9:0]) begin
        image_1_343 <= io_pixelVal_in_1_7;
      end else if (10'h157 == _T_34[9:0]) begin
        image_1_343 <= io_pixelVal_in_1_6;
      end else if (10'h157 == _T_31[9:0]) begin
        image_1_343 <= io_pixelVal_in_1_5;
      end else if (10'h157 == _T_28[9:0]) begin
        image_1_343 <= io_pixelVal_in_1_4;
      end else if (10'h157 == _T_25[9:0]) begin
        image_1_343 <= io_pixelVal_in_1_3;
      end else if (10'h157 == _T_22[9:0]) begin
        image_1_343 <= io_pixelVal_in_1_2;
      end else if (10'h157 == _T_19[9:0]) begin
        image_1_343 <= io_pixelVal_in_1_1;
      end else if (10'h157 == _T_15[9:0]) begin
        image_1_343 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_344 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h158 == _T_37[9:0]) begin
        image_1_344 <= io_pixelVal_in_1_7;
      end else if (10'h158 == _T_34[9:0]) begin
        image_1_344 <= io_pixelVal_in_1_6;
      end else if (10'h158 == _T_31[9:0]) begin
        image_1_344 <= io_pixelVal_in_1_5;
      end else if (10'h158 == _T_28[9:0]) begin
        image_1_344 <= io_pixelVal_in_1_4;
      end else if (10'h158 == _T_25[9:0]) begin
        image_1_344 <= io_pixelVal_in_1_3;
      end else if (10'h158 == _T_22[9:0]) begin
        image_1_344 <= io_pixelVal_in_1_2;
      end else if (10'h158 == _T_19[9:0]) begin
        image_1_344 <= io_pixelVal_in_1_1;
      end else if (10'h158 == _T_15[9:0]) begin
        image_1_344 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_345 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h159 == _T_37[9:0]) begin
        image_1_345 <= io_pixelVal_in_1_7;
      end else if (10'h159 == _T_34[9:0]) begin
        image_1_345 <= io_pixelVal_in_1_6;
      end else if (10'h159 == _T_31[9:0]) begin
        image_1_345 <= io_pixelVal_in_1_5;
      end else if (10'h159 == _T_28[9:0]) begin
        image_1_345 <= io_pixelVal_in_1_4;
      end else if (10'h159 == _T_25[9:0]) begin
        image_1_345 <= io_pixelVal_in_1_3;
      end else if (10'h159 == _T_22[9:0]) begin
        image_1_345 <= io_pixelVal_in_1_2;
      end else if (10'h159 == _T_19[9:0]) begin
        image_1_345 <= io_pixelVal_in_1_1;
      end else if (10'h159 == _T_15[9:0]) begin
        image_1_345 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_346 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15a == _T_37[9:0]) begin
        image_1_346 <= io_pixelVal_in_1_7;
      end else if (10'h15a == _T_34[9:0]) begin
        image_1_346 <= io_pixelVal_in_1_6;
      end else if (10'h15a == _T_31[9:0]) begin
        image_1_346 <= io_pixelVal_in_1_5;
      end else if (10'h15a == _T_28[9:0]) begin
        image_1_346 <= io_pixelVal_in_1_4;
      end else if (10'h15a == _T_25[9:0]) begin
        image_1_346 <= io_pixelVal_in_1_3;
      end else if (10'h15a == _T_22[9:0]) begin
        image_1_346 <= io_pixelVal_in_1_2;
      end else if (10'h15a == _T_19[9:0]) begin
        image_1_346 <= io_pixelVal_in_1_1;
      end else if (10'h15a == _T_15[9:0]) begin
        image_1_346 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_347 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15b == _T_37[9:0]) begin
        image_1_347 <= io_pixelVal_in_1_7;
      end else if (10'h15b == _T_34[9:0]) begin
        image_1_347 <= io_pixelVal_in_1_6;
      end else if (10'h15b == _T_31[9:0]) begin
        image_1_347 <= io_pixelVal_in_1_5;
      end else if (10'h15b == _T_28[9:0]) begin
        image_1_347 <= io_pixelVal_in_1_4;
      end else if (10'h15b == _T_25[9:0]) begin
        image_1_347 <= io_pixelVal_in_1_3;
      end else if (10'h15b == _T_22[9:0]) begin
        image_1_347 <= io_pixelVal_in_1_2;
      end else if (10'h15b == _T_19[9:0]) begin
        image_1_347 <= io_pixelVal_in_1_1;
      end else if (10'h15b == _T_15[9:0]) begin
        image_1_347 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_348 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15c == _T_37[9:0]) begin
        image_1_348 <= io_pixelVal_in_1_7;
      end else if (10'h15c == _T_34[9:0]) begin
        image_1_348 <= io_pixelVal_in_1_6;
      end else if (10'h15c == _T_31[9:0]) begin
        image_1_348 <= io_pixelVal_in_1_5;
      end else if (10'h15c == _T_28[9:0]) begin
        image_1_348 <= io_pixelVal_in_1_4;
      end else if (10'h15c == _T_25[9:0]) begin
        image_1_348 <= io_pixelVal_in_1_3;
      end else if (10'h15c == _T_22[9:0]) begin
        image_1_348 <= io_pixelVal_in_1_2;
      end else if (10'h15c == _T_19[9:0]) begin
        image_1_348 <= io_pixelVal_in_1_1;
      end else if (10'h15c == _T_15[9:0]) begin
        image_1_348 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_349 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15d == _T_37[9:0]) begin
        image_1_349 <= io_pixelVal_in_1_7;
      end else if (10'h15d == _T_34[9:0]) begin
        image_1_349 <= io_pixelVal_in_1_6;
      end else if (10'h15d == _T_31[9:0]) begin
        image_1_349 <= io_pixelVal_in_1_5;
      end else if (10'h15d == _T_28[9:0]) begin
        image_1_349 <= io_pixelVal_in_1_4;
      end else if (10'h15d == _T_25[9:0]) begin
        image_1_349 <= io_pixelVal_in_1_3;
      end else if (10'h15d == _T_22[9:0]) begin
        image_1_349 <= io_pixelVal_in_1_2;
      end else if (10'h15d == _T_19[9:0]) begin
        image_1_349 <= io_pixelVal_in_1_1;
      end else if (10'h15d == _T_15[9:0]) begin
        image_1_349 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_350 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15e == _T_37[9:0]) begin
        image_1_350 <= io_pixelVal_in_1_7;
      end else if (10'h15e == _T_34[9:0]) begin
        image_1_350 <= io_pixelVal_in_1_6;
      end else if (10'h15e == _T_31[9:0]) begin
        image_1_350 <= io_pixelVal_in_1_5;
      end else if (10'h15e == _T_28[9:0]) begin
        image_1_350 <= io_pixelVal_in_1_4;
      end else if (10'h15e == _T_25[9:0]) begin
        image_1_350 <= io_pixelVal_in_1_3;
      end else if (10'h15e == _T_22[9:0]) begin
        image_1_350 <= io_pixelVal_in_1_2;
      end else if (10'h15e == _T_19[9:0]) begin
        image_1_350 <= io_pixelVal_in_1_1;
      end else if (10'h15e == _T_15[9:0]) begin
        image_1_350 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_351 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15f == _T_37[9:0]) begin
        image_1_351 <= io_pixelVal_in_1_7;
      end else if (10'h15f == _T_34[9:0]) begin
        image_1_351 <= io_pixelVal_in_1_6;
      end else if (10'h15f == _T_31[9:0]) begin
        image_1_351 <= io_pixelVal_in_1_5;
      end else if (10'h15f == _T_28[9:0]) begin
        image_1_351 <= io_pixelVal_in_1_4;
      end else if (10'h15f == _T_25[9:0]) begin
        image_1_351 <= io_pixelVal_in_1_3;
      end else if (10'h15f == _T_22[9:0]) begin
        image_1_351 <= io_pixelVal_in_1_2;
      end else if (10'h15f == _T_19[9:0]) begin
        image_1_351 <= io_pixelVal_in_1_1;
      end else if (10'h15f == _T_15[9:0]) begin
        image_1_351 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_352 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h160 == _T_37[9:0]) begin
        image_1_352 <= io_pixelVal_in_1_7;
      end else if (10'h160 == _T_34[9:0]) begin
        image_1_352 <= io_pixelVal_in_1_6;
      end else if (10'h160 == _T_31[9:0]) begin
        image_1_352 <= io_pixelVal_in_1_5;
      end else if (10'h160 == _T_28[9:0]) begin
        image_1_352 <= io_pixelVal_in_1_4;
      end else if (10'h160 == _T_25[9:0]) begin
        image_1_352 <= io_pixelVal_in_1_3;
      end else if (10'h160 == _T_22[9:0]) begin
        image_1_352 <= io_pixelVal_in_1_2;
      end else if (10'h160 == _T_19[9:0]) begin
        image_1_352 <= io_pixelVal_in_1_1;
      end else if (10'h160 == _T_15[9:0]) begin
        image_1_352 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_353 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h161 == _T_37[9:0]) begin
        image_1_353 <= io_pixelVal_in_1_7;
      end else if (10'h161 == _T_34[9:0]) begin
        image_1_353 <= io_pixelVal_in_1_6;
      end else if (10'h161 == _T_31[9:0]) begin
        image_1_353 <= io_pixelVal_in_1_5;
      end else if (10'h161 == _T_28[9:0]) begin
        image_1_353 <= io_pixelVal_in_1_4;
      end else if (10'h161 == _T_25[9:0]) begin
        image_1_353 <= io_pixelVal_in_1_3;
      end else if (10'h161 == _T_22[9:0]) begin
        image_1_353 <= io_pixelVal_in_1_2;
      end else if (10'h161 == _T_19[9:0]) begin
        image_1_353 <= io_pixelVal_in_1_1;
      end else if (10'h161 == _T_15[9:0]) begin
        image_1_353 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_354 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h162 == _T_37[9:0]) begin
        image_1_354 <= io_pixelVal_in_1_7;
      end else if (10'h162 == _T_34[9:0]) begin
        image_1_354 <= io_pixelVal_in_1_6;
      end else if (10'h162 == _T_31[9:0]) begin
        image_1_354 <= io_pixelVal_in_1_5;
      end else if (10'h162 == _T_28[9:0]) begin
        image_1_354 <= io_pixelVal_in_1_4;
      end else if (10'h162 == _T_25[9:0]) begin
        image_1_354 <= io_pixelVal_in_1_3;
      end else if (10'h162 == _T_22[9:0]) begin
        image_1_354 <= io_pixelVal_in_1_2;
      end else if (10'h162 == _T_19[9:0]) begin
        image_1_354 <= io_pixelVal_in_1_1;
      end else if (10'h162 == _T_15[9:0]) begin
        image_1_354 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_355 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h163 == _T_37[9:0]) begin
        image_1_355 <= io_pixelVal_in_1_7;
      end else if (10'h163 == _T_34[9:0]) begin
        image_1_355 <= io_pixelVal_in_1_6;
      end else if (10'h163 == _T_31[9:0]) begin
        image_1_355 <= io_pixelVal_in_1_5;
      end else if (10'h163 == _T_28[9:0]) begin
        image_1_355 <= io_pixelVal_in_1_4;
      end else if (10'h163 == _T_25[9:0]) begin
        image_1_355 <= io_pixelVal_in_1_3;
      end else if (10'h163 == _T_22[9:0]) begin
        image_1_355 <= io_pixelVal_in_1_2;
      end else if (10'h163 == _T_19[9:0]) begin
        image_1_355 <= io_pixelVal_in_1_1;
      end else if (10'h163 == _T_15[9:0]) begin
        image_1_355 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_356 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h164 == _T_37[9:0]) begin
        image_1_356 <= io_pixelVal_in_1_7;
      end else if (10'h164 == _T_34[9:0]) begin
        image_1_356 <= io_pixelVal_in_1_6;
      end else if (10'h164 == _T_31[9:0]) begin
        image_1_356 <= io_pixelVal_in_1_5;
      end else if (10'h164 == _T_28[9:0]) begin
        image_1_356 <= io_pixelVal_in_1_4;
      end else if (10'h164 == _T_25[9:0]) begin
        image_1_356 <= io_pixelVal_in_1_3;
      end else if (10'h164 == _T_22[9:0]) begin
        image_1_356 <= io_pixelVal_in_1_2;
      end else if (10'h164 == _T_19[9:0]) begin
        image_1_356 <= io_pixelVal_in_1_1;
      end else if (10'h164 == _T_15[9:0]) begin
        image_1_356 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_357 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h165 == _T_37[9:0]) begin
        image_1_357 <= io_pixelVal_in_1_7;
      end else if (10'h165 == _T_34[9:0]) begin
        image_1_357 <= io_pixelVal_in_1_6;
      end else if (10'h165 == _T_31[9:0]) begin
        image_1_357 <= io_pixelVal_in_1_5;
      end else if (10'h165 == _T_28[9:0]) begin
        image_1_357 <= io_pixelVal_in_1_4;
      end else if (10'h165 == _T_25[9:0]) begin
        image_1_357 <= io_pixelVal_in_1_3;
      end else if (10'h165 == _T_22[9:0]) begin
        image_1_357 <= io_pixelVal_in_1_2;
      end else if (10'h165 == _T_19[9:0]) begin
        image_1_357 <= io_pixelVal_in_1_1;
      end else if (10'h165 == _T_15[9:0]) begin
        image_1_357 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_358 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h166 == _T_37[9:0]) begin
        image_1_358 <= io_pixelVal_in_1_7;
      end else if (10'h166 == _T_34[9:0]) begin
        image_1_358 <= io_pixelVal_in_1_6;
      end else if (10'h166 == _T_31[9:0]) begin
        image_1_358 <= io_pixelVal_in_1_5;
      end else if (10'h166 == _T_28[9:0]) begin
        image_1_358 <= io_pixelVal_in_1_4;
      end else if (10'h166 == _T_25[9:0]) begin
        image_1_358 <= io_pixelVal_in_1_3;
      end else if (10'h166 == _T_22[9:0]) begin
        image_1_358 <= io_pixelVal_in_1_2;
      end else if (10'h166 == _T_19[9:0]) begin
        image_1_358 <= io_pixelVal_in_1_1;
      end else if (10'h166 == _T_15[9:0]) begin
        image_1_358 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_359 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h167 == _T_37[9:0]) begin
        image_1_359 <= io_pixelVal_in_1_7;
      end else if (10'h167 == _T_34[9:0]) begin
        image_1_359 <= io_pixelVal_in_1_6;
      end else if (10'h167 == _T_31[9:0]) begin
        image_1_359 <= io_pixelVal_in_1_5;
      end else if (10'h167 == _T_28[9:0]) begin
        image_1_359 <= io_pixelVal_in_1_4;
      end else if (10'h167 == _T_25[9:0]) begin
        image_1_359 <= io_pixelVal_in_1_3;
      end else if (10'h167 == _T_22[9:0]) begin
        image_1_359 <= io_pixelVal_in_1_2;
      end else if (10'h167 == _T_19[9:0]) begin
        image_1_359 <= io_pixelVal_in_1_1;
      end else if (10'h167 == _T_15[9:0]) begin
        image_1_359 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_360 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h168 == _T_37[9:0]) begin
        image_1_360 <= io_pixelVal_in_1_7;
      end else if (10'h168 == _T_34[9:0]) begin
        image_1_360 <= io_pixelVal_in_1_6;
      end else if (10'h168 == _T_31[9:0]) begin
        image_1_360 <= io_pixelVal_in_1_5;
      end else if (10'h168 == _T_28[9:0]) begin
        image_1_360 <= io_pixelVal_in_1_4;
      end else if (10'h168 == _T_25[9:0]) begin
        image_1_360 <= io_pixelVal_in_1_3;
      end else if (10'h168 == _T_22[9:0]) begin
        image_1_360 <= io_pixelVal_in_1_2;
      end else if (10'h168 == _T_19[9:0]) begin
        image_1_360 <= io_pixelVal_in_1_1;
      end else if (10'h168 == _T_15[9:0]) begin
        image_1_360 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_361 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h169 == _T_37[9:0]) begin
        image_1_361 <= io_pixelVal_in_1_7;
      end else if (10'h169 == _T_34[9:0]) begin
        image_1_361 <= io_pixelVal_in_1_6;
      end else if (10'h169 == _T_31[9:0]) begin
        image_1_361 <= io_pixelVal_in_1_5;
      end else if (10'h169 == _T_28[9:0]) begin
        image_1_361 <= io_pixelVal_in_1_4;
      end else if (10'h169 == _T_25[9:0]) begin
        image_1_361 <= io_pixelVal_in_1_3;
      end else if (10'h169 == _T_22[9:0]) begin
        image_1_361 <= io_pixelVal_in_1_2;
      end else if (10'h169 == _T_19[9:0]) begin
        image_1_361 <= io_pixelVal_in_1_1;
      end else if (10'h169 == _T_15[9:0]) begin
        image_1_361 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_362 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16a == _T_37[9:0]) begin
        image_1_362 <= io_pixelVal_in_1_7;
      end else if (10'h16a == _T_34[9:0]) begin
        image_1_362 <= io_pixelVal_in_1_6;
      end else if (10'h16a == _T_31[9:0]) begin
        image_1_362 <= io_pixelVal_in_1_5;
      end else if (10'h16a == _T_28[9:0]) begin
        image_1_362 <= io_pixelVal_in_1_4;
      end else if (10'h16a == _T_25[9:0]) begin
        image_1_362 <= io_pixelVal_in_1_3;
      end else if (10'h16a == _T_22[9:0]) begin
        image_1_362 <= io_pixelVal_in_1_2;
      end else if (10'h16a == _T_19[9:0]) begin
        image_1_362 <= io_pixelVal_in_1_1;
      end else if (10'h16a == _T_15[9:0]) begin
        image_1_362 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_363 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16b == _T_37[9:0]) begin
        image_1_363 <= io_pixelVal_in_1_7;
      end else if (10'h16b == _T_34[9:0]) begin
        image_1_363 <= io_pixelVal_in_1_6;
      end else if (10'h16b == _T_31[9:0]) begin
        image_1_363 <= io_pixelVal_in_1_5;
      end else if (10'h16b == _T_28[9:0]) begin
        image_1_363 <= io_pixelVal_in_1_4;
      end else if (10'h16b == _T_25[9:0]) begin
        image_1_363 <= io_pixelVal_in_1_3;
      end else if (10'h16b == _T_22[9:0]) begin
        image_1_363 <= io_pixelVal_in_1_2;
      end else if (10'h16b == _T_19[9:0]) begin
        image_1_363 <= io_pixelVal_in_1_1;
      end else if (10'h16b == _T_15[9:0]) begin
        image_1_363 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_364 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16c == _T_37[9:0]) begin
        image_1_364 <= io_pixelVal_in_1_7;
      end else if (10'h16c == _T_34[9:0]) begin
        image_1_364 <= io_pixelVal_in_1_6;
      end else if (10'h16c == _T_31[9:0]) begin
        image_1_364 <= io_pixelVal_in_1_5;
      end else if (10'h16c == _T_28[9:0]) begin
        image_1_364 <= io_pixelVal_in_1_4;
      end else if (10'h16c == _T_25[9:0]) begin
        image_1_364 <= io_pixelVal_in_1_3;
      end else if (10'h16c == _T_22[9:0]) begin
        image_1_364 <= io_pixelVal_in_1_2;
      end else if (10'h16c == _T_19[9:0]) begin
        image_1_364 <= io_pixelVal_in_1_1;
      end else if (10'h16c == _T_15[9:0]) begin
        image_1_364 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_365 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16d == _T_37[9:0]) begin
        image_1_365 <= io_pixelVal_in_1_7;
      end else if (10'h16d == _T_34[9:0]) begin
        image_1_365 <= io_pixelVal_in_1_6;
      end else if (10'h16d == _T_31[9:0]) begin
        image_1_365 <= io_pixelVal_in_1_5;
      end else if (10'h16d == _T_28[9:0]) begin
        image_1_365 <= io_pixelVal_in_1_4;
      end else if (10'h16d == _T_25[9:0]) begin
        image_1_365 <= io_pixelVal_in_1_3;
      end else if (10'h16d == _T_22[9:0]) begin
        image_1_365 <= io_pixelVal_in_1_2;
      end else if (10'h16d == _T_19[9:0]) begin
        image_1_365 <= io_pixelVal_in_1_1;
      end else if (10'h16d == _T_15[9:0]) begin
        image_1_365 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_366 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16e == _T_37[9:0]) begin
        image_1_366 <= io_pixelVal_in_1_7;
      end else if (10'h16e == _T_34[9:0]) begin
        image_1_366 <= io_pixelVal_in_1_6;
      end else if (10'h16e == _T_31[9:0]) begin
        image_1_366 <= io_pixelVal_in_1_5;
      end else if (10'h16e == _T_28[9:0]) begin
        image_1_366 <= io_pixelVal_in_1_4;
      end else if (10'h16e == _T_25[9:0]) begin
        image_1_366 <= io_pixelVal_in_1_3;
      end else if (10'h16e == _T_22[9:0]) begin
        image_1_366 <= io_pixelVal_in_1_2;
      end else if (10'h16e == _T_19[9:0]) begin
        image_1_366 <= io_pixelVal_in_1_1;
      end else if (10'h16e == _T_15[9:0]) begin
        image_1_366 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_367 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16f == _T_37[9:0]) begin
        image_1_367 <= io_pixelVal_in_1_7;
      end else if (10'h16f == _T_34[9:0]) begin
        image_1_367 <= io_pixelVal_in_1_6;
      end else if (10'h16f == _T_31[9:0]) begin
        image_1_367 <= io_pixelVal_in_1_5;
      end else if (10'h16f == _T_28[9:0]) begin
        image_1_367 <= io_pixelVal_in_1_4;
      end else if (10'h16f == _T_25[9:0]) begin
        image_1_367 <= io_pixelVal_in_1_3;
      end else if (10'h16f == _T_22[9:0]) begin
        image_1_367 <= io_pixelVal_in_1_2;
      end else if (10'h16f == _T_19[9:0]) begin
        image_1_367 <= io_pixelVal_in_1_1;
      end else if (10'h16f == _T_15[9:0]) begin
        image_1_367 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_368 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h170 == _T_37[9:0]) begin
        image_1_368 <= io_pixelVal_in_1_7;
      end else if (10'h170 == _T_34[9:0]) begin
        image_1_368 <= io_pixelVal_in_1_6;
      end else if (10'h170 == _T_31[9:0]) begin
        image_1_368 <= io_pixelVal_in_1_5;
      end else if (10'h170 == _T_28[9:0]) begin
        image_1_368 <= io_pixelVal_in_1_4;
      end else if (10'h170 == _T_25[9:0]) begin
        image_1_368 <= io_pixelVal_in_1_3;
      end else if (10'h170 == _T_22[9:0]) begin
        image_1_368 <= io_pixelVal_in_1_2;
      end else if (10'h170 == _T_19[9:0]) begin
        image_1_368 <= io_pixelVal_in_1_1;
      end else if (10'h170 == _T_15[9:0]) begin
        image_1_368 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_369 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h171 == _T_37[9:0]) begin
        image_1_369 <= io_pixelVal_in_1_7;
      end else if (10'h171 == _T_34[9:0]) begin
        image_1_369 <= io_pixelVal_in_1_6;
      end else if (10'h171 == _T_31[9:0]) begin
        image_1_369 <= io_pixelVal_in_1_5;
      end else if (10'h171 == _T_28[9:0]) begin
        image_1_369 <= io_pixelVal_in_1_4;
      end else if (10'h171 == _T_25[9:0]) begin
        image_1_369 <= io_pixelVal_in_1_3;
      end else if (10'h171 == _T_22[9:0]) begin
        image_1_369 <= io_pixelVal_in_1_2;
      end else if (10'h171 == _T_19[9:0]) begin
        image_1_369 <= io_pixelVal_in_1_1;
      end else if (10'h171 == _T_15[9:0]) begin
        image_1_369 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_370 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h172 == _T_37[9:0]) begin
        image_1_370 <= io_pixelVal_in_1_7;
      end else if (10'h172 == _T_34[9:0]) begin
        image_1_370 <= io_pixelVal_in_1_6;
      end else if (10'h172 == _T_31[9:0]) begin
        image_1_370 <= io_pixelVal_in_1_5;
      end else if (10'h172 == _T_28[9:0]) begin
        image_1_370 <= io_pixelVal_in_1_4;
      end else if (10'h172 == _T_25[9:0]) begin
        image_1_370 <= io_pixelVal_in_1_3;
      end else if (10'h172 == _T_22[9:0]) begin
        image_1_370 <= io_pixelVal_in_1_2;
      end else if (10'h172 == _T_19[9:0]) begin
        image_1_370 <= io_pixelVal_in_1_1;
      end else if (10'h172 == _T_15[9:0]) begin
        image_1_370 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_371 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h173 == _T_37[9:0]) begin
        image_1_371 <= io_pixelVal_in_1_7;
      end else if (10'h173 == _T_34[9:0]) begin
        image_1_371 <= io_pixelVal_in_1_6;
      end else if (10'h173 == _T_31[9:0]) begin
        image_1_371 <= io_pixelVal_in_1_5;
      end else if (10'h173 == _T_28[9:0]) begin
        image_1_371 <= io_pixelVal_in_1_4;
      end else if (10'h173 == _T_25[9:0]) begin
        image_1_371 <= io_pixelVal_in_1_3;
      end else if (10'h173 == _T_22[9:0]) begin
        image_1_371 <= io_pixelVal_in_1_2;
      end else if (10'h173 == _T_19[9:0]) begin
        image_1_371 <= io_pixelVal_in_1_1;
      end else if (10'h173 == _T_15[9:0]) begin
        image_1_371 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_372 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h174 == _T_37[9:0]) begin
        image_1_372 <= io_pixelVal_in_1_7;
      end else if (10'h174 == _T_34[9:0]) begin
        image_1_372 <= io_pixelVal_in_1_6;
      end else if (10'h174 == _T_31[9:0]) begin
        image_1_372 <= io_pixelVal_in_1_5;
      end else if (10'h174 == _T_28[9:0]) begin
        image_1_372 <= io_pixelVal_in_1_4;
      end else if (10'h174 == _T_25[9:0]) begin
        image_1_372 <= io_pixelVal_in_1_3;
      end else if (10'h174 == _T_22[9:0]) begin
        image_1_372 <= io_pixelVal_in_1_2;
      end else if (10'h174 == _T_19[9:0]) begin
        image_1_372 <= io_pixelVal_in_1_1;
      end else if (10'h174 == _T_15[9:0]) begin
        image_1_372 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_373 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h175 == _T_37[9:0]) begin
        image_1_373 <= io_pixelVal_in_1_7;
      end else if (10'h175 == _T_34[9:0]) begin
        image_1_373 <= io_pixelVal_in_1_6;
      end else if (10'h175 == _T_31[9:0]) begin
        image_1_373 <= io_pixelVal_in_1_5;
      end else if (10'h175 == _T_28[9:0]) begin
        image_1_373 <= io_pixelVal_in_1_4;
      end else if (10'h175 == _T_25[9:0]) begin
        image_1_373 <= io_pixelVal_in_1_3;
      end else if (10'h175 == _T_22[9:0]) begin
        image_1_373 <= io_pixelVal_in_1_2;
      end else if (10'h175 == _T_19[9:0]) begin
        image_1_373 <= io_pixelVal_in_1_1;
      end else if (10'h175 == _T_15[9:0]) begin
        image_1_373 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_374 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h176 == _T_37[9:0]) begin
        image_1_374 <= io_pixelVal_in_1_7;
      end else if (10'h176 == _T_34[9:0]) begin
        image_1_374 <= io_pixelVal_in_1_6;
      end else if (10'h176 == _T_31[9:0]) begin
        image_1_374 <= io_pixelVal_in_1_5;
      end else if (10'h176 == _T_28[9:0]) begin
        image_1_374 <= io_pixelVal_in_1_4;
      end else if (10'h176 == _T_25[9:0]) begin
        image_1_374 <= io_pixelVal_in_1_3;
      end else if (10'h176 == _T_22[9:0]) begin
        image_1_374 <= io_pixelVal_in_1_2;
      end else if (10'h176 == _T_19[9:0]) begin
        image_1_374 <= io_pixelVal_in_1_1;
      end else if (10'h176 == _T_15[9:0]) begin
        image_1_374 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_375 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h177 == _T_37[9:0]) begin
        image_1_375 <= io_pixelVal_in_1_7;
      end else if (10'h177 == _T_34[9:0]) begin
        image_1_375 <= io_pixelVal_in_1_6;
      end else if (10'h177 == _T_31[9:0]) begin
        image_1_375 <= io_pixelVal_in_1_5;
      end else if (10'h177 == _T_28[9:0]) begin
        image_1_375 <= io_pixelVal_in_1_4;
      end else if (10'h177 == _T_25[9:0]) begin
        image_1_375 <= io_pixelVal_in_1_3;
      end else if (10'h177 == _T_22[9:0]) begin
        image_1_375 <= io_pixelVal_in_1_2;
      end else if (10'h177 == _T_19[9:0]) begin
        image_1_375 <= io_pixelVal_in_1_1;
      end else if (10'h177 == _T_15[9:0]) begin
        image_1_375 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_376 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h178 == _T_37[9:0]) begin
        image_1_376 <= io_pixelVal_in_1_7;
      end else if (10'h178 == _T_34[9:0]) begin
        image_1_376 <= io_pixelVal_in_1_6;
      end else if (10'h178 == _T_31[9:0]) begin
        image_1_376 <= io_pixelVal_in_1_5;
      end else if (10'h178 == _T_28[9:0]) begin
        image_1_376 <= io_pixelVal_in_1_4;
      end else if (10'h178 == _T_25[9:0]) begin
        image_1_376 <= io_pixelVal_in_1_3;
      end else if (10'h178 == _T_22[9:0]) begin
        image_1_376 <= io_pixelVal_in_1_2;
      end else if (10'h178 == _T_19[9:0]) begin
        image_1_376 <= io_pixelVal_in_1_1;
      end else if (10'h178 == _T_15[9:0]) begin
        image_1_376 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_377 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h179 == _T_37[9:0]) begin
        image_1_377 <= io_pixelVal_in_1_7;
      end else if (10'h179 == _T_34[9:0]) begin
        image_1_377 <= io_pixelVal_in_1_6;
      end else if (10'h179 == _T_31[9:0]) begin
        image_1_377 <= io_pixelVal_in_1_5;
      end else if (10'h179 == _T_28[9:0]) begin
        image_1_377 <= io_pixelVal_in_1_4;
      end else if (10'h179 == _T_25[9:0]) begin
        image_1_377 <= io_pixelVal_in_1_3;
      end else if (10'h179 == _T_22[9:0]) begin
        image_1_377 <= io_pixelVal_in_1_2;
      end else if (10'h179 == _T_19[9:0]) begin
        image_1_377 <= io_pixelVal_in_1_1;
      end else if (10'h179 == _T_15[9:0]) begin
        image_1_377 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_378 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17a == _T_37[9:0]) begin
        image_1_378 <= io_pixelVal_in_1_7;
      end else if (10'h17a == _T_34[9:0]) begin
        image_1_378 <= io_pixelVal_in_1_6;
      end else if (10'h17a == _T_31[9:0]) begin
        image_1_378 <= io_pixelVal_in_1_5;
      end else if (10'h17a == _T_28[9:0]) begin
        image_1_378 <= io_pixelVal_in_1_4;
      end else if (10'h17a == _T_25[9:0]) begin
        image_1_378 <= io_pixelVal_in_1_3;
      end else if (10'h17a == _T_22[9:0]) begin
        image_1_378 <= io_pixelVal_in_1_2;
      end else if (10'h17a == _T_19[9:0]) begin
        image_1_378 <= io_pixelVal_in_1_1;
      end else if (10'h17a == _T_15[9:0]) begin
        image_1_378 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_379 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17b == _T_37[9:0]) begin
        image_1_379 <= io_pixelVal_in_1_7;
      end else if (10'h17b == _T_34[9:0]) begin
        image_1_379 <= io_pixelVal_in_1_6;
      end else if (10'h17b == _T_31[9:0]) begin
        image_1_379 <= io_pixelVal_in_1_5;
      end else if (10'h17b == _T_28[9:0]) begin
        image_1_379 <= io_pixelVal_in_1_4;
      end else if (10'h17b == _T_25[9:0]) begin
        image_1_379 <= io_pixelVal_in_1_3;
      end else if (10'h17b == _T_22[9:0]) begin
        image_1_379 <= io_pixelVal_in_1_2;
      end else if (10'h17b == _T_19[9:0]) begin
        image_1_379 <= io_pixelVal_in_1_1;
      end else if (10'h17b == _T_15[9:0]) begin
        image_1_379 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_380 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17c == _T_37[9:0]) begin
        image_1_380 <= io_pixelVal_in_1_7;
      end else if (10'h17c == _T_34[9:0]) begin
        image_1_380 <= io_pixelVal_in_1_6;
      end else if (10'h17c == _T_31[9:0]) begin
        image_1_380 <= io_pixelVal_in_1_5;
      end else if (10'h17c == _T_28[9:0]) begin
        image_1_380 <= io_pixelVal_in_1_4;
      end else if (10'h17c == _T_25[9:0]) begin
        image_1_380 <= io_pixelVal_in_1_3;
      end else if (10'h17c == _T_22[9:0]) begin
        image_1_380 <= io_pixelVal_in_1_2;
      end else if (10'h17c == _T_19[9:0]) begin
        image_1_380 <= io_pixelVal_in_1_1;
      end else if (10'h17c == _T_15[9:0]) begin
        image_1_380 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_381 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17d == _T_37[9:0]) begin
        image_1_381 <= io_pixelVal_in_1_7;
      end else if (10'h17d == _T_34[9:0]) begin
        image_1_381 <= io_pixelVal_in_1_6;
      end else if (10'h17d == _T_31[9:0]) begin
        image_1_381 <= io_pixelVal_in_1_5;
      end else if (10'h17d == _T_28[9:0]) begin
        image_1_381 <= io_pixelVal_in_1_4;
      end else if (10'h17d == _T_25[9:0]) begin
        image_1_381 <= io_pixelVal_in_1_3;
      end else if (10'h17d == _T_22[9:0]) begin
        image_1_381 <= io_pixelVal_in_1_2;
      end else if (10'h17d == _T_19[9:0]) begin
        image_1_381 <= io_pixelVal_in_1_1;
      end else if (10'h17d == _T_15[9:0]) begin
        image_1_381 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_382 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17e == _T_37[9:0]) begin
        image_1_382 <= io_pixelVal_in_1_7;
      end else if (10'h17e == _T_34[9:0]) begin
        image_1_382 <= io_pixelVal_in_1_6;
      end else if (10'h17e == _T_31[9:0]) begin
        image_1_382 <= io_pixelVal_in_1_5;
      end else if (10'h17e == _T_28[9:0]) begin
        image_1_382 <= io_pixelVal_in_1_4;
      end else if (10'h17e == _T_25[9:0]) begin
        image_1_382 <= io_pixelVal_in_1_3;
      end else if (10'h17e == _T_22[9:0]) begin
        image_1_382 <= io_pixelVal_in_1_2;
      end else if (10'h17e == _T_19[9:0]) begin
        image_1_382 <= io_pixelVal_in_1_1;
      end else if (10'h17e == _T_15[9:0]) begin
        image_1_382 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_383 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17f == _T_37[9:0]) begin
        image_1_383 <= io_pixelVal_in_1_7;
      end else if (10'h17f == _T_34[9:0]) begin
        image_1_383 <= io_pixelVal_in_1_6;
      end else if (10'h17f == _T_31[9:0]) begin
        image_1_383 <= io_pixelVal_in_1_5;
      end else if (10'h17f == _T_28[9:0]) begin
        image_1_383 <= io_pixelVal_in_1_4;
      end else if (10'h17f == _T_25[9:0]) begin
        image_1_383 <= io_pixelVal_in_1_3;
      end else if (10'h17f == _T_22[9:0]) begin
        image_1_383 <= io_pixelVal_in_1_2;
      end else if (10'h17f == _T_19[9:0]) begin
        image_1_383 <= io_pixelVal_in_1_1;
      end else if (10'h17f == _T_15[9:0]) begin
        image_1_383 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_384 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h180 == _T_37[9:0]) begin
        image_1_384 <= io_pixelVal_in_1_7;
      end else if (10'h180 == _T_34[9:0]) begin
        image_1_384 <= io_pixelVal_in_1_6;
      end else if (10'h180 == _T_31[9:0]) begin
        image_1_384 <= io_pixelVal_in_1_5;
      end else if (10'h180 == _T_28[9:0]) begin
        image_1_384 <= io_pixelVal_in_1_4;
      end else if (10'h180 == _T_25[9:0]) begin
        image_1_384 <= io_pixelVal_in_1_3;
      end else if (10'h180 == _T_22[9:0]) begin
        image_1_384 <= io_pixelVal_in_1_2;
      end else if (10'h180 == _T_19[9:0]) begin
        image_1_384 <= io_pixelVal_in_1_1;
      end else if (10'h180 == _T_15[9:0]) begin
        image_1_384 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_385 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h181 == _T_37[9:0]) begin
        image_1_385 <= io_pixelVal_in_1_7;
      end else if (10'h181 == _T_34[9:0]) begin
        image_1_385 <= io_pixelVal_in_1_6;
      end else if (10'h181 == _T_31[9:0]) begin
        image_1_385 <= io_pixelVal_in_1_5;
      end else if (10'h181 == _T_28[9:0]) begin
        image_1_385 <= io_pixelVal_in_1_4;
      end else if (10'h181 == _T_25[9:0]) begin
        image_1_385 <= io_pixelVal_in_1_3;
      end else if (10'h181 == _T_22[9:0]) begin
        image_1_385 <= io_pixelVal_in_1_2;
      end else if (10'h181 == _T_19[9:0]) begin
        image_1_385 <= io_pixelVal_in_1_1;
      end else if (10'h181 == _T_15[9:0]) begin
        image_1_385 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_386 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h182 == _T_37[9:0]) begin
        image_1_386 <= io_pixelVal_in_1_7;
      end else if (10'h182 == _T_34[9:0]) begin
        image_1_386 <= io_pixelVal_in_1_6;
      end else if (10'h182 == _T_31[9:0]) begin
        image_1_386 <= io_pixelVal_in_1_5;
      end else if (10'h182 == _T_28[9:0]) begin
        image_1_386 <= io_pixelVal_in_1_4;
      end else if (10'h182 == _T_25[9:0]) begin
        image_1_386 <= io_pixelVal_in_1_3;
      end else if (10'h182 == _T_22[9:0]) begin
        image_1_386 <= io_pixelVal_in_1_2;
      end else if (10'h182 == _T_19[9:0]) begin
        image_1_386 <= io_pixelVal_in_1_1;
      end else if (10'h182 == _T_15[9:0]) begin
        image_1_386 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_387 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h183 == _T_37[9:0]) begin
        image_1_387 <= io_pixelVal_in_1_7;
      end else if (10'h183 == _T_34[9:0]) begin
        image_1_387 <= io_pixelVal_in_1_6;
      end else if (10'h183 == _T_31[9:0]) begin
        image_1_387 <= io_pixelVal_in_1_5;
      end else if (10'h183 == _T_28[9:0]) begin
        image_1_387 <= io_pixelVal_in_1_4;
      end else if (10'h183 == _T_25[9:0]) begin
        image_1_387 <= io_pixelVal_in_1_3;
      end else if (10'h183 == _T_22[9:0]) begin
        image_1_387 <= io_pixelVal_in_1_2;
      end else if (10'h183 == _T_19[9:0]) begin
        image_1_387 <= io_pixelVal_in_1_1;
      end else if (10'h183 == _T_15[9:0]) begin
        image_1_387 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_388 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h184 == _T_37[9:0]) begin
        image_1_388 <= io_pixelVal_in_1_7;
      end else if (10'h184 == _T_34[9:0]) begin
        image_1_388 <= io_pixelVal_in_1_6;
      end else if (10'h184 == _T_31[9:0]) begin
        image_1_388 <= io_pixelVal_in_1_5;
      end else if (10'h184 == _T_28[9:0]) begin
        image_1_388 <= io_pixelVal_in_1_4;
      end else if (10'h184 == _T_25[9:0]) begin
        image_1_388 <= io_pixelVal_in_1_3;
      end else if (10'h184 == _T_22[9:0]) begin
        image_1_388 <= io_pixelVal_in_1_2;
      end else if (10'h184 == _T_19[9:0]) begin
        image_1_388 <= io_pixelVal_in_1_1;
      end else if (10'h184 == _T_15[9:0]) begin
        image_1_388 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_389 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h185 == _T_37[9:0]) begin
        image_1_389 <= io_pixelVal_in_1_7;
      end else if (10'h185 == _T_34[9:0]) begin
        image_1_389 <= io_pixelVal_in_1_6;
      end else if (10'h185 == _T_31[9:0]) begin
        image_1_389 <= io_pixelVal_in_1_5;
      end else if (10'h185 == _T_28[9:0]) begin
        image_1_389 <= io_pixelVal_in_1_4;
      end else if (10'h185 == _T_25[9:0]) begin
        image_1_389 <= io_pixelVal_in_1_3;
      end else if (10'h185 == _T_22[9:0]) begin
        image_1_389 <= io_pixelVal_in_1_2;
      end else if (10'h185 == _T_19[9:0]) begin
        image_1_389 <= io_pixelVal_in_1_1;
      end else if (10'h185 == _T_15[9:0]) begin
        image_1_389 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_390 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h186 == _T_37[9:0]) begin
        image_1_390 <= io_pixelVal_in_1_7;
      end else if (10'h186 == _T_34[9:0]) begin
        image_1_390 <= io_pixelVal_in_1_6;
      end else if (10'h186 == _T_31[9:0]) begin
        image_1_390 <= io_pixelVal_in_1_5;
      end else if (10'h186 == _T_28[9:0]) begin
        image_1_390 <= io_pixelVal_in_1_4;
      end else if (10'h186 == _T_25[9:0]) begin
        image_1_390 <= io_pixelVal_in_1_3;
      end else if (10'h186 == _T_22[9:0]) begin
        image_1_390 <= io_pixelVal_in_1_2;
      end else if (10'h186 == _T_19[9:0]) begin
        image_1_390 <= io_pixelVal_in_1_1;
      end else if (10'h186 == _T_15[9:0]) begin
        image_1_390 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_391 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h187 == _T_37[9:0]) begin
        image_1_391 <= io_pixelVal_in_1_7;
      end else if (10'h187 == _T_34[9:0]) begin
        image_1_391 <= io_pixelVal_in_1_6;
      end else if (10'h187 == _T_31[9:0]) begin
        image_1_391 <= io_pixelVal_in_1_5;
      end else if (10'h187 == _T_28[9:0]) begin
        image_1_391 <= io_pixelVal_in_1_4;
      end else if (10'h187 == _T_25[9:0]) begin
        image_1_391 <= io_pixelVal_in_1_3;
      end else if (10'h187 == _T_22[9:0]) begin
        image_1_391 <= io_pixelVal_in_1_2;
      end else if (10'h187 == _T_19[9:0]) begin
        image_1_391 <= io_pixelVal_in_1_1;
      end else if (10'h187 == _T_15[9:0]) begin
        image_1_391 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_392 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h188 == _T_37[9:0]) begin
        image_1_392 <= io_pixelVal_in_1_7;
      end else if (10'h188 == _T_34[9:0]) begin
        image_1_392 <= io_pixelVal_in_1_6;
      end else if (10'h188 == _T_31[9:0]) begin
        image_1_392 <= io_pixelVal_in_1_5;
      end else if (10'h188 == _T_28[9:0]) begin
        image_1_392 <= io_pixelVal_in_1_4;
      end else if (10'h188 == _T_25[9:0]) begin
        image_1_392 <= io_pixelVal_in_1_3;
      end else if (10'h188 == _T_22[9:0]) begin
        image_1_392 <= io_pixelVal_in_1_2;
      end else if (10'h188 == _T_19[9:0]) begin
        image_1_392 <= io_pixelVal_in_1_1;
      end else if (10'h188 == _T_15[9:0]) begin
        image_1_392 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_393 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h189 == _T_37[9:0]) begin
        image_1_393 <= io_pixelVal_in_1_7;
      end else if (10'h189 == _T_34[9:0]) begin
        image_1_393 <= io_pixelVal_in_1_6;
      end else if (10'h189 == _T_31[9:0]) begin
        image_1_393 <= io_pixelVal_in_1_5;
      end else if (10'h189 == _T_28[9:0]) begin
        image_1_393 <= io_pixelVal_in_1_4;
      end else if (10'h189 == _T_25[9:0]) begin
        image_1_393 <= io_pixelVal_in_1_3;
      end else if (10'h189 == _T_22[9:0]) begin
        image_1_393 <= io_pixelVal_in_1_2;
      end else if (10'h189 == _T_19[9:0]) begin
        image_1_393 <= io_pixelVal_in_1_1;
      end else if (10'h189 == _T_15[9:0]) begin
        image_1_393 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_394 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18a == _T_37[9:0]) begin
        image_1_394 <= io_pixelVal_in_1_7;
      end else if (10'h18a == _T_34[9:0]) begin
        image_1_394 <= io_pixelVal_in_1_6;
      end else if (10'h18a == _T_31[9:0]) begin
        image_1_394 <= io_pixelVal_in_1_5;
      end else if (10'h18a == _T_28[9:0]) begin
        image_1_394 <= io_pixelVal_in_1_4;
      end else if (10'h18a == _T_25[9:0]) begin
        image_1_394 <= io_pixelVal_in_1_3;
      end else if (10'h18a == _T_22[9:0]) begin
        image_1_394 <= io_pixelVal_in_1_2;
      end else if (10'h18a == _T_19[9:0]) begin
        image_1_394 <= io_pixelVal_in_1_1;
      end else if (10'h18a == _T_15[9:0]) begin
        image_1_394 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_395 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18b == _T_37[9:0]) begin
        image_1_395 <= io_pixelVal_in_1_7;
      end else if (10'h18b == _T_34[9:0]) begin
        image_1_395 <= io_pixelVal_in_1_6;
      end else if (10'h18b == _T_31[9:0]) begin
        image_1_395 <= io_pixelVal_in_1_5;
      end else if (10'h18b == _T_28[9:0]) begin
        image_1_395 <= io_pixelVal_in_1_4;
      end else if (10'h18b == _T_25[9:0]) begin
        image_1_395 <= io_pixelVal_in_1_3;
      end else if (10'h18b == _T_22[9:0]) begin
        image_1_395 <= io_pixelVal_in_1_2;
      end else if (10'h18b == _T_19[9:0]) begin
        image_1_395 <= io_pixelVal_in_1_1;
      end else if (10'h18b == _T_15[9:0]) begin
        image_1_395 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_396 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18c == _T_37[9:0]) begin
        image_1_396 <= io_pixelVal_in_1_7;
      end else if (10'h18c == _T_34[9:0]) begin
        image_1_396 <= io_pixelVal_in_1_6;
      end else if (10'h18c == _T_31[9:0]) begin
        image_1_396 <= io_pixelVal_in_1_5;
      end else if (10'h18c == _T_28[9:0]) begin
        image_1_396 <= io_pixelVal_in_1_4;
      end else if (10'h18c == _T_25[9:0]) begin
        image_1_396 <= io_pixelVal_in_1_3;
      end else if (10'h18c == _T_22[9:0]) begin
        image_1_396 <= io_pixelVal_in_1_2;
      end else if (10'h18c == _T_19[9:0]) begin
        image_1_396 <= io_pixelVal_in_1_1;
      end else if (10'h18c == _T_15[9:0]) begin
        image_1_396 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_397 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18d == _T_37[9:0]) begin
        image_1_397 <= io_pixelVal_in_1_7;
      end else if (10'h18d == _T_34[9:0]) begin
        image_1_397 <= io_pixelVal_in_1_6;
      end else if (10'h18d == _T_31[9:0]) begin
        image_1_397 <= io_pixelVal_in_1_5;
      end else if (10'h18d == _T_28[9:0]) begin
        image_1_397 <= io_pixelVal_in_1_4;
      end else if (10'h18d == _T_25[9:0]) begin
        image_1_397 <= io_pixelVal_in_1_3;
      end else if (10'h18d == _T_22[9:0]) begin
        image_1_397 <= io_pixelVal_in_1_2;
      end else if (10'h18d == _T_19[9:0]) begin
        image_1_397 <= io_pixelVal_in_1_1;
      end else if (10'h18d == _T_15[9:0]) begin
        image_1_397 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_398 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18e == _T_37[9:0]) begin
        image_1_398 <= io_pixelVal_in_1_7;
      end else if (10'h18e == _T_34[9:0]) begin
        image_1_398 <= io_pixelVal_in_1_6;
      end else if (10'h18e == _T_31[9:0]) begin
        image_1_398 <= io_pixelVal_in_1_5;
      end else if (10'h18e == _T_28[9:0]) begin
        image_1_398 <= io_pixelVal_in_1_4;
      end else if (10'h18e == _T_25[9:0]) begin
        image_1_398 <= io_pixelVal_in_1_3;
      end else if (10'h18e == _T_22[9:0]) begin
        image_1_398 <= io_pixelVal_in_1_2;
      end else if (10'h18e == _T_19[9:0]) begin
        image_1_398 <= io_pixelVal_in_1_1;
      end else if (10'h18e == _T_15[9:0]) begin
        image_1_398 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_399 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18f == _T_37[9:0]) begin
        image_1_399 <= io_pixelVal_in_1_7;
      end else if (10'h18f == _T_34[9:0]) begin
        image_1_399 <= io_pixelVal_in_1_6;
      end else if (10'h18f == _T_31[9:0]) begin
        image_1_399 <= io_pixelVal_in_1_5;
      end else if (10'h18f == _T_28[9:0]) begin
        image_1_399 <= io_pixelVal_in_1_4;
      end else if (10'h18f == _T_25[9:0]) begin
        image_1_399 <= io_pixelVal_in_1_3;
      end else if (10'h18f == _T_22[9:0]) begin
        image_1_399 <= io_pixelVal_in_1_2;
      end else if (10'h18f == _T_19[9:0]) begin
        image_1_399 <= io_pixelVal_in_1_1;
      end else if (10'h18f == _T_15[9:0]) begin
        image_1_399 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_400 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h190 == _T_37[9:0]) begin
        image_1_400 <= io_pixelVal_in_1_7;
      end else if (10'h190 == _T_34[9:0]) begin
        image_1_400 <= io_pixelVal_in_1_6;
      end else if (10'h190 == _T_31[9:0]) begin
        image_1_400 <= io_pixelVal_in_1_5;
      end else if (10'h190 == _T_28[9:0]) begin
        image_1_400 <= io_pixelVal_in_1_4;
      end else if (10'h190 == _T_25[9:0]) begin
        image_1_400 <= io_pixelVal_in_1_3;
      end else if (10'h190 == _T_22[9:0]) begin
        image_1_400 <= io_pixelVal_in_1_2;
      end else if (10'h190 == _T_19[9:0]) begin
        image_1_400 <= io_pixelVal_in_1_1;
      end else if (10'h190 == _T_15[9:0]) begin
        image_1_400 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_401 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h191 == _T_37[9:0]) begin
        image_1_401 <= io_pixelVal_in_1_7;
      end else if (10'h191 == _T_34[9:0]) begin
        image_1_401 <= io_pixelVal_in_1_6;
      end else if (10'h191 == _T_31[9:0]) begin
        image_1_401 <= io_pixelVal_in_1_5;
      end else if (10'h191 == _T_28[9:0]) begin
        image_1_401 <= io_pixelVal_in_1_4;
      end else if (10'h191 == _T_25[9:0]) begin
        image_1_401 <= io_pixelVal_in_1_3;
      end else if (10'h191 == _T_22[9:0]) begin
        image_1_401 <= io_pixelVal_in_1_2;
      end else if (10'h191 == _T_19[9:0]) begin
        image_1_401 <= io_pixelVal_in_1_1;
      end else if (10'h191 == _T_15[9:0]) begin
        image_1_401 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_402 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h192 == _T_37[9:0]) begin
        image_1_402 <= io_pixelVal_in_1_7;
      end else if (10'h192 == _T_34[9:0]) begin
        image_1_402 <= io_pixelVal_in_1_6;
      end else if (10'h192 == _T_31[9:0]) begin
        image_1_402 <= io_pixelVal_in_1_5;
      end else if (10'h192 == _T_28[9:0]) begin
        image_1_402 <= io_pixelVal_in_1_4;
      end else if (10'h192 == _T_25[9:0]) begin
        image_1_402 <= io_pixelVal_in_1_3;
      end else if (10'h192 == _T_22[9:0]) begin
        image_1_402 <= io_pixelVal_in_1_2;
      end else if (10'h192 == _T_19[9:0]) begin
        image_1_402 <= io_pixelVal_in_1_1;
      end else if (10'h192 == _T_15[9:0]) begin
        image_1_402 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_403 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h193 == _T_37[9:0]) begin
        image_1_403 <= io_pixelVal_in_1_7;
      end else if (10'h193 == _T_34[9:0]) begin
        image_1_403 <= io_pixelVal_in_1_6;
      end else if (10'h193 == _T_31[9:0]) begin
        image_1_403 <= io_pixelVal_in_1_5;
      end else if (10'h193 == _T_28[9:0]) begin
        image_1_403 <= io_pixelVal_in_1_4;
      end else if (10'h193 == _T_25[9:0]) begin
        image_1_403 <= io_pixelVal_in_1_3;
      end else if (10'h193 == _T_22[9:0]) begin
        image_1_403 <= io_pixelVal_in_1_2;
      end else if (10'h193 == _T_19[9:0]) begin
        image_1_403 <= io_pixelVal_in_1_1;
      end else if (10'h193 == _T_15[9:0]) begin
        image_1_403 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_404 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h194 == _T_37[9:0]) begin
        image_1_404 <= io_pixelVal_in_1_7;
      end else if (10'h194 == _T_34[9:0]) begin
        image_1_404 <= io_pixelVal_in_1_6;
      end else if (10'h194 == _T_31[9:0]) begin
        image_1_404 <= io_pixelVal_in_1_5;
      end else if (10'h194 == _T_28[9:0]) begin
        image_1_404 <= io_pixelVal_in_1_4;
      end else if (10'h194 == _T_25[9:0]) begin
        image_1_404 <= io_pixelVal_in_1_3;
      end else if (10'h194 == _T_22[9:0]) begin
        image_1_404 <= io_pixelVal_in_1_2;
      end else if (10'h194 == _T_19[9:0]) begin
        image_1_404 <= io_pixelVal_in_1_1;
      end else if (10'h194 == _T_15[9:0]) begin
        image_1_404 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_405 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h195 == _T_37[9:0]) begin
        image_1_405 <= io_pixelVal_in_1_7;
      end else if (10'h195 == _T_34[9:0]) begin
        image_1_405 <= io_pixelVal_in_1_6;
      end else if (10'h195 == _T_31[9:0]) begin
        image_1_405 <= io_pixelVal_in_1_5;
      end else if (10'h195 == _T_28[9:0]) begin
        image_1_405 <= io_pixelVal_in_1_4;
      end else if (10'h195 == _T_25[9:0]) begin
        image_1_405 <= io_pixelVal_in_1_3;
      end else if (10'h195 == _T_22[9:0]) begin
        image_1_405 <= io_pixelVal_in_1_2;
      end else if (10'h195 == _T_19[9:0]) begin
        image_1_405 <= io_pixelVal_in_1_1;
      end else if (10'h195 == _T_15[9:0]) begin
        image_1_405 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_406 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h196 == _T_37[9:0]) begin
        image_1_406 <= io_pixelVal_in_1_7;
      end else if (10'h196 == _T_34[9:0]) begin
        image_1_406 <= io_pixelVal_in_1_6;
      end else if (10'h196 == _T_31[9:0]) begin
        image_1_406 <= io_pixelVal_in_1_5;
      end else if (10'h196 == _T_28[9:0]) begin
        image_1_406 <= io_pixelVal_in_1_4;
      end else if (10'h196 == _T_25[9:0]) begin
        image_1_406 <= io_pixelVal_in_1_3;
      end else if (10'h196 == _T_22[9:0]) begin
        image_1_406 <= io_pixelVal_in_1_2;
      end else if (10'h196 == _T_19[9:0]) begin
        image_1_406 <= io_pixelVal_in_1_1;
      end else if (10'h196 == _T_15[9:0]) begin
        image_1_406 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_407 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h197 == _T_37[9:0]) begin
        image_1_407 <= io_pixelVal_in_1_7;
      end else if (10'h197 == _T_34[9:0]) begin
        image_1_407 <= io_pixelVal_in_1_6;
      end else if (10'h197 == _T_31[9:0]) begin
        image_1_407 <= io_pixelVal_in_1_5;
      end else if (10'h197 == _T_28[9:0]) begin
        image_1_407 <= io_pixelVal_in_1_4;
      end else if (10'h197 == _T_25[9:0]) begin
        image_1_407 <= io_pixelVal_in_1_3;
      end else if (10'h197 == _T_22[9:0]) begin
        image_1_407 <= io_pixelVal_in_1_2;
      end else if (10'h197 == _T_19[9:0]) begin
        image_1_407 <= io_pixelVal_in_1_1;
      end else if (10'h197 == _T_15[9:0]) begin
        image_1_407 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_408 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h198 == _T_37[9:0]) begin
        image_1_408 <= io_pixelVal_in_1_7;
      end else if (10'h198 == _T_34[9:0]) begin
        image_1_408 <= io_pixelVal_in_1_6;
      end else if (10'h198 == _T_31[9:0]) begin
        image_1_408 <= io_pixelVal_in_1_5;
      end else if (10'h198 == _T_28[9:0]) begin
        image_1_408 <= io_pixelVal_in_1_4;
      end else if (10'h198 == _T_25[9:0]) begin
        image_1_408 <= io_pixelVal_in_1_3;
      end else if (10'h198 == _T_22[9:0]) begin
        image_1_408 <= io_pixelVal_in_1_2;
      end else if (10'h198 == _T_19[9:0]) begin
        image_1_408 <= io_pixelVal_in_1_1;
      end else if (10'h198 == _T_15[9:0]) begin
        image_1_408 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_409 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h199 == _T_37[9:0]) begin
        image_1_409 <= io_pixelVal_in_1_7;
      end else if (10'h199 == _T_34[9:0]) begin
        image_1_409 <= io_pixelVal_in_1_6;
      end else if (10'h199 == _T_31[9:0]) begin
        image_1_409 <= io_pixelVal_in_1_5;
      end else if (10'h199 == _T_28[9:0]) begin
        image_1_409 <= io_pixelVal_in_1_4;
      end else if (10'h199 == _T_25[9:0]) begin
        image_1_409 <= io_pixelVal_in_1_3;
      end else if (10'h199 == _T_22[9:0]) begin
        image_1_409 <= io_pixelVal_in_1_2;
      end else if (10'h199 == _T_19[9:0]) begin
        image_1_409 <= io_pixelVal_in_1_1;
      end else if (10'h199 == _T_15[9:0]) begin
        image_1_409 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_410 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19a == _T_37[9:0]) begin
        image_1_410 <= io_pixelVal_in_1_7;
      end else if (10'h19a == _T_34[9:0]) begin
        image_1_410 <= io_pixelVal_in_1_6;
      end else if (10'h19a == _T_31[9:0]) begin
        image_1_410 <= io_pixelVal_in_1_5;
      end else if (10'h19a == _T_28[9:0]) begin
        image_1_410 <= io_pixelVal_in_1_4;
      end else if (10'h19a == _T_25[9:0]) begin
        image_1_410 <= io_pixelVal_in_1_3;
      end else if (10'h19a == _T_22[9:0]) begin
        image_1_410 <= io_pixelVal_in_1_2;
      end else if (10'h19a == _T_19[9:0]) begin
        image_1_410 <= io_pixelVal_in_1_1;
      end else if (10'h19a == _T_15[9:0]) begin
        image_1_410 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_411 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19b == _T_37[9:0]) begin
        image_1_411 <= io_pixelVal_in_1_7;
      end else if (10'h19b == _T_34[9:0]) begin
        image_1_411 <= io_pixelVal_in_1_6;
      end else if (10'h19b == _T_31[9:0]) begin
        image_1_411 <= io_pixelVal_in_1_5;
      end else if (10'h19b == _T_28[9:0]) begin
        image_1_411 <= io_pixelVal_in_1_4;
      end else if (10'h19b == _T_25[9:0]) begin
        image_1_411 <= io_pixelVal_in_1_3;
      end else if (10'h19b == _T_22[9:0]) begin
        image_1_411 <= io_pixelVal_in_1_2;
      end else if (10'h19b == _T_19[9:0]) begin
        image_1_411 <= io_pixelVal_in_1_1;
      end else if (10'h19b == _T_15[9:0]) begin
        image_1_411 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_412 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19c == _T_37[9:0]) begin
        image_1_412 <= io_pixelVal_in_1_7;
      end else if (10'h19c == _T_34[9:0]) begin
        image_1_412 <= io_pixelVal_in_1_6;
      end else if (10'h19c == _T_31[9:0]) begin
        image_1_412 <= io_pixelVal_in_1_5;
      end else if (10'h19c == _T_28[9:0]) begin
        image_1_412 <= io_pixelVal_in_1_4;
      end else if (10'h19c == _T_25[9:0]) begin
        image_1_412 <= io_pixelVal_in_1_3;
      end else if (10'h19c == _T_22[9:0]) begin
        image_1_412 <= io_pixelVal_in_1_2;
      end else if (10'h19c == _T_19[9:0]) begin
        image_1_412 <= io_pixelVal_in_1_1;
      end else if (10'h19c == _T_15[9:0]) begin
        image_1_412 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_413 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19d == _T_37[9:0]) begin
        image_1_413 <= io_pixelVal_in_1_7;
      end else if (10'h19d == _T_34[9:0]) begin
        image_1_413 <= io_pixelVal_in_1_6;
      end else if (10'h19d == _T_31[9:0]) begin
        image_1_413 <= io_pixelVal_in_1_5;
      end else if (10'h19d == _T_28[9:0]) begin
        image_1_413 <= io_pixelVal_in_1_4;
      end else if (10'h19d == _T_25[9:0]) begin
        image_1_413 <= io_pixelVal_in_1_3;
      end else if (10'h19d == _T_22[9:0]) begin
        image_1_413 <= io_pixelVal_in_1_2;
      end else if (10'h19d == _T_19[9:0]) begin
        image_1_413 <= io_pixelVal_in_1_1;
      end else if (10'h19d == _T_15[9:0]) begin
        image_1_413 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_414 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19e == _T_37[9:0]) begin
        image_1_414 <= io_pixelVal_in_1_7;
      end else if (10'h19e == _T_34[9:0]) begin
        image_1_414 <= io_pixelVal_in_1_6;
      end else if (10'h19e == _T_31[9:0]) begin
        image_1_414 <= io_pixelVal_in_1_5;
      end else if (10'h19e == _T_28[9:0]) begin
        image_1_414 <= io_pixelVal_in_1_4;
      end else if (10'h19e == _T_25[9:0]) begin
        image_1_414 <= io_pixelVal_in_1_3;
      end else if (10'h19e == _T_22[9:0]) begin
        image_1_414 <= io_pixelVal_in_1_2;
      end else if (10'h19e == _T_19[9:0]) begin
        image_1_414 <= io_pixelVal_in_1_1;
      end else if (10'h19e == _T_15[9:0]) begin
        image_1_414 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_415 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19f == _T_37[9:0]) begin
        image_1_415 <= io_pixelVal_in_1_7;
      end else if (10'h19f == _T_34[9:0]) begin
        image_1_415 <= io_pixelVal_in_1_6;
      end else if (10'h19f == _T_31[9:0]) begin
        image_1_415 <= io_pixelVal_in_1_5;
      end else if (10'h19f == _T_28[9:0]) begin
        image_1_415 <= io_pixelVal_in_1_4;
      end else if (10'h19f == _T_25[9:0]) begin
        image_1_415 <= io_pixelVal_in_1_3;
      end else if (10'h19f == _T_22[9:0]) begin
        image_1_415 <= io_pixelVal_in_1_2;
      end else if (10'h19f == _T_19[9:0]) begin
        image_1_415 <= io_pixelVal_in_1_1;
      end else if (10'h19f == _T_15[9:0]) begin
        image_1_415 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_416 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a0 == _T_37[9:0]) begin
        image_1_416 <= io_pixelVal_in_1_7;
      end else if (10'h1a0 == _T_34[9:0]) begin
        image_1_416 <= io_pixelVal_in_1_6;
      end else if (10'h1a0 == _T_31[9:0]) begin
        image_1_416 <= io_pixelVal_in_1_5;
      end else if (10'h1a0 == _T_28[9:0]) begin
        image_1_416 <= io_pixelVal_in_1_4;
      end else if (10'h1a0 == _T_25[9:0]) begin
        image_1_416 <= io_pixelVal_in_1_3;
      end else if (10'h1a0 == _T_22[9:0]) begin
        image_1_416 <= io_pixelVal_in_1_2;
      end else if (10'h1a0 == _T_19[9:0]) begin
        image_1_416 <= io_pixelVal_in_1_1;
      end else if (10'h1a0 == _T_15[9:0]) begin
        image_1_416 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_417 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a1 == _T_37[9:0]) begin
        image_1_417 <= io_pixelVal_in_1_7;
      end else if (10'h1a1 == _T_34[9:0]) begin
        image_1_417 <= io_pixelVal_in_1_6;
      end else if (10'h1a1 == _T_31[9:0]) begin
        image_1_417 <= io_pixelVal_in_1_5;
      end else if (10'h1a1 == _T_28[9:0]) begin
        image_1_417 <= io_pixelVal_in_1_4;
      end else if (10'h1a1 == _T_25[9:0]) begin
        image_1_417 <= io_pixelVal_in_1_3;
      end else if (10'h1a1 == _T_22[9:0]) begin
        image_1_417 <= io_pixelVal_in_1_2;
      end else if (10'h1a1 == _T_19[9:0]) begin
        image_1_417 <= io_pixelVal_in_1_1;
      end else if (10'h1a1 == _T_15[9:0]) begin
        image_1_417 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_418 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a2 == _T_37[9:0]) begin
        image_1_418 <= io_pixelVal_in_1_7;
      end else if (10'h1a2 == _T_34[9:0]) begin
        image_1_418 <= io_pixelVal_in_1_6;
      end else if (10'h1a2 == _T_31[9:0]) begin
        image_1_418 <= io_pixelVal_in_1_5;
      end else if (10'h1a2 == _T_28[9:0]) begin
        image_1_418 <= io_pixelVal_in_1_4;
      end else if (10'h1a2 == _T_25[9:0]) begin
        image_1_418 <= io_pixelVal_in_1_3;
      end else if (10'h1a2 == _T_22[9:0]) begin
        image_1_418 <= io_pixelVal_in_1_2;
      end else if (10'h1a2 == _T_19[9:0]) begin
        image_1_418 <= io_pixelVal_in_1_1;
      end else if (10'h1a2 == _T_15[9:0]) begin
        image_1_418 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_419 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a3 == _T_37[9:0]) begin
        image_1_419 <= io_pixelVal_in_1_7;
      end else if (10'h1a3 == _T_34[9:0]) begin
        image_1_419 <= io_pixelVal_in_1_6;
      end else if (10'h1a3 == _T_31[9:0]) begin
        image_1_419 <= io_pixelVal_in_1_5;
      end else if (10'h1a3 == _T_28[9:0]) begin
        image_1_419 <= io_pixelVal_in_1_4;
      end else if (10'h1a3 == _T_25[9:0]) begin
        image_1_419 <= io_pixelVal_in_1_3;
      end else if (10'h1a3 == _T_22[9:0]) begin
        image_1_419 <= io_pixelVal_in_1_2;
      end else if (10'h1a3 == _T_19[9:0]) begin
        image_1_419 <= io_pixelVal_in_1_1;
      end else if (10'h1a3 == _T_15[9:0]) begin
        image_1_419 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_420 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a4 == _T_37[9:0]) begin
        image_1_420 <= io_pixelVal_in_1_7;
      end else if (10'h1a4 == _T_34[9:0]) begin
        image_1_420 <= io_pixelVal_in_1_6;
      end else if (10'h1a4 == _T_31[9:0]) begin
        image_1_420 <= io_pixelVal_in_1_5;
      end else if (10'h1a4 == _T_28[9:0]) begin
        image_1_420 <= io_pixelVal_in_1_4;
      end else if (10'h1a4 == _T_25[9:0]) begin
        image_1_420 <= io_pixelVal_in_1_3;
      end else if (10'h1a4 == _T_22[9:0]) begin
        image_1_420 <= io_pixelVal_in_1_2;
      end else if (10'h1a4 == _T_19[9:0]) begin
        image_1_420 <= io_pixelVal_in_1_1;
      end else if (10'h1a4 == _T_15[9:0]) begin
        image_1_420 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_421 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a5 == _T_37[9:0]) begin
        image_1_421 <= io_pixelVal_in_1_7;
      end else if (10'h1a5 == _T_34[9:0]) begin
        image_1_421 <= io_pixelVal_in_1_6;
      end else if (10'h1a5 == _T_31[9:0]) begin
        image_1_421 <= io_pixelVal_in_1_5;
      end else if (10'h1a5 == _T_28[9:0]) begin
        image_1_421 <= io_pixelVal_in_1_4;
      end else if (10'h1a5 == _T_25[9:0]) begin
        image_1_421 <= io_pixelVal_in_1_3;
      end else if (10'h1a5 == _T_22[9:0]) begin
        image_1_421 <= io_pixelVal_in_1_2;
      end else if (10'h1a5 == _T_19[9:0]) begin
        image_1_421 <= io_pixelVal_in_1_1;
      end else if (10'h1a5 == _T_15[9:0]) begin
        image_1_421 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_422 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a6 == _T_37[9:0]) begin
        image_1_422 <= io_pixelVal_in_1_7;
      end else if (10'h1a6 == _T_34[9:0]) begin
        image_1_422 <= io_pixelVal_in_1_6;
      end else if (10'h1a6 == _T_31[9:0]) begin
        image_1_422 <= io_pixelVal_in_1_5;
      end else if (10'h1a6 == _T_28[9:0]) begin
        image_1_422 <= io_pixelVal_in_1_4;
      end else if (10'h1a6 == _T_25[9:0]) begin
        image_1_422 <= io_pixelVal_in_1_3;
      end else if (10'h1a6 == _T_22[9:0]) begin
        image_1_422 <= io_pixelVal_in_1_2;
      end else if (10'h1a6 == _T_19[9:0]) begin
        image_1_422 <= io_pixelVal_in_1_1;
      end else if (10'h1a6 == _T_15[9:0]) begin
        image_1_422 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_423 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a7 == _T_37[9:0]) begin
        image_1_423 <= io_pixelVal_in_1_7;
      end else if (10'h1a7 == _T_34[9:0]) begin
        image_1_423 <= io_pixelVal_in_1_6;
      end else if (10'h1a7 == _T_31[9:0]) begin
        image_1_423 <= io_pixelVal_in_1_5;
      end else if (10'h1a7 == _T_28[9:0]) begin
        image_1_423 <= io_pixelVal_in_1_4;
      end else if (10'h1a7 == _T_25[9:0]) begin
        image_1_423 <= io_pixelVal_in_1_3;
      end else if (10'h1a7 == _T_22[9:0]) begin
        image_1_423 <= io_pixelVal_in_1_2;
      end else if (10'h1a7 == _T_19[9:0]) begin
        image_1_423 <= io_pixelVal_in_1_1;
      end else if (10'h1a7 == _T_15[9:0]) begin
        image_1_423 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_424 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a8 == _T_37[9:0]) begin
        image_1_424 <= io_pixelVal_in_1_7;
      end else if (10'h1a8 == _T_34[9:0]) begin
        image_1_424 <= io_pixelVal_in_1_6;
      end else if (10'h1a8 == _T_31[9:0]) begin
        image_1_424 <= io_pixelVal_in_1_5;
      end else if (10'h1a8 == _T_28[9:0]) begin
        image_1_424 <= io_pixelVal_in_1_4;
      end else if (10'h1a8 == _T_25[9:0]) begin
        image_1_424 <= io_pixelVal_in_1_3;
      end else if (10'h1a8 == _T_22[9:0]) begin
        image_1_424 <= io_pixelVal_in_1_2;
      end else if (10'h1a8 == _T_19[9:0]) begin
        image_1_424 <= io_pixelVal_in_1_1;
      end else if (10'h1a8 == _T_15[9:0]) begin
        image_1_424 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_425 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a9 == _T_37[9:0]) begin
        image_1_425 <= io_pixelVal_in_1_7;
      end else if (10'h1a9 == _T_34[9:0]) begin
        image_1_425 <= io_pixelVal_in_1_6;
      end else if (10'h1a9 == _T_31[9:0]) begin
        image_1_425 <= io_pixelVal_in_1_5;
      end else if (10'h1a9 == _T_28[9:0]) begin
        image_1_425 <= io_pixelVal_in_1_4;
      end else if (10'h1a9 == _T_25[9:0]) begin
        image_1_425 <= io_pixelVal_in_1_3;
      end else if (10'h1a9 == _T_22[9:0]) begin
        image_1_425 <= io_pixelVal_in_1_2;
      end else if (10'h1a9 == _T_19[9:0]) begin
        image_1_425 <= io_pixelVal_in_1_1;
      end else if (10'h1a9 == _T_15[9:0]) begin
        image_1_425 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_426 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1aa == _T_37[9:0]) begin
        image_1_426 <= io_pixelVal_in_1_7;
      end else if (10'h1aa == _T_34[9:0]) begin
        image_1_426 <= io_pixelVal_in_1_6;
      end else if (10'h1aa == _T_31[9:0]) begin
        image_1_426 <= io_pixelVal_in_1_5;
      end else if (10'h1aa == _T_28[9:0]) begin
        image_1_426 <= io_pixelVal_in_1_4;
      end else if (10'h1aa == _T_25[9:0]) begin
        image_1_426 <= io_pixelVal_in_1_3;
      end else if (10'h1aa == _T_22[9:0]) begin
        image_1_426 <= io_pixelVal_in_1_2;
      end else if (10'h1aa == _T_19[9:0]) begin
        image_1_426 <= io_pixelVal_in_1_1;
      end else if (10'h1aa == _T_15[9:0]) begin
        image_1_426 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_427 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ab == _T_37[9:0]) begin
        image_1_427 <= io_pixelVal_in_1_7;
      end else if (10'h1ab == _T_34[9:0]) begin
        image_1_427 <= io_pixelVal_in_1_6;
      end else if (10'h1ab == _T_31[9:0]) begin
        image_1_427 <= io_pixelVal_in_1_5;
      end else if (10'h1ab == _T_28[9:0]) begin
        image_1_427 <= io_pixelVal_in_1_4;
      end else if (10'h1ab == _T_25[9:0]) begin
        image_1_427 <= io_pixelVal_in_1_3;
      end else if (10'h1ab == _T_22[9:0]) begin
        image_1_427 <= io_pixelVal_in_1_2;
      end else if (10'h1ab == _T_19[9:0]) begin
        image_1_427 <= io_pixelVal_in_1_1;
      end else if (10'h1ab == _T_15[9:0]) begin
        image_1_427 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_428 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ac == _T_37[9:0]) begin
        image_1_428 <= io_pixelVal_in_1_7;
      end else if (10'h1ac == _T_34[9:0]) begin
        image_1_428 <= io_pixelVal_in_1_6;
      end else if (10'h1ac == _T_31[9:0]) begin
        image_1_428 <= io_pixelVal_in_1_5;
      end else if (10'h1ac == _T_28[9:0]) begin
        image_1_428 <= io_pixelVal_in_1_4;
      end else if (10'h1ac == _T_25[9:0]) begin
        image_1_428 <= io_pixelVal_in_1_3;
      end else if (10'h1ac == _T_22[9:0]) begin
        image_1_428 <= io_pixelVal_in_1_2;
      end else if (10'h1ac == _T_19[9:0]) begin
        image_1_428 <= io_pixelVal_in_1_1;
      end else if (10'h1ac == _T_15[9:0]) begin
        image_1_428 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_429 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ad == _T_37[9:0]) begin
        image_1_429 <= io_pixelVal_in_1_7;
      end else if (10'h1ad == _T_34[9:0]) begin
        image_1_429 <= io_pixelVal_in_1_6;
      end else if (10'h1ad == _T_31[9:0]) begin
        image_1_429 <= io_pixelVal_in_1_5;
      end else if (10'h1ad == _T_28[9:0]) begin
        image_1_429 <= io_pixelVal_in_1_4;
      end else if (10'h1ad == _T_25[9:0]) begin
        image_1_429 <= io_pixelVal_in_1_3;
      end else if (10'h1ad == _T_22[9:0]) begin
        image_1_429 <= io_pixelVal_in_1_2;
      end else if (10'h1ad == _T_19[9:0]) begin
        image_1_429 <= io_pixelVal_in_1_1;
      end else if (10'h1ad == _T_15[9:0]) begin
        image_1_429 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_430 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ae == _T_37[9:0]) begin
        image_1_430 <= io_pixelVal_in_1_7;
      end else if (10'h1ae == _T_34[9:0]) begin
        image_1_430 <= io_pixelVal_in_1_6;
      end else if (10'h1ae == _T_31[9:0]) begin
        image_1_430 <= io_pixelVal_in_1_5;
      end else if (10'h1ae == _T_28[9:0]) begin
        image_1_430 <= io_pixelVal_in_1_4;
      end else if (10'h1ae == _T_25[9:0]) begin
        image_1_430 <= io_pixelVal_in_1_3;
      end else if (10'h1ae == _T_22[9:0]) begin
        image_1_430 <= io_pixelVal_in_1_2;
      end else if (10'h1ae == _T_19[9:0]) begin
        image_1_430 <= io_pixelVal_in_1_1;
      end else if (10'h1ae == _T_15[9:0]) begin
        image_1_430 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_431 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1af == _T_37[9:0]) begin
        image_1_431 <= io_pixelVal_in_1_7;
      end else if (10'h1af == _T_34[9:0]) begin
        image_1_431 <= io_pixelVal_in_1_6;
      end else if (10'h1af == _T_31[9:0]) begin
        image_1_431 <= io_pixelVal_in_1_5;
      end else if (10'h1af == _T_28[9:0]) begin
        image_1_431 <= io_pixelVal_in_1_4;
      end else if (10'h1af == _T_25[9:0]) begin
        image_1_431 <= io_pixelVal_in_1_3;
      end else if (10'h1af == _T_22[9:0]) begin
        image_1_431 <= io_pixelVal_in_1_2;
      end else if (10'h1af == _T_19[9:0]) begin
        image_1_431 <= io_pixelVal_in_1_1;
      end else if (10'h1af == _T_15[9:0]) begin
        image_1_431 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_432 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b0 == _T_37[9:0]) begin
        image_1_432 <= io_pixelVal_in_1_7;
      end else if (10'h1b0 == _T_34[9:0]) begin
        image_1_432 <= io_pixelVal_in_1_6;
      end else if (10'h1b0 == _T_31[9:0]) begin
        image_1_432 <= io_pixelVal_in_1_5;
      end else if (10'h1b0 == _T_28[9:0]) begin
        image_1_432 <= io_pixelVal_in_1_4;
      end else if (10'h1b0 == _T_25[9:0]) begin
        image_1_432 <= io_pixelVal_in_1_3;
      end else if (10'h1b0 == _T_22[9:0]) begin
        image_1_432 <= io_pixelVal_in_1_2;
      end else if (10'h1b0 == _T_19[9:0]) begin
        image_1_432 <= io_pixelVal_in_1_1;
      end else if (10'h1b0 == _T_15[9:0]) begin
        image_1_432 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_433 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b1 == _T_37[9:0]) begin
        image_1_433 <= io_pixelVal_in_1_7;
      end else if (10'h1b1 == _T_34[9:0]) begin
        image_1_433 <= io_pixelVal_in_1_6;
      end else if (10'h1b1 == _T_31[9:0]) begin
        image_1_433 <= io_pixelVal_in_1_5;
      end else if (10'h1b1 == _T_28[9:0]) begin
        image_1_433 <= io_pixelVal_in_1_4;
      end else if (10'h1b1 == _T_25[9:0]) begin
        image_1_433 <= io_pixelVal_in_1_3;
      end else if (10'h1b1 == _T_22[9:0]) begin
        image_1_433 <= io_pixelVal_in_1_2;
      end else if (10'h1b1 == _T_19[9:0]) begin
        image_1_433 <= io_pixelVal_in_1_1;
      end else if (10'h1b1 == _T_15[9:0]) begin
        image_1_433 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_434 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b2 == _T_37[9:0]) begin
        image_1_434 <= io_pixelVal_in_1_7;
      end else if (10'h1b2 == _T_34[9:0]) begin
        image_1_434 <= io_pixelVal_in_1_6;
      end else if (10'h1b2 == _T_31[9:0]) begin
        image_1_434 <= io_pixelVal_in_1_5;
      end else if (10'h1b2 == _T_28[9:0]) begin
        image_1_434 <= io_pixelVal_in_1_4;
      end else if (10'h1b2 == _T_25[9:0]) begin
        image_1_434 <= io_pixelVal_in_1_3;
      end else if (10'h1b2 == _T_22[9:0]) begin
        image_1_434 <= io_pixelVal_in_1_2;
      end else if (10'h1b2 == _T_19[9:0]) begin
        image_1_434 <= io_pixelVal_in_1_1;
      end else if (10'h1b2 == _T_15[9:0]) begin
        image_1_434 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_435 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b3 == _T_37[9:0]) begin
        image_1_435 <= io_pixelVal_in_1_7;
      end else if (10'h1b3 == _T_34[9:0]) begin
        image_1_435 <= io_pixelVal_in_1_6;
      end else if (10'h1b3 == _T_31[9:0]) begin
        image_1_435 <= io_pixelVal_in_1_5;
      end else if (10'h1b3 == _T_28[9:0]) begin
        image_1_435 <= io_pixelVal_in_1_4;
      end else if (10'h1b3 == _T_25[9:0]) begin
        image_1_435 <= io_pixelVal_in_1_3;
      end else if (10'h1b3 == _T_22[9:0]) begin
        image_1_435 <= io_pixelVal_in_1_2;
      end else if (10'h1b3 == _T_19[9:0]) begin
        image_1_435 <= io_pixelVal_in_1_1;
      end else if (10'h1b3 == _T_15[9:0]) begin
        image_1_435 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_436 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b4 == _T_37[9:0]) begin
        image_1_436 <= io_pixelVal_in_1_7;
      end else if (10'h1b4 == _T_34[9:0]) begin
        image_1_436 <= io_pixelVal_in_1_6;
      end else if (10'h1b4 == _T_31[9:0]) begin
        image_1_436 <= io_pixelVal_in_1_5;
      end else if (10'h1b4 == _T_28[9:0]) begin
        image_1_436 <= io_pixelVal_in_1_4;
      end else if (10'h1b4 == _T_25[9:0]) begin
        image_1_436 <= io_pixelVal_in_1_3;
      end else if (10'h1b4 == _T_22[9:0]) begin
        image_1_436 <= io_pixelVal_in_1_2;
      end else if (10'h1b4 == _T_19[9:0]) begin
        image_1_436 <= io_pixelVal_in_1_1;
      end else if (10'h1b4 == _T_15[9:0]) begin
        image_1_436 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_437 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b5 == _T_37[9:0]) begin
        image_1_437 <= io_pixelVal_in_1_7;
      end else if (10'h1b5 == _T_34[9:0]) begin
        image_1_437 <= io_pixelVal_in_1_6;
      end else if (10'h1b5 == _T_31[9:0]) begin
        image_1_437 <= io_pixelVal_in_1_5;
      end else if (10'h1b5 == _T_28[9:0]) begin
        image_1_437 <= io_pixelVal_in_1_4;
      end else if (10'h1b5 == _T_25[9:0]) begin
        image_1_437 <= io_pixelVal_in_1_3;
      end else if (10'h1b5 == _T_22[9:0]) begin
        image_1_437 <= io_pixelVal_in_1_2;
      end else if (10'h1b5 == _T_19[9:0]) begin
        image_1_437 <= io_pixelVal_in_1_1;
      end else if (10'h1b5 == _T_15[9:0]) begin
        image_1_437 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_438 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b6 == _T_37[9:0]) begin
        image_1_438 <= io_pixelVal_in_1_7;
      end else if (10'h1b6 == _T_34[9:0]) begin
        image_1_438 <= io_pixelVal_in_1_6;
      end else if (10'h1b6 == _T_31[9:0]) begin
        image_1_438 <= io_pixelVal_in_1_5;
      end else if (10'h1b6 == _T_28[9:0]) begin
        image_1_438 <= io_pixelVal_in_1_4;
      end else if (10'h1b6 == _T_25[9:0]) begin
        image_1_438 <= io_pixelVal_in_1_3;
      end else if (10'h1b6 == _T_22[9:0]) begin
        image_1_438 <= io_pixelVal_in_1_2;
      end else if (10'h1b6 == _T_19[9:0]) begin
        image_1_438 <= io_pixelVal_in_1_1;
      end else if (10'h1b6 == _T_15[9:0]) begin
        image_1_438 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_439 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b7 == _T_37[9:0]) begin
        image_1_439 <= io_pixelVal_in_1_7;
      end else if (10'h1b7 == _T_34[9:0]) begin
        image_1_439 <= io_pixelVal_in_1_6;
      end else if (10'h1b7 == _T_31[9:0]) begin
        image_1_439 <= io_pixelVal_in_1_5;
      end else if (10'h1b7 == _T_28[9:0]) begin
        image_1_439 <= io_pixelVal_in_1_4;
      end else if (10'h1b7 == _T_25[9:0]) begin
        image_1_439 <= io_pixelVal_in_1_3;
      end else if (10'h1b7 == _T_22[9:0]) begin
        image_1_439 <= io_pixelVal_in_1_2;
      end else if (10'h1b7 == _T_19[9:0]) begin
        image_1_439 <= io_pixelVal_in_1_1;
      end else if (10'h1b7 == _T_15[9:0]) begin
        image_1_439 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_440 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b8 == _T_37[9:0]) begin
        image_1_440 <= io_pixelVal_in_1_7;
      end else if (10'h1b8 == _T_34[9:0]) begin
        image_1_440 <= io_pixelVal_in_1_6;
      end else if (10'h1b8 == _T_31[9:0]) begin
        image_1_440 <= io_pixelVal_in_1_5;
      end else if (10'h1b8 == _T_28[9:0]) begin
        image_1_440 <= io_pixelVal_in_1_4;
      end else if (10'h1b8 == _T_25[9:0]) begin
        image_1_440 <= io_pixelVal_in_1_3;
      end else if (10'h1b8 == _T_22[9:0]) begin
        image_1_440 <= io_pixelVal_in_1_2;
      end else if (10'h1b8 == _T_19[9:0]) begin
        image_1_440 <= io_pixelVal_in_1_1;
      end else if (10'h1b8 == _T_15[9:0]) begin
        image_1_440 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_441 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b9 == _T_37[9:0]) begin
        image_1_441 <= io_pixelVal_in_1_7;
      end else if (10'h1b9 == _T_34[9:0]) begin
        image_1_441 <= io_pixelVal_in_1_6;
      end else if (10'h1b9 == _T_31[9:0]) begin
        image_1_441 <= io_pixelVal_in_1_5;
      end else if (10'h1b9 == _T_28[9:0]) begin
        image_1_441 <= io_pixelVal_in_1_4;
      end else if (10'h1b9 == _T_25[9:0]) begin
        image_1_441 <= io_pixelVal_in_1_3;
      end else if (10'h1b9 == _T_22[9:0]) begin
        image_1_441 <= io_pixelVal_in_1_2;
      end else if (10'h1b9 == _T_19[9:0]) begin
        image_1_441 <= io_pixelVal_in_1_1;
      end else if (10'h1b9 == _T_15[9:0]) begin
        image_1_441 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_442 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ba == _T_37[9:0]) begin
        image_1_442 <= io_pixelVal_in_1_7;
      end else if (10'h1ba == _T_34[9:0]) begin
        image_1_442 <= io_pixelVal_in_1_6;
      end else if (10'h1ba == _T_31[9:0]) begin
        image_1_442 <= io_pixelVal_in_1_5;
      end else if (10'h1ba == _T_28[9:0]) begin
        image_1_442 <= io_pixelVal_in_1_4;
      end else if (10'h1ba == _T_25[9:0]) begin
        image_1_442 <= io_pixelVal_in_1_3;
      end else if (10'h1ba == _T_22[9:0]) begin
        image_1_442 <= io_pixelVal_in_1_2;
      end else if (10'h1ba == _T_19[9:0]) begin
        image_1_442 <= io_pixelVal_in_1_1;
      end else if (10'h1ba == _T_15[9:0]) begin
        image_1_442 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_443 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1bb == _T_37[9:0]) begin
        image_1_443 <= io_pixelVal_in_1_7;
      end else if (10'h1bb == _T_34[9:0]) begin
        image_1_443 <= io_pixelVal_in_1_6;
      end else if (10'h1bb == _T_31[9:0]) begin
        image_1_443 <= io_pixelVal_in_1_5;
      end else if (10'h1bb == _T_28[9:0]) begin
        image_1_443 <= io_pixelVal_in_1_4;
      end else if (10'h1bb == _T_25[9:0]) begin
        image_1_443 <= io_pixelVal_in_1_3;
      end else if (10'h1bb == _T_22[9:0]) begin
        image_1_443 <= io_pixelVal_in_1_2;
      end else if (10'h1bb == _T_19[9:0]) begin
        image_1_443 <= io_pixelVal_in_1_1;
      end else if (10'h1bb == _T_15[9:0]) begin
        image_1_443 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_444 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1bc == _T_37[9:0]) begin
        image_1_444 <= io_pixelVal_in_1_7;
      end else if (10'h1bc == _T_34[9:0]) begin
        image_1_444 <= io_pixelVal_in_1_6;
      end else if (10'h1bc == _T_31[9:0]) begin
        image_1_444 <= io_pixelVal_in_1_5;
      end else if (10'h1bc == _T_28[9:0]) begin
        image_1_444 <= io_pixelVal_in_1_4;
      end else if (10'h1bc == _T_25[9:0]) begin
        image_1_444 <= io_pixelVal_in_1_3;
      end else if (10'h1bc == _T_22[9:0]) begin
        image_1_444 <= io_pixelVal_in_1_2;
      end else if (10'h1bc == _T_19[9:0]) begin
        image_1_444 <= io_pixelVal_in_1_1;
      end else if (10'h1bc == _T_15[9:0]) begin
        image_1_444 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_445 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1bd == _T_37[9:0]) begin
        image_1_445 <= io_pixelVal_in_1_7;
      end else if (10'h1bd == _T_34[9:0]) begin
        image_1_445 <= io_pixelVal_in_1_6;
      end else if (10'h1bd == _T_31[9:0]) begin
        image_1_445 <= io_pixelVal_in_1_5;
      end else if (10'h1bd == _T_28[9:0]) begin
        image_1_445 <= io_pixelVal_in_1_4;
      end else if (10'h1bd == _T_25[9:0]) begin
        image_1_445 <= io_pixelVal_in_1_3;
      end else if (10'h1bd == _T_22[9:0]) begin
        image_1_445 <= io_pixelVal_in_1_2;
      end else if (10'h1bd == _T_19[9:0]) begin
        image_1_445 <= io_pixelVal_in_1_1;
      end else if (10'h1bd == _T_15[9:0]) begin
        image_1_445 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_446 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1be == _T_37[9:0]) begin
        image_1_446 <= io_pixelVal_in_1_7;
      end else if (10'h1be == _T_34[9:0]) begin
        image_1_446 <= io_pixelVal_in_1_6;
      end else if (10'h1be == _T_31[9:0]) begin
        image_1_446 <= io_pixelVal_in_1_5;
      end else if (10'h1be == _T_28[9:0]) begin
        image_1_446 <= io_pixelVal_in_1_4;
      end else if (10'h1be == _T_25[9:0]) begin
        image_1_446 <= io_pixelVal_in_1_3;
      end else if (10'h1be == _T_22[9:0]) begin
        image_1_446 <= io_pixelVal_in_1_2;
      end else if (10'h1be == _T_19[9:0]) begin
        image_1_446 <= io_pixelVal_in_1_1;
      end else if (10'h1be == _T_15[9:0]) begin
        image_1_446 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_447 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1bf == _T_37[9:0]) begin
        image_1_447 <= io_pixelVal_in_1_7;
      end else if (10'h1bf == _T_34[9:0]) begin
        image_1_447 <= io_pixelVal_in_1_6;
      end else if (10'h1bf == _T_31[9:0]) begin
        image_1_447 <= io_pixelVal_in_1_5;
      end else if (10'h1bf == _T_28[9:0]) begin
        image_1_447 <= io_pixelVal_in_1_4;
      end else if (10'h1bf == _T_25[9:0]) begin
        image_1_447 <= io_pixelVal_in_1_3;
      end else if (10'h1bf == _T_22[9:0]) begin
        image_1_447 <= io_pixelVal_in_1_2;
      end else if (10'h1bf == _T_19[9:0]) begin
        image_1_447 <= io_pixelVal_in_1_1;
      end else if (10'h1bf == _T_15[9:0]) begin
        image_1_447 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_448 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c0 == _T_37[9:0]) begin
        image_1_448 <= io_pixelVal_in_1_7;
      end else if (10'h1c0 == _T_34[9:0]) begin
        image_1_448 <= io_pixelVal_in_1_6;
      end else if (10'h1c0 == _T_31[9:0]) begin
        image_1_448 <= io_pixelVal_in_1_5;
      end else if (10'h1c0 == _T_28[9:0]) begin
        image_1_448 <= io_pixelVal_in_1_4;
      end else if (10'h1c0 == _T_25[9:0]) begin
        image_1_448 <= io_pixelVal_in_1_3;
      end else if (10'h1c0 == _T_22[9:0]) begin
        image_1_448 <= io_pixelVal_in_1_2;
      end else if (10'h1c0 == _T_19[9:0]) begin
        image_1_448 <= io_pixelVal_in_1_1;
      end else if (10'h1c0 == _T_15[9:0]) begin
        image_1_448 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_449 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c1 == _T_37[9:0]) begin
        image_1_449 <= io_pixelVal_in_1_7;
      end else if (10'h1c1 == _T_34[9:0]) begin
        image_1_449 <= io_pixelVal_in_1_6;
      end else if (10'h1c1 == _T_31[9:0]) begin
        image_1_449 <= io_pixelVal_in_1_5;
      end else if (10'h1c1 == _T_28[9:0]) begin
        image_1_449 <= io_pixelVal_in_1_4;
      end else if (10'h1c1 == _T_25[9:0]) begin
        image_1_449 <= io_pixelVal_in_1_3;
      end else if (10'h1c1 == _T_22[9:0]) begin
        image_1_449 <= io_pixelVal_in_1_2;
      end else if (10'h1c1 == _T_19[9:0]) begin
        image_1_449 <= io_pixelVal_in_1_1;
      end else if (10'h1c1 == _T_15[9:0]) begin
        image_1_449 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_450 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c2 == _T_37[9:0]) begin
        image_1_450 <= io_pixelVal_in_1_7;
      end else if (10'h1c2 == _T_34[9:0]) begin
        image_1_450 <= io_pixelVal_in_1_6;
      end else if (10'h1c2 == _T_31[9:0]) begin
        image_1_450 <= io_pixelVal_in_1_5;
      end else if (10'h1c2 == _T_28[9:0]) begin
        image_1_450 <= io_pixelVal_in_1_4;
      end else if (10'h1c2 == _T_25[9:0]) begin
        image_1_450 <= io_pixelVal_in_1_3;
      end else if (10'h1c2 == _T_22[9:0]) begin
        image_1_450 <= io_pixelVal_in_1_2;
      end else if (10'h1c2 == _T_19[9:0]) begin
        image_1_450 <= io_pixelVal_in_1_1;
      end else if (10'h1c2 == _T_15[9:0]) begin
        image_1_450 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_451 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c3 == _T_37[9:0]) begin
        image_1_451 <= io_pixelVal_in_1_7;
      end else if (10'h1c3 == _T_34[9:0]) begin
        image_1_451 <= io_pixelVal_in_1_6;
      end else if (10'h1c3 == _T_31[9:0]) begin
        image_1_451 <= io_pixelVal_in_1_5;
      end else if (10'h1c3 == _T_28[9:0]) begin
        image_1_451 <= io_pixelVal_in_1_4;
      end else if (10'h1c3 == _T_25[9:0]) begin
        image_1_451 <= io_pixelVal_in_1_3;
      end else if (10'h1c3 == _T_22[9:0]) begin
        image_1_451 <= io_pixelVal_in_1_2;
      end else if (10'h1c3 == _T_19[9:0]) begin
        image_1_451 <= io_pixelVal_in_1_1;
      end else if (10'h1c3 == _T_15[9:0]) begin
        image_1_451 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_452 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c4 == _T_37[9:0]) begin
        image_1_452 <= io_pixelVal_in_1_7;
      end else if (10'h1c4 == _T_34[9:0]) begin
        image_1_452 <= io_pixelVal_in_1_6;
      end else if (10'h1c4 == _T_31[9:0]) begin
        image_1_452 <= io_pixelVal_in_1_5;
      end else if (10'h1c4 == _T_28[9:0]) begin
        image_1_452 <= io_pixelVal_in_1_4;
      end else if (10'h1c4 == _T_25[9:0]) begin
        image_1_452 <= io_pixelVal_in_1_3;
      end else if (10'h1c4 == _T_22[9:0]) begin
        image_1_452 <= io_pixelVal_in_1_2;
      end else if (10'h1c4 == _T_19[9:0]) begin
        image_1_452 <= io_pixelVal_in_1_1;
      end else if (10'h1c4 == _T_15[9:0]) begin
        image_1_452 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_453 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c5 == _T_37[9:0]) begin
        image_1_453 <= io_pixelVal_in_1_7;
      end else if (10'h1c5 == _T_34[9:0]) begin
        image_1_453 <= io_pixelVal_in_1_6;
      end else if (10'h1c5 == _T_31[9:0]) begin
        image_1_453 <= io_pixelVal_in_1_5;
      end else if (10'h1c5 == _T_28[9:0]) begin
        image_1_453 <= io_pixelVal_in_1_4;
      end else if (10'h1c5 == _T_25[9:0]) begin
        image_1_453 <= io_pixelVal_in_1_3;
      end else if (10'h1c5 == _T_22[9:0]) begin
        image_1_453 <= io_pixelVal_in_1_2;
      end else if (10'h1c5 == _T_19[9:0]) begin
        image_1_453 <= io_pixelVal_in_1_1;
      end else if (10'h1c5 == _T_15[9:0]) begin
        image_1_453 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_454 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c6 == _T_37[9:0]) begin
        image_1_454 <= io_pixelVal_in_1_7;
      end else if (10'h1c6 == _T_34[9:0]) begin
        image_1_454 <= io_pixelVal_in_1_6;
      end else if (10'h1c6 == _T_31[9:0]) begin
        image_1_454 <= io_pixelVal_in_1_5;
      end else if (10'h1c6 == _T_28[9:0]) begin
        image_1_454 <= io_pixelVal_in_1_4;
      end else if (10'h1c6 == _T_25[9:0]) begin
        image_1_454 <= io_pixelVal_in_1_3;
      end else if (10'h1c6 == _T_22[9:0]) begin
        image_1_454 <= io_pixelVal_in_1_2;
      end else if (10'h1c6 == _T_19[9:0]) begin
        image_1_454 <= io_pixelVal_in_1_1;
      end else if (10'h1c6 == _T_15[9:0]) begin
        image_1_454 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_455 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c7 == _T_37[9:0]) begin
        image_1_455 <= io_pixelVal_in_1_7;
      end else if (10'h1c7 == _T_34[9:0]) begin
        image_1_455 <= io_pixelVal_in_1_6;
      end else if (10'h1c7 == _T_31[9:0]) begin
        image_1_455 <= io_pixelVal_in_1_5;
      end else if (10'h1c7 == _T_28[9:0]) begin
        image_1_455 <= io_pixelVal_in_1_4;
      end else if (10'h1c7 == _T_25[9:0]) begin
        image_1_455 <= io_pixelVal_in_1_3;
      end else if (10'h1c7 == _T_22[9:0]) begin
        image_1_455 <= io_pixelVal_in_1_2;
      end else if (10'h1c7 == _T_19[9:0]) begin
        image_1_455 <= io_pixelVal_in_1_1;
      end else if (10'h1c7 == _T_15[9:0]) begin
        image_1_455 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_456 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c8 == _T_37[9:0]) begin
        image_1_456 <= io_pixelVal_in_1_7;
      end else if (10'h1c8 == _T_34[9:0]) begin
        image_1_456 <= io_pixelVal_in_1_6;
      end else if (10'h1c8 == _T_31[9:0]) begin
        image_1_456 <= io_pixelVal_in_1_5;
      end else if (10'h1c8 == _T_28[9:0]) begin
        image_1_456 <= io_pixelVal_in_1_4;
      end else if (10'h1c8 == _T_25[9:0]) begin
        image_1_456 <= io_pixelVal_in_1_3;
      end else if (10'h1c8 == _T_22[9:0]) begin
        image_1_456 <= io_pixelVal_in_1_2;
      end else if (10'h1c8 == _T_19[9:0]) begin
        image_1_456 <= io_pixelVal_in_1_1;
      end else if (10'h1c8 == _T_15[9:0]) begin
        image_1_456 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_457 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c9 == _T_37[9:0]) begin
        image_1_457 <= io_pixelVal_in_1_7;
      end else if (10'h1c9 == _T_34[9:0]) begin
        image_1_457 <= io_pixelVal_in_1_6;
      end else if (10'h1c9 == _T_31[9:0]) begin
        image_1_457 <= io_pixelVal_in_1_5;
      end else if (10'h1c9 == _T_28[9:0]) begin
        image_1_457 <= io_pixelVal_in_1_4;
      end else if (10'h1c9 == _T_25[9:0]) begin
        image_1_457 <= io_pixelVal_in_1_3;
      end else if (10'h1c9 == _T_22[9:0]) begin
        image_1_457 <= io_pixelVal_in_1_2;
      end else if (10'h1c9 == _T_19[9:0]) begin
        image_1_457 <= io_pixelVal_in_1_1;
      end else if (10'h1c9 == _T_15[9:0]) begin
        image_1_457 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_458 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ca == _T_37[9:0]) begin
        image_1_458 <= io_pixelVal_in_1_7;
      end else if (10'h1ca == _T_34[9:0]) begin
        image_1_458 <= io_pixelVal_in_1_6;
      end else if (10'h1ca == _T_31[9:0]) begin
        image_1_458 <= io_pixelVal_in_1_5;
      end else if (10'h1ca == _T_28[9:0]) begin
        image_1_458 <= io_pixelVal_in_1_4;
      end else if (10'h1ca == _T_25[9:0]) begin
        image_1_458 <= io_pixelVal_in_1_3;
      end else if (10'h1ca == _T_22[9:0]) begin
        image_1_458 <= io_pixelVal_in_1_2;
      end else if (10'h1ca == _T_19[9:0]) begin
        image_1_458 <= io_pixelVal_in_1_1;
      end else if (10'h1ca == _T_15[9:0]) begin
        image_1_458 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_459 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1cb == _T_37[9:0]) begin
        image_1_459 <= io_pixelVal_in_1_7;
      end else if (10'h1cb == _T_34[9:0]) begin
        image_1_459 <= io_pixelVal_in_1_6;
      end else if (10'h1cb == _T_31[9:0]) begin
        image_1_459 <= io_pixelVal_in_1_5;
      end else if (10'h1cb == _T_28[9:0]) begin
        image_1_459 <= io_pixelVal_in_1_4;
      end else if (10'h1cb == _T_25[9:0]) begin
        image_1_459 <= io_pixelVal_in_1_3;
      end else if (10'h1cb == _T_22[9:0]) begin
        image_1_459 <= io_pixelVal_in_1_2;
      end else if (10'h1cb == _T_19[9:0]) begin
        image_1_459 <= io_pixelVal_in_1_1;
      end else if (10'h1cb == _T_15[9:0]) begin
        image_1_459 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_460 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1cc == _T_37[9:0]) begin
        image_1_460 <= io_pixelVal_in_1_7;
      end else if (10'h1cc == _T_34[9:0]) begin
        image_1_460 <= io_pixelVal_in_1_6;
      end else if (10'h1cc == _T_31[9:0]) begin
        image_1_460 <= io_pixelVal_in_1_5;
      end else if (10'h1cc == _T_28[9:0]) begin
        image_1_460 <= io_pixelVal_in_1_4;
      end else if (10'h1cc == _T_25[9:0]) begin
        image_1_460 <= io_pixelVal_in_1_3;
      end else if (10'h1cc == _T_22[9:0]) begin
        image_1_460 <= io_pixelVal_in_1_2;
      end else if (10'h1cc == _T_19[9:0]) begin
        image_1_460 <= io_pixelVal_in_1_1;
      end else if (10'h1cc == _T_15[9:0]) begin
        image_1_460 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_461 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1cd == _T_37[9:0]) begin
        image_1_461 <= io_pixelVal_in_1_7;
      end else if (10'h1cd == _T_34[9:0]) begin
        image_1_461 <= io_pixelVal_in_1_6;
      end else if (10'h1cd == _T_31[9:0]) begin
        image_1_461 <= io_pixelVal_in_1_5;
      end else if (10'h1cd == _T_28[9:0]) begin
        image_1_461 <= io_pixelVal_in_1_4;
      end else if (10'h1cd == _T_25[9:0]) begin
        image_1_461 <= io_pixelVal_in_1_3;
      end else if (10'h1cd == _T_22[9:0]) begin
        image_1_461 <= io_pixelVal_in_1_2;
      end else if (10'h1cd == _T_19[9:0]) begin
        image_1_461 <= io_pixelVal_in_1_1;
      end else if (10'h1cd == _T_15[9:0]) begin
        image_1_461 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_462 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ce == _T_37[9:0]) begin
        image_1_462 <= io_pixelVal_in_1_7;
      end else if (10'h1ce == _T_34[9:0]) begin
        image_1_462 <= io_pixelVal_in_1_6;
      end else if (10'h1ce == _T_31[9:0]) begin
        image_1_462 <= io_pixelVal_in_1_5;
      end else if (10'h1ce == _T_28[9:0]) begin
        image_1_462 <= io_pixelVal_in_1_4;
      end else if (10'h1ce == _T_25[9:0]) begin
        image_1_462 <= io_pixelVal_in_1_3;
      end else if (10'h1ce == _T_22[9:0]) begin
        image_1_462 <= io_pixelVal_in_1_2;
      end else if (10'h1ce == _T_19[9:0]) begin
        image_1_462 <= io_pixelVal_in_1_1;
      end else if (10'h1ce == _T_15[9:0]) begin
        image_1_462 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_463 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1cf == _T_37[9:0]) begin
        image_1_463 <= io_pixelVal_in_1_7;
      end else if (10'h1cf == _T_34[9:0]) begin
        image_1_463 <= io_pixelVal_in_1_6;
      end else if (10'h1cf == _T_31[9:0]) begin
        image_1_463 <= io_pixelVal_in_1_5;
      end else if (10'h1cf == _T_28[9:0]) begin
        image_1_463 <= io_pixelVal_in_1_4;
      end else if (10'h1cf == _T_25[9:0]) begin
        image_1_463 <= io_pixelVal_in_1_3;
      end else if (10'h1cf == _T_22[9:0]) begin
        image_1_463 <= io_pixelVal_in_1_2;
      end else if (10'h1cf == _T_19[9:0]) begin
        image_1_463 <= io_pixelVal_in_1_1;
      end else if (10'h1cf == _T_15[9:0]) begin
        image_1_463 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_464 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d0 == _T_37[9:0]) begin
        image_1_464 <= io_pixelVal_in_1_7;
      end else if (10'h1d0 == _T_34[9:0]) begin
        image_1_464 <= io_pixelVal_in_1_6;
      end else if (10'h1d0 == _T_31[9:0]) begin
        image_1_464 <= io_pixelVal_in_1_5;
      end else if (10'h1d0 == _T_28[9:0]) begin
        image_1_464 <= io_pixelVal_in_1_4;
      end else if (10'h1d0 == _T_25[9:0]) begin
        image_1_464 <= io_pixelVal_in_1_3;
      end else if (10'h1d0 == _T_22[9:0]) begin
        image_1_464 <= io_pixelVal_in_1_2;
      end else if (10'h1d0 == _T_19[9:0]) begin
        image_1_464 <= io_pixelVal_in_1_1;
      end else if (10'h1d0 == _T_15[9:0]) begin
        image_1_464 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_465 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d1 == _T_37[9:0]) begin
        image_1_465 <= io_pixelVal_in_1_7;
      end else if (10'h1d1 == _T_34[9:0]) begin
        image_1_465 <= io_pixelVal_in_1_6;
      end else if (10'h1d1 == _T_31[9:0]) begin
        image_1_465 <= io_pixelVal_in_1_5;
      end else if (10'h1d1 == _T_28[9:0]) begin
        image_1_465 <= io_pixelVal_in_1_4;
      end else if (10'h1d1 == _T_25[9:0]) begin
        image_1_465 <= io_pixelVal_in_1_3;
      end else if (10'h1d1 == _T_22[9:0]) begin
        image_1_465 <= io_pixelVal_in_1_2;
      end else if (10'h1d1 == _T_19[9:0]) begin
        image_1_465 <= io_pixelVal_in_1_1;
      end else if (10'h1d1 == _T_15[9:0]) begin
        image_1_465 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_466 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d2 == _T_37[9:0]) begin
        image_1_466 <= io_pixelVal_in_1_7;
      end else if (10'h1d2 == _T_34[9:0]) begin
        image_1_466 <= io_pixelVal_in_1_6;
      end else if (10'h1d2 == _T_31[9:0]) begin
        image_1_466 <= io_pixelVal_in_1_5;
      end else if (10'h1d2 == _T_28[9:0]) begin
        image_1_466 <= io_pixelVal_in_1_4;
      end else if (10'h1d2 == _T_25[9:0]) begin
        image_1_466 <= io_pixelVal_in_1_3;
      end else if (10'h1d2 == _T_22[9:0]) begin
        image_1_466 <= io_pixelVal_in_1_2;
      end else if (10'h1d2 == _T_19[9:0]) begin
        image_1_466 <= io_pixelVal_in_1_1;
      end else if (10'h1d2 == _T_15[9:0]) begin
        image_1_466 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_467 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d3 == _T_37[9:0]) begin
        image_1_467 <= io_pixelVal_in_1_7;
      end else if (10'h1d3 == _T_34[9:0]) begin
        image_1_467 <= io_pixelVal_in_1_6;
      end else if (10'h1d3 == _T_31[9:0]) begin
        image_1_467 <= io_pixelVal_in_1_5;
      end else if (10'h1d3 == _T_28[9:0]) begin
        image_1_467 <= io_pixelVal_in_1_4;
      end else if (10'h1d3 == _T_25[9:0]) begin
        image_1_467 <= io_pixelVal_in_1_3;
      end else if (10'h1d3 == _T_22[9:0]) begin
        image_1_467 <= io_pixelVal_in_1_2;
      end else if (10'h1d3 == _T_19[9:0]) begin
        image_1_467 <= io_pixelVal_in_1_1;
      end else if (10'h1d3 == _T_15[9:0]) begin
        image_1_467 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_468 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d4 == _T_37[9:0]) begin
        image_1_468 <= io_pixelVal_in_1_7;
      end else if (10'h1d4 == _T_34[9:0]) begin
        image_1_468 <= io_pixelVal_in_1_6;
      end else if (10'h1d4 == _T_31[9:0]) begin
        image_1_468 <= io_pixelVal_in_1_5;
      end else if (10'h1d4 == _T_28[9:0]) begin
        image_1_468 <= io_pixelVal_in_1_4;
      end else if (10'h1d4 == _T_25[9:0]) begin
        image_1_468 <= io_pixelVal_in_1_3;
      end else if (10'h1d4 == _T_22[9:0]) begin
        image_1_468 <= io_pixelVal_in_1_2;
      end else if (10'h1d4 == _T_19[9:0]) begin
        image_1_468 <= io_pixelVal_in_1_1;
      end else if (10'h1d4 == _T_15[9:0]) begin
        image_1_468 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_469 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d5 == _T_37[9:0]) begin
        image_1_469 <= io_pixelVal_in_1_7;
      end else if (10'h1d5 == _T_34[9:0]) begin
        image_1_469 <= io_pixelVal_in_1_6;
      end else if (10'h1d5 == _T_31[9:0]) begin
        image_1_469 <= io_pixelVal_in_1_5;
      end else if (10'h1d5 == _T_28[9:0]) begin
        image_1_469 <= io_pixelVal_in_1_4;
      end else if (10'h1d5 == _T_25[9:0]) begin
        image_1_469 <= io_pixelVal_in_1_3;
      end else if (10'h1d5 == _T_22[9:0]) begin
        image_1_469 <= io_pixelVal_in_1_2;
      end else if (10'h1d5 == _T_19[9:0]) begin
        image_1_469 <= io_pixelVal_in_1_1;
      end else if (10'h1d5 == _T_15[9:0]) begin
        image_1_469 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_470 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d6 == _T_37[9:0]) begin
        image_1_470 <= io_pixelVal_in_1_7;
      end else if (10'h1d6 == _T_34[9:0]) begin
        image_1_470 <= io_pixelVal_in_1_6;
      end else if (10'h1d6 == _T_31[9:0]) begin
        image_1_470 <= io_pixelVal_in_1_5;
      end else if (10'h1d6 == _T_28[9:0]) begin
        image_1_470 <= io_pixelVal_in_1_4;
      end else if (10'h1d6 == _T_25[9:0]) begin
        image_1_470 <= io_pixelVal_in_1_3;
      end else if (10'h1d6 == _T_22[9:0]) begin
        image_1_470 <= io_pixelVal_in_1_2;
      end else if (10'h1d6 == _T_19[9:0]) begin
        image_1_470 <= io_pixelVal_in_1_1;
      end else if (10'h1d6 == _T_15[9:0]) begin
        image_1_470 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_471 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d7 == _T_37[9:0]) begin
        image_1_471 <= io_pixelVal_in_1_7;
      end else if (10'h1d7 == _T_34[9:0]) begin
        image_1_471 <= io_pixelVal_in_1_6;
      end else if (10'h1d7 == _T_31[9:0]) begin
        image_1_471 <= io_pixelVal_in_1_5;
      end else if (10'h1d7 == _T_28[9:0]) begin
        image_1_471 <= io_pixelVal_in_1_4;
      end else if (10'h1d7 == _T_25[9:0]) begin
        image_1_471 <= io_pixelVal_in_1_3;
      end else if (10'h1d7 == _T_22[9:0]) begin
        image_1_471 <= io_pixelVal_in_1_2;
      end else if (10'h1d7 == _T_19[9:0]) begin
        image_1_471 <= io_pixelVal_in_1_1;
      end else if (10'h1d7 == _T_15[9:0]) begin
        image_1_471 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_472 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d8 == _T_37[9:0]) begin
        image_1_472 <= io_pixelVal_in_1_7;
      end else if (10'h1d8 == _T_34[9:0]) begin
        image_1_472 <= io_pixelVal_in_1_6;
      end else if (10'h1d8 == _T_31[9:0]) begin
        image_1_472 <= io_pixelVal_in_1_5;
      end else if (10'h1d8 == _T_28[9:0]) begin
        image_1_472 <= io_pixelVal_in_1_4;
      end else if (10'h1d8 == _T_25[9:0]) begin
        image_1_472 <= io_pixelVal_in_1_3;
      end else if (10'h1d8 == _T_22[9:0]) begin
        image_1_472 <= io_pixelVal_in_1_2;
      end else if (10'h1d8 == _T_19[9:0]) begin
        image_1_472 <= io_pixelVal_in_1_1;
      end else if (10'h1d8 == _T_15[9:0]) begin
        image_1_472 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_473 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d9 == _T_37[9:0]) begin
        image_1_473 <= io_pixelVal_in_1_7;
      end else if (10'h1d9 == _T_34[9:0]) begin
        image_1_473 <= io_pixelVal_in_1_6;
      end else if (10'h1d9 == _T_31[9:0]) begin
        image_1_473 <= io_pixelVal_in_1_5;
      end else if (10'h1d9 == _T_28[9:0]) begin
        image_1_473 <= io_pixelVal_in_1_4;
      end else if (10'h1d9 == _T_25[9:0]) begin
        image_1_473 <= io_pixelVal_in_1_3;
      end else if (10'h1d9 == _T_22[9:0]) begin
        image_1_473 <= io_pixelVal_in_1_2;
      end else if (10'h1d9 == _T_19[9:0]) begin
        image_1_473 <= io_pixelVal_in_1_1;
      end else if (10'h1d9 == _T_15[9:0]) begin
        image_1_473 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_474 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1da == _T_37[9:0]) begin
        image_1_474 <= io_pixelVal_in_1_7;
      end else if (10'h1da == _T_34[9:0]) begin
        image_1_474 <= io_pixelVal_in_1_6;
      end else if (10'h1da == _T_31[9:0]) begin
        image_1_474 <= io_pixelVal_in_1_5;
      end else if (10'h1da == _T_28[9:0]) begin
        image_1_474 <= io_pixelVal_in_1_4;
      end else if (10'h1da == _T_25[9:0]) begin
        image_1_474 <= io_pixelVal_in_1_3;
      end else if (10'h1da == _T_22[9:0]) begin
        image_1_474 <= io_pixelVal_in_1_2;
      end else if (10'h1da == _T_19[9:0]) begin
        image_1_474 <= io_pixelVal_in_1_1;
      end else if (10'h1da == _T_15[9:0]) begin
        image_1_474 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_475 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1db == _T_37[9:0]) begin
        image_1_475 <= io_pixelVal_in_1_7;
      end else if (10'h1db == _T_34[9:0]) begin
        image_1_475 <= io_pixelVal_in_1_6;
      end else if (10'h1db == _T_31[9:0]) begin
        image_1_475 <= io_pixelVal_in_1_5;
      end else if (10'h1db == _T_28[9:0]) begin
        image_1_475 <= io_pixelVal_in_1_4;
      end else if (10'h1db == _T_25[9:0]) begin
        image_1_475 <= io_pixelVal_in_1_3;
      end else if (10'h1db == _T_22[9:0]) begin
        image_1_475 <= io_pixelVal_in_1_2;
      end else if (10'h1db == _T_19[9:0]) begin
        image_1_475 <= io_pixelVal_in_1_1;
      end else if (10'h1db == _T_15[9:0]) begin
        image_1_475 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_476 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1dc == _T_37[9:0]) begin
        image_1_476 <= io_pixelVal_in_1_7;
      end else if (10'h1dc == _T_34[9:0]) begin
        image_1_476 <= io_pixelVal_in_1_6;
      end else if (10'h1dc == _T_31[9:0]) begin
        image_1_476 <= io_pixelVal_in_1_5;
      end else if (10'h1dc == _T_28[9:0]) begin
        image_1_476 <= io_pixelVal_in_1_4;
      end else if (10'h1dc == _T_25[9:0]) begin
        image_1_476 <= io_pixelVal_in_1_3;
      end else if (10'h1dc == _T_22[9:0]) begin
        image_1_476 <= io_pixelVal_in_1_2;
      end else if (10'h1dc == _T_19[9:0]) begin
        image_1_476 <= io_pixelVal_in_1_1;
      end else if (10'h1dc == _T_15[9:0]) begin
        image_1_476 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_477 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1dd == _T_37[9:0]) begin
        image_1_477 <= io_pixelVal_in_1_7;
      end else if (10'h1dd == _T_34[9:0]) begin
        image_1_477 <= io_pixelVal_in_1_6;
      end else if (10'h1dd == _T_31[9:0]) begin
        image_1_477 <= io_pixelVal_in_1_5;
      end else if (10'h1dd == _T_28[9:0]) begin
        image_1_477 <= io_pixelVal_in_1_4;
      end else if (10'h1dd == _T_25[9:0]) begin
        image_1_477 <= io_pixelVal_in_1_3;
      end else if (10'h1dd == _T_22[9:0]) begin
        image_1_477 <= io_pixelVal_in_1_2;
      end else if (10'h1dd == _T_19[9:0]) begin
        image_1_477 <= io_pixelVal_in_1_1;
      end else if (10'h1dd == _T_15[9:0]) begin
        image_1_477 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_478 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1de == _T_37[9:0]) begin
        image_1_478 <= io_pixelVal_in_1_7;
      end else if (10'h1de == _T_34[9:0]) begin
        image_1_478 <= io_pixelVal_in_1_6;
      end else if (10'h1de == _T_31[9:0]) begin
        image_1_478 <= io_pixelVal_in_1_5;
      end else if (10'h1de == _T_28[9:0]) begin
        image_1_478 <= io_pixelVal_in_1_4;
      end else if (10'h1de == _T_25[9:0]) begin
        image_1_478 <= io_pixelVal_in_1_3;
      end else if (10'h1de == _T_22[9:0]) begin
        image_1_478 <= io_pixelVal_in_1_2;
      end else if (10'h1de == _T_19[9:0]) begin
        image_1_478 <= io_pixelVal_in_1_1;
      end else if (10'h1de == _T_15[9:0]) begin
        image_1_478 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_479 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1df == _T_37[9:0]) begin
        image_1_479 <= io_pixelVal_in_1_7;
      end else if (10'h1df == _T_34[9:0]) begin
        image_1_479 <= io_pixelVal_in_1_6;
      end else if (10'h1df == _T_31[9:0]) begin
        image_1_479 <= io_pixelVal_in_1_5;
      end else if (10'h1df == _T_28[9:0]) begin
        image_1_479 <= io_pixelVal_in_1_4;
      end else if (10'h1df == _T_25[9:0]) begin
        image_1_479 <= io_pixelVal_in_1_3;
      end else if (10'h1df == _T_22[9:0]) begin
        image_1_479 <= io_pixelVal_in_1_2;
      end else if (10'h1df == _T_19[9:0]) begin
        image_1_479 <= io_pixelVal_in_1_1;
      end else if (10'h1df == _T_15[9:0]) begin
        image_1_479 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_480 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e0 == _T_37[9:0]) begin
        image_1_480 <= io_pixelVal_in_1_7;
      end else if (10'h1e0 == _T_34[9:0]) begin
        image_1_480 <= io_pixelVal_in_1_6;
      end else if (10'h1e0 == _T_31[9:0]) begin
        image_1_480 <= io_pixelVal_in_1_5;
      end else if (10'h1e0 == _T_28[9:0]) begin
        image_1_480 <= io_pixelVal_in_1_4;
      end else if (10'h1e0 == _T_25[9:0]) begin
        image_1_480 <= io_pixelVal_in_1_3;
      end else if (10'h1e0 == _T_22[9:0]) begin
        image_1_480 <= io_pixelVal_in_1_2;
      end else if (10'h1e0 == _T_19[9:0]) begin
        image_1_480 <= io_pixelVal_in_1_1;
      end else if (10'h1e0 == _T_15[9:0]) begin
        image_1_480 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_481 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e1 == _T_37[9:0]) begin
        image_1_481 <= io_pixelVal_in_1_7;
      end else if (10'h1e1 == _T_34[9:0]) begin
        image_1_481 <= io_pixelVal_in_1_6;
      end else if (10'h1e1 == _T_31[9:0]) begin
        image_1_481 <= io_pixelVal_in_1_5;
      end else if (10'h1e1 == _T_28[9:0]) begin
        image_1_481 <= io_pixelVal_in_1_4;
      end else if (10'h1e1 == _T_25[9:0]) begin
        image_1_481 <= io_pixelVal_in_1_3;
      end else if (10'h1e1 == _T_22[9:0]) begin
        image_1_481 <= io_pixelVal_in_1_2;
      end else if (10'h1e1 == _T_19[9:0]) begin
        image_1_481 <= io_pixelVal_in_1_1;
      end else if (10'h1e1 == _T_15[9:0]) begin
        image_1_481 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_482 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e2 == _T_37[9:0]) begin
        image_1_482 <= io_pixelVal_in_1_7;
      end else if (10'h1e2 == _T_34[9:0]) begin
        image_1_482 <= io_pixelVal_in_1_6;
      end else if (10'h1e2 == _T_31[9:0]) begin
        image_1_482 <= io_pixelVal_in_1_5;
      end else if (10'h1e2 == _T_28[9:0]) begin
        image_1_482 <= io_pixelVal_in_1_4;
      end else if (10'h1e2 == _T_25[9:0]) begin
        image_1_482 <= io_pixelVal_in_1_3;
      end else if (10'h1e2 == _T_22[9:0]) begin
        image_1_482 <= io_pixelVal_in_1_2;
      end else if (10'h1e2 == _T_19[9:0]) begin
        image_1_482 <= io_pixelVal_in_1_1;
      end else if (10'h1e2 == _T_15[9:0]) begin
        image_1_482 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_483 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e3 == _T_37[9:0]) begin
        image_1_483 <= io_pixelVal_in_1_7;
      end else if (10'h1e3 == _T_34[9:0]) begin
        image_1_483 <= io_pixelVal_in_1_6;
      end else if (10'h1e3 == _T_31[9:0]) begin
        image_1_483 <= io_pixelVal_in_1_5;
      end else if (10'h1e3 == _T_28[9:0]) begin
        image_1_483 <= io_pixelVal_in_1_4;
      end else if (10'h1e3 == _T_25[9:0]) begin
        image_1_483 <= io_pixelVal_in_1_3;
      end else if (10'h1e3 == _T_22[9:0]) begin
        image_1_483 <= io_pixelVal_in_1_2;
      end else if (10'h1e3 == _T_19[9:0]) begin
        image_1_483 <= io_pixelVal_in_1_1;
      end else if (10'h1e3 == _T_15[9:0]) begin
        image_1_483 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_484 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e4 == _T_37[9:0]) begin
        image_1_484 <= io_pixelVal_in_1_7;
      end else if (10'h1e4 == _T_34[9:0]) begin
        image_1_484 <= io_pixelVal_in_1_6;
      end else if (10'h1e4 == _T_31[9:0]) begin
        image_1_484 <= io_pixelVal_in_1_5;
      end else if (10'h1e4 == _T_28[9:0]) begin
        image_1_484 <= io_pixelVal_in_1_4;
      end else if (10'h1e4 == _T_25[9:0]) begin
        image_1_484 <= io_pixelVal_in_1_3;
      end else if (10'h1e4 == _T_22[9:0]) begin
        image_1_484 <= io_pixelVal_in_1_2;
      end else if (10'h1e4 == _T_19[9:0]) begin
        image_1_484 <= io_pixelVal_in_1_1;
      end else if (10'h1e4 == _T_15[9:0]) begin
        image_1_484 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_485 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e5 == _T_37[9:0]) begin
        image_1_485 <= io_pixelVal_in_1_7;
      end else if (10'h1e5 == _T_34[9:0]) begin
        image_1_485 <= io_pixelVal_in_1_6;
      end else if (10'h1e5 == _T_31[9:0]) begin
        image_1_485 <= io_pixelVal_in_1_5;
      end else if (10'h1e5 == _T_28[9:0]) begin
        image_1_485 <= io_pixelVal_in_1_4;
      end else if (10'h1e5 == _T_25[9:0]) begin
        image_1_485 <= io_pixelVal_in_1_3;
      end else if (10'h1e5 == _T_22[9:0]) begin
        image_1_485 <= io_pixelVal_in_1_2;
      end else if (10'h1e5 == _T_19[9:0]) begin
        image_1_485 <= io_pixelVal_in_1_1;
      end else if (10'h1e5 == _T_15[9:0]) begin
        image_1_485 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_486 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e6 == _T_37[9:0]) begin
        image_1_486 <= io_pixelVal_in_1_7;
      end else if (10'h1e6 == _T_34[9:0]) begin
        image_1_486 <= io_pixelVal_in_1_6;
      end else if (10'h1e6 == _T_31[9:0]) begin
        image_1_486 <= io_pixelVal_in_1_5;
      end else if (10'h1e6 == _T_28[9:0]) begin
        image_1_486 <= io_pixelVal_in_1_4;
      end else if (10'h1e6 == _T_25[9:0]) begin
        image_1_486 <= io_pixelVal_in_1_3;
      end else if (10'h1e6 == _T_22[9:0]) begin
        image_1_486 <= io_pixelVal_in_1_2;
      end else if (10'h1e6 == _T_19[9:0]) begin
        image_1_486 <= io_pixelVal_in_1_1;
      end else if (10'h1e6 == _T_15[9:0]) begin
        image_1_486 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_487 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e7 == _T_37[9:0]) begin
        image_1_487 <= io_pixelVal_in_1_7;
      end else if (10'h1e7 == _T_34[9:0]) begin
        image_1_487 <= io_pixelVal_in_1_6;
      end else if (10'h1e7 == _T_31[9:0]) begin
        image_1_487 <= io_pixelVal_in_1_5;
      end else if (10'h1e7 == _T_28[9:0]) begin
        image_1_487 <= io_pixelVal_in_1_4;
      end else if (10'h1e7 == _T_25[9:0]) begin
        image_1_487 <= io_pixelVal_in_1_3;
      end else if (10'h1e7 == _T_22[9:0]) begin
        image_1_487 <= io_pixelVal_in_1_2;
      end else if (10'h1e7 == _T_19[9:0]) begin
        image_1_487 <= io_pixelVal_in_1_1;
      end else if (10'h1e7 == _T_15[9:0]) begin
        image_1_487 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_488 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e8 == _T_37[9:0]) begin
        image_1_488 <= io_pixelVal_in_1_7;
      end else if (10'h1e8 == _T_34[9:0]) begin
        image_1_488 <= io_pixelVal_in_1_6;
      end else if (10'h1e8 == _T_31[9:0]) begin
        image_1_488 <= io_pixelVal_in_1_5;
      end else if (10'h1e8 == _T_28[9:0]) begin
        image_1_488 <= io_pixelVal_in_1_4;
      end else if (10'h1e8 == _T_25[9:0]) begin
        image_1_488 <= io_pixelVal_in_1_3;
      end else if (10'h1e8 == _T_22[9:0]) begin
        image_1_488 <= io_pixelVal_in_1_2;
      end else if (10'h1e8 == _T_19[9:0]) begin
        image_1_488 <= io_pixelVal_in_1_1;
      end else if (10'h1e8 == _T_15[9:0]) begin
        image_1_488 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_489 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e9 == _T_37[9:0]) begin
        image_1_489 <= io_pixelVal_in_1_7;
      end else if (10'h1e9 == _T_34[9:0]) begin
        image_1_489 <= io_pixelVal_in_1_6;
      end else if (10'h1e9 == _T_31[9:0]) begin
        image_1_489 <= io_pixelVal_in_1_5;
      end else if (10'h1e9 == _T_28[9:0]) begin
        image_1_489 <= io_pixelVal_in_1_4;
      end else if (10'h1e9 == _T_25[9:0]) begin
        image_1_489 <= io_pixelVal_in_1_3;
      end else if (10'h1e9 == _T_22[9:0]) begin
        image_1_489 <= io_pixelVal_in_1_2;
      end else if (10'h1e9 == _T_19[9:0]) begin
        image_1_489 <= io_pixelVal_in_1_1;
      end else if (10'h1e9 == _T_15[9:0]) begin
        image_1_489 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_490 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ea == _T_37[9:0]) begin
        image_1_490 <= io_pixelVal_in_1_7;
      end else if (10'h1ea == _T_34[9:0]) begin
        image_1_490 <= io_pixelVal_in_1_6;
      end else if (10'h1ea == _T_31[9:0]) begin
        image_1_490 <= io_pixelVal_in_1_5;
      end else if (10'h1ea == _T_28[9:0]) begin
        image_1_490 <= io_pixelVal_in_1_4;
      end else if (10'h1ea == _T_25[9:0]) begin
        image_1_490 <= io_pixelVal_in_1_3;
      end else if (10'h1ea == _T_22[9:0]) begin
        image_1_490 <= io_pixelVal_in_1_2;
      end else if (10'h1ea == _T_19[9:0]) begin
        image_1_490 <= io_pixelVal_in_1_1;
      end else if (10'h1ea == _T_15[9:0]) begin
        image_1_490 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_491 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1eb == _T_37[9:0]) begin
        image_1_491 <= io_pixelVal_in_1_7;
      end else if (10'h1eb == _T_34[9:0]) begin
        image_1_491 <= io_pixelVal_in_1_6;
      end else if (10'h1eb == _T_31[9:0]) begin
        image_1_491 <= io_pixelVal_in_1_5;
      end else if (10'h1eb == _T_28[9:0]) begin
        image_1_491 <= io_pixelVal_in_1_4;
      end else if (10'h1eb == _T_25[9:0]) begin
        image_1_491 <= io_pixelVal_in_1_3;
      end else if (10'h1eb == _T_22[9:0]) begin
        image_1_491 <= io_pixelVal_in_1_2;
      end else if (10'h1eb == _T_19[9:0]) begin
        image_1_491 <= io_pixelVal_in_1_1;
      end else if (10'h1eb == _T_15[9:0]) begin
        image_1_491 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_492 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ec == _T_37[9:0]) begin
        image_1_492 <= io_pixelVal_in_1_7;
      end else if (10'h1ec == _T_34[9:0]) begin
        image_1_492 <= io_pixelVal_in_1_6;
      end else if (10'h1ec == _T_31[9:0]) begin
        image_1_492 <= io_pixelVal_in_1_5;
      end else if (10'h1ec == _T_28[9:0]) begin
        image_1_492 <= io_pixelVal_in_1_4;
      end else if (10'h1ec == _T_25[9:0]) begin
        image_1_492 <= io_pixelVal_in_1_3;
      end else if (10'h1ec == _T_22[9:0]) begin
        image_1_492 <= io_pixelVal_in_1_2;
      end else if (10'h1ec == _T_19[9:0]) begin
        image_1_492 <= io_pixelVal_in_1_1;
      end else if (10'h1ec == _T_15[9:0]) begin
        image_1_492 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_493 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ed == _T_37[9:0]) begin
        image_1_493 <= io_pixelVal_in_1_7;
      end else if (10'h1ed == _T_34[9:0]) begin
        image_1_493 <= io_pixelVal_in_1_6;
      end else if (10'h1ed == _T_31[9:0]) begin
        image_1_493 <= io_pixelVal_in_1_5;
      end else if (10'h1ed == _T_28[9:0]) begin
        image_1_493 <= io_pixelVal_in_1_4;
      end else if (10'h1ed == _T_25[9:0]) begin
        image_1_493 <= io_pixelVal_in_1_3;
      end else if (10'h1ed == _T_22[9:0]) begin
        image_1_493 <= io_pixelVal_in_1_2;
      end else if (10'h1ed == _T_19[9:0]) begin
        image_1_493 <= io_pixelVal_in_1_1;
      end else if (10'h1ed == _T_15[9:0]) begin
        image_1_493 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_494 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ee == _T_37[9:0]) begin
        image_1_494 <= io_pixelVal_in_1_7;
      end else if (10'h1ee == _T_34[9:0]) begin
        image_1_494 <= io_pixelVal_in_1_6;
      end else if (10'h1ee == _T_31[9:0]) begin
        image_1_494 <= io_pixelVal_in_1_5;
      end else if (10'h1ee == _T_28[9:0]) begin
        image_1_494 <= io_pixelVal_in_1_4;
      end else if (10'h1ee == _T_25[9:0]) begin
        image_1_494 <= io_pixelVal_in_1_3;
      end else if (10'h1ee == _T_22[9:0]) begin
        image_1_494 <= io_pixelVal_in_1_2;
      end else if (10'h1ee == _T_19[9:0]) begin
        image_1_494 <= io_pixelVal_in_1_1;
      end else if (10'h1ee == _T_15[9:0]) begin
        image_1_494 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_495 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ef == _T_37[9:0]) begin
        image_1_495 <= io_pixelVal_in_1_7;
      end else if (10'h1ef == _T_34[9:0]) begin
        image_1_495 <= io_pixelVal_in_1_6;
      end else if (10'h1ef == _T_31[9:0]) begin
        image_1_495 <= io_pixelVal_in_1_5;
      end else if (10'h1ef == _T_28[9:0]) begin
        image_1_495 <= io_pixelVal_in_1_4;
      end else if (10'h1ef == _T_25[9:0]) begin
        image_1_495 <= io_pixelVal_in_1_3;
      end else if (10'h1ef == _T_22[9:0]) begin
        image_1_495 <= io_pixelVal_in_1_2;
      end else if (10'h1ef == _T_19[9:0]) begin
        image_1_495 <= io_pixelVal_in_1_1;
      end else if (10'h1ef == _T_15[9:0]) begin
        image_1_495 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_496 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f0 == _T_37[9:0]) begin
        image_1_496 <= io_pixelVal_in_1_7;
      end else if (10'h1f0 == _T_34[9:0]) begin
        image_1_496 <= io_pixelVal_in_1_6;
      end else if (10'h1f0 == _T_31[9:0]) begin
        image_1_496 <= io_pixelVal_in_1_5;
      end else if (10'h1f0 == _T_28[9:0]) begin
        image_1_496 <= io_pixelVal_in_1_4;
      end else if (10'h1f0 == _T_25[9:0]) begin
        image_1_496 <= io_pixelVal_in_1_3;
      end else if (10'h1f0 == _T_22[9:0]) begin
        image_1_496 <= io_pixelVal_in_1_2;
      end else if (10'h1f0 == _T_19[9:0]) begin
        image_1_496 <= io_pixelVal_in_1_1;
      end else if (10'h1f0 == _T_15[9:0]) begin
        image_1_496 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_497 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f1 == _T_37[9:0]) begin
        image_1_497 <= io_pixelVal_in_1_7;
      end else if (10'h1f1 == _T_34[9:0]) begin
        image_1_497 <= io_pixelVal_in_1_6;
      end else if (10'h1f1 == _T_31[9:0]) begin
        image_1_497 <= io_pixelVal_in_1_5;
      end else if (10'h1f1 == _T_28[9:0]) begin
        image_1_497 <= io_pixelVal_in_1_4;
      end else if (10'h1f1 == _T_25[9:0]) begin
        image_1_497 <= io_pixelVal_in_1_3;
      end else if (10'h1f1 == _T_22[9:0]) begin
        image_1_497 <= io_pixelVal_in_1_2;
      end else if (10'h1f1 == _T_19[9:0]) begin
        image_1_497 <= io_pixelVal_in_1_1;
      end else if (10'h1f1 == _T_15[9:0]) begin
        image_1_497 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_498 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f2 == _T_37[9:0]) begin
        image_1_498 <= io_pixelVal_in_1_7;
      end else if (10'h1f2 == _T_34[9:0]) begin
        image_1_498 <= io_pixelVal_in_1_6;
      end else if (10'h1f2 == _T_31[9:0]) begin
        image_1_498 <= io_pixelVal_in_1_5;
      end else if (10'h1f2 == _T_28[9:0]) begin
        image_1_498 <= io_pixelVal_in_1_4;
      end else if (10'h1f2 == _T_25[9:0]) begin
        image_1_498 <= io_pixelVal_in_1_3;
      end else if (10'h1f2 == _T_22[9:0]) begin
        image_1_498 <= io_pixelVal_in_1_2;
      end else if (10'h1f2 == _T_19[9:0]) begin
        image_1_498 <= io_pixelVal_in_1_1;
      end else if (10'h1f2 == _T_15[9:0]) begin
        image_1_498 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_499 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f3 == _T_37[9:0]) begin
        image_1_499 <= io_pixelVal_in_1_7;
      end else if (10'h1f3 == _T_34[9:0]) begin
        image_1_499 <= io_pixelVal_in_1_6;
      end else if (10'h1f3 == _T_31[9:0]) begin
        image_1_499 <= io_pixelVal_in_1_5;
      end else if (10'h1f3 == _T_28[9:0]) begin
        image_1_499 <= io_pixelVal_in_1_4;
      end else if (10'h1f3 == _T_25[9:0]) begin
        image_1_499 <= io_pixelVal_in_1_3;
      end else if (10'h1f3 == _T_22[9:0]) begin
        image_1_499 <= io_pixelVal_in_1_2;
      end else if (10'h1f3 == _T_19[9:0]) begin
        image_1_499 <= io_pixelVal_in_1_1;
      end else if (10'h1f3 == _T_15[9:0]) begin
        image_1_499 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_500 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f4 == _T_37[9:0]) begin
        image_1_500 <= io_pixelVal_in_1_7;
      end else if (10'h1f4 == _T_34[9:0]) begin
        image_1_500 <= io_pixelVal_in_1_6;
      end else if (10'h1f4 == _T_31[9:0]) begin
        image_1_500 <= io_pixelVal_in_1_5;
      end else if (10'h1f4 == _T_28[9:0]) begin
        image_1_500 <= io_pixelVal_in_1_4;
      end else if (10'h1f4 == _T_25[9:0]) begin
        image_1_500 <= io_pixelVal_in_1_3;
      end else if (10'h1f4 == _T_22[9:0]) begin
        image_1_500 <= io_pixelVal_in_1_2;
      end else if (10'h1f4 == _T_19[9:0]) begin
        image_1_500 <= io_pixelVal_in_1_1;
      end else if (10'h1f4 == _T_15[9:0]) begin
        image_1_500 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_501 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f5 == _T_37[9:0]) begin
        image_1_501 <= io_pixelVal_in_1_7;
      end else if (10'h1f5 == _T_34[9:0]) begin
        image_1_501 <= io_pixelVal_in_1_6;
      end else if (10'h1f5 == _T_31[9:0]) begin
        image_1_501 <= io_pixelVal_in_1_5;
      end else if (10'h1f5 == _T_28[9:0]) begin
        image_1_501 <= io_pixelVal_in_1_4;
      end else if (10'h1f5 == _T_25[9:0]) begin
        image_1_501 <= io_pixelVal_in_1_3;
      end else if (10'h1f5 == _T_22[9:0]) begin
        image_1_501 <= io_pixelVal_in_1_2;
      end else if (10'h1f5 == _T_19[9:0]) begin
        image_1_501 <= io_pixelVal_in_1_1;
      end else if (10'h1f5 == _T_15[9:0]) begin
        image_1_501 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_502 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f6 == _T_37[9:0]) begin
        image_1_502 <= io_pixelVal_in_1_7;
      end else if (10'h1f6 == _T_34[9:0]) begin
        image_1_502 <= io_pixelVal_in_1_6;
      end else if (10'h1f6 == _T_31[9:0]) begin
        image_1_502 <= io_pixelVal_in_1_5;
      end else if (10'h1f6 == _T_28[9:0]) begin
        image_1_502 <= io_pixelVal_in_1_4;
      end else if (10'h1f6 == _T_25[9:0]) begin
        image_1_502 <= io_pixelVal_in_1_3;
      end else if (10'h1f6 == _T_22[9:0]) begin
        image_1_502 <= io_pixelVal_in_1_2;
      end else if (10'h1f6 == _T_19[9:0]) begin
        image_1_502 <= io_pixelVal_in_1_1;
      end else if (10'h1f6 == _T_15[9:0]) begin
        image_1_502 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_503 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f7 == _T_37[9:0]) begin
        image_1_503 <= io_pixelVal_in_1_7;
      end else if (10'h1f7 == _T_34[9:0]) begin
        image_1_503 <= io_pixelVal_in_1_6;
      end else if (10'h1f7 == _T_31[9:0]) begin
        image_1_503 <= io_pixelVal_in_1_5;
      end else if (10'h1f7 == _T_28[9:0]) begin
        image_1_503 <= io_pixelVal_in_1_4;
      end else if (10'h1f7 == _T_25[9:0]) begin
        image_1_503 <= io_pixelVal_in_1_3;
      end else if (10'h1f7 == _T_22[9:0]) begin
        image_1_503 <= io_pixelVal_in_1_2;
      end else if (10'h1f7 == _T_19[9:0]) begin
        image_1_503 <= io_pixelVal_in_1_1;
      end else if (10'h1f7 == _T_15[9:0]) begin
        image_1_503 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_504 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f8 == _T_37[9:0]) begin
        image_1_504 <= io_pixelVal_in_1_7;
      end else if (10'h1f8 == _T_34[9:0]) begin
        image_1_504 <= io_pixelVal_in_1_6;
      end else if (10'h1f8 == _T_31[9:0]) begin
        image_1_504 <= io_pixelVal_in_1_5;
      end else if (10'h1f8 == _T_28[9:0]) begin
        image_1_504 <= io_pixelVal_in_1_4;
      end else if (10'h1f8 == _T_25[9:0]) begin
        image_1_504 <= io_pixelVal_in_1_3;
      end else if (10'h1f8 == _T_22[9:0]) begin
        image_1_504 <= io_pixelVal_in_1_2;
      end else if (10'h1f8 == _T_19[9:0]) begin
        image_1_504 <= io_pixelVal_in_1_1;
      end else if (10'h1f8 == _T_15[9:0]) begin
        image_1_504 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_505 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f9 == _T_37[9:0]) begin
        image_1_505 <= io_pixelVal_in_1_7;
      end else if (10'h1f9 == _T_34[9:0]) begin
        image_1_505 <= io_pixelVal_in_1_6;
      end else if (10'h1f9 == _T_31[9:0]) begin
        image_1_505 <= io_pixelVal_in_1_5;
      end else if (10'h1f9 == _T_28[9:0]) begin
        image_1_505 <= io_pixelVal_in_1_4;
      end else if (10'h1f9 == _T_25[9:0]) begin
        image_1_505 <= io_pixelVal_in_1_3;
      end else if (10'h1f9 == _T_22[9:0]) begin
        image_1_505 <= io_pixelVal_in_1_2;
      end else if (10'h1f9 == _T_19[9:0]) begin
        image_1_505 <= io_pixelVal_in_1_1;
      end else if (10'h1f9 == _T_15[9:0]) begin
        image_1_505 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_506 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1fa == _T_37[9:0]) begin
        image_1_506 <= io_pixelVal_in_1_7;
      end else if (10'h1fa == _T_34[9:0]) begin
        image_1_506 <= io_pixelVal_in_1_6;
      end else if (10'h1fa == _T_31[9:0]) begin
        image_1_506 <= io_pixelVal_in_1_5;
      end else if (10'h1fa == _T_28[9:0]) begin
        image_1_506 <= io_pixelVal_in_1_4;
      end else if (10'h1fa == _T_25[9:0]) begin
        image_1_506 <= io_pixelVal_in_1_3;
      end else if (10'h1fa == _T_22[9:0]) begin
        image_1_506 <= io_pixelVal_in_1_2;
      end else if (10'h1fa == _T_19[9:0]) begin
        image_1_506 <= io_pixelVal_in_1_1;
      end else if (10'h1fa == _T_15[9:0]) begin
        image_1_506 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_507 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1fb == _T_37[9:0]) begin
        image_1_507 <= io_pixelVal_in_1_7;
      end else if (10'h1fb == _T_34[9:0]) begin
        image_1_507 <= io_pixelVal_in_1_6;
      end else if (10'h1fb == _T_31[9:0]) begin
        image_1_507 <= io_pixelVal_in_1_5;
      end else if (10'h1fb == _T_28[9:0]) begin
        image_1_507 <= io_pixelVal_in_1_4;
      end else if (10'h1fb == _T_25[9:0]) begin
        image_1_507 <= io_pixelVal_in_1_3;
      end else if (10'h1fb == _T_22[9:0]) begin
        image_1_507 <= io_pixelVal_in_1_2;
      end else if (10'h1fb == _T_19[9:0]) begin
        image_1_507 <= io_pixelVal_in_1_1;
      end else if (10'h1fb == _T_15[9:0]) begin
        image_1_507 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_508 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1fc == _T_37[9:0]) begin
        image_1_508 <= io_pixelVal_in_1_7;
      end else if (10'h1fc == _T_34[9:0]) begin
        image_1_508 <= io_pixelVal_in_1_6;
      end else if (10'h1fc == _T_31[9:0]) begin
        image_1_508 <= io_pixelVal_in_1_5;
      end else if (10'h1fc == _T_28[9:0]) begin
        image_1_508 <= io_pixelVal_in_1_4;
      end else if (10'h1fc == _T_25[9:0]) begin
        image_1_508 <= io_pixelVal_in_1_3;
      end else if (10'h1fc == _T_22[9:0]) begin
        image_1_508 <= io_pixelVal_in_1_2;
      end else if (10'h1fc == _T_19[9:0]) begin
        image_1_508 <= io_pixelVal_in_1_1;
      end else if (10'h1fc == _T_15[9:0]) begin
        image_1_508 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_509 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1fd == _T_37[9:0]) begin
        image_1_509 <= io_pixelVal_in_1_7;
      end else if (10'h1fd == _T_34[9:0]) begin
        image_1_509 <= io_pixelVal_in_1_6;
      end else if (10'h1fd == _T_31[9:0]) begin
        image_1_509 <= io_pixelVal_in_1_5;
      end else if (10'h1fd == _T_28[9:0]) begin
        image_1_509 <= io_pixelVal_in_1_4;
      end else if (10'h1fd == _T_25[9:0]) begin
        image_1_509 <= io_pixelVal_in_1_3;
      end else if (10'h1fd == _T_22[9:0]) begin
        image_1_509 <= io_pixelVal_in_1_2;
      end else if (10'h1fd == _T_19[9:0]) begin
        image_1_509 <= io_pixelVal_in_1_1;
      end else if (10'h1fd == _T_15[9:0]) begin
        image_1_509 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_510 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1fe == _T_37[9:0]) begin
        image_1_510 <= io_pixelVal_in_1_7;
      end else if (10'h1fe == _T_34[9:0]) begin
        image_1_510 <= io_pixelVal_in_1_6;
      end else if (10'h1fe == _T_31[9:0]) begin
        image_1_510 <= io_pixelVal_in_1_5;
      end else if (10'h1fe == _T_28[9:0]) begin
        image_1_510 <= io_pixelVal_in_1_4;
      end else if (10'h1fe == _T_25[9:0]) begin
        image_1_510 <= io_pixelVal_in_1_3;
      end else if (10'h1fe == _T_22[9:0]) begin
        image_1_510 <= io_pixelVal_in_1_2;
      end else if (10'h1fe == _T_19[9:0]) begin
        image_1_510 <= io_pixelVal_in_1_1;
      end else if (10'h1fe == _T_15[9:0]) begin
        image_1_510 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_511 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ff == _T_37[9:0]) begin
        image_1_511 <= io_pixelVal_in_1_7;
      end else if (10'h1ff == _T_34[9:0]) begin
        image_1_511 <= io_pixelVal_in_1_6;
      end else if (10'h1ff == _T_31[9:0]) begin
        image_1_511 <= io_pixelVal_in_1_5;
      end else if (10'h1ff == _T_28[9:0]) begin
        image_1_511 <= io_pixelVal_in_1_4;
      end else if (10'h1ff == _T_25[9:0]) begin
        image_1_511 <= io_pixelVal_in_1_3;
      end else if (10'h1ff == _T_22[9:0]) begin
        image_1_511 <= io_pixelVal_in_1_2;
      end else if (10'h1ff == _T_19[9:0]) begin
        image_1_511 <= io_pixelVal_in_1_1;
      end else if (10'h1ff == _T_15[9:0]) begin
        image_1_511 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_512 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h200 == _T_37[9:0]) begin
        image_1_512 <= io_pixelVal_in_1_7;
      end else if (10'h200 == _T_34[9:0]) begin
        image_1_512 <= io_pixelVal_in_1_6;
      end else if (10'h200 == _T_31[9:0]) begin
        image_1_512 <= io_pixelVal_in_1_5;
      end else if (10'h200 == _T_28[9:0]) begin
        image_1_512 <= io_pixelVal_in_1_4;
      end else if (10'h200 == _T_25[9:0]) begin
        image_1_512 <= io_pixelVal_in_1_3;
      end else if (10'h200 == _T_22[9:0]) begin
        image_1_512 <= io_pixelVal_in_1_2;
      end else if (10'h200 == _T_19[9:0]) begin
        image_1_512 <= io_pixelVal_in_1_1;
      end else if (10'h200 == _T_15[9:0]) begin
        image_1_512 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_513 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h201 == _T_37[9:0]) begin
        image_1_513 <= io_pixelVal_in_1_7;
      end else if (10'h201 == _T_34[9:0]) begin
        image_1_513 <= io_pixelVal_in_1_6;
      end else if (10'h201 == _T_31[9:0]) begin
        image_1_513 <= io_pixelVal_in_1_5;
      end else if (10'h201 == _T_28[9:0]) begin
        image_1_513 <= io_pixelVal_in_1_4;
      end else if (10'h201 == _T_25[9:0]) begin
        image_1_513 <= io_pixelVal_in_1_3;
      end else if (10'h201 == _T_22[9:0]) begin
        image_1_513 <= io_pixelVal_in_1_2;
      end else if (10'h201 == _T_19[9:0]) begin
        image_1_513 <= io_pixelVal_in_1_1;
      end else if (10'h201 == _T_15[9:0]) begin
        image_1_513 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_514 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h202 == _T_37[9:0]) begin
        image_1_514 <= io_pixelVal_in_1_7;
      end else if (10'h202 == _T_34[9:0]) begin
        image_1_514 <= io_pixelVal_in_1_6;
      end else if (10'h202 == _T_31[9:0]) begin
        image_1_514 <= io_pixelVal_in_1_5;
      end else if (10'h202 == _T_28[9:0]) begin
        image_1_514 <= io_pixelVal_in_1_4;
      end else if (10'h202 == _T_25[9:0]) begin
        image_1_514 <= io_pixelVal_in_1_3;
      end else if (10'h202 == _T_22[9:0]) begin
        image_1_514 <= io_pixelVal_in_1_2;
      end else if (10'h202 == _T_19[9:0]) begin
        image_1_514 <= io_pixelVal_in_1_1;
      end else if (10'h202 == _T_15[9:0]) begin
        image_1_514 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_515 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h203 == _T_37[9:0]) begin
        image_1_515 <= io_pixelVal_in_1_7;
      end else if (10'h203 == _T_34[9:0]) begin
        image_1_515 <= io_pixelVal_in_1_6;
      end else if (10'h203 == _T_31[9:0]) begin
        image_1_515 <= io_pixelVal_in_1_5;
      end else if (10'h203 == _T_28[9:0]) begin
        image_1_515 <= io_pixelVal_in_1_4;
      end else if (10'h203 == _T_25[9:0]) begin
        image_1_515 <= io_pixelVal_in_1_3;
      end else if (10'h203 == _T_22[9:0]) begin
        image_1_515 <= io_pixelVal_in_1_2;
      end else if (10'h203 == _T_19[9:0]) begin
        image_1_515 <= io_pixelVal_in_1_1;
      end else if (10'h203 == _T_15[9:0]) begin
        image_1_515 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_516 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h204 == _T_37[9:0]) begin
        image_1_516 <= io_pixelVal_in_1_7;
      end else if (10'h204 == _T_34[9:0]) begin
        image_1_516 <= io_pixelVal_in_1_6;
      end else if (10'h204 == _T_31[9:0]) begin
        image_1_516 <= io_pixelVal_in_1_5;
      end else if (10'h204 == _T_28[9:0]) begin
        image_1_516 <= io_pixelVal_in_1_4;
      end else if (10'h204 == _T_25[9:0]) begin
        image_1_516 <= io_pixelVal_in_1_3;
      end else if (10'h204 == _T_22[9:0]) begin
        image_1_516 <= io_pixelVal_in_1_2;
      end else if (10'h204 == _T_19[9:0]) begin
        image_1_516 <= io_pixelVal_in_1_1;
      end else if (10'h204 == _T_15[9:0]) begin
        image_1_516 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_517 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h205 == _T_37[9:0]) begin
        image_1_517 <= io_pixelVal_in_1_7;
      end else if (10'h205 == _T_34[9:0]) begin
        image_1_517 <= io_pixelVal_in_1_6;
      end else if (10'h205 == _T_31[9:0]) begin
        image_1_517 <= io_pixelVal_in_1_5;
      end else if (10'h205 == _T_28[9:0]) begin
        image_1_517 <= io_pixelVal_in_1_4;
      end else if (10'h205 == _T_25[9:0]) begin
        image_1_517 <= io_pixelVal_in_1_3;
      end else if (10'h205 == _T_22[9:0]) begin
        image_1_517 <= io_pixelVal_in_1_2;
      end else if (10'h205 == _T_19[9:0]) begin
        image_1_517 <= io_pixelVal_in_1_1;
      end else if (10'h205 == _T_15[9:0]) begin
        image_1_517 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_518 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h206 == _T_37[9:0]) begin
        image_1_518 <= io_pixelVal_in_1_7;
      end else if (10'h206 == _T_34[9:0]) begin
        image_1_518 <= io_pixelVal_in_1_6;
      end else if (10'h206 == _T_31[9:0]) begin
        image_1_518 <= io_pixelVal_in_1_5;
      end else if (10'h206 == _T_28[9:0]) begin
        image_1_518 <= io_pixelVal_in_1_4;
      end else if (10'h206 == _T_25[9:0]) begin
        image_1_518 <= io_pixelVal_in_1_3;
      end else if (10'h206 == _T_22[9:0]) begin
        image_1_518 <= io_pixelVal_in_1_2;
      end else if (10'h206 == _T_19[9:0]) begin
        image_1_518 <= io_pixelVal_in_1_1;
      end else if (10'h206 == _T_15[9:0]) begin
        image_1_518 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_519 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h207 == _T_37[9:0]) begin
        image_1_519 <= io_pixelVal_in_1_7;
      end else if (10'h207 == _T_34[9:0]) begin
        image_1_519 <= io_pixelVal_in_1_6;
      end else if (10'h207 == _T_31[9:0]) begin
        image_1_519 <= io_pixelVal_in_1_5;
      end else if (10'h207 == _T_28[9:0]) begin
        image_1_519 <= io_pixelVal_in_1_4;
      end else if (10'h207 == _T_25[9:0]) begin
        image_1_519 <= io_pixelVal_in_1_3;
      end else if (10'h207 == _T_22[9:0]) begin
        image_1_519 <= io_pixelVal_in_1_2;
      end else if (10'h207 == _T_19[9:0]) begin
        image_1_519 <= io_pixelVal_in_1_1;
      end else if (10'h207 == _T_15[9:0]) begin
        image_1_519 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_520 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h208 == _T_37[9:0]) begin
        image_1_520 <= io_pixelVal_in_1_7;
      end else if (10'h208 == _T_34[9:0]) begin
        image_1_520 <= io_pixelVal_in_1_6;
      end else if (10'h208 == _T_31[9:0]) begin
        image_1_520 <= io_pixelVal_in_1_5;
      end else if (10'h208 == _T_28[9:0]) begin
        image_1_520 <= io_pixelVal_in_1_4;
      end else if (10'h208 == _T_25[9:0]) begin
        image_1_520 <= io_pixelVal_in_1_3;
      end else if (10'h208 == _T_22[9:0]) begin
        image_1_520 <= io_pixelVal_in_1_2;
      end else if (10'h208 == _T_19[9:0]) begin
        image_1_520 <= io_pixelVal_in_1_1;
      end else if (10'h208 == _T_15[9:0]) begin
        image_1_520 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_521 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h209 == _T_37[9:0]) begin
        image_1_521 <= io_pixelVal_in_1_7;
      end else if (10'h209 == _T_34[9:0]) begin
        image_1_521 <= io_pixelVal_in_1_6;
      end else if (10'h209 == _T_31[9:0]) begin
        image_1_521 <= io_pixelVal_in_1_5;
      end else if (10'h209 == _T_28[9:0]) begin
        image_1_521 <= io_pixelVal_in_1_4;
      end else if (10'h209 == _T_25[9:0]) begin
        image_1_521 <= io_pixelVal_in_1_3;
      end else if (10'h209 == _T_22[9:0]) begin
        image_1_521 <= io_pixelVal_in_1_2;
      end else if (10'h209 == _T_19[9:0]) begin
        image_1_521 <= io_pixelVal_in_1_1;
      end else if (10'h209 == _T_15[9:0]) begin
        image_1_521 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_522 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20a == _T_37[9:0]) begin
        image_1_522 <= io_pixelVal_in_1_7;
      end else if (10'h20a == _T_34[9:0]) begin
        image_1_522 <= io_pixelVal_in_1_6;
      end else if (10'h20a == _T_31[9:0]) begin
        image_1_522 <= io_pixelVal_in_1_5;
      end else if (10'h20a == _T_28[9:0]) begin
        image_1_522 <= io_pixelVal_in_1_4;
      end else if (10'h20a == _T_25[9:0]) begin
        image_1_522 <= io_pixelVal_in_1_3;
      end else if (10'h20a == _T_22[9:0]) begin
        image_1_522 <= io_pixelVal_in_1_2;
      end else if (10'h20a == _T_19[9:0]) begin
        image_1_522 <= io_pixelVal_in_1_1;
      end else if (10'h20a == _T_15[9:0]) begin
        image_1_522 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_523 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20b == _T_37[9:0]) begin
        image_1_523 <= io_pixelVal_in_1_7;
      end else if (10'h20b == _T_34[9:0]) begin
        image_1_523 <= io_pixelVal_in_1_6;
      end else if (10'h20b == _T_31[9:0]) begin
        image_1_523 <= io_pixelVal_in_1_5;
      end else if (10'h20b == _T_28[9:0]) begin
        image_1_523 <= io_pixelVal_in_1_4;
      end else if (10'h20b == _T_25[9:0]) begin
        image_1_523 <= io_pixelVal_in_1_3;
      end else if (10'h20b == _T_22[9:0]) begin
        image_1_523 <= io_pixelVal_in_1_2;
      end else if (10'h20b == _T_19[9:0]) begin
        image_1_523 <= io_pixelVal_in_1_1;
      end else if (10'h20b == _T_15[9:0]) begin
        image_1_523 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_524 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20c == _T_37[9:0]) begin
        image_1_524 <= io_pixelVal_in_1_7;
      end else if (10'h20c == _T_34[9:0]) begin
        image_1_524 <= io_pixelVal_in_1_6;
      end else if (10'h20c == _T_31[9:0]) begin
        image_1_524 <= io_pixelVal_in_1_5;
      end else if (10'h20c == _T_28[9:0]) begin
        image_1_524 <= io_pixelVal_in_1_4;
      end else if (10'h20c == _T_25[9:0]) begin
        image_1_524 <= io_pixelVal_in_1_3;
      end else if (10'h20c == _T_22[9:0]) begin
        image_1_524 <= io_pixelVal_in_1_2;
      end else if (10'h20c == _T_19[9:0]) begin
        image_1_524 <= io_pixelVal_in_1_1;
      end else if (10'h20c == _T_15[9:0]) begin
        image_1_524 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_525 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20d == _T_37[9:0]) begin
        image_1_525 <= io_pixelVal_in_1_7;
      end else if (10'h20d == _T_34[9:0]) begin
        image_1_525 <= io_pixelVal_in_1_6;
      end else if (10'h20d == _T_31[9:0]) begin
        image_1_525 <= io_pixelVal_in_1_5;
      end else if (10'h20d == _T_28[9:0]) begin
        image_1_525 <= io_pixelVal_in_1_4;
      end else if (10'h20d == _T_25[9:0]) begin
        image_1_525 <= io_pixelVal_in_1_3;
      end else if (10'h20d == _T_22[9:0]) begin
        image_1_525 <= io_pixelVal_in_1_2;
      end else if (10'h20d == _T_19[9:0]) begin
        image_1_525 <= io_pixelVal_in_1_1;
      end else if (10'h20d == _T_15[9:0]) begin
        image_1_525 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_526 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20e == _T_37[9:0]) begin
        image_1_526 <= io_pixelVal_in_1_7;
      end else if (10'h20e == _T_34[9:0]) begin
        image_1_526 <= io_pixelVal_in_1_6;
      end else if (10'h20e == _T_31[9:0]) begin
        image_1_526 <= io_pixelVal_in_1_5;
      end else if (10'h20e == _T_28[9:0]) begin
        image_1_526 <= io_pixelVal_in_1_4;
      end else if (10'h20e == _T_25[9:0]) begin
        image_1_526 <= io_pixelVal_in_1_3;
      end else if (10'h20e == _T_22[9:0]) begin
        image_1_526 <= io_pixelVal_in_1_2;
      end else if (10'h20e == _T_19[9:0]) begin
        image_1_526 <= io_pixelVal_in_1_1;
      end else if (10'h20e == _T_15[9:0]) begin
        image_1_526 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_527 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20f == _T_37[9:0]) begin
        image_1_527 <= io_pixelVal_in_1_7;
      end else if (10'h20f == _T_34[9:0]) begin
        image_1_527 <= io_pixelVal_in_1_6;
      end else if (10'h20f == _T_31[9:0]) begin
        image_1_527 <= io_pixelVal_in_1_5;
      end else if (10'h20f == _T_28[9:0]) begin
        image_1_527 <= io_pixelVal_in_1_4;
      end else if (10'h20f == _T_25[9:0]) begin
        image_1_527 <= io_pixelVal_in_1_3;
      end else if (10'h20f == _T_22[9:0]) begin
        image_1_527 <= io_pixelVal_in_1_2;
      end else if (10'h20f == _T_19[9:0]) begin
        image_1_527 <= io_pixelVal_in_1_1;
      end else if (10'h20f == _T_15[9:0]) begin
        image_1_527 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_528 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h210 == _T_37[9:0]) begin
        image_1_528 <= io_pixelVal_in_1_7;
      end else if (10'h210 == _T_34[9:0]) begin
        image_1_528 <= io_pixelVal_in_1_6;
      end else if (10'h210 == _T_31[9:0]) begin
        image_1_528 <= io_pixelVal_in_1_5;
      end else if (10'h210 == _T_28[9:0]) begin
        image_1_528 <= io_pixelVal_in_1_4;
      end else if (10'h210 == _T_25[9:0]) begin
        image_1_528 <= io_pixelVal_in_1_3;
      end else if (10'h210 == _T_22[9:0]) begin
        image_1_528 <= io_pixelVal_in_1_2;
      end else if (10'h210 == _T_19[9:0]) begin
        image_1_528 <= io_pixelVal_in_1_1;
      end else if (10'h210 == _T_15[9:0]) begin
        image_1_528 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_529 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h211 == _T_37[9:0]) begin
        image_1_529 <= io_pixelVal_in_1_7;
      end else if (10'h211 == _T_34[9:0]) begin
        image_1_529 <= io_pixelVal_in_1_6;
      end else if (10'h211 == _T_31[9:0]) begin
        image_1_529 <= io_pixelVal_in_1_5;
      end else if (10'h211 == _T_28[9:0]) begin
        image_1_529 <= io_pixelVal_in_1_4;
      end else if (10'h211 == _T_25[9:0]) begin
        image_1_529 <= io_pixelVal_in_1_3;
      end else if (10'h211 == _T_22[9:0]) begin
        image_1_529 <= io_pixelVal_in_1_2;
      end else if (10'h211 == _T_19[9:0]) begin
        image_1_529 <= io_pixelVal_in_1_1;
      end else if (10'h211 == _T_15[9:0]) begin
        image_1_529 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_530 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h212 == _T_37[9:0]) begin
        image_1_530 <= io_pixelVal_in_1_7;
      end else if (10'h212 == _T_34[9:0]) begin
        image_1_530 <= io_pixelVal_in_1_6;
      end else if (10'h212 == _T_31[9:0]) begin
        image_1_530 <= io_pixelVal_in_1_5;
      end else if (10'h212 == _T_28[9:0]) begin
        image_1_530 <= io_pixelVal_in_1_4;
      end else if (10'h212 == _T_25[9:0]) begin
        image_1_530 <= io_pixelVal_in_1_3;
      end else if (10'h212 == _T_22[9:0]) begin
        image_1_530 <= io_pixelVal_in_1_2;
      end else if (10'h212 == _T_19[9:0]) begin
        image_1_530 <= io_pixelVal_in_1_1;
      end else if (10'h212 == _T_15[9:0]) begin
        image_1_530 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_531 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h213 == _T_37[9:0]) begin
        image_1_531 <= io_pixelVal_in_1_7;
      end else if (10'h213 == _T_34[9:0]) begin
        image_1_531 <= io_pixelVal_in_1_6;
      end else if (10'h213 == _T_31[9:0]) begin
        image_1_531 <= io_pixelVal_in_1_5;
      end else if (10'h213 == _T_28[9:0]) begin
        image_1_531 <= io_pixelVal_in_1_4;
      end else if (10'h213 == _T_25[9:0]) begin
        image_1_531 <= io_pixelVal_in_1_3;
      end else if (10'h213 == _T_22[9:0]) begin
        image_1_531 <= io_pixelVal_in_1_2;
      end else if (10'h213 == _T_19[9:0]) begin
        image_1_531 <= io_pixelVal_in_1_1;
      end else if (10'h213 == _T_15[9:0]) begin
        image_1_531 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_532 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h214 == _T_37[9:0]) begin
        image_1_532 <= io_pixelVal_in_1_7;
      end else if (10'h214 == _T_34[9:0]) begin
        image_1_532 <= io_pixelVal_in_1_6;
      end else if (10'h214 == _T_31[9:0]) begin
        image_1_532 <= io_pixelVal_in_1_5;
      end else if (10'h214 == _T_28[9:0]) begin
        image_1_532 <= io_pixelVal_in_1_4;
      end else if (10'h214 == _T_25[9:0]) begin
        image_1_532 <= io_pixelVal_in_1_3;
      end else if (10'h214 == _T_22[9:0]) begin
        image_1_532 <= io_pixelVal_in_1_2;
      end else if (10'h214 == _T_19[9:0]) begin
        image_1_532 <= io_pixelVal_in_1_1;
      end else if (10'h214 == _T_15[9:0]) begin
        image_1_532 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_533 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h215 == _T_37[9:0]) begin
        image_1_533 <= io_pixelVal_in_1_7;
      end else if (10'h215 == _T_34[9:0]) begin
        image_1_533 <= io_pixelVal_in_1_6;
      end else if (10'h215 == _T_31[9:0]) begin
        image_1_533 <= io_pixelVal_in_1_5;
      end else if (10'h215 == _T_28[9:0]) begin
        image_1_533 <= io_pixelVal_in_1_4;
      end else if (10'h215 == _T_25[9:0]) begin
        image_1_533 <= io_pixelVal_in_1_3;
      end else if (10'h215 == _T_22[9:0]) begin
        image_1_533 <= io_pixelVal_in_1_2;
      end else if (10'h215 == _T_19[9:0]) begin
        image_1_533 <= io_pixelVal_in_1_1;
      end else if (10'h215 == _T_15[9:0]) begin
        image_1_533 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_534 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h216 == _T_37[9:0]) begin
        image_1_534 <= io_pixelVal_in_1_7;
      end else if (10'h216 == _T_34[9:0]) begin
        image_1_534 <= io_pixelVal_in_1_6;
      end else if (10'h216 == _T_31[9:0]) begin
        image_1_534 <= io_pixelVal_in_1_5;
      end else if (10'h216 == _T_28[9:0]) begin
        image_1_534 <= io_pixelVal_in_1_4;
      end else if (10'h216 == _T_25[9:0]) begin
        image_1_534 <= io_pixelVal_in_1_3;
      end else if (10'h216 == _T_22[9:0]) begin
        image_1_534 <= io_pixelVal_in_1_2;
      end else if (10'h216 == _T_19[9:0]) begin
        image_1_534 <= io_pixelVal_in_1_1;
      end else if (10'h216 == _T_15[9:0]) begin
        image_1_534 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_535 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h217 == _T_37[9:0]) begin
        image_1_535 <= io_pixelVal_in_1_7;
      end else if (10'h217 == _T_34[9:0]) begin
        image_1_535 <= io_pixelVal_in_1_6;
      end else if (10'h217 == _T_31[9:0]) begin
        image_1_535 <= io_pixelVal_in_1_5;
      end else if (10'h217 == _T_28[9:0]) begin
        image_1_535 <= io_pixelVal_in_1_4;
      end else if (10'h217 == _T_25[9:0]) begin
        image_1_535 <= io_pixelVal_in_1_3;
      end else if (10'h217 == _T_22[9:0]) begin
        image_1_535 <= io_pixelVal_in_1_2;
      end else if (10'h217 == _T_19[9:0]) begin
        image_1_535 <= io_pixelVal_in_1_1;
      end else if (10'h217 == _T_15[9:0]) begin
        image_1_535 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_536 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h218 == _T_37[9:0]) begin
        image_1_536 <= io_pixelVal_in_1_7;
      end else if (10'h218 == _T_34[9:0]) begin
        image_1_536 <= io_pixelVal_in_1_6;
      end else if (10'h218 == _T_31[9:0]) begin
        image_1_536 <= io_pixelVal_in_1_5;
      end else if (10'h218 == _T_28[9:0]) begin
        image_1_536 <= io_pixelVal_in_1_4;
      end else if (10'h218 == _T_25[9:0]) begin
        image_1_536 <= io_pixelVal_in_1_3;
      end else if (10'h218 == _T_22[9:0]) begin
        image_1_536 <= io_pixelVal_in_1_2;
      end else if (10'h218 == _T_19[9:0]) begin
        image_1_536 <= io_pixelVal_in_1_1;
      end else if (10'h218 == _T_15[9:0]) begin
        image_1_536 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_537 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h219 == _T_37[9:0]) begin
        image_1_537 <= io_pixelVal_in_1_7;
      end else if (10'h219 == _T_34[9:0]) begin
        image_1_537 <= io_pixelVal_in_1_6;
      end else if (10'h219 == _T_31[9:0]) begin
        image_1_537 <= io_pixelVal_in_1_5;
      end else if (10'h219 == _T_28[9:0]) begin
        image_1_537 <= io_pixelVal_in_1_4;
      end else if (10'h219 == _T_25[9:0]) begin
        image_1_537 <= io_pixelVal_in_1_3;
      end else if (10'h219 == _T_22[9:0]) begin
        image_1_537 <= io_pixelVal_in_1_2;
      end else if (10'h219 == _T_19[9:0]) begin
        image_1_537 <= io_pixelVal_in_1_1;
      end else if (10'h219 == _T_15[9:0]) begin
        image_1_537 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_538 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21a == _T_37[9:0]) begin
        image_1_538 <= io_pixelVal_in_1_7;
      end else if (10'h21a == _T_34[9:0]) begin
        image_1_538 <= io_pixelVal_in_1_6;
      end else if (10'h21a == _T_31[9:0]) begin
        image_1_538 <= io_pixelVal_in_1_5;
      end else if (10'h21a == _T_28[9:0]) begin
        image_1_538 <= io_pixelVal_in_1_4;
      end else if (10'h21a == _T_25[9:0]) begin
        image_1_538 <= io_pixelVal_in_1_3;
      end else if (10'h21a == _T_22[9:0]) begin
        image_1_538 <= io_pixelVal_in_1_2;
      end else if (10'h21a == _T_19[9:0]) begin
        image_1_538 <= io_pixelVal_in_1_1;
      end else if (10'h21a == _T_15[9:0]) begin
        image_1_538 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_539 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21b == _T_37[9:0]) begin
        image_1_539 <= io_pixelVal_in_1_7;
      end else if (10'h21b == _T_34[9:0]) begin
        image_1_539 <= io_pixelVal_in_1_6;
      end else if (10'h21b == _T_31[9:0]) begin
        image_1_539 <= io_pixelVal_in_1_5;
      end else if (10'h21b == _T_28[9:0]) begin
        image_1_539 <= io_pixelVal_in_1_4;
      end else if (10'h21b == _T_25[9:0]) begin
        image_1_539 <= io_pixelVal_in_1_3;
      end else if (10'h21b == _T_22[9:0]) begin
        image_1_539 <= io_pixelVal_in_1_2;
      end else if (10'h21b == _T_19[9:0]) begin
        image_1_539 <= io_pixelVal_in_1_1;
      end else if (10'h21b == _T_15[9:0]) begin
        image_1_539 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_540 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21c == _T_37[9:0]) begin
        image_1_540 <= io_pixelVal_in_1_7;
      end else if (10'h21c == _T_34[9:0]) begin
        image_1_540 <= io_pixelVal_in_1_6;
      end else if (10'h21c == _T_31[9:0]) begin
        image_1_540 <= io_pixelVal_in_1_5;
      end else if (10'h21c == _T_28[9:0]) begin
        image_1_540 <= io_pixelVal_in_1_4;
      end else if (10'h21c == _T_25[9:0]) begin
        image_1_540 <= io_pixelVal_in_1_3;
      end else if (10'h21c == _T_22[9:0]) begin
        image_1_540 <= io_pixelVal_in_1_2;
      end else if (10'h21c == _T_19[9:0]) begin
        image_1_540 <= io_pixelVal_in_1_1;
      end else if (10'h21c == _T_15[9:0]) begin
        image_1_540 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_541 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21d == _T_37[9:0]) begin
        image_1_541 <= io_pixelVal_in_1_7;
      end else if (10'h21d == _T_34[9:0]) begin
        image_1_541 <= io_pixelVal_in_1_6;
      end else if (10'h21d == _T_31[9:0]) begin
        image_1_541 <= io_pixelVal_in_1_5;
      end else if (10'h21d == _T_28[9:0]) begin
        image_1_541 <= io_pixelVal_in_1_4;
      end else if (10'h21d == _T_25[9:0]) begin
        image_1_541 <= io_pixelVal_in_1_3;
      end else if (10'h21d == _T_22[9:0]) begin
        image_1_541 <= io_pixelVal_in_1_2;
      end else if (10'h21d == _T_19[9:0]) begin
        image_1_541 <= io_pixelVal_in_1_1;
      end else if (10'h21d == _T_15[9:0]) begin
        image_1_541 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_542 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21e == _T_37[9:0]) begin
        image_1_542 <= io_pixelVal_in_1_7;
      end else if (10'h21e == _T_34[9:0]) begin
        image_1_542 <= io_pixelVal_in_1_6;
      end else if (10'h21e == _T_31[9:0]) begin
        image_1_542 <= io_pixelVal_in_1_5;
      end else if (10'h21e == _T_28[9:0]) begin
        image_1_542 <= io_pixelVal_in_1_4;
      end else if (10'h21e == _T_25[9:0]) begin
        image_1_542 <= io_pixelVal_in_1_3;
      end else if (10'h21e == _T_22[9:0]) begin
        image_1_542 <= io_pixelVal_in_1_2;
      end else if (10'h21e == _T_19[9:0]) begin
        image_1_542 <= io_pixelVal_in_1_1;
      end else if (10'h21e == _T_15[9:0]) begin
        image_1_542 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_543 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21f == _T_37[9:0]) begin
        image_1_543 <= io_pixelVal_in_1_7;
      end else if (10'h21f == _T_34[9:0]) begin
        image_1_543 <= io_pixelVal_in_1_6;
      end else if (10'h21f == _T_31[9:0]) begin
        image_1_543 <= io_pixelVal_in_1_5;
      end else if (10'h21f == _T_28[9:0]) begin
        image_1_543 <= io_pixelVal_in_1_4;
      end else if (10'h21f == _T_25[9:0]) begin
        image_1_543 <= io_pixelVal_in_1_3;
      end else if (10'h21f == _T_22[9:0]) begin
        image_1_543 <= io_pixelVal_in_1_2;
      end else if (10'h21f == _T_19[9:0]) begin
        image_1_543 <= io_pixelVal_in_1_1;
      end else if (10'h21f == _T_15[9:0]) begin
        image_1_543 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_544 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h220 == _T_37[9:0]) begin
        image_1_544 <= io_pixelVal_in_1_7;
      end else if (10'h220 == _T_34[9:0]) begin
        image_1_544 <= io_pixelVal_in_1_6;
      end else if (10'h220 == _T_31[9:0]) begin
        image_1_544 <= io_pixelVal_in_1_5;
      end else if (10'h220 == _T_28[9:0]) begin
        image_1_544 <= io_pixelVal_in_1_4;
      end else if (10'h220 == _T_25[9:0]) begin
        image_1_544 <= io_pixelVal_in_1_3;
      end else if (10'h220 == _T_22[9:0]) begin
        image_1_544 <= io_pixelVal_in_1_2;
      end else if (10'h220 == _T_19[9:0]) begin
        image_1_544 <= io_pixelVal_in_1_1;
      end else if (10'h220 == _T_15[9:0]) begin
        image_1_544 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_545 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h221 == _T_37[9:0]) begin
        image_1_545 <= io_pixelVal_in_1_7;
      end else if (10'h221 == _T_34[9:0]) begin
        image_1_545 <= io_pixelVal_in_1_6;
      end else if (10'h221 == _T_31[9:0]) begin
        image_1_545 <= io_pixelVal_in_1_5;
      end else if (10'h221 == _T_28[9:0]) begin
        image_1_545 <= io_pixelVal_in_1_4;
      end else if (10'h221 == _T_25[9:0]) begin
        image_1_545 <= io_pixelVal_in_1_3;
      end else if (10'h221 == _T_22[9:0]) begin
        image_1_545 <= io_pixelVal_in_1_2;
      end else if (10'h221 == _T_19[9:0]) begin
        image_1_545 <= io_pixelVal_in_1_1;
      end else if (10'h221 == _T_15[9:0]) begin
        image_1_545 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_546 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h222 == _T_37[9:0]) begin
        image_1_546 <= io_pixelVal_in_1_7;
      end else if (10'h222 == _T_34[9:0]) begin
        image_1_546 <= io_pixelVal_in_1_6;
      end else if (10'h222 == _T_31[9:0]) begin
        image_1_546 <= io_pixelVal_in_1_5;
      end else if (10'h222 == _T_28[9:0]) begin
        image_1_546 <= io_pixelVal_in_1_4;
      end else if (10'h222 == _T_25[9:0]) begin
        image_1_546 <= io_pixelVal_in_1_3;
      end else if (10'h222 == _T_22[9:0]) begin
        image_1_546 <= io_pixelVal_in_1_2;
      end else if (10'h222 == _T_19[9:0]) begin
        image_1_546 <= io_pixelVal_in_1_1;
      end else if (10'h222 == _T_15[9:0]) begin
        image_1_546 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_547 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h223 == _T_37[9:0]) begin
        image_1_547 <= io_pixelVal_in_1_7;
      end else if (10'h223 == _T_34[9:0]) begin
        image_1_547 <= io_pixelVal_in_1_6;
      end else if (10'h223 == _T_31[9:0]) begin
        image_1_547 <= io_pixelVal_in_1_5;
      end else if (10'h223 == _T_28[9:0]) begin
        image_1_547 <= io_pixelVal_in_1_4;
      end else if (10'h223 == _T_25[9:0]) begin
        image_1_547 <= io_pixelVal_in_1_3;
      end else if (10'h223 == _T_22[9:0]) begin
        image_1_547 <= io_pixelVal_in_1_2;
      end else if (10'h223 == _T_19[9:0]) begin
        image_1_547 <= io_pixelVal_in_1_1;
      end else if (10'h223 == _T_15[9:0]) begin
        image_1_547 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_548 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h224 == _T_37[9:0]) begin
        image_1_548 <= io_pixelVal_in_1_7;
      end else if (10'h224 == _T_34[9:0]) begin
        image_1_548 <= io_pixelVal_in_1_6;
      end else if (10'h224 == _T_31[9:0]) begin
        image_1_548 <= io_pixelVal_in_1_5;
      end else if (10'h224 == _T_28[9:0]) begin
        image_1_548 <= io_pixelVal_in_1_4;
      end else if (10'h224 == _T_25[9:0]) begin
        image_1_548 <= io_pixelVal_in_1_3;
      end else if (10'h224 == _T_22[9:0]) begin
        image_1_548 <= io_pixelVal_in_1_2;
      end else if (10'h224 == _T_19[9:0]) begin
        image_1_548 <= io_pixelVal_in_1_1;
      end else if (10'h224 == _T_15[9:0]) begin
        image_1_548 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_549 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h225 == _T_37[9:0]) begin
        image_1_549 <= io_pixelVal_in_1_7;
      end else if (10'h225 == _T_34[9:0]) begin
        image_1_549 <= io_pixelVal_in_1_6;
      end else if (10'h225 == _T_31[9:0]) begin
        image_1_549 <= io_pixelVal_in_1_5;
      end else if (10'h225 == _T_28[9:0]) begin
        image_1_549 <= io_pixelVal_in_1_4;
      end else if (10'h225 == _T_25[9:0]) begin
        image_1_549 <= io_pixelVal_in_1_3;
      end else if (10'h225 == _T_22[9:0]) begin
        image_1_549 <= io_pixelVal_in_1_2;
      end else if (10'h225 == _T_19[9:0]) begin
        image_1_549 <= io_pixelVal_in_1_1;
      end else if (10'h225 == _T_15[9:0]) begin
        image_1_549 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_550 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h226 == _T_37[9:0]) begin
        image_1_550 <= io_pixelVal_in_1_7;
      end else if (10'h226 == _T_34[9:0]) begin
        image_1_550 <= io_pixelVal_in_1_6;
      end else if (10'h226 == _T_31[9:0]) begin
        image_1_550 <= io_pixelVal_in_1_5;
      end else if (10'h226 == _T_28[9:0]) begin
        image_1_550 <= io_pixelVal_in_1_4;
      end else if (10'h226 == _T_25[9:0]) begin
        image_1_550 <= io_pixelVal_in_1_3;
      end else if (10'h226 == _T_22[9:0]) begin
        image_1_550 <= io_pixelVal_in_1_2;
      end else if (10'h226 == _T_19[9:0]) begin
        image_1_550 <= io_pixelVal_in_1_1;
      end else if (10'h226 == _T_15[9:0]) begin
        image_1_550 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_551 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h227 == _T_37[9:0]) begin
        image_1_551 <= io_pixelVal_in_1_7;
      end else if (10'h227 == _T_34[9:0]) begin
        image_1_551 <= io_pixelVal_in_1_6;
      end else if (10'h227 == _T_31[9:0]) begin
        image_1_551 <= io_pixelVal_in_1_5;
      end else if (10'h227 == _T_28[9:0]) begin
        image_1_551 <= io_pixelVal_in_1_4;
      end else if (10'h227 == _T_25[9:0]) begin
        image_1_551 <= io_pixelVal_in_1_3;
      end else if (10'h227 == _T_22[9:0]) begin
        image_1_551 <= io_pixelVal_in_1_2;
      end else if (10'h227 == _T_19[9:0]) begin
        image_1_551 <= io_pixelVal_in_1_1;
      end else if (10'h227 == _T_15[9:0]) begin
        image_1_551 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_552 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h228 == _T_37[9:0]) begin
        image_1_552 <= io_pixelVal_in_1_7;
      end else if (10'h228 == _T_34[9:0]) begin
        image_1_552 <= io_pixelVal_in_1_6;
      end else if (10'h228 == _T_31[9:0]) begin
        image_1_552 <= io_pixelVal_in_1_5;
      end else if (10'h228 == _T_28[9:0]) begin
        image_1_552 <= io_pixelVal_in_1_4;
      end else if (10'h228 == _T_25[9:0]) begin
        image_1_552 <= io_pixelVal_in_1_3;
      end else if (10'h228 == _T_22[9:0]) begin
        image_1_552 <= io_pixelVal_in_1_2;
      end else if (10'h228 == _T_19[9:0]) begin
        image_1_552 <= io_pixelVal_in_1_1;
      end else if (10'h228 == _T_15[9:0]) begin
        image_1_552 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_553 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h229 == _T_37[9:0]) begin
        image_1_553 <= io_pixelVal_in_1_7;
      end else if (10'h229 == _T_34[9:0]) begin
        image_1_553 <= io_pixelVal_in_1_6;
      end else if (10'h229 == _T_31[9:0]) begin
        image_1_553 <= io_pixelVal_in_1_5;
      end else if (10'h229 == _T_28[9:0]) begin
        image_1_553 <= io_pixelVal_in_1_4;
      end else if (10'h229 == _T_25[9:0]) begin
        image_1_553 <= io_pixelVal_in_1_3;
      end else if (10'h229 == _T_22[9:0]) begin
        image_1_553 <= io_pixelVal_in_1_2;
      end else if (10'h229 == _T_19[9:0]) begin
        image_1_553 <= io_pixelVal_in_1_1;
      end else if (10'h229 == _T_15[9:0]) begin
        image_1_553 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_554 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22a == _T_37[9:0]) begin
        image_1_554 <= io_pixelVal_in_1_7;
      end else if (10'h22a == _T_34[9:0]) begin
        image_1_554 <= io_pixelVal_in_1_6;
      end else if (10'h22a == _T_31[9:0]) begin
        image_1_554 <= io_pixelVal_in_1_5;
      end else if (10'h22a == _T_28[9:0]) begin
        image_1_554 <= io_pixelVal_in_1_4;
      end else if (10'h22a == _T_25[9:0]) begin
        image_1_554 <= io_pixelVal_in_1_3;
      end else if (10'h22a == _T_22[9:0]) begin
        image_1_554 <= io_pixelVal_in_1_2;
      end else if (10'h22a == _T_19[9:0]) begin
        image_1_554 <= io_pixelVal_in_1_1;
      end else if (10'h22a == _T_15[9:0]) begin
        image_1_554 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_555 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22b == _T_37[9:0]) begin
        image_1_555 <= io_pixelVal_in_1_7;
      end else if (10'h22b == _T_34[9:0]) begin
        image_1_555 <= io_pixelVal_in_1_6;
      end else if (10'h22b == _T_31[9:0]) begin
        image_1_555 <= io_pixelVal_in_1_5;
      end else if (10'h22b == _T_28[9:0]) begin
        image_1_555 <= io_pixelVal_in_1_4;
      end else if (10'h22b == _T_25[9:0]) begin
        image_1_555 <= io_pixelVal_in_1_3;
      end else if (10'h22b == _T_22[9:0]) begin
        image_1_555 <= io_pixelVal_in_1_2;
      end else if (10'h22b == _T_19[9:0]) begin
        image_1_555 <= io_pixelVal_in_1_1;
      end else if (10'h22b == _T_15[9:0]) begin
        image_1_555 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_556 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22c == _T_37[9:0]) begin
        image_1_556 <= io_pixelVal_in_1_7;
      end else if (10'h22c == _T_34[9:0]) begin
        image_1_556 <= io_pixelVal_in_1_6;
      end else if (10'h22c == _T_31[9:0]) begin
        image_1_556 <= io_pixelVal_in_1_5;
      end else if (10'h22c == _T_28[9:0]) begin
        image_1_556 <= io_pixelVal_in_1_4;
      end else if (10'h22c == _T_25[9:0]) begin
        image_1_556 <= io_pixelVal_in_1_3;
      end else if (10'h22c == _T_22[9:0]) begin
        image_1_556 <= io_pixelVal_in_1_2;
      end else if (10'h22c == _T_19[9:0]) begin
        image_1_556 <= io_pixelVal_in_1_1;
      end else if (10'h22c == _T_15[9:0]) begin
        image_1_556 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_557 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22d == _T_37[9:0]) begin
        image_1_557 <= io_pixelVal_in_1_7;
      end else if (10'h22d == _T_34[9:0]) begin
        image_1_557 <= io_pixelVal_in_1_6;
      end else if (10'h22d == _T_31[9:0]) begin
        image_1_557 <= io_pixelVal_in_1_5;
      end else if (10'h22d == _T_28[9:0]) begin
        image_1_557 <= io_pixelVal_in_1_4;
      end else if (10'h22d == _T_25[9:0]) begin
        image_1_557 <= io_pixelVal_in_1_3;
      end else if (10'h22d == _T_22[9:0]) begin
        image_1_557 <= io_pixelVal_in_1_2;
      end else if (10'h22d == _T_19[9:0]) begin
        image_1_557 <= io_pixelVal_in_1_1;
      end else if (10'h22d == _T_15[9:0]) begin
        image_1_557 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_558 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22e == _T_37[9:0]) begin
        image_1_558 <= io_pixelVal_in_1_7;
      end else if (10'h22e == _T_34[9:0]) begin
        image_1_558 <= io_pixelVal_in_1_6;
      end else if (10'h22e == _T_31[9:0]) begin
        image_1_558 <= io_pixelVal_in_1_5;
      end else if (10'h22e == _T_28[9:0]) begin
        image_1_558 <= io_pixelVal_in_1_4;
      end else if (10'h22e == _T_25[9:0]) begin
        image_1_558 <= io_pixelVal_in_1_3;
      end else if (10'h22e == _T_22[9:0]) begin
        image_1_558 <= io_pixelVal_in_1_2;
      end else if (10'h22e == _T_19[9:0]) begin
        image_1_558 <= io_pixelVal_in_1_1;
      end else if (10'h22e == _T_15[9:0]) begin
        image_1_558 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_559 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22f == _T_37[9:0]) begin
        image_1_559 <= io_pixelVal_in_1_7;
      end else if (10'h22f == _T_34[9:0]) begin
        image_1_559 <= io_pixelVal_in_1_6;
      end else if (10'h22f == _T_31[9:0]) begin
        image_1_559 <= io_pixelVal_in_1_5;
      end else if (10'h22f == _T_28[9:0]) begin
        image_1_559 <= io_pixelVal_in_1_4;
      end else if (10'h22f == _T_25[9:0]) begin
        image_1_559 <= io_pixelVal_in_1_3;
      end else if (10'h22f == _T_22[9:0]) begin
        image_1_559 <= io_pixelVal_in_1_2;
      end else if (10'h22f == _T_19[9:0]) begin
        image_1_559 <= io_pixelVal_in_1_1;
      end else if (10'h22f == _T_15[9:0]) begin
        image_1_559 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_560 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h230 == _T_37[9:0]) begin
        image_1_560 <= io_pixelVal_in_1_7;
      end else if (10'h230 == _T_34[9:0]) begin
        image_1_560 <= io_pixelVal_in_1_6;
      end else if (10'h230 == _T_31[9:0]) begin
        image_1_560 <= io_pixelVal_in_1_5;
      end else if (10'h230 == _T_28[9:0]) begin
        image_1_560 <= io_pixelVal_in_1_4;
      end else if (10'h230 == _T_25[9:0]) begin
        image_1_560 <= io_pixelVal_in_1_3;
      end else if (10'h230 == _T_22[9:0]) begin
        image_1_560 <= io_pixelVal_in_1_2;
      end else if (10'h230 == _T_19[9:0]) begin
        image_1_560 <= io_pixelVal_in_1_1;
      end else if (10'h230 == _T_15[9:0]) begin
        image_1_560 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_561 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h231 == _T_37[9:0]) begin
        image_1_561 <= io_pixelVal_in_1_7;
      end else if (10'h231 == _T_34[9:0]) begin
        image_1_561 <= io_pixelVal_in_1_6;
      end else if (10'h231 == _T_31[9:0]) begin
        image_1_561 <= io_pixelVal_in_1_5;
      end else if (10'h231 == _T_28[9:0]) begin
        image_1_561 <= io_pixelVal_in_1_4;
      end else if (10'h231 == _T_25[9:0]) begin
        image_1_561 <= io_pixelVal_in_1_3;
      end else if (10'h231 == _T_22[9:0]) begin
        image_1_561 <= io_pixelVal_in_1_2;
      end else if (10'h231 == _T_19[9:0]) begin
        image_1_561 <= io_pixelVal_in_1_1;
      end else if (10'h231 == _T_15[9:0]) begin
        image_1_561 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_562 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h232 == _T_37[9:0]) begin
        image_1_562 <= io_pixelVal_in_1_7;
      end else if (10'h232 == _T_34[9:0]) begin
        image_1_562 <= io_pixelVal_in_1_6;
      end else if (10'h232 == _T_31[9:0]) begin
        image_1_562 <= io_pixelVal_in_1_5;
      end else if (10'h232 == _T_28[9:0]) begin
        image_1_562 <= io_pixelVal_in_1_4;
      end else if (10'h232 == _T_25[9:0]) begin
        image_1_562 <= io_pixelVal_in_1_3;
      end else if (10'h232 == _T_22[9:0]) begin
        image_1_562 <= io_pixelVal_in_1_2;
      end else if (10'h232 == _T_19[9:0]) begin
        image_1_562 <= io_pixelVal_in_1_1;
      end else if (10'h232 == _T_15[9:0]) begin
        image_1_562 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_563 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h233 == _T_37[9:0]) begin
        image_1_563 <= io_pixelVal_in_1_7;
      end else if (10'h233 == _T_34[9:0]) begin
        image_1_563 <= io_pixelVal_in_1_6;
      end else if (10'h233 == _T_31[9:0]) begin
        image_1_563 <= io_pixelVal_in_1_5;
      end else if (10'h233 == _T_28[9:0]) begin
        image_1_563 <= io_pixelVal_in_1_4;
      end else if (10'h233 == _T_25[9:0]) begin
        image_1_563 <= io_pixelVal_in_1_3;
      end else if (10'h233 == _T_22[9:0]) begin
        image_1_563 <= io_pixelVal_in_1_2;
      end else if (10'h233 == _T_19[9:0]) begin
        image_1_563 <= io_pixelVal_in_1_1;
      end else if (10'h233 == _T_15[9:0]) begin
        image_1_563 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_564 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h234 == _T_37[9:0]) begin
        image_1_564 <= io_pixelVal_in_1_7;
      end else if (10'h234 == _T_34[9:0]) begin
        image_1_564 <= io_pixelVal_in_1_6;
      end else if (10'h234 == _T_31[9:0]) begin
        image_1_564 <= io_pixelVal_in_1_5;
      end else if (10'h234 == _T_28[9:0]) begin
        image_1_564 <= io_pixelVal_in_1_4;
      end else if (10'h234 == _T_25[9:0]) begin
        image_1_564 <= io_pixelVal_in_1_3;
      end else if (10'h234 == _T_22[9:0]) begin
        image_1_564 <= io_pixelVal_in_1_2;
      end else if (10'h234 == _T_19[9:0]) begin
        image_1_564 <= io_pixelVal_in_1_1;
      end else if (10'h234 == _T_15[9:0]) begin
        image_1_564 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_565 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h235 == _T_37[9:0]) begin
        image_1_565 <= io_pixelVal_in_1_7;
      end else if (10'h235 == _T_34[9:0]) begin
        image_1_565 <= io_pixelVal_in_1_6;
      end else if (10'h235 == _T_31[9:0]) begin
        image_1_565 <= io_pixelVal_in_1_5;
      end else if (10'h235 == _T_28[9:0]) begin
        image_1_565 <= io_pixelVal_in_1_4;
      end else if (10'h235 == _T_25[9:0]) begin
        image_1_565 <= io_pixelVal_in_1_3;
      end else if (10'h235 == _T_22[9:0]) begin
        image_1_565 <= io_pixelVal_in_1_2;
      end else if (10'h235 == _T_19[9:0]) begin
        image_1_565 <= io_pixelVal_in_1_1;
      end else if (10'h235 == _T_15[9:0]) begin
        image_1_565 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_566 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h236 == _T_37[9:0]) begin
        image_1_566 <= io_pixelVal_in_1_7;
      end else if (10'h236 == _T_34[9:0]) begin
        image_1_566 <= io_pixelVal_in_1_6;
      end else if (10'h236 == _T_31[9:0]) begin
        image_1_566 <= io_pixelVal_in_1_5;
      end else if (10'h236 == _T_28[9:0]) begin
        image_1_566 <= io_pixelVal_in_1_4;
      end else if (10'h236 == _T_25[9:0]) begin
        image_1_566 <= io_pixelVal_in_1_3;
      end else if (10'h236 == _T_22[9:0]) begin
        image_1_566 <= io_pixelVal_in_1_2;
      end else if (10'h236 == _T_19[9:0]) begin
        image_1_566 <= io_pixelVal_in_1_1;
      end else if (10'h236 == _T_15[9:0]) begin
        image_1_566 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_567 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h237 == _T_37[9:0]) begin
        image_1_567 <= io_pixelVal_in_1_7;
      end else if (10'h237 == _T_34[9:0]) begin
        image_1_567 <= io_pixelVal_in_1_6;
      end else if (10'h237 == _T_31[9:0]) begin
        image_1_567 <= io_pixelVal_in_1_5;
      end else if (10'h237 == _T_28[9:0]) begin
        image_1_567 <= io_pixelVal_in_1_4;
      end else if (10'h237 == _T_25[9:0]) begin
        image_1_567 <= io_pixelVal_in_1_3;
      end else if (10'h237 == _T_22[9:0]) begin
        image_1_567 <= io_pixelVal_in_1_2;
      end else if (10'h237 == _T_19[9:0]) begin
        image_1_567 <= io_pixelVal_in_1_1;
      end else if (10'h237 == _T_15[9:0]) begin
        image_1_567 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_568 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h238 == _T_37[9:0]) begin
        image_1_568 <= io_pixelVal_in_1_7;
      end else if (10'h238 == _T_34[9:0]) begin
        image_1_568 <= io_pixelVal_in_1_6;
      end else if (10'h238 == _T_31[9:0]) begin
        image_1_568 <= io_pixelVal_in_1_5;
      end else if (10'h238 == _T_28[9:0]) begin
        image_1_568 <= io_pixelVal_in_1_4;
      end else if (10'h238 == _T_25[9:0]) begin
        image_1_568 <= io_pixelVal_in_1_3;
      end else if (10'h238 == _T_22[9:0]) begin
        image_1_568 <= io_pixelVal_in_1_2;
      end else if (10'h238 == _T_19[9:0]) begin
        image_1_568 <= io_pixelVal_in_1_1;
      end else if (10'h238 == _T_15[9:0]) begin
        image_1_568 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_569 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h239 == _T_37[9:0]) begin
        image_1_569 <= io_pixelVal_in_1_7;
      end else if (10'h239 == _T_34[9:0]) begin
        image_1_569 <= io_pixelVal_in_1_6;
      end else if (10'h239 == _T_31[9:0]) begin
        image_1_569 <= io_pixelVal_in_1_5;
      end else if (10'h239 == _T_28[9:0]) begin
        image_1_569 <= io_pixelVal_in_1_4;
      end else if (10'h239 == _T_25[9:0]) begin
        image_1_569 <= io_pixelVal_in_1_3;
      end else if (10'h239 == _T_22[9:0]) begin
        image_1_569 <= io_pixelVal_in_1_2;
      end else if (10'h239 == _T_19[9:0]) begin
        image_1_569 <= io_pixelVal_in_1_1;
      end else if (10'h239 == _T_15[9:0]) begin
        image_1_569 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_570 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23a == _T_37[9:0]) begin
        image_1_570 <= io_pixelVal_in_1_7;
      end else if (10'h23a == _T_34[9:0]) begin
        image_1_570 <= io_pixelVal_in_1_6;
      end else if (10'h23a == _T_31[9:0]) begin
        image_1_570 <= io_pixelVal_in_1_5;
      end else if (10'h23a == _T_28[9:0]) begin
        image_1_570 <= io_pixelVal_in_1_4;
      end else if (10'h23a == _T_25[9:0]) begin
        image_1_570 <= io_pixelVal_in_1_3;
      end else if (10'h23a == _T_22[9:0]) begin
        image_1_570 <= io_pixelVal_in_1_2;
      end else if (10'h23a == _T_19[9:0]) begin
        image_1_570 <= io_pixelVal_in_1_1;
      end else if (10'h23a == _T_15[9:0]) begin
        image_1_570 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_571 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23b == _T_37[9:0]) begin
        image_1_571 <= io_pixelVal_in_1_7;
      end else if (10'h23b == _T_34[9:0]) begin
        image_1_571 <= io_pixelVal_in_1_6;
      end else if (10'h23b == _T_31[9:0]) begin
        image_1_571 <= io_pixelVal_in_1_5;
      end else if (10'h23b == _T_28[9:0]) begin
        image_1_571 <= io_pixelVal_in_1_4;
      end else if (10'h23b == _T_25[9:0]) begin
        image_1_571 <= io_pixelVal_in_1_3;
      end else if (10'h23b == _T_22[9:0]) begin
        image_1_571 <= io_pixelVal_in_1_2;
      end else if (10'h23b == _T_19[9:0]) begin
        image_1_571 <= io_pixelVal_in_1_1;
      end else if (10'h23b == _T_15[9:0]) begin
        image_1_571 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_572 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23c == _T_37[9:0]) begin
        image_1_572 <= io_pixelVal_in_1_7;
      end else if (10'h23c == _T_34[9:0]) begin
        image_1_572 <= io_pixelVal_in_1_6;
      end else if (10'h23c == _T_31[9:0]) begin
        image_1_572 <= io_pixelVal_in_1_5;
      end else if (10'h23c == _T_28[9:0]) begin
        image_1_572 <= io_pixelVal_in_1_4;
      end else if (10'h23c == _T_25[9:0]) begin
        image_1_572 <= io_pixelVal_in_1_3;
      end else if (10'h23c == _T_22[9:0]) begin
        image_1_572 <= io_pixelVal_in_1_2;
      end else if (10'h23c == _T_19[9:0]) begin
        image_1_572 <= io_pixelVal_in_1_1;
      end else if (10'h23c == _T_15[9:0]) begin
        image_1_572 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_573 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23d == _T_37[9:0]) begin
        image_1_573 <= io_pixelVal_in_1_7;
      end else if (10'h23d == _T_34[9:0]) begin
        image_1_573 <= io_pixelVal_in_1_6;
      end else if (10'h23d == _T_31[9:0]) begin
        image_1_573 <= io_pixelVal_in_1_5;
      end else if (10'h23d == _T_28[9:0]) begin
        image_1_573 <= io_pixelVal_in_1_4;
      end else if (10'h23d == _T_25[9:0]) begin
        image_1_573 <= io_pixelVal_in_1_3;
      end else if (10'h23d == _T_22[9:0]) begin
        image_1_573 <= io_pixelVal_in_1_2;
      end else if (10'h23d == _T_19[9:0]) begin
        image_1_573 <= io_pixelVal_in_1_1;
      end else if (10'h23d == _T_15[9:0]) begin
        image_1_573 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_574 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23e == _T_37[9:0]) begin
        image_1_574 <= io_pixelVal_in_1_7;
      end else if (10'h23e == _T_34[9:0]) begin
        image_1_574 <= io_pixelVal_in_1_6;
      end else if (10'h23e == _T_31[9:0]) begin
        image_1_574 <= io_pixelVal_in_1_5;
      end else if (10'h23e == _T_28[9:0]) begin
        image_1_574 <= io_pixelVal_in_1_4;
      end else if (10'h23e == _T_25[9:0]) begin
        image_1_574 <= io_pixelVal_in_1_3;
      end else if (10'h23e == _T_22[9:0]) begin
        image_1_574 <= io_pixelVal_in_1_2;
      end else if (10'h23e == _T_19[9:0]) begin
        image_1_574 <= io_pixelVal_in_1_1;
      end else if (10'h23e == _T_15[9:0]) begin
        image_1_574 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_575 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23f == _T_37[9:0]) begin
        image_1_575 <= io_pixelVal_in_1_7;
      end else if (10'h23f == _T_34[9:0]) begin
        image_1_575 <= io_pixelVal_in_1_6;
      end else if (10'h23f == _T_31[9:0]) begin
        image_1_575 <= io_pixelVal_in_1_5;
      end else if (10'h23f == _T_28[9:0]) begin
        image_1_575 <= io_pixelVal_in_1_4;
      end else if (10'h23f == _T_25[9:0]) begin
        image_1_575 <= io_pixelVal_in_1_3;
      end else if (10'h23f == _T_22[9:0]) begin
        image_1_575 <= io_pixelVal_in_1_2;
      end else if (10'h23f == _T_19[9:0]) begin
        image_1_575 <= io_pixelVal_in_1_1;
      end else if (10'h23f == _T_15[9:0]) begin
        image_1_575 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_2_0 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h0 == _T_37[9:0]) begin
        image_2_0 <= io_pixelVal_in_2_7;
      end else if (10'h0 == _T_34[9:0]) begin
        image_2_0 <= io_pixelVal_in_2_6;
      end else if (10'h0 == _T_31[9:0]) begin
        image_2_0 <= io_pixelVal_in_2_5;
      end else if (10'h0 == _T_28[9:0]) begin
        image_2_0 <= io_pixelVal_in_2_4;
      end else if (10'h0 == _T_25[9:0]) begin
        image_2_0 <= io_pixelVal_in_2_3;
      end else if (10'h0 == _T_22[9:0]) begin
        image_2_0 <= io_pixelVal_in_2_2;
      end else if (10'h0 == _T_19[9:0]) begin
        image_2_0 <= io_pixelVal_in_2_1;
      end else if (10'h0 == _T_15[9:0]) begin
        image_2_0 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_1 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1 == _T_37[9:0]) begin
        image_2_1 <= io_pixelVal_in_2_7;
      end else if (10'h1 == _T_34[9:0]) begin
        image_2_1 <= io_pixelVal_in_2_6;
      end else if (10'h1 == _T_31[9:0]) begin
        image_2_1 <= io_pixelVal_in_2_5;
      end else if (10'h1 == _T_28[9:0]) begin
        image_2_1 <= io_pixelVal_in_2_4;
      end else if (10'h1 == _T_25[9:0]) begin
        image_2_1 <= io_pixelVal_in_2_3;
      end else if (10'h1 == _T_22[9:0]) begin
        image_2_1 <= io_pixelVal_in_2_2;
      end else if (10'h1 == _T_19[9:0]) begin
        image_2_1 <= io_pixelVal_in_2_1;
      end else if (10'h1 == _T_15[9:0]) begin
        image_2_1 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_2 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2 == _T_37[9:0]) begin
        image_2_2 <= io_pixelVal_in_2_7;
      end else if (10'h2 == _T_34[9:0]) begin
        image_2_2 <= io_pixelVal_in_2_6;
      end else if (10'h2 == _T_31[9:0]) begin
        image_2_2 <= io_pixelVal_in_2_5;
      end else if (10'h2 == _T_28[9:0]) begin
        image_2_2 <= io_pixelVal_in_2_4;
      end else if (10'h2 == _T_25[9:0]) begin
        image_2_2 <= io_pixelVal_in_2_3;
      end else if (10'h2 == _T_22[9:0]) begin
        image_2_2 <= io_pixelVal_in_2_2;
      end else if (10'h2 == _T_19[9:0]) begin
        image_2_2 <= io_pixelVal_in_2_1;
      end else if (10'h2 == _T_15[9:0]) begin
        image_2_2 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_3 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3 == _T_37[9:0]) begin
        image_2_3 <= io_pixelVal_in_2_7;
      end else if (10'h3 == _T_34[9:0]) begin
        image_2_3 <= io_pixelVal_in_2_6;
      end else if (10'h3 == _T_31[9:0]) begin
        image_2_3 <= io_pixelVal_in_2_5;
      end else if (10'h3 == _T_28[9:0]) begin
        image_2_3 <= io_pixelVal_in_2_4;
      end else if (10'h3 == _T_25[9:0]) begin
        image_2_3 <= io_pixelVal_in_2_3;
      end else if (10'h3 == _T_22[9:0]) begin
        image_2_3 <= io_pixelVal_in_2_2;
      end else if (10'h3 == _T_19[9:0]) begin
        image_2_3 <= io_pixelVal_in_2_1;
      end else if (10'h3 == _T_15[9:0]) begin
        image_2_3 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_4 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4 == _T_37[9:0]) begin
        image_2_4 <= io_pixelVal_in_2_7;
      end else if (10'h4 == _T_34[9:0]) begin
        image_2_4 <= io_pixelVal_in_2_6;
      end else if (10'h4 == _T_31[9:0]) begin
        image_2_4 <= io_pixelVal_in_2_5;
      end else if (10'h4 == _T_28[9:0]) begin
        image_2_4 <= io_pixelVal_in_2_4;
      end else if (10'h4 == _T_25[9:0]) begin
        image_2_4 <= io_pixelVal_in_2_3;
      end else if (10'h4 == _T_22[9:0]) begin
        image_2_4 <= io_pixelVal_in_2_2;
      end else if (10'h4 == _T_19[9:0]) begin
        image_2_4 <= io_pixelVal_in_2_1;
      end else if (10'h4 == _T_15[9:0]) begin
        image_2_4 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_5 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5 == _T_37[9:0]) begin
        image_2_5 <= io_pixelVal_in_2_7;
      end else if (10'h5 == _T_34[9:0]) begin
        image_2_5 <= io_pixelVal_in_2_6;
      end else if (10'h5 == _T_31[9:0]) begin
        image_2_5 <= io_pixelVal_in_2_5;
      end else if (10'h5 == _T_28[9:0]) begin
        image_2_5 <= io_pixelVal_in_2_4;
      end else if (10'h5 == _T_25[9:0]) begin
        image_2_5 <= io_pixelVal_in_2_3;
      end else if (10'h5 == _T_22[9:0]) begin
        image_2_5 <= io_pixelVal_in_2_2;
      end else if (10'h5 == _T_19[9:0]) begin
        image_2_5 <= io_pixelVal_in_2_1;
      end else if (10'h5 == _T_15[9:0]) begin
        image_2_5 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_6 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6 == _T_37[9:0]) begin
        image_2_6 <= io_pixelVal_in_2_7;
      end else if (10'h6 == _T_34[9:0]) begin
        image_2_6 <= io_pixelVal_in_2_6;
      end else if (10'h6 == _T_31[9:0]) begin
        image_2_6 <= io_pixelVal_in_2_5;
      end else if (10'h6 == _T_28[9:0]) begin
        image_2_6 <= io_pixelVal_in_2_4;
      end else if (10'h6 == _T_25[9:0]) begin
        image_2_6 <= io_pixelVal_in_2_3;
      end else if (10'h6 == _T_22[9:0]) begin
        image_2_6 <= io_pixelVal_in_2_2;
      end else if (10'h6 == _T_19[9:0]) begin
        image_2_6 <= io_pixelVal_in_2_1;
      end else if (10'h6 == _T_15[9:0]) begin
        image_2_6 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_7 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7 == _T_37[9:0]) begin
        image_2_7 <= io_pixelVal_in_2_7;
      end else if (10'h7 == _T_34[9:0]) begin
        image_2_7 <= io_pixelVal_in_2_6;
      end else if (10'h7 == _T_31[9:0]) begin
        image_2_7 <= io_pixelVal_in_2_5;
      end else if (10'h7 == _T_28[9:0]) begin
        image_2_7 <= io_pixelVal_in_2_4;
      end else if (10'h7 == _T_25[9:0]) begin
        image_2_7 <= io_pixelVal_in_2_3;
      end else if (10'h7 == _T_22[9:0]) begin
        image_2_7 <= io_pixelVal_in_2_2;
      end else if (10'h7 == _T_19[9:0]) begin
        image_2_7 <= io_pixelVal_in_2_1;
      end else if (10'h7 == _T_15[9:0]) begin
        image_2_7 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_8 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8 == _T_37[9:0]) begin
        image_2_8 <= io_pixelVal_in_2_7;
      end else if (10'h8 == _T_34[9:0]) begin
        image_2_8 <= io_pixelVal_in_2_6;
      end else if (10'h8 == _T_31[9:0]) begin
        image_2_8 <= io_pixelVal_in_2_5;
      end else if (10'h8 == _T_28[9:0]) begin
        image_2_8 <= io_pixelVal_in_2_4;
      end else if (10'h8 == _T_25[9:0]) begin
        image_2_8 <= io_pixelVal_in_2_3;
      end else if (10'h8 == _T_22[9:0]) begin
        image_2_8 <= io_pixelVal_in_2_2;
      end else if (10'h8 == _T_19[9:0]) begin
        image_2_8 <= io_pixelVal_in_2_1;
      end else if (10'h8 == _T_15[9:0]) begin
        image_2_8 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_9 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9 == _T_37[9:0]) begin
        image_2_9 <= io_pixelVal_in_2_7;
      end else if (10'h9 == _T_34[9:0]) begin
        image_2_9 <= io_pixelVal_in_2_6;
      end else if (10'h9 == _T_31[9:0]) begin
        image_2_9 <= io_pixelVal_in_2_5;
      end else if (10'h9 == _T_28[9:0]) begin
        image_2_9 <= io_pixelVal_in_2_4;
      end else if (10'h9 == _T_25[9:0]) begin
        image_2_9 <= io_pixelVal_in_2_3;
      end else if (10'h9 == _T_22[9:0]) begin
        image_2_9 <= io_pixelVal_in_2_2;
      end else if (10'h9 == _T_19[9:0]) begin
        image_2_9 <= io_pixelVal_in_2_1;
      end else if (10'h9 == _T_15[9:0]) begin
        image_2_9 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_10 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha == _T_37[9:0]) begin
        image_2_10 <= io_pixelVal_in_2_7;
      end else if (10'ha == _T_34[9:0]) begin
        image_2_10 <= io_pixelVal_in_2_6;
      end else if (10'ha == _T_31[9:0]) begin
        image_2_10 <= io_pixelVal_in_2_5;
      end else if (10'ha == _T_28[9:0]) begin
        image_2_10 <= io_pixelVal_in_2_4;
      end else if (10'ha == _T_25[9:0]) begin
        image_2_10 <= io_pixelVal_in_2_3;
      end else if (10'ha == _T_22[9:0]) begin
        image_2_10 <= io_pixelVal_in_2_2;
      end else if (10'ha == _T_19[9:0]) begin
        image_2_10 <= io_pixelVal_in_2_1;
      end else if (10'ha == _T_15[9:0]) begin
        image_2_10 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_11 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb == _T_37[9:0]) begin
        image_2_11 <= io_pixelVal_in_2_7;
      end else if (10'hb == _T_34[9:0]) begin
        image_2_11 <= io_pixelVal_in_2_6;
      end else if (10'hb == _T_31[9:0]) begin
        image_2_11 <= io_pixelVal_in_2_5;
      end else if (10'hb == _T_28[9:0]) begin
        image_2_11 <= io_pixelVal_in_2_4;
      end else if (10'hb == _T_25[9:0]) begin
        image_2_11 <= io_pixelVal_in_2_3;
      end else if (10'hb == _T_22[9:0]) begin
        image_2_11 <= io_pixelVal_in_2_2;
      end else if (10'hb == _T_19[9:0]) begin
        image_2_11 <= io_pixelVal_in_2_1;
      end else if (10'hb == _T_15[9:0]) begin
        image_2_11 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_12 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc == _T_37[9:0]) begin
        image_2_12 <= io_pixelVal_in_2_7;
      end else if (10'hc == _T_34[9:0]) begin
        image_2_12 <= io_pixelVal_in_2_6;
      end else if (10'hc == _T_31[9:0]) begin
        image_2_12 <= io_pixelVal_in_2_5;
      end else if (10'hc == _T_28[9:0]) begin
        image_2_12 <= io_pixelVal_in_2_4;
      end else if (10'hc == _T_25[9:0]) begin
        image_2_12 <= io_pixelVal_in_2_3;
      end else if (10'hc == _T_22[9:0]) begin
        image_2_12 <= io_pixelVal_in_2_2;
      end else if (10'hc == _T_19[9:0]) begin
        image_2_12 <= io_pixelVal_in_2_1;
      end else if (10'hc == _T_15[9:0]) begin
        image_2_12 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_13 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd == _T_37[9:0]) begin
        image_2_13 <= io_pixelVal_in_2_7;
      end else if (10'hd == _T_34[9:0]) begin
        image_2_13 <= io_pixelVal_in_2_6;
      end else if (10'hd == _T_31[9:0]) begin
        image_2_13 <= io_pixelVal_in_2_5;
      end else if (10'hd == _T_28[9:0]) begin
        image_2_13 <= io_pixelVal_in_2_4;
      end else if (10'hd == _T_25[9:0]) begin
        image_2_13 <= io_pixelVal_in_2_3;
      end else if (10'hd == _T_22[9:0]) begin
        image_2_13 <= io_pixelVal_in_2_2;
      end else if (10'hd == _T_19[9:0]) begin
        image_2_13 <= io_pixelVal_in_2_1;
      end else if (10'hd == _T_15[9:0]) begin
        image_2_13 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_14 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he == _T_37[9:0]) begin
        image_2_14 <= io_pixelVal_in_2_7;
      end else if (10'he == _T_34[9:0]) begin
        image_2_14 <= io_pixelVal_in_2_6;
      end else if (10'he == _T_31[9:0]) begin
        image_2_14 <= io_pixelVal_in_2_5;
      end else if (10'he == _T_28[9:0]) begin
        image_2_14 <= io_pixelVal_in_2_4;
      end else if (10'he == _T_25[9:0]) begin
        image_2_14 <= io_pixelVal_in_2_3;
      end else if (10'he == _T_22[9:0]) begin
        image_2_14 <= io_pixelVal_in_2_2;
      end else if (10'he == _T_19[9:0]) begin
        image_2_14 <= io_pixelVal_in_2_1;
      end else if (10'he == _T_15[9:0]) begin
        image_2_14 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_15 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf == _T_37[9:0]) begin
        image_2_15 <= io_pixelVal_in_2_7;
      end else if (10'hf == _T_34[9:0]) begin
        image_2_15 <= io_pixelVal_in_2_6;
      end else if (10'hf == _T_31[9:0]) begin
        image_2_15 <= io_pixelVal_in_2_5;
      end else if (10'hf == _T_28[9:0]) begin
        image_2_15 <= io_pixelVal_in_2_4;
      end else if (10'hf == _T_25[9:0]) begin
        image_2_15 <= io_pixelVal_in_2_3;
      end else if (10'hf == _T_22[9:0]) begin
        image_2_15 <= io_pixelVal_in_2_2;
      end else if (10'hf == _T_19[9:0]) begin
        image_2_15 <= io_pixelVal_in_2_1;
      end else if (10'hf == _T_15[9:0]) begin
        image_2_15 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_16 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10 == _T_37[9:0]) begin
        image_2_16 <= io_pixelVal_in_2_7;
      end else if (10'h10 == _T_34[9:0]) begin
        image_2_16 <= io_pixelVal_in_2_6;
      end else if (10'h10 == _T_31[9:0]) begin
        image_2_16 <= io_pixelVal_in_2_5;
      end else if (10'h10 == _T_28[9:0]) begin
        image_2_16 <= io_pixelVal_in_2_4;
      end else if (10'h10 == _T_25[9:0]) begin
        image_2_16 <= io_pixelVal_in_2_3;
      end else if (10'h10 == _T_22[9:0]) begin
        image_2_16 <= io_pixelVal_in_2_2;
      end else if (10'h10 == _T_19[9:0]) begin
        image_2_16 <= io_pixelVal_in_2_1;
      end else if (10'h10 == _T_15[9:0]) begin
        image_2_16 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_17 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11 == _T_37[9:0]) begin
        image_2_17 <= io_pixelVal_in_2_7;
      end else if (10'h11 == _T_34[9:0]) begin
        image_2_17 <= io_pixelVal_in_2_6;
      end else if (10'h11 == _T_31[9:0]) begin
        image_2_17 <= io_pixelVal_in_2_5;
      end else if (10'h11 == _T_28[9:0]) begin
        image_2_17 <= io_pixelVal_in_2_4;
      end else if (10'h11 == _T_25[9:0]) begin
        image_2_17 <= io_pixelVal_in_2_3;
      end else if (10'h11 == _T_22[9:0]) begin
        image_2_17 <= io_pixelVal_in_2_2;
      end else if (10'h11 == _T_19[9:0]) begin
        image_2_17 <= io_pixelVal_in_2_1;
      end else if (10'h11 == _T_15[9:0]) begin
        image_2_17 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_18 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12 == _T_37[9:0]) begin
        image_2_18 <= io_pixelVal_in_2_7;
      end else if (10'h12 == _T_34[9:0]) begin
        image_2_18 <= io_pixelVal_in_2_6;
      end else if (10'h12 == _T_31[9:0]) begin
        image_2_18 <= io_pixelVal_in_2_5;
      end else if (10'h12 == _T_28[9:0]) begin
        image_2_18 <= io_pixelVal_in_2_4;
      end else if (10'h12 == _T_25[9:0]) begin
        image_2_18 <= io_pixelVal_in_2_3;
      end else if (10'h12 == _T_22[9:0]) begin
        image_2_18 <= io_pixelVal_in_2_2;
      end else if (10'h12 == _T_19[9:0]) begin
        image_2_18 <= io_pixelVal_in_2_1;
      end else if (10'h12 == _T_15[9:0]) begin
        image_2_18 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_19 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13 == _T_37[9:0]) begin
        image_2_19 <= io_pixelVal_in_2_7;
      end else if (10'h13 == _T_34[9:0]) begin
        image_2_19 <= io_pixelVal_in_2_6;
      end else if (10'h13 == _T_31[9:0]) begin
        image_2_19 <= io_pixelVal_in_2_5;
      end else if (10'h13 == _T_28[9:0]) begin
        image_2_19 <= io_pixelVal_in_2_4;
      end else if (10'h13 == _T_25[9:0]) begin
        image_2_19 <= io_pixelVal_in_2_3;
      end else if (10'h13 == _T_22[9:0]) begin
        image_2_19 <= io_pixelVal_in_2_2;
      end else if (10'h13 == _T_19[9:0]) begin
        image_2_19 <= io_pixelVal_in_2_1;
      end else if (10'h13 == _T_15[9:0]) begin
        image_2_19 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_20 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14 == _T_37[9:0]) begin
        image_2_20 <= io_pixelVal_in_2_7;
      end else if (10'h14 == _T_34[9:0]) begin
        image_2_20 <= io_pixelVal_in_2_6;
      end else if (10'h14 == _T_31[9:0]) begin
        image_2_20 <= io_pixelVal_in_2_5;
      end else if (10'h14 == _T_28[9:0]) begin
        image_2_20 <= io_pixelVal_in_2_4;
      end else if (10'h14 == _T_25[9:0]) begin
        image_2_20 <= io_pixelVal_in_2_3;
      end else if (10'h14 == _T_22[9:0]) begin
        image_2_20 <= io_pixelVal_in_2_2;
      end else if (10'h14 == _T_19[9:0]) begin
        image_2_20 <= io_pixelVal_in_2_1;
      end else if (10'h14 == _T_15[9:0]) begin
        image_2_20 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_21 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15 == _T_37[9:0]) begin
        image_2_21 <= io_pixelVal_in_2_7;
      end else if (10'h15 == _T_34[9:0]) begin
        image_2_21 <= io_pixelVal_in_2_6;
      end else if (10'h15 == _T_31[9:0]) begin
        image_2_21 <= io_pixelVal_in_2_5;
      end else if (10'h15 == _T_28[9:0]) begin
        image_2_21 <= io_pixelVal_in_2_4;
      end else if (10'h15 == _T_25[9:0]) begin
        image_2_21 <= io_pixelVal_in_2_3;
      end else if (10'h15 == _T_22[9:0]) begin
        image_2_21 <= io_pixelVal_in_2_2;
      end else if (10'h15 == _T_19[9:0]) begin
        image_2_21 <= io_pixelVal_in_2_1;
      end else if (10'h15 == _T_15[9:0]) begin
        image_2_21 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_22 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16 == _T_37[9:0]) begin
        image_2_22 <= io_pixelVal_in_2_7;
      end else if (10'h16 == _T_34[9:0]) begin
        image_2_22 <= io_pixelVal_in_2_6;
      end else if (10'h16 == _T_31[9:0]) begin
        image_2_22 <= io_pixelVal_in_2_5;
      end else if (10'h16 == _T_28[9:0]) begin
        image_2_22 <= io_pixelVal_in_2_4;
      end else if (10'h16 == _T_25[9:0]) begin
        image_2_22 <= io_pixelVal_in_2_3;
      end else if (10'h16 == _T_22[9:0]) begin
        image_2_22 <= io_pixelVal_in_2_2;
      end else if (10'h16 == _T_19[9:0]) begin
        image_2_22 <= io_pixelVal_in_2_1;
      end else if (10'h16 == _T_15[9:0]) begin
        image_2_22 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_23 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17 == _T_37[9:0]) begin
        image_2_23 <= io_pixelVal_in_2_7;
      end else if (10'h17 == _T_34[9:0]) begin
        image_2_23 <= io_pixelVal_in_2_6;
      end else if (10'h17 == _T_31[9:0]) begin
        image_2_23 <= io_pixelVal_in_2_5;
      end else if (10'h17 == _T_28[9:0]) begin
        image_2_23 <= io_pixelVal_in_2_4;
      end else if (10'h17 == _T_25[9:0]) begin
        image_2_23 <= io_pixelVal_in_2_3;
      end else if (10'h17 == _T_22[9:0]) begin
        image_2_23 <= io_pixelVal_in_2_2;
      end else if (10'h17 == _T_19[9:0]) begin
        image_2_23 <= io_pixelVal_in_2_1;
      end else if (10'h17 == _T_15[9:0]) begin
        image_2_23 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_24 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18 == _T_37[9:0]) begin
        image_2_24 <= io_pixelVal_in_2_7;
      end else if (10'h18 == _T_34[9:0]) begin
        image_2_24 <= io_pixelVal_in_2_6;
      end else if (10'h18 == _T_31[9:0]) begin
        image_2_24 <= io_pixelVal_in_2_5;
      end else if (10'h18 == _T_28[9:0]) begin
        image_2_24 <= io_pixelVal_in_2_4;
      end else if (10'h18 == _T_25[9:0]) begin
        image_2_24 <= io_pixelVal_in_2_3;
      end else if (10'h18 == _T_22[9:0]) begin
        image_2_24 <= io_pixelVal_in_2_2;
      end else if (10'h18 == _T_19[9:0]) begin
        image_2_24 <= io_pixelVal_in_2_1;
      end else if (10'h18 == _T_15[9:0]) begin
        image_2_24 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_25 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19 == _T_37[9:0]) begin
        image_2_25 <= io_pixelVal_in_2_7;
      end else if (10'h19 == _T_34[9:0]) begin
        image_2_25 <= io_pixelVal_in_2_6;
      end else if (10'h19 == _T_31[9:0]) begin
        image_2_25 <= io_pixelVal_in_2_5;
      end else if (10'h19 == _T_28[9:0]) begin
        image_2_25 <= io_pixelVal_in_2_4;
      end else if (10'h19 == _T_25[9:0]) begin
        image_2_25 <= io_pixelVal_in_2_3;
      end else if (10'h19 == _T_22[9:0]) begin
        image_2_25 <= io_pixelVal_in_2_2;
      end else if (10'h19 == _T_19[9:0]) begin
        image_2_25 <= io_pixelVal_in_2_1;
      end else if (10'h19 == _T_15[9:0]) begin
        image_2_25 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_26 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a == _T_37[9:0]) begin
        image_2_26 <= io_pixelVal_in_2_7;
      end else if (10'h1a == _T_34[9:0]) begin
        image_2_26 <= io_pixelVal_in_2_6;
      end else if (10'h1a == _T_31[9:0]) begin
        image_2_26 <= io_pixelVal_in_2_5;
      end else if (10'h1a == _T_28[9:0]) begin
        image_2_26 <= io_pixelVal_in_2_4;
      end else if (10'h1a == _T_25[9:0]) begin
        image_2_26 <= io_pixelVal_in_2_3;
      end else if (10'h1a == _T_22[9:0]) begin
        image_2_26 <= io_pixelVal_in_2_2;
      end else if (10'h1a == _T_19[9:0]) begin
        image_2_26 <= io_pixelVal_in_2_1;
      end else if (10'h1a == _T_15[9:0]) begin
        image_2_26 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_27 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b == _T_37[9:0]) begin
        image_2_27 <= io_pixelVal_in_2_7;
      end else if (10'h1b == _T_34[9:0]) begin
        image_2_27 <= io_pixelVal_in_2_6;
      end else if (10'h1b == _T_31[9:0]) begin
        image_2_27 <= io_pixelVal_in_2_5;
      end else if (10'h1b == _T_28[9:0]) begin
        image_2_27 <= io_pixelVal_in_2_4;
      end else if (10'h1b == _T_25[9:0]) begin
        image_2_27 <= io_pixelVal_in_2_3;
      end else if (10'h1b == _T_22[9:0]) begin
        image_2_27 <= io_pixelVal_in_2_2;
      end else if (10'h1b == _T_19[9:0]) begin
        image_2_27 <= io_pixelVal_in_2_1;
      end else if (10'h1b == _T_15[9:0]) begin
        image_2_27 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_28 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c == _T_37[9:0]) begin
        image_2_28 <= io_pixelVal_in_2_7;
      end else if (10'h1c == _T_34[9:0]) begin
        image_2_28 <= io_pixelVal_in_2_6;
      end else if (10'h1c == _T_31[9:0]) begin
        image_2_28 <= io_pixelVal_in_2_5;
      end else if (10'h1c == _T_28[9:0]) begin
        image_2_28 <= io_pixelVal_in_2_4;
      end else if (10'h1c == _T_25[9:0]) begin
        image_2_28 <= io_pixelVal_in_2_3;
      end else if (10'h1c == _T_22[9:0]) begin
        image_2_28 <= io_pixelVal_in_2_2;
      end else if (10'h1c == _T_19[9:0]) begin
        image_2_28 <= io_pixelVal_in_2_1;
      end else if (10'h1c == _T_15[9:0]) begin
        image_2_28 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_29 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d == _T_37[9:0]) begin
        image_2_29 <= io_pixelVal_in_2_7;
      end else if (10'h1d == _T_34[9:0]) begin
        image_2_29 <= io_pixelVal_in_2_6;
      end else if (10'h1d == _T_31[9:0]) begin
        image_2_29 <= io_pixelVal_in_2_5;
      end else if (10'h1d == _T_28[9:0]) begin
        image_2_29 <= io_pixelVal_in_2_4;
      end else if (10'h1d == _T_25[9:0]) begin
        image_2_29 <= io_pixelVal_in_2_3;
      end else if (10'h1d == _T_22[9:0]) begin
        image_2_29 <= io_pixelVal_in_2_2;
      end else if (10'h1d == _T_19[9:0]) begin
        image_2_29 <= io_pixelVal_in_2_1;
      end else if (10'h1d == _T_15[9:0]) begin
        image_2_29 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_30 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e == _T_37[9:0]) begin
        image_2_30 <= io_pixelVal_in_2_7;
      end else if (10'h1e == _T_34[9:0]) begin
        image_2_30 <= io_pixelVal_in_2_6;
      end else if (10'h1e == _T_31[9:0]) begin
        image_2_30 <= io_pixelVal_in_2_5;
      end else if (10'h1e == _T_28[9:0]) begin
        image_2_30 <= io_pixelVal_in_2_4;
      end else if (10'h1e == _T_25[9:0]) begin
        image_2_30 <= io_pixelVal_in_2_3;
      end else if (10'h1e == _T_22[9:0]) begin
        image_2_30 <= io_pixelVal_in_2_2;
      end else if (10'h1e == _T_19[9:0]) begin
        image_2_30 <= io_pixelVal_in_2_1;
      end else if (10'h1e == _T_15[9:0]) begin
        image_2_30 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_31 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f == _T_37[9:0]) begin
        image_2_31 <= io_pixelVal_in_2_7;
      end else if (10'h1f == _T_34[9:0]) begin
        image_2_31 <= io_pixelVal_in_2_6;
      end else if (10'h1f == _T_31[9:0]) begin
        image_2_31 <= io_pixelVal_in_2_5;
      end else if (10'h1f == _T_28[9:0]) begin
        image_2_31 <= io_pixelVal_in_2_4;
      end else if (10'h1f == _T_25[9:0]) begin
        image_2_31 <= io_pixelVal_in_2_3;
      end else if (10'h1f == _T_22[9:0]) begin
        image_2_31 <= io_pixelVal_in_2_2;
      end else if (10'h1f == _T_19[9:0]) begin
        image_2_31 <= io_pixelVal_in_2_1;
      end else if (10'h1f == _T_15[9:0]) begin
        image_2_31 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_32 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20 == _T_37[9:0]) begin
        image_2_32 <= io_pixelVal_in_2_7;
      end else if (10'h20 == _T_34[9:0]) begin
        image_2_32 <= io_pixelVal_in_2_6;
      end else if (10'h20 == _T_31[9:0]) begin
        image_2_32 <= io_pixelVal_in_2_5;
      end else if (10'h20 == _T_28[9:0]) begin
        image_2_32 <= io_pixelVal_in_2_4;
      end else if (10'h20 == _T_25[9:0]) begin
        image_2_32 <= io_pixelVal_in_2_3;
      end else if (10'h20 == _T_22[9:0]) begin
        image_2_32 <= io_pixelVal_in_2_2;
      end else if (10'h20 == _T_19[9:0]) begin
        image_2_32 <= io_pixelVal_in_2_1;
      end else if (10'h20 == _T_15[9:0]) begin
        image_2_32 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_33 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21 == _T_37[9:0]) begin
        image_2_33 <= io_pixelVal_in_2_7;
      end else if (10'h21 == _T_34[9:0]) begin
        image_2_33 <= io_pixelVal_in_2_6;
      end else if (10'h21 == _T_31[9:0]) begin
        image_2_33 <= io_pixelVal_in_2_5;
      end else if (10'h21 == _T_28[9:0]) begin
        image_2_33 <= io_pixelVal_in_2_4;
      end else if (10'h21 == _T_25[9:0]) begin
        image_2_33 <= io_pixelVal_in_2_3;
      end else if (10'h21 == _T_22[9:0]) begin
        image_2_33 <= io_pixelVal_in_2_2;
      end else if (10'h21 == _T_19[9:0]) begin
        image_2_33 <= io_pixelVal_in_2_1;
      end else if (10'h21 == _T_15[9:0]) begin
        image_2_33 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_34 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22 == _T_37[9:0]) begin
        image_2_34 <= io_pixelVal_in_2_7;
      end else if (10'h22 == _T_34[9:0]) begin
        image_2_34 <= io_pixelVal_in_2_6;
      end else if (10'h22 == _T_31[9:0]) begin
        image_2_34 <= io_pixelVal_in_2_5;
      end else if (10'h22 == _T_28[9:0]) begin
        image_2_34 <= io_pixelVal_in_2_4;
      end else if (10'h22 == _T_25[9:0]) begin
        image_2_34 <= io_pixelVal_in_2_3;
      end else if (10'h22 == _T_22[9:0]) begin
        image_2_34 <= io_pixelVal_in_2_2;
      end else if (10'h22 == _T_19[9:0]) begin
        image_2_34 <= io_pixelVal_in_2_1;
      end else if (10'h22 == _T_15[9:0]) begin
        image_2_34 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_35 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23 == _T_37[9:0]) begin
        image_2_35 <= io_pixelVal_in_2_7;
      end else if (10'h23 == _T_34[9:0]) begin
        image_2_35 <= io_pixelVal_in_2_6;
      end else if (10'h23 == _T_31[9:0]) begin
        image_2_35 <= io_pixelVal_in_2_5;
      end else if (10'h23 == _T_28[9:0]) begin
        image_2_35 <= io_pixelVal_in_2_4;
      end else if (10'h23 == _T_25[9:0]) begin
        image_2_35 <= io_pixelVal_in_2_3;
      end else if (10'h23 == _T_22[9:0]) begin
        image_2_35 <= io_pixelVal_in_2_2;
      end else if (10'h23 == _T_19[9:0]) begin
        image_2_35 <= io_pixelVal_in_2_1;
      end else if (10'h23 == _T_15[9:0]) begin
        image_2_35 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_36 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h24 == _T_37[9:0]) begin
        image_2_36 <= io_pixelVal_in_2_7;
      end else if (10'h24 == _T_34[9:0]) begin
        image_2_36 <= io_pixelVal_in_2_6;
      end else if (10'h24 == _T_31[9:0]) begin
        image_2_36 <= io_pixelVal_in_2_5;
      end else if (10'h24 == _T_28[9:0]) begin
        image_2_36 <= io_pixelVal_in_2_4;
      end else if (10'h24 == _T_25[9:0]) begin
        image_2_36 <= io_pixelVal_in_2_3;
      end else if (10'h24 == _T_22[9:0]) begin
        image_2_36 <= io_pixelVal_in_2_2;
      end else if (10'h24 == _T_19[9:0]) begin
        image_2_36 <= io_pixelVal_in_2_1;
      end else if (10'h24 == _T_15[9:0]) begin
        image_2_36 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_37 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h25 == _T_37[9:0]) begin
        image_2_37 <= io_pixelVal_in_2_7;
      end else if (10'h25 == _T_34[9:0]) begin
        image_2_37 <= io_pixelVal_in_2_6;
      end else if (10'h25 == _T_31[9:0]) begin
        image_2_37 <= io_pixelVal_in_2_5;
      end else if (10'h25 == _T_28[9:0]) begin
        image_2_37 <= io_pixelVal_in_2_4;
      end else if (10'h25 == _T_25[9:0]) begin
        image_2_37 <= io_pixelVal_in_2_3;
      end else if (10'h25 == _T_22[9:0]) begin
        image_2_37 <= io_pixelVal_in_2_2;
      end else if (10'h25 == _T_19[9:0]) begin
        image_2_37 <= io_pixelVal_in_2_1;
      end else if (10'h25 == _T_15[9:0]) begin
        image_2_37 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_38 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h26 == _T_37[9:0]) begin
        image_2_38 <= io_pixelVal_in_2_7;
      end else if (10'h26 == _T_34[9:0]) begin
        image_2_38 <= io_pixelVal_in_2_6;
      end else if (10'h26 == _T_31[9:0]) begin
        image_2_38 <= io_pixelVal_in_2_5;
      end else if (10'h26 == _T_28[9:0]) begin
        image_2_38 <= io_pixelVal_in_2_4;
      end else if (10'h26 == _T_25[9:0]) begin
        image_2_38 <= io_pixelVal_in_2_3;
      end else if (10'h26 == _T_22[9:0]) begin
        image_2_38 <= io_pixelVal_in_2_2;
      end else if (10'h26 == _T_19[9:0]) begin
        image_2_38 <= io_pixelVal_in_2_1;
      end else if (10'h26 == _T_15[9:0]) begin
        image_2_38 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_39 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h27 == _T_37[9:0]) begin
        image_2_39 <= io_pixelVal_in_2_7;
      end else if (10'h27 == _T_34[9:0]) begin
        image_2_39 <= io_pixelVal_in_2_6;
      end else if (10'h27 == _T_31[9:0]) begin
        image_2_39 <= io_pixelVal_in_2_5;
      end else if (10'h27 == _T_28[9:0]) begin
        image_2_39 <= io_pixelVal_in_2_4;
      end else if (10'h27 == _T_25[9:0]) begin
        image_2_39 <= io_pixelVal_in_2_3;
      end else if (10'h27 == _T_22[9:0]) begin
        image_2_39 <= io_pixelVal_in_2_2;
      end else if (10'h27 == _T_19[9:0]) begin
        image_2_39 <= io_pixelVal_in_2_1;
      end else if (10'h27 == _T_15[9:0]) begin
        image_2_39 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_40 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h28 == _T_37[9:0]) begin
        image_2_40 <= io_pixelVal_in_2_7;
      end else if (10'h28 == _T_34[9:0]) begin
        image_2_40 <= io_pixelVal_in_2_6;
      end else if (10'h28 == _T_31[9:0]) begin
        image_2_40 <= io_pixelVal_in_2_5;
      end else if (10'h28 == _T_28[9:0]) begin
        image_2_40 <= io_pixelVal_in_2_4;
      end else if (10'h28 == _T_25[9:0]) begin
        image_2_40 <= io_pixelVal_in_2_3;
      end else if (10'h28 == _T_22[9:0]) begin
        image_2_40 <= io_pixelVal_in_2_2;
      end else if (10'h28 == _T_19[9:0]) begin
        image_2_40 <= io_pixelVal_in_2_1;
      end else if (10'h28 == _T_15[9:0]) begin
        image_2_40 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_41 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h29 == _T_37[9:0]) begin
        image_2_41 <= io_pixelVal_in_2_7;
      end else if (10'h29 == _T_34[9:0]) begin
        image_2_41 <= io_pixelVal_in_2_6;
      end else if (10'h29 == _T_31[9:0]) begin
        image_2_41 <= io_pixelVal_in_2_5;
      end else if (10'h29 == _T_28[9:0]) begin
        image_2_41 <= io_pixelVal_in_2_4;
      end else if (10'h29 == _T_25[9:0]) begin
        image_2_41 <= io_pixelVal_in_2_3;
      end else if (10'h29 == _T_22[9:0]) begin
        image_2_41 <= io_pixelVal_in_2_2;
      end else if (10'h29 == _T_19[9:0]) begin
        image_2_41 <= io_pixelVal_in_2_1;
      end else if (10'h29 == _T_15[9:0]) begin
        image_2_41 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_42 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2a == _T_37[9:0]) begin
        image_2_42 <= io_pixelVal_in_2_7;
      end else if (10'h2a == _T_34[9:0]) begin
        image_2_42 <= io_pixelVal_in_2_6;
      end else if (10'h2a == _T_31[9:0]) begin
        image_2_42 <= io_pixelVal_in_2_5;
      end else if (10'h2a == _T_28[9:0]) begin
        image_2_42 <= io_pixelVal_in_2_4;
      end else if (10'h2a == _T_25[9:0]) begin
        image_2_42 <= io_pixelVal_in_2_3;
      end else if (10'h2a == _T_22[9:0]) begin
        image_2_42 <= io_pixelVal_in_2_2;
      end else if (10'h2a == _T_19[9:0]) begin
        image_2_42 <= io_pixelVal_in_2_1;
      end else if (10'h2a == _T_15[9:0]) begin
        image_2_42 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_43 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2b == _T_37[9:0]) begin
        image_2_43 <= io_pixelVal_in_2_7;
      end else if (10'h2b == _T_34[9:0]) begin
        image_2_43 <= io_pixelVal_in_2_6;
      end else if (10'h2b == _T_31[9:0]) begin
        image_2_43 <= io_pixelVal_in_2_5;
      end else if (10'h2b == _T_28[9:0]) begin
        image_2_43 <= io_pixelVal_in_2_4;
      end else if (10'h2b == _T_25[9:0]) begin
        image_2_43 <= io_pixelVal_in_2_3;
      end else if (10'h2b == _T_22[9:0]) begin
        image_2_43 <= io_pixelVal_in_2_2;
      end else if (10'h2b == _T_19[9:0]) begin
        image_2_43 <= io_pixelVal_in_2_1;
      end else if (10'h2b == _T_15[9:0]) begin
        image_2_43 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_44 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2c == _T_37[9:0]) begin
        image_2_44 <= io_pixelVal_in_2_7;
      end else if (10'h2c == _T_34[9:0]) begin
        image_2_44 <= io_pixelVal_in_2_6;
      end else if (10'h2c == _T_31[9:0]) begin
        image_2_44 <= io_pixelVal_in_2_5;
      end else if (10'h2c == _T_28[9:0]) begin
        image_2_44 <= io_pixelVal_in_2_4;
      end else if (10'h2c == _T_25[9:0]) begin
        image_2_44 <= io_pixelVal_in_2_3;
      end else if (10'h2c == _T_22[9:0]) begin
        image_2_44 <= io_pixelVal_in_2_2;
      end else if (10'h2c == _T_19[9:0]) begin
        image_2_44 <= io_pixelVal_in_2_1;
      end else if (10'h2c == _T_15[9:0]) begin
        image_2_44 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_45 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2d == _T_37[9:0]) begin
        image_2_45 <= io_pixelVal_in_2_7;
      end else if (10'h2d == _T_34[9:0]) begin
        image_2_45 <= io_pixelVal_in_2_6;
      end else if (10'h2d == _T_31[9:0]) begin
        image_2_45 <= io_pixelVal_in_2_5;
      end else if (10'h2d == _T_28[9:0]) begin
        image_2_45 <= io_pixelVal_in_2_4;
      end else if (10'h2d == _T_25[9:0]) begin
        image_2_45 <= io_pixelVal_in_2_3;
      end else if (10'h2d == _T_22[9:0]) begin
        image_2_45 <= io_pixelVal_in_2_2;
      end else if (10'h2d == _T_19[9:0]) begin
        image_2_45 <= io_pixelVal_in_2_1;
      end else if (10'h2d == _T_15[9:0]) begin
        image_2_45 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_46 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2e == _T_37[9:0]) begin
        image_2_46 <= io_pixelVal_in_2_7;
      end else if (10'h2e == _T_34[9:0]) begin
        image_2_46 <= io_pixelVal_in_2_6;
      end else if (10'h2e == _T_31[9:0]) begin
        image_2_46 <= io_pixelVal_in_2_5;
      end else if (10'h2e == _T_28[9:0]) begin
        image_2_46 <= io_pixelVal_in_2_4;
      end else if (10'h2e == _T_25[9:0]) begin
        image_2_46 <= io_pixelVal_in_2_3;
      end else if (10'h2e == _T_22[9:0]) begin
        image_2_46 <= io_pixelVal_in_2_2;
      end else if (10'h2e == _T_19[9:0]) begin
        image_2_46 <= io_pixelVal_in_2_1;
      end else if (10'h2e == _T_15[9:0]) begin
        image_2_46 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_47 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2f == _T_37[9:0]) begin
        image_2_47 <= io_pixelVal_in_2_7;
      end else if (10'h2f == _T_34[9:0]) begin
        image_2_47 <= io_pixelVal_in_2_6;
      end else if (10'h2f == _T_31[9:0]) begin
        image_2_47 <= io_pixelVal_in_2_5;
      end else if (10'h2f == _T_28[9:0]) begin
        image_2_47 <= io_pixelVal_in_2_4;
      end else if (10'h2f == _T_25[9:0]) begin
        image_2_47 <= io_pixelVal_in_2_3;
      end else if (10'h2f == _T_22[9:0]) begin
        image_2_47 <= io_pixelVal_in_2_2;
      end else if (10'h2f == _T_19[9:0]) begin
        image_2_47 <= io_pixelVal_in_2_1;
      end else if (10'h2f == _T_15[9:0]) begin
        image_2_47 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_48 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h30 == _T_37[9:0]) begin
        image_2_48 <= io_pixelVal_in_2_7;
      end else if (10'h30 == _T_34[9:0]) begin
        image_2_48 <= io_pixelVal_in_2_6;
      end else if (10'h30 == _T_31[9:0]) begin
        image_2_48 <= io_pixelVal_in_2_5;
      end else if (10'h30 == _T_28[9:0]) begin
        image_2_48 <= io_pixelVal_in_2_4;
      end else if (10'h30 == _T_25[9:0]) begin
        image_2_48 <= io_pixelVal_in_2_3;
      end else if (10'h30 == _T_22[9:0]) begin
        image_2_48 <= io_pixelVal_in_2_2;
      end else if (10'h30 == _T_19[9:0]) begin
        image_2_48 <= io_pixelVal_in_2_1;
      end else if (10'h30 == _T_15[9:0]) begin
        image_2_48 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_49 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h31 == _T_37[9:0]) begin
        image_2_49 <= io_pixelVal_in_2_7;
      end else if (10'h31 == _T_34[9:0]) begin
        image_2_49 <= io_pixelVal_in_2_6;
      end else if (10'h31 == _T_31[9:0]) begin
        image_2_49 <= io_pixelVal_in_2_5;
      end else if (10'h31 == _T_28[9:0]) begin
        image_2_49 <= io_pixelVal_in_2_4;
      end else if (10'h31 == _T_25[9:0]) begin
        image_2_49 <= io_pixelVal_in_2_3;
      end else if (10'h31 == _T_22[9:0]) begin
        image_2_49 <= io_pixelVal_in_2_2;
      end else if (10'h31 == _T_19[9:0]) begin
        image_2_49 <= io_pixelVal_in_2_1;
      end else if (10'h31 == _T_15[9:0]) begin
        image_2_49 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_50 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h32 == _T_37[9:0]) begin
        image_2_50 <= io_pixelVal_in_2_7;
      end else if (10'h32 == _T_34[9:0]) begin
        image_2_50 <= io_pixelVal_in_2_6;
      end else if (10'h32 == _T_31[9:0]) begin
        image_2_50 <= io_pixelVal_in_2_5;
      end else if (10'h32 == _T_28[9:0]) begin
        image_2_50 <= io_pixelVal_in_2_4;
      end else if (10'h32 == _T_25[9:0]) begin
        image_2_50 <= io_pixelVal_in_2_3;
      end else if (10'h32 == _T_22[9:0]) begin
        image_2_50 <= io_pixelVal_in_2_2;
      end else if (10'h32 == _T_19[9:0]) begin
        image_2_50 <= io_pixelVal_in_2_1;
      end else if (10'h32 == _T_15[9:0]) begin
        image_2_50 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_51 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h33 == _T_37[9:0]) begin
        image_2_51 <= io_pixelVal_in_2_7;
      end else if (10'h33 == _T_34[9:0]) begin
        image_2_51 <= io_pixelVal_in_2_6;
      end else if (10'h33 == _T_31[9:0]) begin
        image_2_51 <= io_pixelVal_in_2_5;
      end else if (10'h33 == _T_28[9:0]) begin
        image_2_51 <= io_pixelVal_in_2_4;
      end else if (10'h33 == _T_25[9:0]) begin
        image_2_51 <= io_pixelVal_in_2_3;
      end else if (10'h33 == _T_22[9:0]) begin
        image_2_51 <= io_pixelVal_in_2_2;
      end else if (10'h33 == _T_19[9:0]) begin
        image_2_51 <= io_pixelVal_in_2_1;
      end else if (10'h33 == _T_15[9:0]) begin
        image_2_51 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_52 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h34 == _T_37[9:0]) begin
        image_2_52 <= io_pixelVal_in_2_7;
      end else if (10'h34 == _T_34[9:0]) begin
        image_2_52 <= io_pixelVal_in_2_6;
      end else if (10'h34 == _T_31[9:0]) begin
        image_2_52 <= io_pixelVal_in_2_5;
      end else if (10'h34 == _T_28[9:0]) begin
        image_2_52 <= io_pixelVal_in_2_4;
      end else if (10'h34 == _T_25[9:0]) begin
        image_2_52 <= io_pixelVal_in_2_3;
      end else if (10'h34 == _T_22[9:0]) begin
        image_2_52 <= io_pixelVal_in_2_2;
      end else if (10'h34 == _T_19[9:0]) begin
        image_2_52 <= io_pixelVal_in_2_1;
      end else if (10'h34 == _T_15[9:0]) begin
        image_2_52 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_53 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h35 == _T_37[9:0]) begin
        image_2_53 <= io_pixelVal_in_2_7;
      end else if (10'h35 == _T_34[9:0]) begin
        image_2_53 <= io_pixelVal_in_2_6;
      end else if (10'h35 == _T_31[9:0]) begin
        image_2_53 <= io_pixelVal_in_2_5;
      end else if (10'h35 == _T_28[9:0]) begin
        image_2_53 <= io_pixelVal_in_2_4;
      end else if (10'h35 == _T_25[9:0]) begin
        image_2_53 <= io_pixelVal_in_2_3;
      end else if (10'h35 == _T_22[9:0]) begin
        image_2_53 <= io_pixelVal_in_2_2;
      end else if (10'h35 == _T_19[9:0]) begin
        image_2_53 <= io_pixelVal_in_2_1;
      end else if (10'h35 == _T_15[9:0]) begin
        image_2_53 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_54 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h36 == _T_37[9:0]) begin
        image_2_54 <= io_pixelVal_in_2_7;
      end else if (10'h36 == _T_34[9:0]) begin
        image_2_54 <= io_pixelVal_in_2_6;
      end else if (10'h36 == _T_31[9:0]) begin
        image_2_54 <= io_pixelVal_in_2_5;
      end else if (10'h36 == _T_28[9:0]) begin
        image_2_54 <= io_pixelVal_in_2_4;
      end else if (10'h36 == _T_25[9:0]) begin
        image_2_54 <= io_pixelVal_in_2_3;
      end else if (10'h36 == _T_22[9:0]) begin
        image_2_54 <= io_pixelVal_in_2_2;
      end else if (10'h36 == _T_19[9:0]) begin
        image_2_54 <= io_pixelVal_in_2_1;
      end else if (10'h36 == _T_15[9:0]) begin
        image_2_54 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_55 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h37 == _T_37[9:0]) begin
        image_2_55 <= io_pixelVal_in_2_7;
      end else if (10'h37 == _T_34[9:0]) begin
        image_2_55 <= io_pixelVal_in_2_6;
      end else if (10'h37 == _T_31[9:0]) begin
        image_2_55 <= io_pixelVal_in_2_5;
      end else if (10'h37 == _T_28[9:0]) begin
        image_2_55 <= io_pixelVal_in_2_4;
      end else if (10'h37 == _T_25[9:0]) begin
        image_2_55 <= io_pixelVal_in_2_3;
      end else if (10'h37 == _T_22[9:0]) begin
        image_2_55 <= io_pixelVal_in_2_2;
      end else if (10'h37 == _T_19[9:0]) begin
        image_2_55 <= io_pixelVal_in_2_1;
      end else if (10'h37 == _T_15[9:0]) begin
        image_2_55 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_56 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h38 == _T_37[9:0]) begin
        image_2_56 <= io_pixelVal_in_2_7;
      end else if (10'h38 == _T_34[9:0]) begin
        image_2_56 <= io_pixelVal_in_2_6;
      end else if (10'h38 == _T_31[9:0]) begin
        image_2_56 <= io_pixelVal_in_2_5;
      end else if (10'h38 == _T_28[9:0]) begin
        image_2_56 <= io_pixelVal_in_2_4;
      end else if (10'h38 == _T_25[9:0]) begin
        image_2_56 <= io_pixelVal_in_2_3;
      end else if (10'h38 == _T_22[9:0]) begin
        image_2_56 <= io_pixelVal_in_2_2;
      end else if (10'h38 == _T_19[9:0]) begin
        image_2_56 <= io_pixelVal_in_2_1;
      end else if (10'h38 == _T_15[9:0]) begin
        image_2_56 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_57 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h39 == _T_37[9:0]) begin
        image_2_57 <= io_pixelVal_in_2_7;
      end else if (10'h39 == _T_34[9:0]) begin
        image_2_57 <= io_pixelVal_in_2_6;
      end else if (10'h39 == _T_31[9:0]) begin
        image_2_57 <= io_pixelVal_in_2_5;
      end else if (10'h39 == _T_28[9:0]) begin
        image_2_57 <= io_pixelVal_in_2_4;
      end else if (10'h39 == _T_25[9:0]) begin
        image_2_57 <= io_pixelVal_in_2_3;
      end else if (10'h39 == _T_22[9:0]) begin
        image_2_57 <= io_pixelVal_in_2_2;
      end else if (10'h39 == _T_19[9:0]) begin
        image_2_57 <= io_pixelVal_in_2_1;
      end else if (10'h39 == _T_15[9:0]) begin
        image_2_57 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_58 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3a == _T_37[9:0]) begin
        image_2_58 <= io_pixelVal_in_2_7;
      end else if (10'h3a == _T_34[9:0]) begin
        image_2_58 <= io_pixelVal_in_2_6;
      end else if (10'h3a == _T_31[9:0]) begin
        image_2_58 <= io_pixelVal_in_2_5;
      end else if (10'h3a == _T_28[9:0]) begin
        image_2_58 <= io_pixelVal_in_2_4;
      end else if (10'h3a == _T_25[9:0]) begin
        image_2_58 <= io_pixelVal_in_2_3;
      end else if (10'h3a == _T_22[9:0]) begin
        image_2_58 <= io_pixelVal_in_2_2;
      end else if (10'h3a == _T_19[9:0]) begin
        image_2_58 <= io_pixelVal_in_2_1;
      end else if (10'h3a == _T_15[9:0]) begin
        image_2_58 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_59 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3b == _T_37[9:0]) begin
        image_2_59 <= io_pixelVal_in_2_7;
      end else if (10'h3b == _T_34[9:0]) begin
        image_2_59 <= io_pixelVal_in_2_6;
      end else if (10'h3b == _T_31[9:0]) begin
        image_2_59 <= io_pixelVal_in_2_5;
      end else if (10'h3b == _T_28[9:0]) begin
        image_2_59 <= io_pixelVal_in_2_4;
      end else if (10'h3b == _T_25[9:0]) begin
        image_2_59 <= io_pixelVal_in_2_3;
      end else if (10'h3b == _T_22[9:0]) begin
        image_2_59 <= io_pixelVal_in_2_2;
      end else if (10'h3b == _T_19[9:0]) begin
        image_2_59 <= io_pixelVal_in_2_1;
      end else if (10'h3b == _T_15[9:0]) begin
        image_2_59 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_60 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3c == _T_37[9:0]) begin
        image_2_60 <= io_pixelVal_in_2_7;
      end else if (10'h3c == _T_34[9:0]) begin
        image_2_60 <= io_pixelVal_in_2_6;
      end else if (10'h3c == _T_31[9:0]) begin
        image_2_60 <= io_pixelVal_in_2_5;
      end else if (10'h3c == _T_28[9:0]) begin
        image_2_60 <= io_pixelVal_in_2_4;
      end else if (10'h3c == _T_25[9:0]) begin
        image_2_60 <= io_pixelVal_in_2_3;
      end else if (10'h3c == _T_22[9:0]) begin
        image_2_60 <= io_pixelVal_in_2_2;
      end else if (10'h3c == _T_19[9:0]) begin
        image_2_60 <= io_pixelVal_in_2_1;
      end else if (10'h3c == _T_15[9:0]) begin
        image_2_60 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_61 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3d == _T_37[9:0]) begin
        image_2_61 <= io_pixelVal_in_2_7;
      end else if (10'h3d == _T_34[9:0]) begin
        image_2_61 <= io_pixelVal_in_2_6;
      end else if (10'h3d == _T_31[9:0]) begin
        image_2_61 <= io_pixelVal_in_2_5;
      end else if (10'h3d == _T_28[9:0]) begin
        image_2_61 <= io_pixelVal_in_2_4;
      end else if (10'h3d == _T_25[9:0]) begin
        image_2_61 <= io_pixelVal_in_2_3;
      end else if (10'h3d == _T_22[9:0]) begin
        image_2_61 <= io_pixelVal_in_2_2;
      end else if (10'h3d == _T_19[9:0]) begin
        image_2_61 <= io_pixelVal_in_2_1;
      end else if (10'h3d == _T_15[9:0]) begin
        image_2_61 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_62 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3e == _T_37[9:0]) begin
        image_2_62 <= io_pixelVal_in_2_7;
      end else if (10'h3e == _T_34[9:0]) begin
        image_2_62 <= io_pixelVal_in_2_6;
      end else if (10'h3e == _T_31[9:0]) begin
        image_2_62 <= io_pixelVal_in_2_5;
      end else if (10'h3e == _T_28[9:0]) begin
        image_2_62 <= io_pixelVal_in_2_4;
      end else if (10'h3e == _T_25[9:0]) begin
        image_2_62 <= io_pixelVal_in_2_3;
      end else if (10'h3e == _T_22[9:0]) begin
        image_2_62 <= io_pixelVal_in_2_2;
      end else if (10'h3e == _T_19[9:0]) begin
        image_2_62 <= io_pixelVal_in_2_1;
      end else if (10'h3e == _T_15[9:0]) begin
        image_2_62 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_63 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3f == _T_37[9:0]) begin
        image_2_63 <= io_pixelVal_in_2_7;
      end else if (10'h3f == _T_34[9:0]) begin
        image_2_63 <= io_pixelVal_in_2_6;
      end else if (10'h3f == _T_31[9:0]) begin
        image_2_63 <= io_pixelVal_in_2_5;
      end else if (10'h3f == _T_28[9:0]) begin
        image_2_63 <= io_pixelVal_in_2_4;
      end else if (10'h3f == _T_25[9:0]) begin
        image_2_63 <= io_pixelVal_in_2_3;
      end else if (10'h3f == _T_22[9:0]) begin
        image_2_63 <= io_pixelVal_in_2_2;
      end else if (10'h3f == _T_19[9:0]) begin
        image_2_63 <= io_pixelVal_in_2_1;
      end else if (10'h3f == _T_15[9:0]) begin
        image_2_63 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_64 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h40 == _T_37[9:0]) begin
        image_2_64 <= io_pixelVal_in_2_7;
      end else if (10'h40 == _T_34[9:0]) begin
        image_2_64 <= io_pixelVal_in_2_6;
      end else if (10'h40 == _T_31[9:0]) begin
        image_2_64 <= io_pixelVal_in_2_5;
      end else if (10'h40 == _T_28[9:0]) begin
        image_2_64 <= io_pixelVal_in_2_4;
      end else if (10'h40 == _T_25[9:0]) begin
        image_2_64 <= io_pixelVal_in_2_3;
      end else if (10'h40 == _T_22[9:0]) begin
        image_2_64 <= io_pixelVal_in_2_2;
      end else if (10'h40 == _T_19[9:0]) begin
        image_2_64 <= io_pixelVal_in_2_1;
      end else if (10'h40 == _T_15[9:0]) begin
        image_2_64 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_65 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h41 == _T_37[9:0]) begin
        image_2_65 <= io_pixelVal_in_2_7;
      end else if (10'h41 == _T_34[9:0]) begin
        image_2_65 <= io_pixelVal_in_2_6;
      end else if (10'h41 == _T_31[9:0]) begin
        image_2_65 <= io_pixelVal_in_2_5;
      end else if (10'h41 == _T_28[9:0]) begin
        image_2_65 <= io_pixelVal_in_2_4;
      end else if (10'h41 == _T_25[9:0]) begin
        image_2_65 <= io_pixelVal_in_2_3;
      end else if (10'h41 == _T_22[9:0]) begin
        image_2_65 <= io_pixelVal_in_2_2;
      end else if (10'h41 == _T_19[9:0]) begin
        image_2_65 <= io_pixelVal_in_2_1;
      end else if (10'h41 == _T_15[9:0]) begin
        image_2_65 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_66 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h42 == _T_37[9:0]) begin
        image_2_66 <= io_pixelVal_in_2_7;
      end else if (10'h42 == _T_34[9:0]) begin
        image_2_66 <= io_pixelVal_in_2_6;
      end else if (10'h42 == _T_31[9:0]) begin
        image_2_66 <= io_pixelVal_in_2_5;
      end else if (10'h42 == _T_28[9:0]) begin
        image_2_66 <= io_pixelVal_in_2_4;
      end else if (10'h42 == _T_25[9:0]) begin
        image_2_66 <= io_pixelVal_in_2_3;
      end else if (10'h42 == _T_22[9:0]) begin
        image_2_66 <= io_pixelVal_in_2_2;
      end else if (10'h42 == _T_19[9:0]) begin
        image_2_66 <= io_pixelVal_in_2_1;
      end else if (10'h42 == _T_15[9:0]) begin
        image_2_66 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_67 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h43 == _T_37[9:0]) begin
        image_2_67 <= io_pixelVal_in_2_7;
      end else if (10'h43 == _T_34[9:0]) begin
        image_2_67 <= io_pixelVal_in_2_6;
      end else if (10'h43 == _T_31[9:0]) begin
        image_2_67 <= io_pixelVal_in_2_5;
      end else if (10'h43 == _T_28[9:0]) begin
        image_2_67 <= io_pixelVal_in_2_4;
      end else if (10'h43 == _T_25[9:0]) begin
        image_2_67 <= io_pixelVal_in_2_3;
      end else if (10'h43 == _T_22[9:0]) begin
        image_2_67 <= io_pixelVal_in_2_2;
      end else if (10'h43 == _T_19[9:0]) begin
        image_2_67 <= io_pixelVal_in_2_1;
      end else if (10'h43 == _T_15[9:0]) begin
        image_2_67 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_68 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h44 == _T_37[9:0]) begin
        image_2_68 <= io_pixelVal_in_2_7;
      end else if (10'h44 == _T_34[9:0]) begin
        image_2_68 <= io_pixelVal_in_2_6;
      end else if (10'h44 == _T_31[9:0]) begin
        image_2_68 <= io_pixelVal_in_2_5;
      end else if (10'h44 == _T_28[9:0]) begin
        image_2_68 <= io_pixelVal_in_2_4;
      end else if (10'h44 == _T_25[9:0]) begin
        image_2_68 <= io_pixelVal_in_2_3;
      end else if (10'h44 == _T_22[9:0]) begin
        image_2_68 <= io_pixelVal_in_2_2;
      end else if (10'h44 == _T_19[9:0]) begin
        image_2_68 <= io_pixelVal_in_2_1;
      end else if (10'h44 == _T_15[9:0]) begin
        image_2_68 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_69 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h45 == _T_37[9:0]) begin
        image_2_69 <= io_pixelVal_in_2_7;
      end else if (10'h45 == _T_34[9:0]) begin
        image_2_69 <= io_pixelVal_in_2_6;
      end else if (10'h45 == _T_31[9:0]) begin
        image_2_69 <= io_pixelVal_in_2_5;
      end else if (10'h45 == _T_28[9:0]) begin
        image_2_69 <= io_pixelVal_in_2_4;
      end else if (10'h45 == _T_25[9:0]) begin
        image_2_69 <= io_pixelVal_in_2_3;
      end else if (10'h45 == _T_22[9:0]) begin
        image_2_69 <= io_pixelVal_in_2_2;
      end else if (10'h45 == _T_19[9:0]) begin
        image_2_69 <= io_pixelVal_in_2_1;
      end else if (10'h45 == _T_15[9:0]) begin
        image_2_69 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_70 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h46 == _T_37[9:0]) begin
        image_2_70 <= io_pixelVal_in_2_7;
      end else if (10'h46 == _T_34[9:0]) begin
        image_2_70 <= io_pixelVal_in_2_6;
      end else if (10'h46 == _T_31[9:0]) begin
        image_2_70 <= io_pixelVal_in_2_5;
      end else if (10'h46 == _T_28[9:0]) begin
        image_2_70 <= io_pixelVal_in_2_4;
      end else if (10'h46 == _T_25[9:0]) begin
        image_2_70 <= io_pixelVal_in_2_3;
      end else if (10'h46 == _T_22[9:0]) begin
        image_2_70 <= io_pixelVal_in_2_2;
      end else if (10'h46 == _T_19[9:0]) begin
        image_2_70 <= io_pixelVal_in_2_1;
      end else if (10'h46 == _T_15[9:0]) begin
        image_2_70 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_71 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h47 == _T_37[9:0]) begin
        image_2_71 <= io_pixelVal_in_2_7;
      end else if (10'h47 == _T_34[9:0]) begin
        image_2_71 <= io_pixelVal_in_2_6;
      end else if (10'h47 == _T_31[9:0]) begin
        image_2_71 <= io_pixelVal_in_2_5;
      end else if (10'h47 == _T_28[9:0]) begin
        image_2_71 <= io_pixelVal_in_2_4;
      end else if (10'h47 == _T_25[9:0]) begin
        image_2_71 <= io_pixelVal_in_2_3;
      end else if (10'h47 == _T_22[9:0]) begin
        image_2_71 <= io_pixelVal_in_2_2;
      end else if (10'h47 == _T_19[9:0]) begin
        image_2_71 <= io_pixelVal_in_2_1;
      end else if (10'h47 == _T_15[9:0]) begin
        image_2_71 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_72 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h48 == _T_37[9:0]) begin
        image_2_72 <= io_pixelVal_in_2_7;
      end else if (10'h48 == _T_34[9:0]) begin
        image_2_72 <= io_pixelVal_in_2_6;
      end else if (10'h48 == _T_31[9:0]) begin
        image_2_72 <= io_pixelVal_in_2_5;
      end else if (10'h48 == _T_28[9:0]) begin
        image_2_72 <= io_pixelVal_in_2_4;
      end else if (10'h48 == _T_25[9:0]) begin
        image_2_72 <= io_pixelVal_in_2_3;
      end else if (10'h48 == _T_22[9:0]) begin
        image_2_72 <= io_pixelVal_in_2_2;
      end else if (10'h48 == _T_19[9:0]) begin
        image_2_72 <= io_pixelVal_in_2_1;
      end else if (10'h48 == _T_15[9:0]) begin
        image_2_72 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_73 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h49 == _T_37[9:0]) begin
        image_2_73 <= io_pixelVal_in_2_7;
      end else if (10'h49 == _T_34[9:0]) begin
        image_2_73 <= io_pixelVal_in_2_6;
      end else if (10'h49 == _T_31[9:0]) begin
        image_2_73 <= io_pixelVal_in_2_5;
      end else if (10'h49 == _T_28[9:0]) begin
        image_2_73 <= io_pixelVal_in_2_4;
      end else if (10'h49 == _T_25[9:0]) begin
        image_2_73 <= io_pixelVal_in_2_3;
      end else if (10'h49 == _T_22[9:0]) begin
        image_2_73 <= io_pixelVal_in_2_2;
      end else if (10'h49 == _T_19[9:0]) begin
        image_2_73 <= io_pixelVal_in_2_1;
      end else if (10'h49 == _T_15[9:0]) begin
        image_2_73 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_74 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4a == _T_37[9:0]) begin
        image_2_74 <= io_pixelVal_in_2_7;
      end else if (10'h4a == _T_34[9:0]) begin
        image_2_74 <= io_pixelVal_in_2_6;
      end else if (10'h4a == _T_31[9:0]) begin
        image_2_74 <= io_pixelVal_in_2_5;
      end else if (10'h4a == _T_28[9:0]) begin
        image_2_74 <= io_pixelVal_in_2_4;
      end else if (10'h4a == _T_25[9:0]) begin
        image_2_74 <= io_pixelVal_in_2_3;
      end else if (10'h4a == _T_22[9:0]) begin
        image_2_74 <= io_pixelVal_in_2_2;
      end else if (10'h4a == _T_19[9:0]) begin
        image_2_74 <= io_pixelVal_in_2_1;
      end else if (10'h4a == _T_15[9:0]) begin
        image_2_74 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_75 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4b == _T_37[9:0]) begin
        image_2_75 <= io_pixelVal_in_2_7;
      end else if (10'h4b == _T_34[9:0]) begin
        image_2_75 <= io_pixelVal_in_2_6;
      end else if (10'h4b == _T_31[9:0]) begin
        image_2_75 <= io_pixelVal_in_2_5;
      end else if (10'h4b == _T_28[9:0]) begin
        image_2_75 <= io_pixelVal_in_2_4;
      end else if (10'h4b == _T_25[9:0]) begin
        image_2_75 <= io_pixelVal_in_2_3;
      end else if (10'h4b == _T_22[9:0]) begin
        image_2_75 <= io_pixelVal_in_2_2;
      end else if (10'h4b == _T_19[9:0]) begin
        image_2_75 <= io_pixelVal_in_2_1;
      end else if (10'h4b == _T_15[9:0]) begin
        image_2_75 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_76 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4c == _T_37[9:0]) begin
        image_2_76 <= io_pixelVal_in_2_7;
      end else if (10'h4c == _T_34[9:0]) begin
        image_2_76 <= io_pixelVal_in_2_6;
      end else if (10'h4c == _T_31[9:0]) begin
        image_2_76 <= io_pixelVal_in_2_5;
      end else if (10'h4c == _T_28[9:0]) begin
        image_2_76 <= io_pixelVal_in_2_4;
      end else if (10'h4c == _T_25[9:0]) begin
        image_2_76 <= io_pixelVal_in_2_3;
      end else if (10'h4c == _T_22[9:0]) begin
        image_2_76 <= io_pixelVal_in_2_2;
      end else if (10'h4c == _T_19[9:0]) begin
        image_2_76 <= io_pixelVal_in_2_1;
      end else if (10'h4c == _T_15[9:0]) begin
        image_2_76 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_77 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4d == _T_37[9:0]) begin
        image_2_77 <= io_pixelVal_in_2_7;
      end else if (10'h4d == _T_34[9:0]) begin
        image_2_77 <= io_pixelVal_in_2_6;
      end else if (10'h4d == _T_31[9:0]) begin
        image_2_77 <= io_pixelVal_in_2_5;
      end else if (10'h4d == _T_28[9:0]) begin
        image_2_77 <= io_pixelVal_in_2_4;
      end else if (10'h4d == _T_25[9:0]) begin
        image_2_77 <= io_pixelVal_in_2_3;
      end else if (10'h4d == _T_22[9:0]) begin
        image_2_77 <= io_pixelVal_in_2_2;
      end else if (10'h4d == _T_19[9:0]) begin
        image_2_77 <= io_pixelVal_in_2_1;
      end else if (10'h4d == _T_15[9:0]) begin
        image_2_77 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_78 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4e == _T_37[9:0]) begin
        image_2_78 <= io_pixelVal_in_2_7;
      end else if (10'h4e == _T_34[9:0]) begin
        image_2_78 <= io_pixelVal_in_2_6;
      end else if (10'h4e == _T_31[9:0]) begin
        image_2_78 <= io_pixelVal_in_2_5;
      end else if (10'h4e == _T_28[9:0]) begin
        image_2_78 <= io_pixelVal_in_2_4;
      end else if (10'h4e == _T_25[9:0]) begin
        image_2_78 <= io_pixelVal_in_2_3;
      end else if (10'h4e == _T_22[9:0]) begin
        image_2_78 <= io_pixelVal_in_2_2;
      end else if (10'h4e == _T_19[9:0]) begin
        image_2_78 <= io_pixelVal_in_2_1;
      end else if (10'h4e == _T_15[9:0]) begin
        image_2_78 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_79 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4f == _T_37[9:0]) begin
        image_2_79 <= io_pixelVal_in_2_7;
      end else if (10'h4f == _T_34[9:0]) begin
        image_2_79 <= io_pixelVal_in_2_6;
      end else if (10'h4f == _T_31[9:0]) begin
        image_2_79 <= io_pixelVal_in_2_5;
      end else if (10'h4f == _T_28[9:0]) begin
        image_2_79 <= io_pixelVal_in_2_4;
      end else if (10'h4f == _T_25[9:0]) begin
        image_2_79 <= io_pixelVal_in_2_3;
      end else if (10'h4f == _T_22[9:0]) begin
        image_2_79 <= io_pixelVal_in_2_2;
      end else if (10'h4f == _T_19[9:0]) begin
        image_2_79 <= io_pixelVal_in_2_1;
      end else if (10'h4f == _T_15[9:0]) begin
        image_2_79 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_80 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h50 == _T_37[9:0]) begin
        image_2_80 <= io_pixelVal_in_2_7;
      end else if (10'h50 == _T_34[9:0]) begin
        image_2_80 <= io_pixelVal_in_2_6;
      end else if (10'h50 == _T_31[9:0]) begin
        image_2_80 <= io_pixelVal_in_2_5;
      end else if (10'h50 == _T_28[9:0]) begin
        image_2_80 <= io_pixelVal_in_2_4;
      end else if (10'h50 == _T_25[9:0]) begin
        image_2_80 <= io_pixelVal_in_2_3;
      end else if (10'h50 == _T_22[9:0]) begin
        image_2_80 <= io_pixelVal_in_2_2;
      end else if (10'h50 == _T_19[9:0]) begin
        image_2_80 <= io_pixelVal_in_2_1;
      end else if (10'h50 == _T_15[9:0]) begin
        image_2_80 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_81 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h51 == _T_37[9:0]) begin
        image_2_81 <= io_pixelVal_in_2_7;
      end else if (10'h51 == _T_34[9:0]) begin
        image_2_81 <= io_pixelVal_in_2_6;
      end else if (10'h51 == _T_31[9:0]) begin
        image_2_81 <= io_pixelVal_in_2_5;
      end else if (10'h51 == _T_28[9:0]) begin
        image_2_81 <= io_pixelVal_in_2_4;
      end else if (10'h51 == _T_25[9:0]) begin
        image_2_81 <= io_pixelVal_in_2_3;
      end else if (10'h51 == _T_22[9:0]) begin
        image_2_81 <= io_pixelVal_in_2_2;
      end else if (10'h51 == _T_19[9:0]) begin
        image_2_81 <= io_pixelVal_in_2_1;
      end else if (10'h51 == _T_15[9:0]) begin
        image_2_81 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_82 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h52 == _T_37[9:0]) begin
        image_2_82 <= io_pixelVal_in_2_7;
      end else if (10'h52 == _T_34[9:0]) begin
        image_2_82 <= io_pixelVal_in_2_6;
      end else if (10'h52 == _T_31[9:0]) begin
        image_2_82 <= io_pixelVal_in_2_5;
      end else if (10'h52 == _T_28[9:0]) begin
        image_2_82 <= io_pixelVal_in_2_4;
      end else if (10'h52 == _T_25[9:0]) begin
        image_2_82 <= io_pixelVal_in_2_3;
      end else if (10'h52 == _T_22[9:0]) begin
        image_2_82 <= io_pixelVal_in_2_2;
      end else if (10'h52 == _T_19[9:0]) begin
        image_2_82 <= io_pixelVal_in_2_1;
      end else if (10'h52 == _T_15[9:0]) begin
        image_2_82 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_83 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h53 == _T_37[9:0]) begin
        image_2_83 <= io_pixelVal_in_2_7;
      end else if (10'h53 == _T_34[9:0]) begin
        image_2_83 <= io_pixelVal_in_2_6;
      end else if (10'h53 == _T_31[9:0]) begin
        image_2_83 <= io_pixelVal_in_2_5;
      end else if (10'h53 == _T_28[9:0]) begin
        image_2_83 <= io_pixelVal_in_2_4;
      end else if (10'h53 == _T_25[9:0]) begin
        image_2_83 <= io_pixelVal_in_2_3;
      end else if (10'h53 == _T_22[9:0]) begin
        image_2_83 <= io_pixelVal_in_2_2;
      end else if (10'h53 == _T_19[9:0]) begin
        image_2_83 <= io_pixelVal_in_2_1;
      end else if (10'h53 == _T_15[9:0]) begin
        image_2_83 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_84 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h54 == _T_37[9:0]) begin
        image_2_84 <= io_pixelVal_in_2_7;
      end else if (10'h54 == _T_34[9:0]) begin
        image_2_84 <= io_pixelVal_in_2_6;
      end else if (10'h54 == _T_31[9:0]) begin
        image_2_84 <= io_pixelVal_in_2_5;
      end else if (10'h54 == _T_28[9:0]) begin
        image_2_84 <= io_pixelVal_in_2_4;
      end else if (10'h54 == _T_25[9:0]) begin
        image_2_84 <= io_pixelVal_in_2_3;
      end else if (10'h54 == _T_22[9:0]) begin
        image_2_84 <= io_pixelVal_in_2_2;
      end else if (10'h54 == _T_19[9:0]) begin
        image_2_84 <= io_pixelVal_in_2_1;
      end else if (10'h54 == _T_15[9:0]) begin
        image_2_84 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_85 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h55 == _T_37[9:0]) begin
        image_2_85 <= io_pixelVal_in_2_7;
      end else if (10'h55 == _T_34[9:0]) begin
        image_2_85 <= io_pixelVal_in_2_6;
      end else if (10'h55 == _T_31[9:0]) begin
        image_2_85 <= io_pixelVal_in_2_5;
      end else if (10'h55 == _T_28[9:0]) begin
        image_2_85 <= io_pixelVal_in_2_4;
      end else if (10'h55 == _T_25[9:0]) begin
        image_2_85 <= io_pixelVal_in_2_3;
      end else if (10'h55 == _T_22[9:0]) begin
        image_2_85 <= io_pixelVal_in_2_2;
      end else if (10'h55 == _T_19[9:0]) begin
        image_2_85 <= io_pixelVal_in_2_1;
      end else if (10'h55 == _T_15[9:0]) begin
        image_2_85 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_86 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h56 == _T_37[9:0]) begin
        image_2_86 <= io_pixelVal_in_2_7;
      end else if (10'h56 == _T_34[9:0]) begin
        image_2_86 <= io_pixelVal_in_2_6;
      end else if (10'h56 == _T_31[9:0]) begin
        image_2_86 <= io_pixelVal_in_2_5;
      end else if (10'h56 == _T_28[9:0]) begin
        image_2_86 <= io_pixelVal_in_2_4;
      end else if (10'h56 == _T_25[9:0]) begin
        image_2_86 <= io_pixelVal_in_2_3;
      end else if (10'h56 == _T_22[9:0]) begin
        image_2_86 <= io_pixelVal_in_2_2;
      end else if (10'h56 == _T_19[9:0]) begin
        image_2_86 <= io_pixelVal_in_2_1;
      end else if (10'h56 == _T_15[9:0]) begin
        image_2_86 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_87 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h57 == _T_37[9:0]) begin
        image_2_87 <= io_pixelVal_in_2_7;
      end else if (10'h57 == _T_34[9:0]) begin
        image_2_87 <= io_pixelVal_in_2_6;
      end else if (10'h57 == _T_31[9:0]) begin
        image_2_87 <= io_pixelVal_in_2_5;
      end else if (10'h57 == _T_28[9:0]) begin
        image_2_87 <= io_pixelVal_in_2_4;
      end else if (10'h57 == _T_25[9:0]) begin
        image_2_87 <= io_pixelVal_in_2_3;
      end else if (10'h57 == _T_22[9:0]) begin
        image_2_87 <= io_pixelVal_in_2_2;
      end else if (10'h57 == _T_19[9:0]) begin
        image_2_87 <= io_pixelVal_in_2_1;
      end else if (10'h57 == _T_15[9:0]) begin
        image_2_87 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_88 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h58 == _T_37[9:0]) begin
        image_2_88 <= io_pixelVal_in_2_7;
      end else if (10'h58 == _T_34[9:0]) begin
        image_2_88 <= io_pixelVal_in_2_6;
      end else if (10'h58 == _T_31[9:0]) begin
        image_2_88 <= io_pixelVal_in_2_5;
      end else if (10'h58 == _T_28[9:0]) begin
        image_2_88 <= io_pixelVal_in_2_4;
      end else if (10'h58 == _T_25[9:0]) begin
        image_2_88 <= io_pixelVal_in_2_3;
      end else if (10'h58 == _T_22[9:0]) begin
        image_2_88 <= io_pixelVal_in_2_2;
      end else if (10'h58 == _T_19[9:0]) begin
        image_2_88 <= io_pixelVal_in_2_1;
      end else if (10'h58 == _T_15[9:0]) begin
        image_2_88 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_89 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h59 == _T_37[9:0]) begin
        image_2_89 <= io_pixelVal_in_2_7;
      end else if (10'h59 == _T_34[9:0]) begin
        image_2_89 <= io_pixelVal_in_2_6;
      end else if (10'h59 == _T_31[9:0]) begin
        image_2_89 <= io_pixelVal_in_2_5;
      end else if (10'h59 == _T_28[9:0]) begin
        image_2_89 <= io_pixelVal_in_2_4;
      end else if (10'h59 == _T_25[9:0]) begin
        image_2_89 <= io_pixelVal_in_2_3;
      end else if (10'h59 == _T_22[9:0]) begin
        image_2_89 <= io_pixelVal_in_2_2;
      end else if (10'h59 == _T_19[9:0]) begin
        image_2_89 <= io_pixelVal_in_2_1;
      end else if (10'h59 == _T_15[9:0]) begin
        image_2_89 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_90 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5a == _T_37[9:0]) begin
        image_2_90 <= io_pixelVal_in_2_7;
      end else if (10'h5a == _T_34[9:0]) begin
        image_2_90 <= io_pixelVal_in_2_6;
      end else if (10'h5a == _T_31[9:0]) begin
        image_2_90 <= io_pixelVal_in_2_5;
      end else if (10'h5a == _T_28[9:0]) begin
        image_2_90 <= io_pixelVal_in_2_4;
      end else if (10'h5a == _T_25[9:0]) begin
        image_2_90 <= io_pixelVal_in_2_3;
      end else if (10'h5a == _T_22[9:0]) begin
        image_2_90 <= io_pixelVal_in_2_2;
      end else if (10'h5a == _T_19[9:0]) begin
        image_2_90 <= io_pixelVal_in_2_1;
      end else if (10'h5a == _T_15[9:0]) begin
        image_2_90 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_91 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5b == _T_37[9:0]) begin
        image_2_91 <= io_pixelVal_in_2_7;
      end else if (10'h5b == _T_34[9:0]) begin
        image_2_91 <= io_pixelVal_in_2_6;
      end else if (10'h5b == _T_31[9:0]) begin
        image_2_91 <= io_pixelVal_in_2_5;
      end else if (10'h5b == _T_28[9:0]) begin
        image_2_91 <= io_pixelVal_in_2_4;
      end else if (10'h5b == _T_25[9:0]) begin
        image_2_91 <= io_pixelVal_in_2_3;
      end else if (10'h5b == _T_22[9:0]) begin
        image_2_91 <= io_pixelVal_in_2_2;
      end else if (10'h5b == _T_19[9:0]) begin
        image_2_91 <= io_pixelVal_in_2_1;
      end else if (10'h5b == _T_15[9:0]) begin
        image_2_91 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_92 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5c == _T_37[9:0]) begin
        image_2_92 <= io_pixelVal_in_2_7;
      end else if (10'h5c == _T_34[9:0]) begin
        image_2_92 <= io_pixelVal_in_2_6;
      end else if (10'h5c == _T_31[9:0]) begin
        image_2_92 <= io_pixelVal_in_2_5;
      end else if (10'h5c == _T_28[9:0]) begin
        image_2_92 <= io_pixelVal_in_2_4;
      end else if (10'h5c == _T_25[9:0]) begin
        image_2_92 <= io_pixelVal_in_2_3;
      end else if (10'h5c == _T_22[9:0]) begin
        image_2_92 <= io_pixelVal_in_2_2;
      end else if (10'h5c == _T_19[9:0]) begin
        image_2_92 <= io_pixelVal_in_2_1;
      end else if (10'h5c == _T_15[9:0]) begin
        image_2_92 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_93 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5d == _T_37[9:0]) begin
        image_2_93 <= io_pixelVal_in_2_7;
      end else if (10'h5d == _T_34[9:0]) begin
        image_2_93 <= io_pixelVal_in_2_6;
      end else if (10'h5d == _T_31[9:0]) begin
        image_2_93 <= io_pixelVal_in_2_5;
      end else if (10'h5d == _T_28[9:0]) begin
        image_2_93 <= io_pixelVal_in_2_4;
      end else if (10'h5d == _T_25[9:0]) begin
        image_2_93 <= io_pixelVal_in_2_3;
      end else if (10'h5d == _T_22[9:0]) begin
        image_2_93 <= io_pixelVal_in_2_2;
      end else if (10'h5d == _T_19[9:0]) begin
        image_2_93 <= io_pixelVal_in_2_1;
      end else if (10'h5d == _T_15[9:0]) begin
        image_2_93 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_94 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5e == _T_37[9:0]) begin
        image_2_94 <= io_pixelVal_in_2_7;
      end else if (10'h5e == _T_34[9:0]) begin
        image_2_94 <= io_pixelVal_in_2_6;
      end else if (10'h5e == _T_31[9:0]) begin
        image_2_94 <= io_pixelVal_in_2_5;
      end else if (10'h5e == _T_28[9:0]) begin
        image_2_94 <= io_pixelVal_in_2_4;
      end else if (10'h5e == _T_25[9:0]) begin
        image_2_94 <= io_pixelVal_in_2_3;
      end else if (10'h5e == _T_22[9:0]) begin
        image_2_94 <= io_pixelVal_in_2_2;
      end else if (10'h5e == _T_19[9:0]) begin
        image_2_94 <= io_pixelVal_in_2_1;
      end else if (10'h5e == _T_15[9:0]) begin
        image_2_94 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_95 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5f == _T_37[9:0]) begin
        image_2_95 <= io_pixelVal_in_2_7;
      end else if (10'h5f == _T_34[9:0]) begin
        image_2_95 <= io_pixelVal_in_2_6;
      end else if (10'h5f == _T_31[9:0]) begin
        image_2_95 <= io_pixelVal_in_2_5;
      end else if (10'h5f == _T_28[9:0]) begin
        image_2_95 <= io_pixelVal_in_2_4;
      end else if (10'h5f == _T_25[9:0]) begin
        image_2_95 <= io_pixelVal_in_2_3;
      end else if (10'h5f == _T_22[9:0]) begin
        image_2_95 <= io_pixelVal_in_2_2;
      end else if (10'h5f == _T_19[9:0]) begin
        image_2_95 <= io_pixelVal_in_2_1;
      end else if (10'h5f == _T_15[9:0]) begin
        image_2_95 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_96 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h60 == _T_37[9:0]) begin
        image_2_96 <= io_pixelVal_in_2_7;
      end else if (10'h60 == _T_34[9:0]) begin
        image_2_96 <= io_pixelVal_in_2_6;
      end else if (10'h60 == _T_31[9:0]) begin
        image_2_96 <= io_pixelVal_in_2_5;
      end else if (10'h60 == _T_28[9:0]) begin
        image_2_96 <= io_pixelVal_in_2_4;
      end else if (10'h60 == _T_25[9:0]) begin
        image_2_96 <= io_pixelVal_in_2_3;
      end else if (10'h60 == _T_22[9:0]) begin
        image_2_96 <= io_pixelVal_in_2_2;
      end else if (10'h60 == _T_19[9:0]) begin
        image_2_96 <= io_pixelVal_in_2_1;
      end else if (10'h60 == _T_15[9:0]) begin
        image_2_96 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_97 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h61 == _T_37[9:0]) begin
        image_2_97 <= io_pixelVal_in_2_7;
      end else if (10'h61 == _T_34[9:0]) begin
        image_2_97 <= io_pixelVal_in_2_6;
      end else if (10'h61 == _T_31[9:0]) begin
        image_2_97 <= io_pixelVal_in_2_5;
      end else if (10'h61 == _T_28[9:0]) begin
        image_2_97 <= io_pixelVal_in_2_4;
      end else if (10'h61 == _T_25[9:0]) begin
        image_2_97 <= io_pixelVal_in_2_3;
      end else if (10'h61 == _T_22[9:0]) begin
        image_2_97 <= io_pixelVal_in_2_2;
      end else if (10'h61 == _T_19[9:0]) begin
        image_2_97 <= io_pixelVal_in_2_1;
      end else if (10'h61 == _T_15[9:0]) begin
        image_2_97 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_98 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h62 == _T_37[9:0]) begin
        image_2_98 <= io_pixelVal_in_2_7;
      end else if (10'h62 == _T_34[9:0]) begin
        image_2_98 <= io_pixelVal_in_2_6;
      end else if (10'h62 == _T_31[9:0]) begin
        image_2_98 <= io_pixelVal_in_2_5;
      end else if (10'h62 == _T_28[9:0]) begin
        image_2_98 <= io_pixelVal_in_2_4;
      end else if (10'h62 == _T_25[9:0]) begin
        image_2_98 <= io_pixelVal_in_2_3;
      end else if (10'h62 == _T_22[9:0]) begin
        image_2_98 <= io_pixelVal_in_2_2;
      end else if (10'h62 == _T_19[9:0]) begin
        image_2_98 <= io_pixelVal_in_2_1;
      end else if (10'h62 == _T_15[9:0]) begin
        image_2_98 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_99 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h63 == _T_37[9:0]) begin
        image_2_99 <= io_pixelVal_in_2_7;
      end else if (10'h63 == _T_34[9:0]) begin
        image_2_99 <= io_pixelVal_in_2_6;
      end else if (10'h63 == _T_31[9:0]) begin
        image_2_99 <= io_pixelVal_in_2_5;
      end else if (10'h63 == _T_28[9:0]) begin
        image_2_99 <= io_pixelVal_in_2_4;
      end else if (10'h63 == _T_25[9:0]) begin
        image_2_99 <= io_pixelVal_in_2_3;
      end else if (10'h63 == _T_22[9:0]) begin
        image_2_99 <= io_pixelVal_in_2_2;
      end else if (10'h63 == _T_19[9:0]) begin
        image_2_99 <= io_pixelVal_in_2_1;
      end else if (10'h63 == _T_15[9:0]) begin
        image_2_99 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_100 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h64 == _T_37[9:0]) begin
        image_2_100 <= io_pixelVal_in_2_7;
      end else if (10'h64 == _T_34[9:0]) begin
        image_2_100 <= io_pixelVal_in_2_6;
      end else if (10'h64 == _T_31[9:0]) begin
        image_2_100 <= io_pixelVal_in_2_5;
      end else if (10'h64 == _T_28[9:0]) begin
        image_2_100 <= io_pixelVal_in_2_4;
      end else if (10'h64 == _T_25[9:0]) begin
        image_2_100 <= io_pixelVal_in_2_3;
      end else if (10'h64 == _T_22[9:0]) begin
        image_2_100 <= io_pixelVal_in_2_2;
      end else if (10'h64 == _T_19[9:0]) begin
        image_2_100 <= io_pixelVal_in_2_1;
      end else if (10'h64 == _T_15[9:0]) begin
        image_2_100 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_101 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h65 == _T_37[9:0]) begin
        image_2_101 <= io_pixelVal_in_2_7;
      end else if (10'h65 == _T_34[9:0]) begin
        image_2_101 <= io_pixelVal_in_2_6;
      end else if (10'h65 == _T_31[9:0]) begin
        image_2_101 <= io_pixelVal_in_2_5;
      end else if (10'h65 == _T_28[9:0]) begin
        image_2_101 <= io_pixelVal_in_2_4;
      end else if (10'h65 == _T_25[9:0]) begin
        image_2_101 <= io_pixelVal_in_2_3;
      end else if (10'h65 == _T_22[9:0]) begin
        image_2_101 <= io_pixelVal_in_2_2;
      end else if (10'h65 == _T_19[9:0]) begin
        image_2_101 <= io_pixelVal_in_2_1;
      end else if (10'h65 == _T_15[9:0]) begin
        image_2_101 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_102 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h66 == _T_37[9:0]) begin
        image_2_102 <= io_pixelVal_in_2_7;
      end else if (10'h66 == _T_34[9:0]) begin
        image_2_102 <= io_pixelVal_in_2_6;
      end else if (10'h66 == _T_31[9:0]) begin
        image_2_102 <= io_pixelVal_in_2_5;
      end else if (10'h66 == _T_28[9:0]) begin
        image_2_102 <= io_pixelVal_in_2_4;
      end else if (10'h66 == _T_25[9:0]) begin
        image_2_102 <= io_pixelVal_in_2_3;
      end else if (10'h66 == _T_22[9:0]) begin
        image_2_102 <= io_pixelVal_in_2_2;
      end else if (10'h66 == _T_19[9:0]) begin
        image_2_102 <= io_pixelVal_in_2_1;
      end else if (10'h66 == _T_15[9:0]) begin
        image_2_102 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_103 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h67 == _T_37[9:0]) begin
        image_2_103 <= io_pixelVal_in_2_7;
      end else if (10'h67 == _T_34[9:0]) begin
        image_2_103 <= io_pixelVal_in_2_6;
      end else if (10'h67 == _T_31[9:0]) begin
        image_2_103 <= io_pixelVal_in_2_5;
      end else if (10'h67 == _T_28[9:0]) begin
        image_2_103 <= io_pixelVal_in_2_4;
      end else if (10'h67 == _T_25[9:0]) begin
        image_2_103 <= io_pixelVal_in_2_3;
      end else if (10'h67 == _T_22[9:0]) begin
        image_2_103 <= io_pixelVal_in_2_2;
      end else if (10'h67 == _T_19[9:0]) begin
        image_2_103 <= io_pixelVal_in_2_1;
      end else if (10'h67 == _T_15[9:0]) begin
        image_2_103 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_104 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h68 == _T_37[9:0]) begin
        image_2_104 <= io_pixelVal_in_2_7;
      end else if (10'h68 == _T_34[9:0]) begin
        image_2_104 <= io_pixelVal_in_2_6;
      end else if (10'h68 == _T_31[9:0]) begin
        image_2_104 <= io_pixelVal_in_2_5;
      end else if (10'h68 == _T_28[9:0]) begin
        image_2_104 <= io_pixelVal_in_2_4;
      end else if (10'h68 == _T_25[9:0]) begin
        image_2_104 <= io_pixelVal_in_2_3;
      end else if (10'h68 == _T_22[9:0]) begin
        image_2_104 <= io_pixelVal_in_2_2;
      end else if (10'h68 == _T_19[9:0]) begin
        image_2_104 <= io_pixelVal_in_2_1;
      end else if (10'h68 == _T_15[9:0]) begin
        image_2_104 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_105 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h69 == _T_37[9:0]) begin
        image_2_105 <= io_pixelVal_in_2_7;
      end else if (10'h69 == _T_34[9:0]) begin
        image_2_105 <= io_pixelVal_in_2_6;
      end else if (10'h69 == _T_31[9:0]) begin
        image_2_105 <= io_pixelVal_in_2_5;
      end else if (10'h69 == _T_28[9:0]) begin
        image_2_105 <= io_pixelVal_in_2_4;
      end else if (10'h69 == _T_25[9:0]) begin
        image_2_105 <= io_pixelVal_in_2_3;
      end else if (10'h69 == _T_22[9:0]) begin
        image_2_105 <= io_pixelVal_in_2_2;
      end else if (10'h69 == _T_19[9:0]) begin
        image_2_105 <= io_pixelVal_in_2_1;
      end else if (10'h69 == _T_15[9:0]) begin
        image_2_105 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_106 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6a == _T_37[9:0]) begin
        image_2_106 <= io_pixelVal_in_2_7;
      end else if (10'h6a == _T_34[9:0]) begin
        image_2_106 <= io_pixelVal_in_2_6;
      end else if (10'h6a == _T_31[9:0]) begin
        image_2_106 <= io_pixelVal_in_2_5;
      end else if (10'h6a == _T_28[9:0]) begin
        image_2_106 <= io_pixelVal_in_2_4;
      end else if (10'h6a == _T_25[9:0]) begin
        image_2_106 <= io_pixelVal_in_2_3;
      end else if (10'h6a == _T_22[9:0]) begin
        image_2_106 <= io_pixelVal_in_2_2;
      end else if (10'h6a == _T_19[9:0]) begin
        image_2_106 <= io_pixelVal_in_2_1;
      end else if (10'h6a == _T_15[9:0]) begin
        image_2_106 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_107 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6b == _T_37[9:0]) begin
        image_2_107 <= io_pixelVal_in_2_7;
      end else if (10'h6b == _T_34[9:0]) begin
        image_2_107 <= io_pixelVal_in_2_6;
      end else if (10'h6b == _T_31[9:0]) begin
        image_2_107 <= io_pixelVal_in_2_5;
      end else if (10'h6b == _T_28[9:0]) begin
        image_2_107 <= io_pixelVal_in_2_4;
      end else if (10'h6b == _T_25[9:0]) begin
        image_2_107 <= io_pixelVal_in_2_3;
      end else if (10'h6b == _T_22[9:0]) begin
        image_2_107 <= io_pixelVal_in_2_2;
      end else if (10'h6b == _T_19[9:0]) begin
        image_2_107 <= io_pixelVal_in_2_1;
      end else if (10'h6b == _T_15[9:0]) begin
        image_2_107 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_108 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6c == _T_37[9:0]) begin
        image_2_108 <= io_pixelVal_in_2_7;
      end else if (10'h6c == _T_34[9:0]) begin
        image_2_108 <= io_pixelVal_in_2_6;
      end else if (10'h6c == _T_31[9:0]) begin
        image_2_108 <= io_pixelVal_in_2_5;
      end else if (10'h6c == _T_28[9:0]) begin
        image_2_108 <= io_pixelVal_in_2_4;
      end else if (10'h6c == _T_25[9:0]) begin
        image_2_108 <= io_pixelVal_in_2_3;
      end else if (10'h6c == _T_22[9:0]) begin
        image_2_108 <= io_pixelVal_in_2_2;
      end else if (10'h6c == _T_19[9:0]) begin
        image_2_108 <= io_pixelVal_in_2_1;
      end else if (10'h6c == _T_15[9:0]) begin
        image_2_108 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_109 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6d == _T_37[9:0]) begin
        image_2_109 <= io_pixelVal_in_2_7;
      end else if (10'h6d == _T_34[9:0]) begin
        image_2_109 <= io_pixelVal_in_2_6;
      end else if (10'h6d == _T_31[9:0]) begin
        image_2_109 <= io_pixelVal_in_2_5;
      end else if (10'h6d == _T_28[9:0]) begin
        image_2_109 <= io_pixelVal_in_2_4;
      end else if (10'h6d == _T_25[9:0]) begin
        image_2_109 <= io_pixelVal_in_2_3;
      end else if (10'h6d == _T_22[9:0]) begin
        image_2_109 <= io_pixelVal_in_2_2;
      end else if (10'h6d == _T_19[9:0]) begin
        image_2_109 <= io_pixelVal_in_2_1;
      end else if (10'h6d == _T_15[9:0]) begin
        image_2_109 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_110 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6e == _T_37[9:0]) begin
        image_2_110 <= io_pixelVal_in_2_7;
      end else if (10'h6e == _T_34[9:0]) begin
        image_2_110 <= io_pixelVal_in_2_6;
      end else if (10'h6e == _T_31[9:0]) begin
        image_2_110 <= io_pixelVal_in_2_5;
      end else if (10'h6e == _T_28[9:0]) begin
        image_2_110 <= io_pixelVal_in_2_4;
      end else if (10'h6e == _T_25[9:0]) begin
        image_2_110 <= io_pixelVal_in_2_3;
      end else if (10'h6e == _T_22[9:0]) begin
        image_2_110 <= io_pixelVal_in_2_2;
      end else if (10'h6e == _T_19[9:0]) begin
        image_2_110 <= io_pixelVal_in_2_1;
      end else if (10'h6e == _T_15[9:0]) begin
        image_2_110 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_111 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6f == _T_37[9:0]) begin
        image_2_111 <= io_pixelVal_in_2_7;
      end else if (10'h6f == _T_34[9:0]) begin
        image_2_111 <= io_pixelVal_in_2_6;
      end else if (10'h6f == _T_31[9:0]) begin
        image_2_111 <= io_pixelVal_in_2_5;
      end else if (10'h6f == _T_28[9:0]) begin
        image_2_111 <= io_pixelVal_in_2_4;
      end else if (10'h6f == _T_25[9:0]) begin
        image_2_111 <= io_pixelVal_in_2_3;
      end else if (10'h6f == _T_22[9:0]) begin
        image_2_111 <= io_pixelVal_in_2_2;
      end else if (10'h6f == _T_19[9:0]) begin
        image_2_111 <= io_pixelVal_in_2_1;
      end else if (10'h6f == _T_15[9:0]) begin
        image_2_111 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_112 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h70 == _T_37[9:0]) begin
        image_2_112 <= io_pixelVal_in_2_7;
      end else if (10'h70 == _T_34[9:0]) begin
        image_2_112 <= io_pixelVal_in_2_6;
      end else if (10'h70 == _T_31[9:0]) begin
        image_2_112 <= io_pixelVal_in_2_5;
      end else if (10'h70 == _T_28[9:0]) begin
        image_2_112 <= io_pixelVal_in_2_4;
      end else if (10'h70 == _T_25[9:0]) begin
        image_2_112 <= io_pixelVal_in_2_3;
      end else if (10'h70 == _T_22[9:0]) begin
        image_2_112 <= io_pixelVal_in_2_2;
      end else if (10'h70 == _T_19[9:0]) begin
        image_2_112 <= io_pixelVal_in_2_1;
      end else if (10'h70 == _T_15[9:0]) begin
        image_2_112 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_113 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h71 == _T_37[9:0]) begin
        image_2_113 <= io_pixelVal_in_2_7;
      end else if (10'h71 == _T_34[9:0]) begin
        image_2_113 <= io_pixelVal_in_2_6;
      end else if (10'h71 == _T_31[9:0]) begin
        image_2_113 <= io_pixelVal_in_2_5;
      end else if (10'h71 == _T_28[9:0]) begin
        image_2_113 <= io_pixelVal_in_2_4;
      end else if (10'h71 == _T_25[9:0]) begin
        image_2_113 <= io_pixelVal_in_2_3;
      end else if (10'h71 == _T_22[9:0]) begin
        image_2_113 <= io_pixelVal_in_2_2;
      end else if (10'h71 == _T_19[9:0]) begin
        image_2_113 <= io_pixelVal_in_2_1;
      end else if (10'h71 == _T_15[9:0]) begin
        image_2_113 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_114 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h72 == _T_37[9:0]) begin
        image_2_114 <= io_pixelVal_in_2_7;
      end else if (10'h72 == _T_34[9:0]) begin
        image_2_114 <= io_pixelVal_in_2_6;
      end else if (10'h72 == _T_31[9:0]) begin
        image_2_114 <= io_pixelVal_in_2_5;
      end else if (10'h72 == _T_28[9:0]) begin
        image_2_114 <= io_pixelVal_in_2_4;
      end else if (10'h72 == _T_25[9:0]) begin
        image_2_114 <= io_pixelVal_in_2_3;
      end else if (10'h72 == _T_22[9:0]) begin
        image_2_114 <= io_pixelVal_in_2_2;
      end else if (10'h72 == _T_19[9:0]) begin
        image_2_114 <= io_pixelVal_in_2_1;
      end else if (10'h72 == _T_15[9:0]) begin
        image_2_114 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_115 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h73 == _T_37[9:0]) begin
        image_2_115 <= io_pixelVal_in_2_7;
      end else if (10'h73 == _T_34[9:0]) begin
        image_2_115 <= io_pixelVal_in_2_6;
      end else if (10'h73 == _T_31[9:0]) begin
        image_2_115 <= io_pixelVal_in_2_5;
      end else if (10'h73 == _T_28[9:0]) begin
        image_2_115 <= io_pixelVal_in_2_4;
      end else if (10'h73 == _T_25[9:0]) begin
        image_2_115 <= io_pixelVal_in_2_3;
      end else if (10'h73 == _T_22[9:0]) begin
        image_2_115 <= io_pixelVal_in_2_2;
      end else if (10'h73 == _T_19[9:0]) begin
        image_2_115 <= io_pixelVal_in_2_1;
      end else if (10'h73 == _T_15[9:0]) begin
        image_2_115 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_116 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h74 == _T_37[9:0]) begin
        image_2_116 <= io_pixelVal_in_2_7;
      end else if (10'h74 == _T_34[9:0]) begin
        image_2_116 <= io_pixelVal_in_2_6;
      end else if (10'h74 == _T_31[9:0]) begin
        image_2_116 <= io_pixelVal_in_2_5;
      end else if (10'h74 == _T_28[9:0]) begin
        image_2_116 <= io_pixelVal_in_2_4;
      end else if (10'h74 == _T_25[9:0]) begin
        image_2_116 <= io_pixelVal_in_2_3;
      end else if (10'h74 == _T_22[9:0]) begin
        image_2_116 <= io_pixelVal_in_2_2;
      end else if (10'h74 == _T_19[9:0]) begin
        image_2_116 <= io_pixelVal_in_2_1;
      end else if (10'h74 == _T_15[9:0]) begin
        image_2_116 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_117 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h75 == _T_37[9:0]) begin
        image_2_117 <= io_pixelVal_in_2_7;
      end else if (10'h75 == _T_34[9:0]) begin
        image_2_117 <= io_pixelVal_in_2_6;
      end else if (10'h75 == _T_31[9:0]) begin
        image_2_117 <= io_pixelVal_in_2_5;
      end else if (10'h75 == _T_28[9:0]) begin
        image_2_117 <= io_pixelVal_in_2_4;
      end else if (10'h75 == _T_25[9:0]) begin
        image_2_117 <= io_pixelVal_in_2_3;
      end else if (10'h75 == _T_22[9:0]) begin
        image_2_117 <= io_pixelVal_in_2_2;
      end else if (10'h75 == _T_19[9:0]) begin
        image_2_117 <= io_pixelVal_in_2_1;
      end else if (10'h75 == _T_15[9:0]) begin
        image_2_117 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_118 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h76 == _T_37[9:0]) begin
        image_2_118 <= io_pixelVal_in_2_7;
      end else if (10'h76 == _T_34[9:0]) begin
        image_2_118 <= io_pixelVal_in_2_6;
      end else if (10'h76 == _T_31[9:0]) begin
        image_2_118 <= io_pixelVal_in_2_5;
      end else if (10'h76 == _T_28[9:0]) begin
        image_2_118 <= io_pixelVal_in_2_4;
      end else if (10'h76 == _T_25[9:0]) begin
        image_2_118 <= io_pixelVal_in_2_3;
      end else if (10'h76 == _T_22[9:0]) begin
        image_2_118 <= io_pixelVal_in_2_2;
      end else if (10'h76 == _T_19[9:0]) begin
        image_2_118 <= io_pixelVal_in_2_1;
      end else if (10'h76 == _T_15[9:0]) begin
        image_2_118 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_119 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h77 == _T_37[9:0]) begin
        image_2_119 <= io_pixelVal_in_2_7;
      end else if (10'h77 == _T_34[9:0]) begin
        image_2_119 <= io_pixelVal_in_2_6;
      end else if (10'h77 == _T_31[9:0]) begin
        image_2_119 <= io_pixelVal_in_2_5;
      end else if (10'h77 == _T_28[9:0]) begin
        image_2_119 <= io_pixelVal_in_2_4;
      end else if (10'h77 == _T_25[9:0]) begin
        image_2_119 <= io_pixelVal_in_2_3;
      end else if (10'h77 == _T_22[9:0]) begin
        image_2_119 <= io_pixelVal_in_2_2;
      end else if (10'h77 == _T_19[9:0]) begin
        image_2_119 <= io_pixelVal_in_2_1;
      end else if (10'h77 == _T_15[9:0]) begin
        image_2_119 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_120 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h78 == _T_37[9:0]) begin
        image_2_120 <= io_pixelVal_in_2_7;
      end else if (10'h78 == _T_34[9:0]) begin
        image_2_120 <= io_pixelVal_in_2_6;
      end else if (10'h78 == _T_31[9:0]) begin
        image_2_120 <= io_pixelVal_in_2_5;
      end else if (10'h78 == _T_28[9:0]) begin
        image_2_120 <= io_pixelVal_in_2_4;
      end else if (10'h78 == _T_25[9:0]) begin
        image_2_120 <= io_pixelVal_in_2_3;
      end else if (10'h78 == _T_22[9:0]) begin
        image_2_120 <= io_pixelVal_in_2_2;
      end else if (10'h78 == _T_19[9:0]) begin
        image_2_120 <= io_pixelVal_in_2_1;
      end else if (10'h78 == _T_15[9:0]) begin
        image_2_120 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_121 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h79 == _T_37[9:0]) begin
        image_2_121 <= io_pixelVal_in_2_7;
      end else if (10'h79 == _T_34[9:0]) begin
        image_2_121 <= io_pixelVal_in_2_6;
      end else if (10'h79 == _T_31[9:0]) begin
        image_2_121 <= io_pixelVal_in_2_5;
      end else if (10'h79 == _T_28[9:0]) begin
        image_2_121 <= io_pixelVal_in_2_4;
      end else if (10'h79 == _T_25[9:0]) begin
        image_2_121 <= io_pixelVal_in_2_3;
      end else if (10'h79 == _T_22[9:0]) begin
        image_2_121 <= io_pixelVal_in_2_2;
      end else if (10'h79 == _T_19[9:0]) begin
        image_2_121 <= io_pixelVal_in_2_1;
      end else if (10'h79 == _T_15[9:0]) begin
        image_2_121 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_122 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7a == _T_37[9:0]) begin
        image_2_122 <= io_pixelVal_in_2_7;
      end else if (10'h7a == _T_34[9:0]) begin
        image_2_122 <= io_pixelVal_in_2_6;
      end else if (10'h7a == _T_31[9:0]) begin
        image_2_122 <= io_pixelVal_in_2_5;
      end else if (10'h7a == _T_28[9:0]) begin
        image_2_122 <= io_pixelVal_in_2_4;
      end else if (10'h7a == _T_25[9:0]) begin
        image_2_122 <= io_pixelVal_in_2_3;
      end else if (10'h7a == _T_22[9:0]) begin
        image_2_122 <= io_pixelVal_in_2_2;
      end else if (10'h7a == _T_19[9:0]) begin
        image_2_122 <= io_pixelVal_in_2_1;
      end else if (10'h7a == _T_15[9:0]) begin
        image_2_122 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_123 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7b == _T_37[9:0]) begin
        image_2_123 <= io_pixelVal_in_2_7;
      end else if (10'h7b == _T_34[9:0]) begin
        image_2_123 <= io_pixelVal_in_2_6;
      end else if (10'h7b == _T_31[9:0]) begin
        image_2_123 <= io_pixelVal_in_2_5;
      end else if (10'h7b == _T_28[9:0]) begin
        image_2_123 <= io_pixelVal_in_2_4;
      end else if (10'h7b == _T_25[9:0]) begin
        image_2_123 <= io_pixelVal_in_2_3;
      end else if (10'h7b == _T_22[9:0]) begin
        image_2_123 <= io_pixelVal_in_2_2;
      end else if (10'h7b == _T_19[9:0]) begin
        image_2_123 <= io_pixelVal_in_2_1;
      end else if (10'h7b == _T_15[9:0]) begin
        image_2_123 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_124 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7c == _T_37[9:0]) begin
        image_2_124 <= io_pixelVal_in_2_7;
      end else if (10'h7c == _T_34[9:0]) begin
        image_2_124 <= io_pixelVal_in_2_6;
      end else if (10'h7c == _T_31[9:0]) begin
        image_2_124 <= io_pixelVal_in_2_5;
      end else if (10'h7c == _T_28[9:0]) begin
        image_2_124 <= io_pixelVal_in_2_4;
      end else if (10'h7c == _T_25[9:0]) begin
        image_2_124 <= io_pixelVal_in_2_3;
      end else if (10'h7c == _T_22[9:0]) begin
        image_2_124 <= io_pixelVal_in_2_2;
      end else if (10'h7c == _T_19[9:0]) begin
        image_2_124 <= io_pixelVal_in_2_1;
      end else if (10'h7c == _T_15[9:0]) begin
        image_2_124 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_125 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7d == _T_37[9:0]) begin
        image_2_125 <= io_pixelVal_in_2_7;
      end else if (10'h7d == _T_34[9:0]) begin
        image_2_125 <= io_pixelVal_in_2_6;
      end else if (10'h7d == _T_31[9:0]) begin
        image_2_125 <= io_pixelVal_in_2_5;
      end else if (10'h7d == _T_28[9:0]) begin
        image_2_125 <= io_pixelVal_in_2_4;
      end else if (10'h7d == _T_25[9:0]) begin
        image_2_125 <= io_pixelVal_in_2_3;
      end else if (10'h7d == _T_22[9:0]) begin
        image_2_125 <= io_pixelVal_in_2_2;
      end else if (10'h7d == _T_19[9:0]) begin
        image_2_125 <= io_pixelVal_in_2_1;
      end else if (10'h7d == _T_15[9:0]) begin
        image_2_125 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_126 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7e == _T_37[9:0]) begin
        image_2_126 <= io_pixelVal_in_2_7;
      end else if (10'h7e == _T_34[9:0]) begin
        image_2_126 <= io_pixelVal_in_2_6;
      end else if (10'h7e == _T_31[9:0]) begin
        image_2_126 <= io_pixelVal_in_2_5;
      end else if (10'h7e == _T_28[9:0]) begin
        image_2_126 <= io_pixelVal_in_2_4;
      end else if (10'h7e == _T_25[9:0]) begin
        image_2_126 <= io_pixelVal_in_2_3;
      end else if (10'h7e == _T_22[9:0]) begin
        image_2_126 <= io_pixelVal_in_2_2;
      end else if (10'h7e == _T_19[9:0]) begin
        image_2_126 <= io_pixelVal_in_2_1;
      end else if (10'h7e == _T_15[9:0]) begin
        image_2_126 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_127 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7f == _T_37[9:0]) begin
        image_2_127 <= io_pixelVal_in_2_7;
      end else if (10'h7f == _T_34[9:0]) begin
        image_2_127 <= io_pixelVal_in_2_6;
      end else if (10'h7f == _T_31[9:0]) begin
        image_2_127 <= io_pixelVal_in_2_5;
      end else if (10'h7f == _T_28[9:0]) begin
        image_2_127 <= io_pixelVal_in_2_4;
      end else if (10'h7f == _T_25[9:0]) begin
        image_2_127 <= io_pixelVal_in_2_3;
      end else if (10'h7f == _T_22[9:0]) begin
        image_2_127 <= io_pixelVal_in_2_2;
      end else if (10'h7f == _T_19[9:0]) begin
        image_2_127 <= io_pixelVal_in_2_1;
      end else if (10'h7f == _T_15[9:0]) begin
        image_2_127 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_128 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h80 == _T_37[9:0]) begin
        image_2_128 <= io_pixelVal_in_2_7;
      end else if (10'h80 == _T_34[9:0]) begin
        image_2_128 <= io_pixelVal_in_2_6;
      end else if (10'h80 == _T_31[9:0]) begin
        image_2_128 <= io_pixelVal_in_2_5;
      end else if (10'h80 == _T_28[9:0]) begin
        image_2_128 <= io_pixelVal_in_2_4;
      end else if (10'h80 == _T_25[9:0]) begin
        image_2_128 <= io_pixelVal_in_2_3;
      end else if (10'h80 == _T_22[9:0]) begin
        image_2_128 <= io_pixelVal_in_2_2;
      end else if (10'h80 == _T_19[9:0]) begin
        image_2_128 <= io_pixelVal_in_2_1;
      end else if (10'h80 == _T_15[9:0]) begin
        image_2_128 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_129 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h81 == _T_37[9:0]) begin
        image_2_129 <= io_pixelVal_in_2_7;
      end else if (10'h81 == _T_34[9:0]) begin
        image_2_129 <= io_pixelVal_in_2_6;
      end else if (10'h81 == _T_31[9:0]) begin
        image_2_129 <= io_pixelVal_in_2_5;
      end else if (10'h81 == _T_28[9:0]) begin
        image_2_129 <= io_pixelVal_in_2_4;
      end else if (10'h81 == _T_25[9:0]) begin
        image_2_129 <= io_pixelVal_in_2_3;
      end else if (10'h81 == _T_22[9:0]) begin
        image_2_129 <= io_pixelVal_in_2_2;
      end else if (10'h81 == _T_19[9:0]) begin
        image_2_129 <= io_pixelVal_in_2_1;
      end else if (10'h81 == _T_15[9:0]) begin
        image_2_129 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_130 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h82 == _T_37[9:0]) begin
        image_2_130 <= io_pixelVal_in_2_7;
      end else if (10'h82 == _T_34[9:0]) begin
        image_2_130 <= io_pixelVal_in_2_6;
      end else if (10'h82 == _T_31[9:0]) begin
        image_2_130 <= io_pixelVal_in_2_5;
      end else if (10'h82 == _T_28[9:0]) begin
        image_2_130 <= io_pixelVal_in_2_4;
      end else if (10'h82 == _T_25[9:0]) begin
        image_2_130 <= io_pixelVal_in_2_3;
      end else if (10'h82 == _T_22[9:0]) begin
        image_2_130 <= io_pixelVal_in_2_2;
      end else if (10'h82 == _T_19[9:0]) begin
        image_2_130 <= io_pixelVal_in_2_1;
      end else if (10'h82 == _T_15[9:0]) begin
        image_2_130 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_131 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h83 == _T_37[9:0]) begin
        image_2_131 <= io_pixelVal_in_2_7;
      end else if (10'h83 == _T_34[9:0]) begin
        image_2_131 <= io_pixelVal_in_2_6;
      end else if (10'h83 == _T_31[9:0]) begin
        image_2_131 <= io_pixelVal_in_2_5;
      end else if (10'h83 == _T_28[9:0]) begin
        image_2_131 <= io_pixelVal_in_2_4;
      end else if (10'h83 == _T_25[9:0]) begin
        image_2_131 <= io_pixelVal_in_2_3;
      end else if (10'h83 == _T_22[9:0]) begin
        image_2_131 <= io_pixelVal_in_2_2;
      end else if (10'h83 == _T_19[9:0]) begin
        image_2_131 <= io_pixelVal_in_2_1;
      end else if (10'h83 == _T_15[9:0]) begin
        image_2_131 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_132 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h84 == _T_37[9:0]) begin
        image_2_132 <= io_pixelVal_in_2_7;
      end else if (10'h84 == _T_34[9:0]) begin
        image_2_132 <= io_pixelVal_in_2_6;
      end else if (10'h84 == _T_31[9:0]) begin
        image_2_132 <= io_pixelVal_in_2_5;
      end else if (10'h84 == _T_28[9:0]) begin
        image_2_132 <= io_pixelVal_in_2_4;
      end else if (10'h84 == _T_25[9:0]) begin
        image_2_132 <= io_pixelVal_in_2_3;
      end else if (10'h84 == _T_22[9:0]) begin
        image_2_132 <= io_pixelVal_in_2_2;
      end else if (10'h84 == _T_19[9:0]) begin
        image_2_132 <= io_pixelVal_in_2_1;
      end else if (10'h84 == _T_15[9:0]) begin
        image_2_132 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_133 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h85 == _T_37[9:0]) begin
        image_2_133 <= io_pixelVal_in_2_7;
      end else if (10'h85 == _T_34[9:0]) begin
        image_2_133 <= io_pixelVal_in_2_6;
      end else if (10'h85 == _T_31[9:0]) begin
        image_2_133 <= io_pixelVal_in_2_5;
      end else if (10'h85 == _T_28[9:0]) begin
        image_2_133 <= io_pixelVal_in_2_4;
      end else if (10'h85 == _T_25[9:0]) begin
        image_2_133 <= io_pixelVal_in_2_3;
      end else if (10'h85 == _T_22[9:0]) begin
        image_2_133 <= io_pixelVal_in_2_2;
      end else if (10'h85 == _T_19[9:0]) begin
        image_2_133 <= io_pixelVal_in_2_1;
      end else if (10'h85 == _T_15[9:0]) begin
        image_2_133 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_134 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h86 == _T_37[9:0]) begin
        image_2_134 <= io_pixelVal_in_2_7;
      end else if (10'h86 == _T_34[9:0]) begin
        image_2_134 <= io_pixelVal_in_2_6;
      end else if (10'h86 == _T_31[9:0]) begin
        image_2_134 <= io_pixelVal_in_2_5;
      end else if (10'h86 == _T_28[9:0]) begin
        image_2_134 <= io_pixelVal_in_2_4;
      end else if (10'h86 == _T_25[9:0]) begin
        image_2_134 <= io_pixelVal_in_2_3;
      end else if (10'h86 == _T_22[9:0]) begin
        image_2_134 <= io_pixelVal_in_2_2;
      end else if (10'h86 == _T_19[9:0]) begin
        image_2_134 <= io_pixelVal_in_2_1;
      end else if (10'h86 == _T_15[9:0]) begin
        image_2_134 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_135 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h87 == _T_37[9:0]) begin
        image_2_135 <= io_pixelVal_in_2_7;
      end else if (10'h87 == _T_34[9:0]) begin
        image_2_135 <= io_pixelVal_in_2_6;
      end else if (10'h87 == _T_31[9:0]) begin
        image_2_135 <= io_pixelVal_in_2_5;
      end else if (10'h87 == _T_28[9:0]) begin
        image_2_135 <= io_pixelVal_in_2_4;
      end else if (10'h87 == _T_25[9:0]) begin
        image_2_135 <= io_pixelVal_in_2_3;
      end else if (10'h87 == _T_22[9:0]) begin
        image_2_135 <= io_pixelVal_in_2_2;
      end else if (10'h87 == _T_19[9:0]) begin
        image_2_135 <= io_pixelVal_in_2_1;
      end else if (10'h87 == _T_15[9:0]) begin
        image_2_135 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_136 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h88 == _T_37[9:0]) begin
        image_2_136 <= io_pixelVal_in_2_7;
      end else if (10'h88 == _T_34[9:0]) begin
        image_2_136 <= io_pixelVal_in_2_6;
      end else if (10'h88 == _T_31[9:0]) begin
        image_2_136 <= io_pixelVal_in_2_5;
      end else if (10'h88 == _T_28[9:0]) begin
        image_2_136 <= io_pixelVal_in_2_4;
      end else if (10'h88 == _T_25[9:0]) begin
        image_2_136 <= io_pixelVal_in_2_3;
      end else if (10'h88 == _T_22[9:0]) begin
        image_2_136 <= io_pixelVal_in_2_2;
      end else if (10'h88 == _T_19[9:0]) begin
        image_2_136 <= io_pixelVal_in_2_1;
      end else if (10'h88 == _T_15[9:0]) begin
        image_2_136 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_137 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h89 == _T_37[9:0]) begin
        image_2_137 <= io_pixelVal_in_2_7;
      end else if (10'h89 == _T_34[9:0]) begin
        image_2_137 <= io_pixelVal_in_2_6;
      end else if (10'h89 == _T_31[9:0]) begin
        image_2_137 <= io_pixelVal_in_2_5;
      end else if (10'h89 == _T_28[9:0]) begin
        image_2_137 <= io_pixelVal_in_2_4;
      end else if (10'h89 == _T_25[9:0]) begin
        image_2_137 <= io_pixelVal_in_2_3;
      end else if (10'h89 == _T_22[9:0]) begin
        image_2_137 <= io_pixelVal_in_2_2;
      end else if (10'h89 == _T_19[9:0]) begin
        image_2_137 <= io_pixelVal_in_2_1;
      end else if (10'h89 == _T_15[9:0]) begin
        image_2_137 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_138 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8a == _T_37[9:0]) begin
        image_2_138 <= io_pixelVal_in_2_7;
      end else if (10'h8a == _T_34[9:0]) begin
        image_2_138 <= io_pixelVal_in_2_6;
      end else if (10'h8a == _T_31[9:0]) begin
        image_2_138 <= io_pixelVal_in_2_5;
      end else if (10'h8a == _T_28[9:0]) begin
        image_2_138 <= io_pixelVal_in_2_4;
      end else if (10'h8a == _T_25[9:0]) begin
        image_2_138 <= io_pixelVal_in_2_3;
      end else if (10'h8a == _T_22[9:0]) begin
        image_2_138 <= io_pixelVal_in_2_2;
      end else if (10'h8a == _T_19[9:0]) begin
        image_2_138 <= io_pixelVal_in_2_1;
      end else if (10'h8a == _T_15[9:0]) begin
        image_2_138 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_139 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8b == _T_37[9:0]) begin
        image_2_139 <= io_pixelVal_in_2_7;
      end else if (10'h8b == _T_34[9:0]) begin
        image_2_139 <= io_pixelVal_in_2_6;
      end else if (10'h8b == _T_31[9:0]) begin
        image_2_139 <= io_pixelVal_in_2_5;
      end else if (10'h8b == _T_28[9:0]) begin
        image_2_139 <= io_pixelVal_in_2_4;
      end else if (10'h8b == _T_25[9:0]) begin
        image_2_139 <= io_pixelVal_in_2_3;
      end else if (10'h8b == _T_22[9:0]) begin
        image_2_139 <= io_pixelVal_in_2_2;
      end else if (10'h8b == _T_19[9:0]) begin
        image_2_139 <= io_pixelVal_in_2_1;
      end else if (10'h8b == _T_15[9:0]) begin
        image_2_139 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_140 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8c == _T_37[9:0]) begin
        image_2_140 <= io_pixelVal_in_2_7;
      end else if (10'h8c == _T_34[9:0]) begin
        image_2_140 <= io_pixelVal_in_2_6;
      end else if (10'h8c == _T_31[9:0]) begin
        image_2_140 <= io_pixelVal_in_2_5;
      end else if (10'h8c == _T_28[9:0]) begin
        image_2_140 <= io_pixelVal_in_2_4;
      end else if (10'h8c == _T_25[9:0]) begin
        image_2_140 <= io_pixelVal_in_2_3;
      end else if (10'h8c == _T_22[9:0]) begin
        image_2_140 <= io_pixelVal_in_2_2;
      end else if (10'h8c == _T_19[9:0]) begin
        image_2_140 <= io_pixelVal_in_2_1;
      end else if (10'h8c == _T_15[9:0]) begin
        image_2_140 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_141 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8d == _T_37[9:0]) begin
        image_2_141 <= io_pixelVal_in_2_7;
      end else if (10'h8d == _T_34[9:0]) begin
        image_2_141 <= io_pixelVal_in_2_6;
      end else if (10'h8d == _T_31[9:0]) begin
        image_2_141 <= io_pixelVal_in_2_5;
      end else if (10'h8d == _T_28[9:0]) begin
        image_2_141 <= io_pixelVal_in_2_4;
      end else if (10'h8d == _T_25[9:0]) begin
        image_2_141 <= io_pixelVal_in_2_3;
      end else if (10'h8d == _T_22[9:0]) begin
        image_2_141 <= io_pixelVal_in_2_2;
      end else if (10'h8d == _T_19[9:0]) begin
        image_2_141 <= io_pixelVal_in_2_1;
      end else if (10'h8d == _T_15[9:0]) begin
        image_2_141 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_142 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8e == _T_37[9:0]) begin
        image_2_142 <= io_pixelVal_in_2_7;
      end else if (10'h8e == _T_34[9:0]) begin
        image_2_142 <= io_pixelVal_in_2_6;
      end else if (10'h8e == _T_31[9:0]) begin
        image_2_142 <= io_pixelVal_in_2_5;
      end else if (10'h8e == _T_28[9:0]) begin
        image_2_142 <= io_pixelVal_in_2_4;
      end else if (10'h8e == _T_25[9:0]) begin
        image_2_142 <= io_pixelVal_in_2_3;
      end else if (10'h8e == _T_22[9:0]) begin
        image_2_142 <= io_pixelVal_in_2_2;
      end else if (10'h8e == _T_19[9:0]) begin
        image_2_142 <= io_pixelVal_in_2_1;
      end else if (10'h8e == _T_15[9:0]) begin
        image_2_142 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_143 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8f == _T_37[9:0]) begin
        image_2_143 <= io_pixelVal_in_2_7;
      end else if (10'h8f == _T_34[9:0]) begin
        image_2_143 <= io_pixelVal_in_2_6;
      end else if (10'h8f == _T_31[9:0]) begin
        image_2_143 <= io_pixelVal_in_2_5;
      end else if (10'h8f == _T_28[9:0]) begin
        image_2_143 <= io_pixelVal_in_2_4;
      end else if (10'h8f == _T_25[9:0]) begin
        image_2_143 <= io_pixelVal_in_2_3;
      end else if (10'h8f == _T_22[9:0]) begin
        image_2_143 <= io_pixelVal_in_2_2;
      end else if (10'h8f == _T_19[9:0]) begin
        image_2_143 <= io_pixelVal_in_2_1;
      end else if (10'h8f == _T_15[9:0]) begin
        image_2_143 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_144 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h90 == _T_37[9:0]) begin
        image_2_144 <= io_pixelVal_in_2_7;
      end else if (10'h90 == _T_34[9:0]) begin
        image_2_144 <= io_pixelVal_in_2_6;
      end else if (10'h90 == _T_31[9:0]) begin
        image_2_144 <= io_pixelVal_in_2_5;
      end else if (10'h90 == _T_28[9:0]) begin
        image_2_144 <= io_pixelVal_in_2_4;
      end else if (10'h90 == _T_25[9:0]) begin
        image_2_144 <= io_pixelVal_in_2_3;
      end else if (10'h90 == _T_22[9:0]) begin
        image_2_144 <= io_pixelVal_in_2_2;
      end else if (10'h90 == _T_19[9:0]) begin
        image_2_144 <= io_pixelVal_in_2_1;
      end else if (10'h90 == _T_15[9:0]) begin
        image_2_144 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_145 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h91 == _T_37[9:0]) begin
        image_2_145 <= io_pixelVal_in_2_7;
      end else if (10'h91 == _T_34[9:0]) begin
        image_2_145 <= io_pixelVal_in_2_6;
      end else if (10'h91 == _T_31[9:0]) begin
        image_2_145 <= io_pixelVal_in_2_5;
      end else if (10'h91 == _T_28[9:0]) begin
        image_2_145 <= io_pixelVal_in_2_4;
      end else if (10'h91 == _T_25[9:0]) begin
        image_2_145 <= io_pixelVal_in_2_3;
      end else if (10'h91 == _T_22[9:0]) begin
        image_2_145 <= io_pixelVal_in_2_2;
      end else if (10'h91 == _T_19[9:0]) begin
        image_2_145 <= io_pixelVal_in_2_1;
      end else if (10'h91 == _T_15[9:0]) begin
        image_2_145 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_146 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h92 == _T_37[9:0]) begin
        image_2_146 <= io_pixelVal_in_2_7;
      end else if (10'h92 == _T_34[9:0]) begin
        image_2_146 <= io_pixelVal_in_2_6;
      end else if (10'h92 == _T_31[9:0]) begin
        image_2_146 <= io_pixelVal_in_2_5;
      end else if (10'h92 == _T_28[9:0]) begin
        image_2_146 <= io_pixelVal_in_2_4;
      end else if (10'h92 == _T_25[9:0]) begin
        image_2_146 <= io_pixelVal_in_2_3;
      end else if (10'h92 == _T_22[9:0]) begin
        image_2_146 <= io_pixelVal_in_2_2;
      end else if (10'h92 == _T_19[9:0]) begin
        image_2_146 <= io_pixelVal_in_2_1;
      end else if (10'h92 == _T_15[9:0]) begin
        image_2_146 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_147 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h93 == _T_37[9:0]) begin
        image_2_147 <= io_pixelVal_in_2_7;
      end else if (10'h93 == _T_34[9:0]) begin
        image_2_147 <= io_pixelVal_in_2_6;
      end else if (10'h93 == _T_31[9:0]) begin
        image_2_147 <= io_pixelVal_in_2_5;
      end else if (10'h93 == _T_28[9:0]) begin
        image_2_147 <= io_pixelVal_in_2_4;
      end else if (10'h93 == _T_25[9:0]) begin
        image_2_147 <= io_pixelVal_in_2_3;
      end else if (10'h93 == _T_22[9:0]) begin
        image_2_147 <= io_pixelVal_in_2_2;
      end else if (10'h93 == _T_19[9:0]) begin
        image_2_147 <= io_pixelVal_in_2_1;
      end else if (10'h93 == _T_15[9:0]) begin
        image_2_147 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_148 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h94 == _T_37[9:0]) begin
        image_2_148 <= io_pixelVal_in_2_7;
      end else if (10'h94 == _T_34[9:0]) begin
        image_2_148 <= io_pixelVal_in_2_6;
      end else if (10'h94 == _T_31[9:0]) begin
        image_2_148 <= io_pixelVal_in_2_5;
      end else if (10'h94 == _T_28[9:0]) begin
        image_2_148 <= io_pixelVal_in_2_4;
      end else if (10'h94 == _T_25[9:0]) begin
        image_2_148 <= io_pixelVal_in_2_3;
      end else if (10'h94 == _T_22[9:0]) begin
        image_2_148 <= io_pixelVal_in_2_2;
      end else if (10'h94 == _T_19[9:0]) begin
        image_2_148 <= io_pixelVal_in_2_1;
      end else if (10'h94 == _T_15[9:0]) begin
        image_2_148 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_149 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h95 == _T_37[9:0]) begin
        image_2_149 <= io_pixelVal_in_2_7;
      end else if (10'h95 == _T_34[9:0]) begin
        image_2_149 <= io_pixelVal_in_2_6;
      end else if (10'h95 == _T_31[9:0]) begin
        image_2_149 <= io_pixelVal_in_2_5;
      end else if (10'h95 == _T_28[9:0]) begin
        image_2_149 <= io_pixelVal_in_2_4;
      end else if (10'h95 == _T_25[9:0]) begin
        image_2_149 <= io_pixelVal_in_2_3;
      end else if (10'h95 == _T_22[9:0]) begin
        image_2_149 <= io_pixelVal_in_2_2;
      end else if (10'h95 == _T_19[9:0]) begin
        image_2_149 <= io_pixelVal_in_2_1;
      end else if (10'h95 == _T_15[9:0]) begin
        image_2_149 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_150 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h96 == _T_37[9:0]) begin
        image_2_150 <= io_pixelVal_in_2_7;
      end else if (10'h96 == _T_34[9:0]) begin
        image_2_150 <= io_pixelVal_in_2_6;
      end else if (10'h96 == _T_31[9:0]) begin
        image_2_150 <= io_pixelVal_in_2_5;
      end else if (10'h96 == _T_28[9:0]) begin
        image_2_150 <= io_pixelVal_in_2_4;
      end else if (10'h96 == _T_25[9:0]) begin
        image_2_150 <= io_pixelVal_in_2_3;
      end else if (10'h96 == _T_22[9:0]) begin
        image_2_150 <= io_pixelVal_in_2_2;
      end else if (10'h96 == _T_19[9:0]) begin
        image_2_150 <= io_pixelVal_in_2_1;
      end else if (10'h96 == _T_15[9:0]) begin
        image_2_150 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_151 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h97 == _T_37[9:0]) begin
        image_2_151 <= io_pixelVal_in_2_7;
      end else if (10'h97 == _T_34[9:0]) begin
        image_2_151 <= io_pixelVal_in_2_6;
      end else if (10'h97 == _T_31[9:0]) begin
        image_2_151 <= io_pixelVal_in_2_5;
      end else if (10'h97 == _T_28[9:0]) begin
        image_2_151 <= io_pixelVal_in_2_4;
      end else if (10'h97 == _T_25[9:0]) begin
        image_2_151 <= io_pixelVal_in_2_3;
      end else if (10'h97 == _T_22[9:0]) begin
        image_2_151 <= io_pixelVal_in_2_2;
      end else if (10'h97 == _T_19[9:0]) begin
        image_2_151 <= io_pixelVal_in_2_1;
      end else if (10'h97 == _T_15[9:0]) begin
        image_2_151 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_152 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h98 == _T_37[9:0]) begin
        image_2_152 <= io_pixelVal_in_2_7;
      end else if (10'h98 == _T_34[9:0]) begin
        image_2_152 <= io_pixelVal_in_2_6;
      end else if (10'h98 == _T_31[9:0]) begin
        image_2_152 <= io_pixelVal_in_2_5;
      end else if (10'h98 == _T_28[9:0]) begin
        image_2_152 <= io_pixelVal_in_2_4;
      end else if (10'h98 == _T_25[9:0]) begin
        image_2_152 <= io_pixelVal_in_2_3;
      end else if (10'h98 == _T_22[9:0]) begin
        image_2_152 <= io_pixelVal_in_2_2;
      end else if (10'h98 == _T_19[9:0]) begin
        image_2_152 <= io_pixelVal_in_2_1;
      end else if (10'h98 == _T_15[9:0]) begin
        image_2_152 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_153 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h99 == _T_37[9:0]) begin
        image_2_153 <= io_pixelVal_in_2_7;
      end else if (10'h99 == _T_34[9:0]) begin
        image_2_153 <= io_pixelVal_in_2_6;
      end else if (10'h99 == _T_31[9:0]) begin
        image_2_153 <= io_pixelVal_in_2_5;
      end else if (10'h99 == _T_28[9:0]) begin
        image_2_153 <= io_pixelVal_in_2_4;
      end else if (10'h99 == _T_25[9:0]) begin
        image_2_153 <= io_pixelVal_in_2_3;
      end else if (10'h99 == _T_22[9:0]) begin
        image_2_153 <= io_pixelVal_in_2_2;
      end else if (10'h99 == _T_19[9:0]) begin
        image_2_153 <= io_pixelVal_in_2_1;
      end else if (10'h99 == _T_15[9:0]) begin
        image_2_153 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_154 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9a == _T_37[9:0]) begin
        image_2_154 <= io_pixelVal_in_2_7;
      end else if (10'h9a == _T_34[9:0]) begin
        image_2_154 <= io_pixelVal_in_2_6;
      end else if (10'h9a == _T_31[9:0]) begin
        image_2_154 <= io_pixelVal_in_2_5;
      end else if (10'h9a == _T_28[9:0]) begin
        image_2_154 <= io_pixelVal_in_2_4;
      end else if (10'h9a == _T_25[9:0]) begin
        image_2_154 <= io_pixelVal_in_2_3;
      end else if (10'h9a == _T_22[9:0]) begin
        image_2_154 <= io_pixelVal_in_2_2;
      end else if (10'h9a == _T_19[9:0]) begin
        image_2_154 <= io_pixelVal_in_2_1;
      end else if (10'h9a == _T_15[9:0]) begin
        image_2_154 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_155 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9b == _T_37[9:0]) begin
        image_2_155 <= io_pixelVal_in_2_7;
      end else if (10'h9b == _T_34[9:0]) begin
        image_2_155 <= io_pixelVal_in_2_6;
      end else if (10'h9b == _T_31[9:0]) begin
        image_2_155 <= io_pixelVal_in_2_5;
      end else if (10'h9b == _T_28[9:0]) begin
        image_2_155 <= io_pixelVal_in_2_4;
      end else if (10'h9b == _T_25[9:0]) begin
        image_2_155 <= io_pixelVal_in_2_3;
      end else if (10'h9b == _T_22[9:0]) begin
        image_2_155 <= io_pixelVal_in_2_2;
      end else if (10'h9b == _T_19[9:0]) begin
        image_2_155 <= io_pixelVal_in_2_1;
      end else if (10'h9b == _T_15[9:0]) begin
        image_2_155 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_156 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9c == _T_37[9:0]) begin
        image_2_156 <= io_pixelVal_in_2_7;
      end else if (10'h9c == _T_34[9:0]) begin
        image_2_156 <= io_pixelVal_in_2_6;
      end else if (10'h9c == _T_31[9:0]) begin
        image_2_156 <= io_pixelVal_in_2_5;
      end else if (10'h9c == _T_28[9:0]) begin
        image_2_156 <= io_pixelVal_in_2_4;
      end else if (10'h9c == _T_25[9:0]) begin
        image_2_156 <= io_pixelVal_in_2_3;
      end else if (10'h9c == _T_22[9:0]) begin
        image_2_156 <= io_pixelVal_in_2_2;
      end else if (10'h9c == _T_19[9:0]) begin
        image_2_156 <= io_pixelVal_in_2_1;
      end else if (10'h9c == _T_15[9:0]) begin
        image_2_156 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_157 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9d == _T_37[9:0]) begin
        image_2_157 <= io_pixelVal_in_2_7;
      end else if (10'h9d == _T_34[9:0]) begin
        image_2_157 <= io_pixelVal_in_2_6;
      end else if (10'h9d == _T_31[9:0]) begin
        image_2_157 <= io_pixelVal_in_2_5;
      end else if (10'h9d == _T_28[9:0]) begin
        image_2_157 <= io_pixelVal_in_2_4;
      end else if (10'h9d == _T_25[9:0]) begin
        image_2_157 <= io_pixelVal_in_2_3;
      end else if (10'h9d == _T_22[9:0]) begin
        image_2_157 <= io_pixelVal_in_2_2;
      end else if (10'h9d == _T_19[9:0]) begin
        image_2_157 <= io_pixelVal_in_2_1;
      end else if (10'h9d == _T_15[9:0]) begin
        image_2_157 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_158 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9e == _T_37[9:0]) begin
        image_2_158 <= io_pixelVal_in_2_7;
      end else if (10'h9e == _T_34[9:0]) begin
        image_2_158 <= io_pixelVal_in_2_6;
      end else if (10'h9e == _T_31[9:0]) begin
        image_2_158 <= io_pixelVal_in_2_5;
      end else if (10'h9e == _T_28[9:0]) begin
        image_2_158 <= io_pixelVal_in_2_4;
      end else if (10'h9e == _T_25[9:0]) begin
        image_2_158 <= io_pixelVal_in_2_3;
      end else if (10'h9e == _T_22[9:0]) begin
        image_2_158 <= io_pixelVal_in_2_2;
      end else if (10'h9e == _T_19[9:0]) begin
        image_2_158 <= io_pixelVal_in_2_1;
      end else if (10'h9e == _T_15[9:0]) begin
        image_2_158 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_159 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9f == _T_37[9:0]) begin
        image_2_159 <= io_pixelVal_in_2_7;
      end else if (10'h9f == _T_34[9:0]) begin
        image_2_159 <= io_pixelVal_in_2_6;
      end else if (10'h9f == _T_31[9:0]) begin
        image_2_159 <= io_pixelVal_in_2_5;
      end else if (10'h9f == _T_28[9:0]) begin
        image_2_159 <= io_pixelVal_in_2_4;
      end else if (10'h9f == _T_25[9:0]) begin
        image_2_159 <= io_pixelVal_in_2_3;
      end else if (10'h9f == _T_22[9:0]) begin
        image_2_159 <= io_pixelVal_in_2_2;
      end else if (10'h9f == _T_19[9:0]) begin
        image_2_159 <= io_pixelVal_in_2_1;
      end else if (10'h9f == _T_15[9:0]) begin
        image_2_159 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_160 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha0 == _T_37[9:0]) begin
        image_2_160 <= io_pixelVal_in_2_7;
      end else if (10'ha0 == _T_34[9:0]) begin
        image_2_160 <= io_pixelVal_in_2_6;
      end else if (10'ha0 == _T_31[9:0]) begin
        image_2_160 <= io_pixelVal_in_2_5;
      end else if (10'ha0 == _T_28[9:0]) begin
        image_2_160 <= io_pixelVal_in_2_4;
      end else if (10'ha0 == _T_25[9:0]) begin
        image_2_160 <= io_pixelVal_in_2_3;
      end else if (10'ha0 == _T_22[9:0]) begin
        image_2_160 <= io_pixelVal_in_2_2;
      end else if (10'ha0 == _T_19[9:0]) begin
        image_2_160 <= io_pixelVal_in_2_1;
      end else if (10'ha0 == _T_15[9:0]) begin
        image_2_160 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_161 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha1 == _T_37[9:0]) begin
        image_2_161 <= io_pixelVal_in_2_7;
      end else if (10'ha1 == _T_34[9:0]) begin
        image_2_161 <= io_pixelVal_in_2_6;
      end else if (10'ha1 == _T_31[9:0]) begin
        image_2_161 <= io_pixelVal_in_2_5;
      end else if (10'ha1 == _T_28[9:0]) begin
        image_2_161 <= io_pixelVal_in_2_4;
      end else if (10'ha1 == _T_25[9:0]) begin
        image_2_161 <= io_pixelVal_in_2_3;
      end else if (10'ha1 == _T_22[9:0]) begin
        image_2_161 <= io_pixelVal_in_2_2;
      end else if (10'ha1 == _T_19[9:0]) begin
        image_2_161 <= io_pixelVal_in_2_1;
      end else if (10'ha1 == _T_15[9:0]) begin
        image_2_161 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_162 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha2 == _T_37[9:0]) begin
        image_2_162 <= io_pixelVal_in_2_7;
      end else if (10'ha2 == _T_34[9:0]) begin
        image_2_162 <= io_pixelVal_in_2_6;
      end else if (10'ha2 == _T_31[9:0]) begin
        image_2_162 <= io_pixelVal_in_2_5;
      end else if (10'ha2 == _T_28[9:0]) begin
        image_2_162 <= io_pixelVal_in_2_4;
      end else if (10'ha2 == _T_25[9:0]) begin
        image_2_162 <= io_pixelVal_in_2_3;
      end else if (10'ha2 == _T_22[9:0]) begin
        image_2_162 <= io_pixelVal_in_2_2;
      end else if (10'ha2 == _T_19[9:0]) begin
        image_2_162 <= io_pixelVal_in_2_1;
      end else if (10'ha2 == _T_15[9:0]) begin
        image_2_162 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_163 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha3 == _T_37[9:0]) begin
        image_2_163 <= io_pixelVal_in_2_7;
      end else if (10'ha3 == _T_34[9:0]) begin
        image_2_163 <= io_pixelVal_in_2_6;
      end else if (10'ha3 == _T_31[9:0]) begin
        image_2_163 <= io_pixelVal_in_2_5;
      end else if (10'ha3 == _T_28[9:0]) begin
        image_2_163 <= io_pixelVal_in_2_4;
      end else if (10'ha3 == _T_25[9:0]) begin
        image_2_163 <= io_pixelVal_in_2_3;
      end else if (10'ha3 == _T_22[9:0]) begin
        image_2_163 <= io_pixelVal_in_2_2;
      end else if (10'ha3 == _T_19[9:0]) begin
        image_2_163 <= io_pixelVal_in_2_1;
      end else if (10'ha3 == _T_15[9:0]) begin
        image_2_163 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_164 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha4 == _T_37[9:0]) begin
        image_2_164 <= io_pixelVal_in_2_7;
      end else if (10'ha4 == _T_34[9:0]) begin
        image_2_164 <= io_pixelVal_in_2_6;
      end else if (10'ha4 == _T_31[9:0]) begin
        image_2_164 <= io_pixelVal_in_2_5;
      end else if (10'ha4 == _T_28[9:0]) begin
        image_2_164 <= io_pixelVal_in_2_4;
      end else if (10'ha4 == _T_25[9:0]) begin
        image_2_164 <= io_pixelVal_in_2_3;
      end else if (10'ha4 == _T_22[9:0]) begin
        image_2_164 <= io_pixelVal_in_2_2;
      end else if (10'ha4 == _T_19[9:0]) begin
        image_2_164 <= io_pixelVal_in_2_1;
      end else if (10'ha4 == _T_15[9:0]) begin
        image_2_164 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_165 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha5 == _T_37[9:0]) begin
        image_2_165 <= io_pixelVal_in_2_7;
      end else if (10'ha5 == _T_34[9:0]) begin
        image_2_165 <= io_pixelVal_in_2_6;
      end else if (10'ha5 == _T_31[9:0]) begin
        image_2_165 <= io_pixelVal_in_2_5;
      end else if (10'ha5 == _T_28[9:0]) begin
        image_2_165 <= io_pixelVal_in_2_4;
      end else if (10'ha5 == _T_25[9:0]) begin
        image_2_165 <= io_pixelVal_in_2_3;
      end else if (10'ha5 == _T_22[9:0]) begin
        image_2_165 <= io_pixelVal_in_2_2;
      end else if (10'ha5 == _T_19[9:0]) begin
        image_2_165 <= io_pixelVal_in_2_1;
      end else if (10'ha5 == _T_15[9:0]) begin
        image_2_165 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_166 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha6 == _T_37[9:0]) begin
        image_2_166 <= io_pixelVal_in_2_7;
      end else if (10'ha6 == _T_34[9:0]) begin
        image_2_166 <= io_pixelVal_in_2_6;
      end else if (10'ha6 == _T_31[9:0]) begin
        image_2_166 <= io_pixelVal_in_2_5;
      end else if (10'ha6 == _T_28[9:0]) begin
        image_2_166 <= io_pixelVal_in_2_4;
      end else if (10'ha6 == _T_25[9:0]) begin
        image_2_166 <= io_pixelVal_in_2_3;
      end else if (10'ha6 == _T_22[9:0]) begin
        image_2_166 <= io_pixelVal_in_2_2;
      end else if (10'ha6 == _T_19[9:0]) begin
        image_2_166 <= io_pixelVal_in_2_1;
      end else if (10'ha6 == _T_15[9:0]) begin
        image_2_166 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_167 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha7 == _T_37[9:0]) begin
        image_2_167 <= io_pixelVal_in_2_7;
      end else if (10'ha7 == _T_34[9:0]) begin
        image_2_167 <= io_pixelVal_in_2_6;
      end else if (10'ha7 == _T_31[9:0]) begin
        image_2_167 <= io_pixelVal_in_2_5;
      end else if (10'ha7 == _T_28[9:0]) begin
        image_2_167 <= io_pixelVal_in_2_4;
      end else if (10'ha7 == _T_25[9:0]) begin
        image_2_167 <= io_pixelVal_in_2_3;
      end else if (10'ha7 == _T_22[9:0]) begin
        image_2_167 <= io_pixelVal_in_2_2;
      end else if (10'ha7 == _T_19[9:0]) begin
        image_2_167 <= io_pixelVal_in_2_1;
      end else if (10'ha7 == _T_15[9:0]) begin
        image_2_167 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_168 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha8 == _T_37[9:0]) begin
        image_2_168 <= io_pixelVal_in_2_7;
      end else if (10'ha8 == _T_34[9:0]) begin
        image_2_168 <= io_pixelVal_in_2_6;
      end else if (10'ha8 == _T_31[9:0]) begin
        image_2_168 <= io_pixelVal_in_2_5;
      end else if (10'ha8 == _T_28[9:0]) begin
        image_2_168 <= io_pixelVal_in_2_4;
      end else if (10'ha8 == _T_25[9:0]) begin
        image_2_168 <= io_pixelVal_in_2_3;
      end else if (10'ha8 == _T_22[9:0]) begin
        image_2_168 <= io_pixelVal_in_2_2;
      end else if (10'ha8 == _T_19[9:0]) begin
        image_2_168 <= io_pixelVal_in_2_1;
      end else if (10'ha8 == _T_15[9:0]) begin
        image_2_168 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_169 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha9 == _T_37[9:0]) begin
        image_2_169 <= io_pixelVal_in_2_7;
      end else if (10'ha9 == _T_34[9:0]) begin
        image_2_169 <= io_pixelVal_in_2_6;
      end else if (10'ha9 == _T_31[9:0]) begin
        image_2_169 <= io_pixelVal_in_2_5;
      end else if (10'ha9 == _T_28[9:0]) begin
        image_2_169 <= io_pixelVal_in_2_4;
      end else if (10'ha9 == _T_25[9:0]) begin
        image_2_169 <= io_pixelVal_in_2_3;
      end else if (10'ha9 == _T_22[9:0]) begin
        image_2_169 <= io_pixelVal_in_2_2;
      end else if (10'ha9 == _T_19[9:0]) begin
        image_2_169 <= io_pixelVal_in_2_1;
      end else if (10'ha9 == _T_15[9:0]) begin
        image_2_169 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_170 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'haa == _T_37[9:0]) begin
        image_2_170 <= io_pixelVal_in_2_7;
      end else if (10'haa == _T_34[9:0]) begin
        image_2_170 <= io_pixelVal_in_2_6;
      end else if (10'haa == _T_31[9:0]) begin
        image_2_170 <= io_pixelVal_in_2_5;
      end else if (10'haa == _T_28[9:0]) begin
        image_2_170 <= io_pixelVal_in_2_4;
      end else if (10'haa == _T_25[9:0]) begin
        image_2_170 <= io_pixelVal_in_2_3;
      end else if (10'haa == _T_22[9:0]) begin
        image_2_170 <= io_pixelVal_in_2_2;
      end else if (10'haa == _T_19[9:0]) begin
        image_2_170 <= io_pixelVal_in_2_1;
      end else if (10'haa == _T_15[9:0]) begin
        image_2_170 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_171 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hab == _T_37[9:0]) begin
        image_2_171 <= io_pixelVal_in_2_7;
      end else if (10'hab == _T_34[9:0]) begin
        image_2_171 <= io_pixelVal_in_2_6;
      end else if (10'hab == _T_31[9:0]) begin
        image_2_171 <= io_pixelVal_in_2_5;
      end else if (10'hab == _T_28[9:0]) begin
        image_2_171 <= io_pixelVal_in_2_4;
      end else if (10'hab == _T_25[9:0]) begin
        image_2_171 <= io_pixelVal_in_2_3;
      end else if (10'hab == _T_22[9:0]) begin
        image_2_171 <= io_pixelVal_in_2_2;
      end else if (10'hab == _T_19[9:0]) begin
        image_2_171 <= io_pixelVal_in_2_1;
      end else if (10'hab == _T_15[9:0]) begin
        image_2_171 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_172 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hac == _T_37[9:0]) begin
        image_2_172 <= io_pixelVal_in_2_7;
      end else if (10'hac == _T_34[9:0]) begin
        image_2_172 <= io_pixelVal_in_2_6;
      end else if (10'hac == _T_31[9:0]) begin
        image_2_172 <= io_pixelVal_in_2_5;
      end else if (10'hac == _T_28[9:0]) begin
        image_2_172 <= io_pixelVal_in_2_4;
      end else if (10'hac == _T_25[9:0]) begin
        image_2_172 <= io_pixelVal_in_2_3;
      end else if (10'hac == _T_22[9:0]) begin
        image_2_172 <= io_pixelVal_in_2_2;
      end else if (10'hac == _T_19[9:0]) begin
        image_2_172 <= io_pixelVal_in_2_1;
      end else if (10'hac == _T_15[9:0]) begin
        image_2_172 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_173 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'had == _T_37[9:0]) begin
        image_2_173 <= io_pixelVal_in_2_7;
      end else if (10'had == _T_34[9:0]) begin
        image_2_173 <= io_pixelVal_in_2_6;
      end else if (10'had == _T_31[9:0]) begin
        image_2_173 <= io_pixelVal_in_2_5;
      end else if (10'had == _T_28[9:0]) begin
        image_2_173 <= io_pixelVal_in_2_4;
      end else if (10'had == _T_25[9:0]) begin
        image_2_173 <= io_pixelVal_in_2_3;
      end else if (10'had == _T_22[9:0]) begin
        image_2_173 <= io_pixelVal_in_2_2;
      end else if (10'had == _T_19[9:0]) begin
        image_2_173 <= io_pixelVal_in_2_1;
      end else if (10'had == _T_15[9:0]) begin
        image_2_173 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_174 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hae == _T_37[9:0]) begin
        image_2_174 <= io_pixelVal_in_2_7;
      end else if (10'hae == _T_34[9:0]) begin
        image_2_174 <= io_pixelVal_in_2_6;
      end else if (10'hae == _T_31[9:0]) begin
        image_2_174 <= io_pixelVal_in_2_5;
      end else if (10'hae == _T_28[9:0]) begin
        image_2_174 <= io_pixelVal_in_2_4;
      end else if (10'hae == _T_25[9:0]) begin
        image_2_174 <= io_pixelVal_in_2_3;
      end else if (10'hae == _T_22[9:0]) begin
        image_2_174 <= io_pixelVal_in_2_2;
      end else if (10'hae == _T_19[9:0]) begin
        image_2_174 <= io_pixelVal_in_2_1;
      end else if (10'hae == _T_15[9:0]) begin
        image_2_174 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_175 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'haf == _T_37[9:0]) begin
        image_2_175 <= io_pixelVal_in_2_7;
      end else if (10'haf == _T_34[9:0]) begin
        image_2_175 <= io_pixelVal_in_2_6;
      end else if (10'haf == _T_31[9:0]) begin
        image_2_175 <= io_pixelVal_in_2_5;
      end else if (10'haf == _T_28[9:0]) begin
        image_2_175 <= io_pixelVal_in_2_4;
      end else if (10'haf == _T_25[9:0]) begin
        image_2_175 <= io_pixelVal_in_2_3;
      end else if (10'haf == _T_22[9:0]) begin
        image_2_175 <= io_pixelVal_in_2_2;
      end else if (10'haf == _T_19[9:0]) begin
        image_2_175 <= io_pixelVal_in_2_1;
      end else if (10'haf == _T_15[9:0]) begin
        image_2_175 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_176 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb0 == _T_37[9:0]) begin
        image_2_176 <= io_pixelVal_in_2_7;
      end else if (10'hb0 == _T_34[9:0]) begin
        image_2_176 <= io_pixelVal_in_2_6;
      end else if (10'hb0 == _T_31[9:0]) begin
        image_2_176 <= io_pixelVal_in_2_5;
      end else if (10'hb0 == _T_28[9:0]) begin
        image_2_176 <= io_pixelVal_in_2_4;
      end else if (10'hb0 == _T_25[9:0]) begin
        image_2_176 <= io_pixelVal_in_2_3;
      end else if (10'hb0 == _T_22[9:0]) begin
        image_2_176 <= io_pixelVal_in_2_2;
      end else if (10'hb0 == _T_19[9:0]) begin
        image_2_176 <= io_pixelVal_in_2_1;
      end else if (10'hb0 == _T_15[9:0]) begin
        image_2_176 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_177 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb1 == _T_37[9:0]) begin
        image_2_177 <= io_pixelVal_in_2_7;
      end else if (10'hb1 == _T_34[9:0]) begin
        image_2_177 <= io_pixelVal_in_2_6;
      end else if (10'hb1 == _T_31[9:0]) begin
        image_2_177 <= io_pixelVal_in_2_5;
      end else if (10'hb1 == _T_28[9:0]) begin
        image_2_177 <= io_pixelVal_in_2_4;
      end else if (10'hb1 == _T_25[9:0]) begin
        image_2_177 <= io_pixelVal_in_2_3;
      end else if (10'hb1 == _T_22[9:0]) begin
        image_2_177 <= io_pixelVal_in_2_2;
      end else if (10'hb1 == _T_19[9:0]) begin
        image_2_177 <= io_pixelVal_in_2_1;
      end else if (10'hb1 == _T_15[9:0]) begin
        image_2_177 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_178 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb2 == _T_37[9:0]) begin
        image_2_178 <= io_pixelVal_in_2_7;
      end else if (10'hb2 == _T_34[9:0]) begin
        image_2_178 <= io_pixelVal_in_2_6;
      end else if (10'hb2 == _T_31[9:0]) begin
        image_2_178 <= io_pixelVal_in_2_5;
      end else if (10'hb2 == _T_28[9:0]) begin
        image_2_178 <= io_pixelVal_in_2_4;
      end else if (10'hb2 == _T_25[9:0]) begin
        image_2_178 <= io_pixelVal_in_2_3;
      end else if (10'hb2 == _T_22[9:0]) begin
        image_2_178 <= io_pixelVal_in_2_2;
      end else if (10'hb2 == _T_19[9:0]) begin
        image_2_178 <= io_pixelVal_in_2_1;
      end else if (10'hb2 == _T_15[9:0]) begin
        image_2_178 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_179 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb3 == _T_37[9:0]) begin
        image_2_179 <= io_pixelVal_in_2_7;
      end else if (10'hb3 == _T_34[9:0]) begin
        image_2_179 <= io_pixelVal_in_2_6;
      end else if (10'hb3 == _T_31[9:0]) begin
        image_2_179 <= io_pixelVal_in_2_5;
      end else if (10'hb3 == _T_28[9:0]) begin
        image_2_179 <= io_pixelVal_in_2_4;
      end else if (10'hb3 == _T_25[9:0]) begin
        image_2_179 <= io_pixelVal_in_2_3;
      end else if (10'hb3 == _T_22[9:0]) begin
        image_2_179 <= io_pixelVal_in_2_2;
      end else if (10'hb3 == _T_19[9:0]) begin
        image_2_179 <= io_pixelVal_in_2_1;
      end else if (10'hb3 == _T_15[9:0]) begin
        image_2_179 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_180 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb4 == _T_37[9:0]) begin
        image_2_180 <= io_pixelVal_in_2_7;
      end else if (10'hb4 == _T_34[9:0]) begin
        image_2_180 <= io_pixelVal_in_2_6;
      end else if (10'hb4 == _T_31[9:0]) begin
        image_2_180 <= io_pixelVal_in_2_5;
      end else if (10'hb4 == _T_28[9:0]) begin
        image_2_180 <= io_pixelVal_in_2_4;
      end else if (10'hb4 == _T_25[9:0]) begin
        image_2_180 <= io_pixelVal_in_2_3;
      end else if (10'hb4 == _T_22[9:0]) begin
        image_2_180 <= io_pixelVal_in_2_2;
      end else if (10'hb4 == _T_19[9:0]) begin
        image_2_180 <= io_pixelVal_in_2_1;
      end else if (10'hb4 == _T_15[9:0]) begin
        image_2_180 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_181 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb5 == _T_37[9:0]) begin
        image_2_181 <= io_pixelVal_in_2_7;
      end else if (10'hb5 == _T_34[9:0]) begin
        image_2_181 <= io_pixelVal_in_2_6;
      end else if (10'hb5 == _T_31[9:0]) begin
        image_2_181 <= io_pixelVal_in_2_5;
      end else if (10'hb5 == _T_28[9:0]) begin
        image_2_181 <= io_pixelVal_in_2_4;
      end else if (10'hb5 == _T_25[9:0]) begin
        image_2_181 <= io_pixelVal_in_2_3;
      end else if (10'hb5 == _T_22[9:0]) begin
        image_2_181 <= io_pixelVal_in_2_2;
      end else if (10'hb5 == _T_19[9:0]) begin
        image_2_181 <= io_pixelVal_in_2_1;
      end else if (10'hb5 == _T_15[9:0]) begin
        image_2_181 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_182 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb6 == _T_37[9:0]) begin
        image_2_182 <= io_pixelVal_in_2_7;
      end else if (10'hb6 == _T_34[9:0]) begin
        image_2_182 <= io_pixelVal_in_2_6;
      end else if (10'hb6 == _T_31[9:0]) begin
        image_2_182 <= io_pixelVal_in_2_5;
      end else if (10'hb6 == _T_28[9:0]) begin
        image_2_182 <= io_pixelVal_in_2_4;
      end else if (10'hb6 == _T_25[9:0]) begin
        image_2_182 <= io_pixelVal_in_2_3;
      end else if (10'hb6 == _T_22[9:0]) begin
        image_2_182 <= io_pixelVal_in_2_2;
      end else if (10'hb6 == _T_19[9:0]) begin
        image_2_182 <= io_pixelVal_in_2_1;
      end else if (10'hb6 == _T_15[9:0]) begin
        image_2_182 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_183 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb7 == _T_37[9:0]) begin
        image_2_183 <= io_pixelVal_in_2_7;
      end else if (10'hb7 == _T_34[9:0]) begin
        image_2_183 <= io_pixelVal_in_2_6;
      end else if (10'hb7 == _T_31[9:0]) begin
        image_2_183 <= io_pixelVal_in_2_5;
      end else if (10'hb7 == _T_28[9:0]) begin
        image_2_183 <= io_pixelVal_in_2_4;
      end else if (10'hb7 == _T_25[9:0]) begin
        image_2_183 <= io_pixelVal_in_2_3;
      end else if (10'hb7 == _T_22[9:0]) begin
        image_2_183 <= io_pixelVal_in_2_2;
      end else if (10'hb7 == _T_19[9:0]) begin
        image_2_183 <= io_pixelVal_in_2_1;
      end else if (10'hb7 == _T_15[9:0]) begin
        image_2_183 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_184 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb8 == _T_37[9:0]) begin
        image_2_184 <= io_pixelVal_in_2_7;
      end else if (10'hb8 == _T_34[9:0]) begin
        image_2_184 <= io_pixelVal_in_2_6;
      end else if (10'hb8 == _T_31[9:0]) begin
        image_2_184 <= io_pixelVal_in_2_5;
      end else if (10'hb8 == _T_28[9:0]) begin
        image_2_184 <= io_pixelVal_in_2_4;
      end else if (10'hb8 == _T_25[9:0]) begin
        image_2_184 <= io_pixelVal_in_2_3;
      end else if (10'hb8 == _T_22[9:0]) begin
        image_2_184 <= io_pixelVal_in_2_2;
      end else if (10'hb8 == _T_19[9:0]) begin
        image_2_184 <= io_pixelVal_in_2_1;
      end else if (10'hb8 == _T_15[9:0]) begin
        image_2_184 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_185 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb9 == _T_37[9:0]) begin
        image_2_185 <= io_pixelVal_in_2_7;
      end else if (10'hb9 == _T_34[9:0]) begin
        image_2_185 <= io_pixelVal_in_2_6;
      end else if (10'hb9 == _T_31[9:0]) begin
        image_2_185 <= io_pixelVal_in_2_5;
      end else if (10'hb9 == _T_28[9:0]) begin
        image_2_185 <= io_pixelVal_in_2_4;
      end else if (10'hb9 == _T_25[9:0]) begin
        image_2_185 <= io_pixelVal_in_2_3;
      end else if (10'hb9 == _T_22[9:0]) begin
        image_2_185 <= io_pixelVal_in_2_2;
      end else if (10'hb9 == _T_19[9:0]) begin
        image_2_185 <= io_pixelVal_in_2_1;
      end else if (10'hb9 == _T_15[9:0]) begin
        image_2_185 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_186 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hba == _T_37[9:0]) begin
        image_2_186 <= io_pixelVal_in_2_7;
      end else if (10'hba == _T_34[9:0]) begin
        image_2_186 <= io_pixelVal_in_2_6;
      end else if (10'hba == _T_31[9:0]) begin
        image_2_186 <= io_pixelVal_in_2_5;
      end else if (10'hba == _T_28[9:0]) begin
        image_2_186 <= io_pixelVal_in_2_4;
      end else if (10'hba == _T_25[9:0]) begin
        image_2_186 <= io_pixelVal_in_2_3;
      end else if (10'hba == _T_22[9:0]) begin
        image_2_186 <= io_pixelVal_in_2_2;
      end else if (10'hba == _T_19[9:0]) begin
        image_2_186 <= io_pixelVal_in_2_1;
      end else if (10'hba == _T_15[9:0]) begin
        image_2_186 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_187 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hbb == _T_37[9:0]) begin
        image_2_187 <= io_pixelVal_in_2_7;
      end else if (10'hbb == _T_34[9:0]) begin
        image_2_187 <= io_pixelVal_in_2_6;
      end else if (10'hbb == _T_31[9:0]) begin
        image_2_187 <= io_pixelVal_in_2_5;
      end else if (10'hbb == _T_28[9:0]) begin
        image_2_187 <= io_pixelVal_in_2_4;
      end else if (10'hbb == _T_25[9:0]) begin
        image_2_187 <= io_pixelVal_in_2_3;
      end else if (10'hbb == _T_22[9:0]) begin
        image_2_187 <= io_pixelVal_in_2_2;
      end else if (10'hbb == _T_19[9:0]) begin
        image_2_187 <= io_pixelVal_in_2_1;
      end else if (10'hbb == _T_15[9:0]) begin
        image_2_187 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_188 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hbc == _T_37[9:0]) begin
        image_2_188 <= io_pixelVal_in_2_7;
      end else if (10'hbc == _T_34[9:0]) begin
        image_2_188 <= io_pixelVal_in_2_6;
      end else if (10'hbc == _T_31[9:0]) begin
        image_2_188 <= io_pixelVal_in_2_5;
      end else if (10'hbc == _T_28[9:0]) begin
        image_2_188 <= io_pixelVal_in_2_4;
      end else if (10'hbc == _T_25[9:0]) begin
        image_2_188 <= io_pixelVal_in_2_3;
      end else if (10'hbc == _T_22[9:0]) begin
        image_2_188 <= io_pixelVal_in_2_2;
      end else if (10'hbc == _T_19[9:0]) begin
        image_2_188 <= io_pixelVal_in_2_1;
      end else if (10'hbc == _T_15[9:0]) begin
        image_2_188 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_189 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hbd == _T_37[9:0]) begin
        image_2_189 <= io_pixelVal_in_2_7;
      end else if (10'hbd == _T_34[9:0]) begin
        image_2_189 <= io_pixelVal_in_2_6;
      end else if (10'hbd == _T_31[9:0]) begin
        image_2_189 <= io_pixelVal_in_2_5;
      end else if (10'hbd == _T_28[9:0]) begin
        image_2_189 <= io_pixelVal_in_2_4;
      end else if (10'hbd == _T_25[9:0]) begin
        image_2_189 <= io_pixelVal_in_2_3;
      end else if (10'hbd == _T_22[9:0]) begin
        image_2_189 <= io_pixelVal_in_2_2;
      end else if (10'hbd == _T_19[9:0]) begin
        image_2_189 <= io_pixelVal_in_2_1;
      end else if (10'hbd == _T_15[9:0]) begin
        image_2_189 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_190 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hbe == _T_37[9:0]) begin
        image_2_190 <= io_pixelVal_in_2_7;
      end else if (10'hbe == _T_34[9:0]) begin
        image_2_190 <= io_pixelVal_in_2_6;
      end else if (10'hbe == _T_31[9:0]) begin
        image_2_190 <= io_pixelVal_in_2_5;
      end else if (10'hbe == _T_28[9:0]) begin
        image_2_190 <= io_pixelVal_in_2_4;
      end else if (10'hbe == _T_25[9:0]) begin
        image_2_190 <= io_pixelVal_in_2_3;
      end else if (10'hbe == _T_22[9:0]) begin
        image_2_190 <= io_pixelVal_in_2_2;
      end else if (10'hbe == _T_19[9:0]) begin
        image_2_190 <= io_pixelVal_in_2_1;
      end else if (10'hbe == _T_15[9:0]) begin
        image_2_190 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_191 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hbf == _T_37[9:0]) begin
        image_2_191 <= io_pixelVal_in_2_7;
      end else if (10'hbf == _T_34[9:0]) begin
        image_2_191 <= io_pixelVal_in_2_6;
      end else if (10'hbf == _T_31[9:0]) begin
        image_2_191 <= io_pixelVal_in_2_5;
      end else if (10'hbf == _T_28[9:0]) begin
        image_2_191 <= io_pixelVal_in_2_4;
      end else if (10'hbf == _T_25[9:0]) begin
        image_2_191 <= io_pixelVal_in_2_3;
      end else if (10'hbf == _T_22[9:0]) begin
        image_2_191 <= io_pixelVal_in_2_2;
      end else if (10'hbf == _T_19[9:0]) begin
        image_2_191 <= io_pixelVal_in_2_1;
      end else if (10'hbf == _T_15[9:0]) begin
        image_2_191 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_192 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc0 == _T_37[9:0]) begin
        image_2_192 <= io_pixelVal_in_2_7;
      end else if (10'hc0 == _T_34[9:0]) begin
        image_2_192 <= io_pixelVal_in_2_6;
      end else if (10'hc0 == _T_31[9:0]) begin
        image_2_192 <= io_pixelVal_in_2_5;
      end else if (10'hc0 == _T_28[9:0]) begin
        image_2_192 <= io_pixelVal_in_2_4;
      end else if (10'hc0 == _T_25[9:0]) begin
        image_2_192 <= io_pixelVal_in_2_3;
      end else if (10'hc0 == _T_22[9:0]) begin
        image_2_192 <= io_pixelVal_in_2_2;
      end else if (10'hc0 == _T_19[9:0]) begin
        image_2_192 <= io_pixelVal_in_2_1;
      end else if (10'hc0 == _T_15[9:0]) begin
        image_2_192 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_193 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc1 == _T_37[9:0]) begin
        image_2_193 <= io_pixelVal_in_2_7;
      end else if (10'hc1 == _T_34[9:0]) begin
        image_2_193 <= io_pixelVal_in_2_6;
      end else if (10'hc1 == _T_31[9:0]) begin
        image_2_193 <= io_pixelVal_in_2_5;
      end else if (10'hc1 == _T_28[9:0]) begin
        image_2_193 <= io_pixelVal_in_2_4;
      end else if (10'hc1 == _T_25[9:0]) begin
        image_2_193 <= io_pixelVal_in_2_3;
      end else if (10'hc1 == _T_22[9:0]) begin
        image_2_193 <= io_pixelVal_in_2_2;
      end else if (10'hc1 == _T_19[9:0]) begin
        image_2_193 <= io_pixelVal_in_2_1;
      end else if (10'hc1 == _T_15[9:0]) begin
        image_2_193 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_194 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc2 == _T_37[9:0]) begin
        image_2_194 <= io_pixelVal_in_2_7;
      end else if (10'hc2 == _T_34[9:0]) begin
        image_2_194 <= io_pixelVal_in_2_6;
      end else if (10'hc2 == _T_31[9:0]) begin
        image_2_194 <= io_pixelVal_in_2_5;
      end else if (10'hc2 == _T_28[9:0]) begin
        image_2_194 <= io_pixelVal_in_2_4;
      end else if (10'hc2 == _T_25[9:0]) begin
        image_2_194 <= io_pixelVal_in_2_3;
      end else if (10'hc2 == _T_22[9:0]) begin
        image_2_194 <= io_pixelVal_in_2_2;
      end else if (10'hc2 == _T_19[9:0]) begin
        image_2_194 <= io_pixelVal_in_2_1;
      end else if (10'hc2 == _T_15[9:0]) begin
        image_2_194 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_195 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc3 == _T_37[9:0]) begin
        image_2_195 <= io_pixelVal_in_2_7;
      end else if (10'hc3 == _T_34[9:0]) begin
        image_2_195 <= io_pixelVal_in_2_6;
      end else if (10'hc3 == _T_31[9:0]) begin
        image_2_195 <= io_pixelVal_in_2_5;
      end else if (10'hc3 == _T_28[9:0]) begin
        image_2_195 <= io_pixelVal_in_2_4;
      end else if (10'hc3 == _T_25[9:0]) begin
        image_2_195 <= io_pixelVal_in_2_3;
      end else if (10'hc3 == _T_22[9:0]) begin
        image_2_195 <= io_pixelVal_in_2_2;
      end else if (10'hc3 == _T_19[9:0]) begin
        image_2_195 <= io_pixelVal_in_2_1;
      end else if (10'hc3 == _T_15[9:0]) begin
        image_2_195 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_196 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc4 == _T_37[9:0]) begin
        image_2_196 <= io_pixelVal_in_2_7;
      end else if (10'hc4 == _T_34[9:0]) begin
        image_2_196 <= io_pixelVal_in_2_6;
      end else if (10'hc4 == _T_31[9:0]) begin
        image_2_196 <= io_pixelVal_in_2_5;
      end else if (10'hc4 == _T_28[9:0]) begin
        image_2_196 <= io_pixelVal_in_2_4;
      end else if (10'hc4 == _T_25[9:0]) begin
        image_2_196 <= io_pixelVal_in_2_3;
      end else if (10'hc4 == _T_22[9:0]) begin
        image_2_196 <= io_pixelVal_in_2_2;
      end else if (10'hc4 == _T_19[9:0]) begin
        image_2_196 <= io_pixelVal_in_2_1;
      end else if (10'hc4 == _T_15[9:0]) begin
        image_2_196 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_197 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc5 == _T_37[9:0]) begin
        image_2_197 <= io_pixelVal_in_2_7;
      end else if (10'hc5 == _T_34[9:0]) begin
        image_2_197 <= io_pixelVal_in_2_6;
      end else if (10'hc5 == _T_31[9:0]) begin
        image_2_197 <= io_pixelVal_in_2_5;
      end else if (10'hc5 == _T_28[9:0]) begin
        image_2_197 <= io_pixelVal_in_2_4;
      end else if (10'hc5 == _T_25[9:0]) begin
        image_2_197 <= io_pixelVal_in_2_3;
      end else if (10'hc5 == _T_22[9:0]) begin
        image_2_197 <= io_pixelVal_in_2_2;
      end else if (10'hc5 == _T_19[9:0]) begin
        image_2_197 <= io_pixelVal_in_2_1;
      end else if (10'hc5 == _T_15[9:0]) begin
        image_2_197 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_198 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc6 == _T_37[9:0]) begin
        image_2_198 <= io_pixelVal_in_2_7;
      end else if (10'hc6 == _T_34[9:0]) begin
        image_2_198 <= io_pixelVal_in_2_6;
      end else if (10'hc6 == _T_31[9:0]) begin
        image_2_198 <= io_pixelVal_in_2_5;
      end else if (10'hc6 == _T_28[9:0]) begin
        image_2_198 <= io_pixelVal_in_2_4;
      end else if (10'hc6 == _T_25[9:0]) begin
        image_2_198 <= io_pixelVal_in_2_3;
      end else if (10'hc6 == _T_22[9:0]) begin
        image_2_198 <= io_pixelVal_in_2_2;
      end else if (10'hc6 == _T_19[9:0]) begin
        image_2_198 <= io_pixelVal_in_2_1;
      end else if (10'hc6 == _T_15[9:0]) begin
        image_2_198 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_199 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc7 == _T_37[9:0]) begin
        image_2_199 <= io_pixelVal_in_2_7;
      end else if (10'hc7 == _T_34[9:0]) begin
        image_2_199 <= io_pixelVal_in_2_6;
      end else if (10'hc7 == _T_31[9:0]) begin
        image_2_199 <= io_pixelVal_in_2_5;
      end else if (10'hc7 == _T_28[9:0]) begin
        image_2_199 <= io_pixelVal_in_2_4;
      end else if (10'hc7 == _T_25[9:0]) begin
        image_2_199 <= io_pixelVal_in_2_3;
      end else if (10'hc7 == _T_22[9:0]) begin
        image_2_199 <= io_pixelVal_in_2_2;
      end else if (10'hc7 == _T_19[9:0]) begin
        image_2_199 <= io_pixelVal_in_2_1;
      end else if (10'hc7 == _T_15[9:0]) begin
        image_2_199 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_200 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc8 == _T_37[9:0]) begin
        image_2_200 <= io_pixelVal_in_2_7;
      end else if (10'hc8 == _T_34[9:0]) begin
        image_2_200 <= io_pixelVal_in_2_6;
      end else if (10'hc8 == _T_31[9:0]) begin
        image_2_200 <= io_pixelVal_in_2_5;
      end else if (10'hc8 == _T_28[9:0]) begin
        image_2_200 <= io_pixelVal_in_2_4;
      end else if (10'hc8 == _T_25[9:0]) begin
        image_2_200 <= io_pixelVal_in_2_3;
      end else if (10'hc8 == _T_22[9:0]) begin
        image_2_200 <= io_pixelVal_in_2_2;
      end else if (10'hc8 == _T_19[9:0]) begin
        image_2_200 <= io_pixelVal_in_2_1;
      end else if (10'hc8 == _T_15[9:0]) begin
        image_2_200 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_201 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc9 == _T_37[9:0]) begin
        image_2_201 <= io_pixelVal_in_2_7;
      end else if (10'hc9 == _T_34[9:0]) begin
        image_2_201 <= io_pixelVal_in_2_6;
      end else if (10'hc9 == _T_31[9:0]) begin
        image_2_201 <= io_pixelVal_in_2_5;
      end else if (10'hc9 == _T_28[9:0]) begin
        image_2_201 <= io_pixelVal_in_2_4;
      end else if (10'hc9 == _T_25[9:0]) begin
        image_2_201 <= io_pixelVal_in_2_3;
      end else if (10'hc9 == _T_22[9:0]) begin
        image_2_201 <= io_pixelVal_in_2_2;
      end else if (10'hc9 == _T_19[9:0]) begin
        image_2_201 <= io_pixelVal_in_2_1;
      end else if (10'hc9 == _T_15[9:0]) begin
        image_2_201 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_202 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hca == _T_37[9:0]) begin
        image_2_202 <= io_pixelVal_in_2_7;
      end else if (10'hca == _T_34[9:0]) begin
        image_2_202 <= io_pixelVal_in_2_6;
      end else if (10'hca == _T_31[9:0]) begin
        image_2_202 <= io_pixelVal_in_2_5;
      end else if (10'hca == _T_28[9:0]) begin
        image_2_202 <= io_pixelVal_in_2_4;
      end else if (10'hca == _T_25[9:0]) begin
        image_2_202 <= io_pixelVal_in_2_3;
      end else if (10'hca == _T_22[9:0]) begin
        image_2_202 <= io_pixelVal_in_2_2;
      end else if (10'hca == _T_19[9:0]) begin
        image_2_202 <= io_pixelVal_in_2_1;
      end else if (10'hca == _T_15[9:0]) begin
        image_2_202 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_203 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hcb == _T_37[9:0]) begin
        image_2_203 <= io_pixelVal_in_2_7;
      end else if (10'hcb == _T_34[9:0]) begin
        image_2_203 <= io_pixelVal_in_2_6;
      end else if (10'hcb == _T_31[9:0]) begin
        image_2_203 <= io_pixelVal_in_2_5;
      end else if (10'hcb == _T_28[9:0]) begin
        image_2_203 <= io_pixelVal_in_2_4;
      end else if (10'hcb == _T_25[9:0]) begin
        image_2_203 <= io_pixelVal_in_2_3;
      end else if (10'hcb == _T_22[9:0]) begin
        image_2_203 <= io_pixelVal_in_2_2;
      end else if (10'hcb == _T_19[9:0]) begin
        image_2_203 <= io_pixelVal_in_2_1;
      end else if (10'hcb == _T_15[9:0]) begin
        image_2_203 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_204 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hcc == _T_37[9:0]) begin
        image_2_204 <= io_pixelVal_in_2_7;
      end else if (10'hcc == _T_34[9:0]) begin
        image_2_204 <= io_pixelVal_in_2_6;
      end else if (10'hcc == _T_31[9:0]) begin
        image_2_204 <= io_pixelVal_in_2_5;
      end else if (10'hcc == _T_28[9:0]) begin
        image_2_204 <= io_pixelVal_in_2_4;
      end else if (10'hcc == _T_25[9:0]) begin
        image_2_204 <= io_pixelVal_in_2_3;
      end else if (10'hcc == _T_22[9:0]) begin
        image_2_204 <= io_pixelVal_in_2_2;
      end else if (10'hcc == _T_19[9:0]) begin
        image_2_204 <= io_pixelVal_in_2_1;
      end else if (10'hcc == _T_15[9:0]) begin
        image_2_204 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_205 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hcd == _T_37[9:0]) begin
        image_2_205 <= io_pixelVal_in_2_7;
      end else if (10'hcd == _T_34[9:0]) begin
        image_2_205 <= io_pixelVal_in_2_6;
      end else if (10'hcd == _T_31[9:0]) begin
        image_2_205 <= io_pixelVal_in_2_5;
      end else if (10'hcd == _T_28[9:0]) begin
        image_2_205 <= io_pixelVal_in_2_4;
      end else if (10'hcd == _T_25[9:0]) begin
        image_2_205 <= io_pixelVal_in_2_3;
      end else if (10'hcd == _T_22[9:0]) begin
        image_2_205 <= io_pixelVal_in_2_2;
      end else if (10'hcd == _T_19[9:0]) begin
        image_2_205 <= io_pixelVal_in_2_1;
      end else if (10'hcd == _T_15[9:0]) begin
        image_2_205 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_206 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hce == _T_37[9:0]) begin
        image_2_206 <= io_pixelVal_in_2_7;
      end else if (10'hce == _T_34[9:0]) begin
        image_2_206 <= io_pixelVal_in_2_6;
      end else if (10'hce == _T_31[9:0]) begin
        image_2_206 <= io_pixelVal_in_2_5;
      end else if (10'hce == _T_28[9:0]) begin
        image_2_206 <= io_pixelVal_in_2_4;
      end else if (10'hce == _T_25[9:0]) begin
        image_2_206 <= io_pixelVal_in_2_3;
      end else if (10'hce == _T_22[9:0]) begin
        image_2_206 <= io_pixelVal_in_2_2;
      end else if (10'hce == _T_19[9:0]) begin
        image_2_206 <= io_pixelVal_in_2_1;
      end else if (10'hce == _T_15[9:0]) begin
        image_2_206 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_207 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hcf == _T_37[9:0]) begin
        image_2_207 <= io_pixelVal_in_2_7;
      end else if (10'hcf == _T_34[9:0]) begin
        image_2_207 <= io_pixelVal_in_2_6;
      end else if (10'hcf == _T_31[9:0]) begin
        image_2_207 <= io_pixelVal_in_2_5;
      end else if (10'hcf == _T_28[9:0]) begin
        image_2_207 <= io_pixelVal_in_2_4;
      end else if (10'hcf == _T_25[9:0]) begin
        image_2_207 <= io_pixelVal_in_2_3;
      end else if (10'hcf == _T_22[9:0]) begin
        image_2_207 <= io_pixelVal_in_2_2;
      end else if (10'hcf == _T_19[9:0]) begin
        image_2_207 <= io_pixelVal_in_2_1;
      end else if (10'hcf == _T_15[9:0]) begin
        image_2_207 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_208 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd0 == _T_37[9:0]) begin
        image_2_208 <= io_pixelVal_in_2_7;
      end else if (10'hd0 == _T_34[9:0]) begin
        image_2_208 <= io_pixelVal_in_2_6;
      end else if (10'hd0 == _T_31[9:0]) begin
        image_2_208 <= io_pixelVal_in_2_5;
      end else if (10'hd0 == _T_28[9:0]) begin
        image_2_208 <= io_pixelVal_in_2_4;
      end else if (10'hd0 == _T_25[9:0]) begin
        image_2_208 <= io_pixelVal_in_2_3;
      end else if (10'hd0 == _T_22[9:0]) begin
        image_2_208 <= io_pixelVal_in_2_2;
      end else if (10'hd0 == _T_19[9:0]) begin
        image_2_208 <= io_pixelVal_in_2_1;
      end else if (10'hd0 == _T_15[9:0]) begin
        image_2_208 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_209 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd1 == _T_37[9:0]) begin
        image_2_209 <= io_pixelVal_in_2_7;
      end else if (10'hd1 == _T_34[9:0]) begin
        image_2_209 <= io_pixelVal_in_2_6;
      end else if (10'hd1 == _T_31[9:0]) begin
        image_2_209 <= io_pixelVal_in_2_5;
      end else if (10'hd1 == _T_28[9:0]) begin
        image_2_209 <= io_pixelVal_in_2_4;
      end else if (10'hd1 == _T_25[9:0]) begin
        image_2_209 <= io_pixelVal_in_2_3;
      end else if (10'hd1 == _T_22[9:0]) begin
        image_2_209 <= io_pixelVal_in_2_2;
      end else if (10'hd1 == _T_19[9:0]) begin
        image_2_209 <= io_pixelVal_in_2_1;
      end else if (10'hd1 == _T_15[9:0]) begin
        image_2_209 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_210 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd2 == _T_37[9:0]) begin
        image_2_210 <= io_pixelVal_in_2_7;
      end else if (10'hd2 == _T_34[9:0]) begin
        image_2_210 <= io_pixelVal_in_2_6;
      end else if (10'hd2 == _T_31[9:0]) begin
        image_2_210 <= io_pixelVal_in_2_5;
      end else if (10'hd2 == _T_28[9:0]) begin
        image_2_210 <= io_pixelVal_in_2_4;
      end else if (10'hd2 == _T_25[9:0]) begin
        image_2_210 <= io_pixelVal_in_2_3;
      end else if (10'hd2 == _T_22[9:0]) begin
        image_2_210 <= io_pixelVal_in_2_2;
      end else if (10'hd2 == _T_19[9:0]) begin
        image_2_210 <= io_pixelVal_in_2_1;
      end else if (10'hd2 == _T_15[9:0]) begin
        image_2_210 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_211 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd3 == _T_37[9:0]) begin
        image_2_211 <= io_pixelVal_in_2_7;
      end else if (10'hd3 == _T_34[9:0]) begin
        image_2_211 <= io_pixelVal_in_2_6;
      end else if (10'hd3 == _T_31[9:0]) begin
        image_2_211 <= io_pixelVal_in_2_5;
      end else if (10'hd3 == _T_28[9:0]) begin
        image_2_211 <= io_pixelVal_in_2_4;
      end else if (10'hd3 == _T_25[9:0]) begin
        image_2_211 <= io_pixelVal_in_2_3;
      end else if (10'hd3 == _T_22[9:0]) begin
        image_2_211 <= io_pixelVal_in_2_2;
      end else if (10'hd3 == _T_19[9:0]) begin
        image_2_211 <= io_pixelVal_in_2_1;
      end else if (10'hd3 == _T_15[9:0]) begin
        image_2_211 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_212 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd4 == _T_37[9:0]) begin
        image_2_212 <= io_pixelVal_in_2_7;
      end else if (10'hd4 == _T_34[9:0]) begin
        image_2_212 <= io_pixelVal_in_2_6;
      end else if (10'hd4 == _T_31[9:0]) begin
        image_2_212 <= io_pixelVal_in_2_5;
      end else if (10'hd4 == _T_28[9:0]) begin
        image_2_212 <= io_pixelVal_in_2_4;
      end else if (10'hd4 == _T_25[9:0]) begin
        image_2_212 <= io_pixelVal_in_2_3;
      end else if (10'hd4 == _T_22[9:0]) begin
        image_2_212 <= io_pixelVal_in_2_2;
      end else if (10'hd4 == _T_19[9:0]) begin
        image_2_212 <= io_pixelVal_in_2_1;
      end else if (10'hd4 == _T_15[9:0]) begin
        image_2_212 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_213 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd5 == _T_37[9:0]) begin
        image_2_213 <= io_pixelVal_in_2_7;
      end else if (10'hd5 == _T_34[9:0]) begin
        image_2_213 <= io_pixelVal_in_2_6;
      end else if (10'hd5 == _T_31[9:0]) begin
        image_2_213 <= io_pixelVal_in_2_5;
      end else if (10'hd5 == _T_28[9:0]) begin
        image_2_213 <= io_pixelVal_in_2_4;
      end else if (10'hd5 == _T_25[9:0]) begin
        image_2_213 <= io_pixelVal_in_2_3;
      end else if (10'hd5 == _T_22[9:0]) begin
        image_2_213 <= io_pixelVal_in_2_2;
      end else if (10'hd5 == _T_19[9:0]) begin
        image_2_213 <= io_pixelVal_in_2_1;
      end else if (10'hd5 == _T_15[9:0]) begin
        image_2_213 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_214 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd6 == _T_37[9:0]) begin
        image_2_214 <= io_pixelVal_in_2_7;
      end else if (10'hd6 == _T_34[9:0]) begin
        image_2_214 <= io_pixelVal_in_2_6;
      end else if (10'hd6 == _T_31[9:0]) begin
        image_2_214 <= io_pixelVal_in_2_5;
      end else if (10'hd6 == _T_28[9:0]) begin
        image_2_214 <= io_pixelVal_in_2_4;
      end else if (10'hd6 == _T_25[9:0]) begin
        image_2_214 <= io_pixelVal_in_2_3;
      end else if (10'hd6 == _T_22[9:0]) begin
        image_2_214 <= io_pixelVal_in_2_2;
      end else if (10'hd6 == _T_19[9:0]) begin
        image_2_214 <= io_pixelVal_in_2_1;
      end else if (10'hd6 == _T_15[9:0]) begin
        image_2_214 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_215 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd7 == _T_37[9:0]) begin
        image_2_215 <= io_pixelVal_in_2_7;
      end else if (10'hd7 == _T_34[9:0]) begin
        image_2_215 <= io_pixelVal_in_2_6;
      end else if (10'hd7 == _T_31[9:0]) begin
        image_2_215 <= io_pixelVal_in_2_5;
      end else if (10'hd7 == _T_28[9:0]) begin
        image_2_215 <= io_pixelVal_in_2_4;
      end else if (10'hd7 == _T_25[9:0]) begin
        image_2_215 <= io_pixelVal_in_2_3;
      end else if (10'hd7 == _T_22[9:0]) begin
        image_2_215 <= io_pixelVal_in_2_2;
      end else if (10'hd7 == _T_19[9:0]) begin
        image_2_215 <= io_pixelVal_in_2_1;
      end else if (10'hd7 == _T_15[9:0]) begin
        image_2_215 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_216 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd8 == _T_37[9:0]) begin
        image_2_216 <= io_pixelVal_in_2_7;
      end else if (10'hd8 == _T_34[9:0]) begin
        image_2_216 <= io_pixelVal_in_2_6;
      end else if (10'hd8 == _T_31[9:0]) begin
        image_2_216 <= io_pixelVal_in_2_5;
      end else if (10'hd8 == _T_28[9:0]) begin
        image_2_216 <= io_pixelVal_in_2_4;
      end else if (10'hd8 == _T_25[9:0]) begin
        image_2_216 <= io_pixelVal_in_2_3;
      end else if (10'hd8 == _T_22[9:0]) begin
        image_2_216 <= io_pixelVal_in_2_2;
      end else if (10'hd8 == _T_19[9:0]) begin
        image_2_216 <= io_pixelVal_in_2_1;
      end else if (10'hd8 == _T_15[9:0]) begin
        image_2_216 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_217 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd9 == _T_37[9:0]) begin
        image_2_217 <= io_pixelVal_in_2_7;
      end else if (10'hd9 == _T_34[9:0]) begin
        image_2_217 <= io_pixelVal_in_2_6;
      end else if (10'hd9 == _T_31[9:0]) begin
        image_2_217 <= io_pixelVal_in_2_5;
      end else if (10'hd9 == _T_28[9:0]) begin
        image_2_217 <= io_pixelVal_in_2_4;
      end else if (10'hd9 == _T_25[9:0]) begin
        image_2_217 <= io_pixelVal_in_2_3;
      end else if (10'hd9 == _T_22[9:0]) begin
        image_2_217 <= io_pixelVal_in_2_2;
      end else if (10'hd9 == _T_19[9:0]) begin
        image_2_217 <= io_pixelVal_in_2_1;
      end else if (10'hd9 == _T_15[9:0]) begin
        image_2_217 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_218 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hda == _T_37[9:0]) begin
        image_2_218 <= io_pixelVal_in_2_7;
      end else if (10'hda == _T_34[9:0]) begin
        image_2_218 <= io_pixelVal_in_2_6;
      end else if (10'hda == _T_31[9:0]) begin
        image_2_218 <= io_pixelVal_in_2_5;
      end else if (10'hda == _T_28[9:0]) begin
        image_2_218 <= io_pixelVal_in_2_4;
      end else if (10'hda == _T_25[9:0]) begin
        image_2_218 <= io_pixelVal_in_2_3;
      end else if (10'hda == _T_22[9:0]) begin
        image_2_218 <= io_pixelVal_in_2_2;
      end else if (10'hda == _T_19[9:0]) begin
        image_2_218 <= io_pixelVal_in_2_1;
      end else if (10'hda == _T_15[9:0]) begin
        image_2_218 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_219 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hdb == _T_37[9:0]) begin
        image_2_219 <= io_pixelVal_in_2_7;
      end else if (10'hdb == _T_34[9:0]) begin
        image_2_219 <= io_pixelVal_in_2_6;
      end else if (10'hdb == _T_31[9:0]) begin
        image_2_219 <= io_pixelVal_in_2_5;
      end else if (10'hdb == _T_28[9:0]) begin
        image_2_219 <= io_pixelVal_in_2_4;
      end else if (10'hdb == _T_25[9:0]) begin
        image_2_219 <= io_pixelVal_in_2_3;
      end else if (10'hdb == _T_22[9:0]) begin
        image_2_219 <= io_pixelVal_in_2_2;
      end else if (10'hdb == _T_19[9:0]) begin
        image_2_219 <= io_pixelVal_in_2_1;
      end else if (10'hdb == _T_15[9:0]) begin
        image_2_219 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_220 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hdc == _T_37[9:0]) begin
        image_2_220 <= io_pixelVal_in_2_7;
      end else if (10'hdc == _T_34[9:0]) begin
        image_2_220 <= io_pixelVal_in_2_6;
      end else if (10'hdc == _T_31[9:0]) begin
        image_2_220 <= io_pixelVal_in_2_5;
      end else if (10'hdc == _T_28[9:0]) begin
        image_2_220 <= io_pixelVal_in_2_4;
      end else if (10'hdc == _T_25[9:0]) begin
        image_2_220 <= io_pixelVal_in_2_3;
      end else if (10'hdc == _T_22[9:0]) begin
        image_2_220 <= io_pixelVal_in_2_2;
      end else if (10'hdc == _T_19[9:0]) begin
        image_2_220 <= io_pixelVal_in_2_1;
      end else if (10'hdc == _T_15[9:0]) begin
        image_2_220 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_221 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hdd == _T_37[9:0]) begin
        image_2_221 <= io_pixelVal_in_2_7;
      end else if (10'hdd == _T_34[9:0]) begin
        image_2_221 <= io_pixelVal_in_2_6;
      end else if (10'hdd == _T_31[9:0]) begin
        image_2_221 <= io_pixelVal_in_2_5;
      end else if (10'hdd == _T_28[9:0]) begin
        image_2_221 <= io_pixelVal_in_2_4;
      end else if (10'hdd == _T_25[9:0]) begin
        image_2_221 <= io_pixelVal_in_2_3;
      end else if (10'hdd == _T_22[9:0]) begin
        image_2_221 <= io_pixelVal_in_2_2;
      end else if (10'hdd == _T_19[9:0]) begin
        image_2_221 <= io_pixelVal_in_2_1;
      end else if (10'hdd == _T_15[9:0]) begin
        image_2_221 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_222 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hde == _T_37[9:0]) begin
        image_2_222 <= io_pixelVal_in_2_7;
      end else if (10'hde == _T_34[9:0]) begin
        image_2_222 <= io_pixelVal_in_2_6;
      end else if (10'hde == _T_31[9:0]) begin
        image_2_222 <= io_pixelVal_in_2_5;
      end else if (10'hde == _T_28[9:0]) begin
        image_2_222 <= io_pixelVal_in_2_4;
      end else if (10'hde == _T_25[9:0]) begin
        image_2_222 <= io_pixelVal_in_2_3;
      end else if (10'hde == _T_22[9:0]) begin
        image_2_222 <= io_pixelVal_in_2_2;
      end else if (10'hde == _T_19[9:0]) begin
        image_2_222 <= io_pixelVal_in_2_1;
      end else if (10'hde == _T_15[9:0]) begin
        image_2_222 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_223 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hdf == _T_37[9:0]) begin
        image_2_223 <= io_pixelVal_in_2_7;
      end else if (10'hdf == _T_34[9:0]) begin
        image_2_223 <= io_pixelVal_in_2_6;
      end else if (10'hdf == _T_31[9:0]) begin
        image_2_223 <= io_pixelVal_in_2_5;
      end else if (10'hdf == _T_28[9:0]) begin
        image_2_223 <= io_pixelVal_in_2_4;
      end else if (10'hdf == _T_25[9:0]) begin
        image_2_223 <= io_pixelVal_in_2_3;
      end else if (10'hdf == _T_22[9:0]) begin
        image_2_223 <= io_pixelVal_in_2_2;
      end else if (10'hdf == _T_19[9:0]) begin
        image_2_223 <= io_pixelVal_in_2_1;
      end else if (10'hdf == _T_15[9:0]) begin
        image_2_223 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_224 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he0 == _T_37[9:0]) begin
        image_2_224 <= io_pixelVal_in_2_7;
      end else if (10'he0 == _T_34[9:0]) begin
        image_2_224 <= io_pixelVal_in_2_6;
      end else if (10'he0 == _T_31[9:0]) begin
        image_2_224 <= io_pixelVal_in_2_5;
      end else if (10'he0 == _T_28[9:0]) begin
        image_2_224 <= io_pixelVal_in_2_4;
      end else if (10'he0 == _T_25[9:0]) begin
        image_2_224 <= io_pixelVal_in_2_3;
      end else if (10'he0 == _T_22[9:0]) begin
        image_2_224 <= io_pixelVal_in_2_2;
      end else if (10'he0 == _T_19[9:0]) begin
        image_2_224 <= io_pixelVal_in_2_1;
      end else if (10'he0 == _T_15[9:0]) begin
        image_2_224 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_225 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he1 == _T_37[9:0]) begin
        image_2_225 <= io_pixelVal_in_2_7;
      end else if (10'he1 == _T_34[9:0]) begin
        image_2_225 <= io_pixelVal_in_2_6;
      end else if (10'he1 == _T_31[9:0]) begin
        image_2_225 <= io_pixelVal_in_2_5;
      end else if (10'he1 == _T_28[9:0]) begin
        image_2_225 <= io_pixelVal_in_2_4;
      end else if (10'he1 == _T_25[9:0]) begin
        image_2_225 <= io_pixelVal_in_2_3;
      end else if (10'he1 == _T_22[9:0]) begin
        image_2_225 <= io_pixelVal_in_2_2;
      end else if (10'he1 == _T_19[9:0]) begin
        image_2_225 <= io_pixelVal_in_2_1;
      end else if (10'he1 == _T_15[9:0]) begin
        image_2_225 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_226 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he2 == _T_37[9:0]) begin
        image_2_226 <= io_pixelVal_in_2_7;
      end else if (10'he2 == _T_34[9:0]) begin
        image_2_226 <= io_pixelVal_in_2_6;
      end else if (10'he2 == _T_31[9:0]) begin
        image_2_226 <= io_pixelVal_in_2_5;
      end else if (10'he2 == _T_28[9:0]) begin
        image_2_226 <= io_pixelVal_in_2_4;
      end else if (10'he2 == _T_25[9:0]) begin
        image_2_226 <= io_pixelVal_in_2_3;
      end else if (10'he2 == _T_22[9:0]) begin
        image_2_226 <= io_pixelVal_in_2_2;
      end else if (10'he2 == _T_19[9:0]) begin
        image_2_226 <= io_pixelVal_in_2_1;
      end else if (10'he2 == _T_15[9:0]) begin
        image_2_226 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_227 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he3 == _T_37[9:0]) begin
        image_2_227 <= io_pixelVal_in_2_7;
      end else if (10'he3 == _T_34[9:0]) begin
        image_2_227 <= io_pixelVal_in_2_6;
      end else if (10'he3 == _T_31[9:0]) begin
        image_2_227 <= io_pixelVal_in_2_5;
      end else if (10'he3 == _T_28[9:0]) begin
        image_2_227 <= io_pixelVal_in_2_4;
      end else if (10'he3 == _T_25[9:0]) begin
        image_2_227 <= io_pixelVal_in_2_3;
      end else if (10'he3 == _T_22[9:0]) begin
        image_2_227 <= io_pixelVal_in_2_2;
      end else if (10'he3 == _T_19[9:0]) begin
        image_2_227 <= io_pixelVal_in_2_1;
      end else if (10'he3 == _T_15[9:0]) begin
        image_2_227 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_228 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he4 == _T_37[9:0]) begin
        image_2_228 <= io_pixelVal_in_2_7;
      end else if (10'he4 == _T_34[9:0]) begin
        image_2_228 <= io_pixelVal_in_2_6;
      end else if (10'he4 == _T_31[9:0]) begin
        image_2_228 <= io_pixelVal_in_2_5;
      end else if (10'he4 == _T_28[9:0]) begin
        image_2_228 <= io_pixelVal_in_2_4;
      end else if (10'he4 == _T_25[9:0]) begin
        image_2_228 <= io_pixelVal_in_2_3;
      end else if (10'he4 == _T_22[9:0]) begin
        image_2_228 <= io_pixelVal_in_2_2;
      end else if (10'he4 == _T_19[9:0]) begin
        image_2_228 <= io_pixelVal_in_2_1;
      end else if (10'he4 == _T_15[9:0]) begin
        image_2_228 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_229 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he5 == _T_37[9:0]) begin
        image_2_229 <= io_pixelVal_in_2_7;
      end else if (10'he5 == _T_34[9:0]) begin
        image_2_229 <= io_pixelVal_in_2_6;
      end else if (10'he5 == _T_31[9:0]) begin
        image_2_229 <= io_pixelVal_in_2_5;
      end else if (10'he5 == _T_28[9:0]) begin
        image_2_229 <= io_pixelVal_in_2_4;
      end else if (10'he5 == _T_25[9:0]) begin
        image_2_229 <= io_pixelVal_in_2_3;
      end else if (10'he5 == _T_22[9:0]) begin
        image_2_229 <= io_pixelVal_in_2_2;
      end else if (10'he5 == _T_19[9:0]) begin
        image_2_229 <= io_pixelVal_in_2_1;
      end else if (10'he5 == _T_15[9:0]) begin
        image_2_229 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_230 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he6 == _T_37[9:0]) begin
        image_2_230 <= io_pixelVal_in_2_7;
      end else if (10'he6 == _T_34[9:0]) begin
        image_2_230 <= io_pixelVal_in_2_6;
      end else if (10'he6 == _T_31[9:0]) begin
        image_2_230 <= io_pixelVal_in_2_5;
      end else if (10'he6 == _T_28[9:0]) begin
        image_2_230 <= io_pixelVal_in_2_4;
      end else if (10'he6 == _T_25[9:0]) begin
        image_2_230 <= io_pixelVal_in_2_3;
      end else if (10'he6 == _T_22[9:0]) begin
        image_2_230 <= io_pixelVal_in_2_2;
      end else if (10'he6 == _T_19[9:0]) begin
        image_2_230 <= io_pixelVal_in_2_1;
      end else if (10'he6 == _T_15[9:0]) begin
        image_2_230 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_231 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he7 == _T_37[9:0]) begin
        image_2_231 <= io_pixelVal_in_2_7;
      end else if (10'he7 == _T_34[9:0]) begin
        image_2_231 <= io_pixelVal_in_2_6;
      end else if (10'he7 == _T_31[9:0]) begin
        image_2_231 <= io_pixelVal_in_2_5;
      end else if (10'he7 == _T_28[9:0]) begin
        image_2_231 <= io_pixelVal_in_2_4;
      end else if (10'he7 == _T_25[9:0]) begin
        image_2_231 <= io_pixelVal_in_2_3;
      end else if (10'he7 == _T_22[9:0]) begin
        image_2_231 <= io_pixelVal_in_2_2;
      end else if (10'he7 == _T_19[9:0]) begin
        image_2_231 <= io_pixelVal_in_2_1;
      end else if (10'he7 == _T_15[9:0]) begin
        image_2_231 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_232 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he8 == _T_37[9:0]) begin
        image_2_232 <= io_pixelVal_in_2_7;
      end else if (10'he8 == _T_34[9:0]) begin
        image_2_232 <= io_pixelVal_in_2_6;
      end else if (10'he8 == _T_31[9:0]) begin
        image_2_232 <= io_pixelVal_in_2_5;
      end else if (10'he8 == _T_28[9:0]) begin
        image_2_232 <= io_pixelVal_in_2_4;
      end else if (10'he8 == _T_25[9:0]) begin
        image_2_232 <= io_pixelVal_in_2_3;
      end else if (10'he8 == _T_22[9:0]) begin
        image_2_232 <= io_pixelVal_in_2_2;
      end else if (10'he8 == _T_19[9:0]) begin
        image_2_232 <= io_pixelVal_in_2_1;
      end else if (10'he8 == _T_15[9:0]) begin
        image_2_232 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_233 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he9 == _T_37[9:0]) begin
        image_2_233 <= io_pixelVal_in_2_7;
      end else if (10'he9 == _T_34[9:0]) begin
        image_2_233 <= io_pixelVal_in_2_6;
      end else if (10'he9 == _T_31[9:0]) begin
        image_2_233 <= io_pixelVal_in_2_5;
      end else if (10'he9 == _T_28[9:0]) begin
        image_2_233 <= io_pixelVal_in_2_4;
      end else if (10'he9 == _T_25[9:0]) begin
        image_2_233 <= io_pixelVal_in_2_3;
      end else if (10'he9 == _T_22[9:0]) begin
        image_2_233 <= io_pixelVal_in_2_2;
      end else if (10'he9 == _T_19[9:0]) begin
        image_2_233 <= io_pixelVal_in_2_1;
      end else if (10'he9 == _T_15[9:0]) begin
        image_2_233 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_234 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hea == _T_37[9:0]) begin
        image_2_234 <= io_pixelVal_in_2_7;
      end else if (10'hea == _T_34[9:0]) begin
        image_2_234 <= io_pixelVal_in_2_6;
      end else if (10'hea == _T_31[9:0]) begin
        image_2_234 <= io_pixelVal_in_2_5;
      end else if (10'hea == _T_28[9:0]) begin
        image_2_234 <= io_pixelVal_in_2_4;
      end else if (10'hea == _T_25[9:0]) begin
        image_2_234 <= io_pixelVal_in_2_3;
      end else if (10'hea == _T_22[9:0]) begin
        image_2_234 <= io_pixelVal_in_2_2;
      end else if (10'hea == _T_19[9:0]) begin
        image_2_234 <= io_pixelVal_in_2_1;
      end else if (10'hea == _T_15[9:0]) begin
        image_2_234 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_235 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'heb == _T_37[9:0]) begin
        image_2_235 <= io_pixelVal_in_2_7;
      end else if (10'heb == _T_34[9:0]) begin
        image_2_235 <= io_pixelVal_in_2_6;
      end else if (10'heb == _T_31[9:0]) begin
        image_2_235 <= io_pixelVal_in_2_5;
      end else if (10'heb == _T_28[9:0]) begin
        image_2_235 <= io_pixelVal_in_2_4;
      end else if (10'heb == _T_25[9:0]) begin
        image_2_235 <= io_pixelVal_in_2_3;
      end else if (10'heb == _T_22[9:0]) begin
        image_2_235 <= io_pixelVal_in_2_2;
      end else if (10'heb == _T_19[9:0]) begin
        image_2_235 <= io_pixelVal_in_2_1;
      end else if (10'heb == _T_15[9:0]) begin
        image_2_235 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_236 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hec == _T_37[9:0]) begin
        image_2_236 <= io_pixelVal_in_2_7;
      end else if (10'hec == _T_34[9:0]) begin
        image_2_236 <= io_pixelVal_in_2_6;
      end else if (10'hec == _T_31[9:0]) begin
        image_2_236 <= io_pixelVal_in_2_5;
      end else if (10'hec == _T_28[9:0]) begin
        image_2_236 <= io_pixelVal_in_2_4;
      end else if (10'hec == _T_25[9:0]) begin
        image_2_236 <= io_pixelVal_in_2_3;
      end else if (10'hec == _T_22[9:0]) begin
        image_2_236 <= io_pixelVal_in_2_2;
      end else if (10'hec == _T_19[9:0]) begin
        image_2_236 <= io_pixelVal_in_2_1;
      end else if (10'hec == _T_15[9:0]) begin
        image_2_236 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_237 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hed == _T_37[9:0]) begin
        image_2_237 <= io_pixelVal_in_2_7;
      end else if (10'hed == _T_34[9:0]) begin
        image_2_237 <= io_pixelVal_in_2_6;
      end else if (10'hed == _T_31[9:0]) begin
        image_2_237 <= io_pixelVal_in_2_5;
      end else if (10'hed == _T_28[9:0]) begin
        image_2_237 <= io_pixelVal_in_2_4;
      end else if (10'hed == _T_25[9:0]) begin
        image_2_237 <= io_pixelVal_in_2_3;
      end else if (10'hed == _T_22[9:0]) begin
        image_2_237 <= io_pixelVal_in_2_2;
      end else if (10'hed == _T_19[9:0]) begin
        image_2_237 <= io_pixelVal_in_2_1;
      end else if (10'hed == _T_15[9:0]) begin
        image_2_237 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_238 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hee == _T_37[9:0]) begin
        image_2_238 <= io_pixelVal_in_2_7;
      end else if (10'hee == _T_34[9:0]) begin
        image_2_238 <= io_pixelVal_in_2_6;
      end else if (10'hee == _T_31[9:0]) begin
        image_2_238 <= io_pixelVal_in_2_5;
      end else if (10'hee == _T_28[9:0]) begin
        image_2_238 <= io_pixelVal_in_2_4;
      end else if (10'hee == _T_25[9:0]) begin
        image_2_238 <= io_pixelVal_in_2_3;
      end else if (10'hee == _T_22[9:0]) begin
        image_2_238 <= io_pixelVal_in_2_2;
      end else if (10'hee == _T_19[9:0]) begin
        image_2_238 <= io_pixelVal_in_2_1;
      end else if (10'hee == _T_15[9:0]) begin
        image_2_238 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_239 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hef == _T_37[9:0]) begin
        image_2_239 <= io_pixelVal_in_2_7;
      end else if (10'hef == _T_34[9:0]) begin
        image_2_239 <= io_pixelVal_in_2_6;
      end else if (10'hef == _T_31[9:0]) begin
        image_2_239 <= io_pixelVal_in_2_5;
      end else if (10'hef == _T_28[9:0]) begin
        image_2_239 <= io_pixelVal_in_2_4;
      end else if (10'hef == _T_25[9:0]) begin
        image_2_239 <= io_pixelVal_in_2_3;
      end else if (10'hef == _T_22[9:0]) begin
        image_2_239 <= io_pixelVal_in_2_2;
      end else if (10'hef == _T_19[9:0]) begin
        image_2_239 <= io_pixelVal_in_2_1;
      end else if (10'hef == _T_15[9:0]) begin
        image_2_239 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_240 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf0 == _T_37[9:0]) begin
        image_2_240 <= io_pixelVal_in_2_7;
      end else if (10'hf0 == _T_34[9:0]) begin
        image_2_240 <= io_pixelVal_in_2_6;
      end else if (10'hf0 == _T_31[9:0]) begin
        image_2_240 <= io_pixelVal_in_2_5;
      end else if (10'hf0 == _T_28[9:0]) begin
        image_2_240 <= io_pixelVal_in_2_4;
      end else if (10'hf0 == _T_25[9:0]) begin
        image_2_240 <= io_pixelVal_in_2_3;
      end else if (10'hf0 == _T_22[9:0]) begin
        image_2_240 <= io_pixelVal_in_2_2;
      end else if (10'hf0 == _T_19[9:0]) begin
        image_2_240 <= io_pixelVal_in_2_1;
      end else if (10'hf0 == _T_15[9:0]) begin
        image_2_240 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_241 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf1 == _T_37[9:0]) begin
        image_2_241 <= io_pixelVal_in_2_7;
      end else if (10'hf1 == _T_34[9:0]) begin
        image_2_241 <= io_pixelVal_in_2_6;
      end else if (10'hf1 == _T_31[9:0]) begin
        image_2_241 <= io_pixelVal_in_2_5;
      end else if (10'hf1 == _T_28[9:0]) begin
        image_2_241 <= io_pixelVal_in_2_4;
      end else if (10'hf1 == _T_25[9:0]) begin
        image_2_241 <= io_pixelVal_in_2_3;
      end else if (10'hf1 == _T_22[9:0]) begin
        image_2_241 <= io_pixelVal_in_2_2;
      end else if (10'hf1 == _T_19[9:0]) begin
        image_2_241 <= io_pixelVal_in_2_1;
      end else if (10'hf1 == _T_15[9:0]) begin
        image_2_241 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_242 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf2 == _T_37[9:0]) begin
        image_2_242 <= io_pixelVal_in_2_7;
      end else if (10'hf2 == _T_34[9:0]) begin
        image_2_242 <= io_pixelVal_in_2_6;
      end else if (10'hf2 == _T_31[9:0]) begin
        image_2_242 <= io_pixelVal_in_2_5;
      end else if (10'hf2 == _T_28[9:0]) begin
        image_2_242 <= io_pixelVal_in_2_4;
      end else if (10'hf2 == _T_25[9:0]) begin
        image_2_242 <= io_pixelVal_in_2_3;
      end else if (10'hf2 == _T_22[9:0]) begin
        image_2_242 <= io_pixelVal_in_2_2;
      end else if (10'hf2 == _T_19[9:0]) begin
        image_2_242 <= io_pixelVal_in_2_1;
      end else if (10'hf2 == _T_15[9:0]) begin
        image_2_242 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_243 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf3 == _T_37[9:0]) begin
        image_2_243 <= io_pixelVal_in_2_7;
      end else if (10'hf3 == _T_34[9:0]) begin
        image_2_243 <= io_pixelVal_in_2_6;
      end else if (10'hf3 == _T_31[9:0]) begin
        image_2_243 <= io_pixelVal_in_2_5;
      end else if (10'hf3 == _T_28[9:0]) begin
        image_2_243 <= io_pixelVal_in_2_4;
      end else if (10'hf3 == _T_25[9:0]) begin
        image_2_243 <= io_pixelVal_in_2_3;
      end else if (10'hf3 == _T_22[9:0]) begin
        image_2_243 <= io_pixelVal_in_2_2;
      end else if (10'hf3 == _T_19[9:0]) begin
        image_2_243 <= io_pixelVal_in_2_1;
      end else if (10'hf3 == _T_15[9:0]) begin
        image_2_243 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_244 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf4 == _T_37[9:0]) begin
        image_2_244 <= io_pixelVal_in_2_7;
      end else if (10'hf4 == _T_34[9:0]) begin
        image_2_244 <= io_pixelVal_in_2_6;
      end else if (10'hf4 == _T_31[9:0]) begin
        image_2_244 <= io_pixelVal_in_2_5;
      end else if (10'hf4 == _T_28[9:0]) begin
        image_2_244 <= io_pixelVal_in_2_4;
      end else if (10'hf4 == _T_25[9:0]) begin
        image_2_244 <= io_pixelVal_in_2_3;
      end else if (10'hf4 == _T_22[9:0]) begin
        image_2_244 <= io_pixelVal_in_2_2;
      end else if (10'hf4 == _T_19[9:0]) begin
        image_2_244 <= io_pixelVal_in_2_1;
      end else if (10'hf4 == _T_15[9:0]) begin
        image_2_244 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_245 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf5 == _T_37[9:0]) begin
        image_2_245 <= io_pixelVal_in_2_7;
      end else if (10'hf5 == _T_34[9:0]) begin
        image_2_245 <= io_pixelVal_in_2_6;
      end else if (10'hf5 == _T_31[9:0]) begin
        image_2_245 <= io_pixelVal_in_2_5;
      end else if (10'hf5 == _T_28[9:0]) begin
        image_2_245 <= io_pixelVal_in_2_4;
      end else if (10'hf5 == _T_25[9:0]) begin
        image_2_245 <= io_pixelVal_in_2_3;
      end else if (10'hf5 == _T_22[9:0]) begin
        image_2_245 <= io_pixelVal_in_2_2;
      end else if (10'hf5 == _T_19[9:0]) begin
        image_2_245 <= io_pixelVal_in_2_1;
      end else if (10'hf5 == _T_15[9:0]) begin
        image_2_245 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_246 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf6 == _T_37[9:0]) begin
        image_2_246 <= io_pixelVal_in_2_7;
      end else if (10'hf6 == _T_34[9:0]) begin
        image_2_246 <= io_pixelVal_in_2_6;
      end else if (10'hf6 == _T_31[9:0]) begin
        image_2_246 <= io_pixelVal_in_2_5;
      end else if (10'hf6 == _T_28[9:0]) begin
        image_2_246 <= io_pixelVal_in_2_4;
      end else if (10'hf6 == _T_25[9:0]) begin
        image_2_246 <= io_pixelVal_in_2_3;
      end else if (10'hf6 == _T_22[9:0]) begin
        image_2_246 <= io_pixelVal_in_2_2;
      end else if (10'hf6 == _T_19[9:0]) begin
        image_2_246 <= io_pixelVal_in_2_1;
      end else if (10'hf6 == _T_15[9:0]) begin
        image_2_246 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_247 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf7 == _T_37[9:0]) begin
        image_2_247 <= io_pixelVal_in_2_7;
      end else if (10'hf7 == _T_34[9:0]) begin
        image_2_247 <= io_pixelVal_in_2_6;
      end else if (10'hf7 == _T_31[9:0]) begin
        image_2_247 <= io_pixelVal_in_2_5;
      end else if (10'hf7 == _T_28[9:0]) begin
        image_2_247 <= io_pixelVal_in_2_4;
      end else if (10'hf7 == _T_25[9:0]) begin
        image_2_247 <= io_pixelVal_in_2_3;
      end else if (10'hf7 == _T_22[9:0]) begin
        image_2_247 <= io_pixelVal_in_2_2;
      end else if (10'hf7 == _T_19[9:0]) begin
        image_2_247 <= io_pixelVal_in_2_1;
      end else if (10'hf7 == _T_15[9:0]) begin
        image_2_247 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_248 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf8 == _T_37[9:0]) begin
        image_2_248 <= io_pixelVal_in_2_7;
      end else if (10'hf8 == _T_34[9:0]) begin
        image_2_248 <= io_pixelVal_in_2_6;
      end else if (10'hf8 == _T_31[9:0]) begin
        image_2_248 <= io_pixelVal_in_2_5;
      end else if (10'hf8 == _T_28[9:0]) begin
        image_2_248 <= io_pixelVal_in_2_4;
      end else if (10'hf8 == _T_25[9:0]) begin
        image_2_248 <= io_pixelVal_in_2_3;
      end else if (10'hf8 == _T_22[9:0]) begin
        image_2_248 <= io_pixelVal_in_2_2;
      end else if (10'hf8 == _T_19[9:0]) begin
        image_2_248 <= io_pixelVal_in_2_1;
      end else if (10'hf8 == _T_15[9:0]) begin
        image_2_248 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_249 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf9 == _T_37[9:0]) begin
        image_2_249 <= io_pixelVal_in_2_7;
      end else if (10'hf9 == _T_34[9:0]) begin
        image_2_249 <= io_pixelVal_in_2_6;
      end else if (10'hf9 == _T_31[9:0]) begin
        image_2_249 <= io_pixelVal_in_2_5;
      end else if (10'hf9 == _T_28[9:0]) begin
        image_2_249 <= io_pixelVal_in_2_4;
      end else if (10'hf9 == _T_25[9:0]) begin
        image_2_249 <= io_pixelVal_in_2_3;
      end else if (10'hf9 == _T_22[9:0]) begin
        image_2_249 <= io_pixelVal_in_2_2;
      end else if (10'hf9 == _T_19[9:0]) begin
        image_2_249 <= io_pixelVal_in_2_1;
      end else if (10'hf9 == _T_15[9:0]) begin
        image_2_249 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_250 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hfa == _T_37[9:0]) begin
        image_2_250 <= io_pixelVal_in_2_7;
      end else if (10'hfa == _T_34[9:0]) begin
        image_2_250 <= io_pixelVal_in_2_6;
      end else if (10'hfa == _T_31[9:0]) begin
        image_2_250 <= io_pixelVal_in_2_5;
      end else if (10'hfa == _T_28[9:0]) begin
        image_2_250 <= io_pixelVal_in_2_4;
      end else if (10'hfa == _T_25[9:0]) begin
        image_2_250 <= io_pixelVal_in_2_3;
      end else if (10'hfa == _T_22[9:0]) begin
        image_2_250 <= io_pixelVal_in_2_2;
      end else if (10'hfa == _T_19[9:0]) begin
        image_2_250 <= io_pixelVal_in_2_1;
      end else if (10'hfa == _T_15[9:0]) begin
        image_2_250 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_251 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hfb == _T_37[9:0]) begin
        image_2_251 <= io_pixelVal_in_2_7;
      end else if (10'hfb == _T_34[9:0]) begin
        image_2_251 <= io_pixelVal_in_2_6;
      end else if (10'hfb == _T_31[9:0]) begin
        image_2_251 <= io_pixelVal_in_2_5;
      end else if (10'hfb == _T_28[9:0]) begin
        image_2_251 <= io_pixelVal_in_2_4;
      end else if (10'hfb == _T_25[9:0]) begin
        image_2_251 <= io_pixelVal_in_2_3;
      end else if (10'hfb == _T_22[9:0]) begin
        image_2_251 <= io_pixelVal_in_2_2;
      end else if (10'hfb == _T_19[9:0]) begin
        image_2_251 <= io_pixelVal_in_2_1;
      end else if (10'hfb == _T_15[9:0]) begin
        image_2_251 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_252 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hfc == _T_37[9:0]) begin
        image_2_252 <= io_pixelVal_in_2_7;
      end else if (10'hfc == _T_34[9:0]) begin
        image_2_252 <= io_pixelVal_in_2_6;
      end else if (10'hfc == _T_31[9:0]) begin
        image_2_252 <= io_pixelVal_in_2_5;
      end else if (10'hfc == _T_28[9:0]) begin
        image_2_252 <= io_pixelVal_in_2_4;
      end else if (10'hfc == _T_25[9:0]) begin
        image_2_252 <= io_pixelVal_in_2_3;
      end else if (10'hfc == _T_22[9:0]) begin
        image_2_252 <= io_pixelVal_in_2_2;
      end else if (10'hfc == _T_19[9:0]) begin
        image_2_252 <= io_pixelVal_in_2_1;
      end else if (10'hfc == _T_15[9:0]) begin
        image_2_252 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_253 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hfd == _T_37[9:0]) begin
        image_2_253 <= io_pixelVal_in_2_7;
      end else if (10'hfd == _T_34[9:0]) begin
        image_2_253 <= io_pixelVal_in_2_6;
      end else if (10'hfd == _T_31[9:0]) begin
        image_2_253 <= io_pixelVal_in_2_5;
      end else if (10'hfd == _T_28[9:0]) begin
        image_2_253 <= io_pixelVal_in_2_4;
      end else if (10'hfd == _T_25[9:0]) begin
        image_2_253 <= io_pixelVal_in_2_3;
      end else if (10'hfd == _T_22[9:0]) begin
        image_2_253 <= io_pixelVal_in_2_2;
      end else if (10'hfd == _T_19[9:0]) begin
        image_2_253 <= io_pixelVal_in_2_1;
      end else if (10'hfd == _T_15[9:0]) begin
        image_2_253 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_254 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hfe == _T_37[9:0]) begin
        image_2_254 <= io_pixelVal_in_2_7;
      end else if (10'hfe == _T_34[9:0]) begin
        image_2_254 <= io_pixelVal_in_2_6;
      end else if (10'hfe == _T_31[9:0]) begin
        image_2_254 <= io_pixelVal_in_2_5;
      end else if (10'hfe == _T_28[9:0]) begin
        image_2_254 <= io_pixelVal_in_2_4;
      end else if (10'hfe == _T_25[9:0]) begin
        image_2_254 <= io_pixelVal_in_2_3;
      end else if (10'hfe == _T_22[9:0]) begin
        image_2_254 <= io_pixelVal_in_2_2;
      end else if (10'hfe == _T_19[9:0]) begin
        image_2_254 <= io_pixelVal_in_2_1;
      end else if (10'hfe == _T_15[9:0]) begin
        image_2_254 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_255 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hff == _T_37[9:0]) begin
        image_2_255 <= io_pixelVal_in_2_7;
      end else if (10'hff == _T_34[9:0]) begin
        image_2_255 <= io_pixelVal_in_2_6;
      end else if (10'hff == _T_31[9:0]) begin
        image_2_255 <= io_pixelVal_in_2_5;
      end else if (10'hff == _T_28[9:0]) begin
        image_2_255 <= io_pixelVal_in_2_4;
      end else if (10'hff == _T_25[9:0]) begin
        image_2_255 <= io_pixelVal_in_2_3;
      end else if (10'hff == _T_22[9:0]) begin
        image_2_255 <= io_pixelVal_in_2_2;
      end else if (10'hff == _T_19[9:0]) begin
        image_2_255 <= io_pixelVal_in_2_1;
      end else if (10'hff == _T_15[9:0]) begin
        image_2_255 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_256 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h100 == _T_37[9:0]) begin
        image_2_256 <= io_pixelVal_in_2_7;
      end else if (10'h100 == _T_34[9:0]) begin
        image_2_256 <= io_pixelVal_in_2_6;
      end else if (10'h100 == _T_31[9:0]) begin
        image_2_256 <= io_pixelVal_in_2_5;
      end else if (10'h100 == _T_28[9:0]) begin
        image_2_256 <= io_pixelVal_in_2_4;
      end else if (10'h100 == _T_25[9:0]) begin
        image_2_256 <= io_pixelVal_in_2_3;
      end else if (10'h100 == _T_22[9:0]) begin
        image_2_256 <= io_pixelVal_in_2_2;
      end else if (10'h100 == _T_19[9:0]) begin
        image_2_256 <= io_pixelVal_in_2_1;
      end else if (10'h100 == _T_15[9:0]) begin
        image_2_256 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_257 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h101 == _T_37[9:0]) begin
        image_2_257 <= io_pixelVal_in_2_7;
      end else if (10'h101 == _T_34[9:0]) begin
        image_2_257 <= io_pixelVal_in_2_6;
      end else if (10'h101 == _T_31[9:0]) begin
        image_2_257 <= io_pixelVal_in_2_5;
      end else if (10'h101 == _T_28[9:0]) begin
        image_2_257 <= io_pixelVal_in_2_4;
      end else if (10'h101 == _T_25[9:0]) begin
        image_2_257 <= io_pixelVal_in_2_3;
      end else if (10'h101 == _T_22[9:0]) begin
        image_2_257 <= io_pixelVal_in_2_2;
      end else if (10'h101 == _T_19[9:0]) begin
        image_2_257 <= io_pixelVal_in_2_1;
      end else if (10'h101 == _T_15[9:0]) begin
        image_2_257 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_258 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h102 == _T_37[9:0]) begin
        image_2_258 <= io_pixelVal_in_2_7;
      end else if (10'h102 == _T_34[9:0]) begin
        image_2_258 <= io_pixelVal_in_2_6;
      end else if (10'h102 == _T_31[9:0]) begin
        image_2_258 <= io_pixelVal_in_2_5;
      end else if (10'h102 == _T_28[9:0]) begin
        image_2_258 <= io_pixelVal_in_2_4;
      end else if (10'h102 == _T_25[9:0]) begin
        image_2_258 <= io_pixelVal_in_2_3;
      end else if (10'h102 == _T_22[9:0]) begin
        image_2_258 <= io_pixelVal_in_2_2;
      end else if (10'h102 == _T_19[9:0]) begin
        image_2_258 <= io_pixelVal_in_2_1;
      end else if (10'h102 == _T_15[9:0]) begin
        image_2_258 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_259 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h103 == _T_37[9:0]) begin
        image_2_259 <= io_pixelVal_in_2_7;
      end else if (10'h103 == _T_34[9:0]) begin
        image_2_259 <= io_pixelVal_in_2_6;
      end else if (10'h103 == _T_31[9:0]) begin
        image_2_259 <= io_pixelVal_in_2_5;
      end else if (10'h103 == _T_28[9:0]) begin
        image_2_259 <= io_pixelVal_in_2_4;
      end else if (10'h103 == _T_25[9:0]) begin
        image_2_259 <= io_pixelVal_in_2_3;
      end else if (10'h103 == _T_22[9:0]) begin
        image_2_259 <= io_pixelVal_in_2_2;
      end else if (10'h103 == _T_19[9:0]) begin
        image_2_259 <= io_pixelVal_in_2_1;
      end else if (10'h103 == _T_15[9:0]) begin
        image_2_259 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_260 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h104 == _T_37[9:0]) begin
        image_2_260 <= io_pixelVal_in_2_7;
      end else if (10'h104 == _T_34[9:0]) begin
        image_2_260 <= io_pixelVal_in_2_6;
      end else if (10'h104 == _T_31[9:0]) begin
        image_2_260 <= io_pixelVal_in_2_5;
      end else if (10'h104 == _T_28[9:0]) begin
        image_2_260 <= io_pixelVal_in_2_4;
      end else if (10'h104 == _T_25[9:0]) begin
        image_2_260 <= io_pixelVal_in_2_3;
      end else if (10'h104 == _T_22[9:0]) begin
        image_2_260 <= io_pixelVal_in_2_2;
      end else if (10'h104 == _T_19[9:0]) begin
        image_2_260 <= io_pixelVal_in_2_1;
      end else if (10'h104 == _T_15[9:0]) begin
        image_2_260 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_261 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h105 == _T_37[9:0]) begin
        image_2_261 <= io_pixelVal_in_2_7;
      end else if (10'h105 == _T_34[9:0]) begin
        image_2_261 <= io_pixelVal_in_2_6;
      end else if (10'h105 == _T_31[9:0]) begin
        image_2_261 <= io_pixelVal_in_2_5;
      end else if (10'h105 == _T_28[9:0]) begin
        image_2_261 <= io_pixelVal_in_2_4;
      end else if (10'h105 == _T_25[9:0]) begin
        image_2_261 <= io_pixelVal_in_2_3;
      end else if (10'h105 == _T_22[9:0]) begin
        image_2_261 <= io_pixelVal_in_2_2;
      end else if (10'h105 == _T_19[9:0]) begin
        image_2_261 <= io_pixelVal_in_2_1;
      end else if (10'h105 == _T_15[9:0]) begin
        image_2_261 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_262 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h106 == _T_37[9:0]) begin
        image_2_262 <= io_pixelVal_in_2_7;
      end else if (10'h106 == _T_34[9:0]) begin
        image_2_262 <= io_pixelVal_in_2_6;
      end else if (10'h106 == _T_31[9:0]) begin
        image_2_262 <= io_pixelVal_in_2_5;
      end else if (10'h106 == _T_28[9:0]) begin
        image_2_262 <= io_pixelVal_in_2_4;
      end else if (10'h106 == _T_25[9:0]) begin
        image_2_262 <= io_pixelVal_in_2_3;
      end else if (10'h106 == _T_22[9:0]) begin
        image_2_262 <= io_pixelVal_in_2_2;
      end else if (10'h106 == _T_19[9:0]) begin
        image_2_262 <= io_pixelVal_in_2_1;
      end else if (10'h106 == _T_15[9:0]) begin
        image_2_262 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_263 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h107 == _T_37[9:0]) begin
        image_2_263 <= io_pixelVal_in_2_7;
      end else if (10'h107 == _T_34[9:0]) begin
        image_2_263 <= io_pixelVal_in_2_6;
      end else if (10'h107 == _T_31[9:0]) begin
        image_2_263 <= io_pixelVal_in_2_5;
      end else if (10'h107 == _T_28[9:0]) begin
        image_2_263 <= io_pixelVal_in_2_4;
      end else if (10'h107 == _T_25[9:0]) begin
        image_2_263 <= io_pixelVal_in_2_3;
      end else if (10'h107 == _T_22[9:0]) begin
        image_2_263 <= io_pixelVal_in_2_2;
      end else if (10'h107 == _T_19[9:0]) begin
        image_2_263 <= io_pixelVal_in_2_1;
      end else if (10'h107 == _T_15[9:0]) begin
        image_2_263 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_264 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h108 == _T_37[9:0]) begin
        image_2_264 <= io_pixelVal_in_2_7;
      end else if (10'h108 == _T_34[9:0]) begin
        image_2_264 <= io_pixelVal_in_2_6;
      end else if (10'h108 == _T_31[9:0]) begin
        image_2_264 <= io_pixelVal_in_2_5;
      end else if (10'h108 == _T_28[9:0]) begin
        image_2_264 <= io_pixelVal_in_2_4;
      end else if (10'h108 == _T_25[9:0]) begin
        image_2_264 <= io_pixelVal_in_2_3;
      end else if (10'h108 == _T_22[9:0]) begin
        image_2_264 <= io_pixelVal_in_2_2;
      end else if (10'h108 == _T_19[9:0]) begin
        image_2_264 <= io_pixelVal_in_2_1;
      end else if (10'h108 == _T_15[9:0]) begin
        image_2_264 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_265 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h109 == _T_37[9:0]) begin
        image_2_265 <= io_pixelVal_in_2_7;
      end else if (10'h109 == _T_34[9:0]) begin
        image_2_265 <= io_pixelVal_in_2_6;
      end else if (10'h109 == _T_31[9:0]) begin
        image_2_265 <= io_pixelVal_in_2_5;
      end else if (10'h109 == _T_28[9:0]) begin
        image_2_265 <= io_pixelVal_in_2_4;
      end else if (10'h109 == _T_25[9:0]) begin
        image_2_265 <= io_pixelVal_in_2_3;
      end else if (10'h109 == _T_22[9:0]) begin
        image_2_265 <= io_pixelVal_in_2_2;
      end else if (10'h109 == _T_19[9:0]) begin
        image_2_265 <= io_pixelVal_in_2_1;
      end else if (10'h109 == _T_15[9:0]) begin
        image_2_265 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_266 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10a == _T_37[9:0]) begin
        image_2_266 <= io_pixelVal_in_2_7;
      end else if (10'h10a == _T_34[9:0]) begin
        image_2_266 <= io_pixelVal_in_2_6;
      end else if (10'h10a == _T_31[9:0]) begin
        image_2_266 <= io_pixelVal_in_2_5;
      end else if (10'h10a == _T_28[9:0]) begin
        image_2_266 <= io_pixelVal_in_2_4;
      end else if (10'h10a == _T_25[9:0]) begin
        image_2_266 <= io_pixelVal_in_2_3;
      end else if (10'h10a == _T_22[9:0]) begin
        image_2_266 <= io_pixelVal_in_2_2;
      end else if (10'h10a == _T_19[9:0]) begin
        image_2_266 <= io_pixelVal_in_2_1;
      end else if (10'h10a == _T_15[9:0]) begin
        image_2_266 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_267 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10b == _T_37[9:0]) begin
        image_2_267 <= io_pixelVal_in_2_7;
      end else if (10'h10b == _T_34[9:0]) begin
        image_2_267 <= io_pixelVal_in_2_6;
      end else if (10'h10b == _T_31[9:0]) begin
        image_2_267 <= io_pixelVal_in_2_5;
      end else if (10'h10b == _T_28[9:0]) begin
        image_2_267 <= io_pixelVal_in_2_4;
      end else if (10'h10b == _T_25[9:0]) begin
        image_2_267 <= io_pixelVal_in_2_3;
      end else if (10'h10b == _T_22[9:0]) begin
        image_2_267 <= io_pixelVal_in_2_2;
      end else if (10'h10b == _T_19[9:0]) begin
        image_2_267 <= io_pixelVal_in_2_1;
      end else if (10'h10b == _T_15[9:0]) begin
        image_2_267 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_268 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10c == _T_37[9:0]) begin
        image_2_268 <= io_pixelVal_in_2_7;
      end else if (10'h10c == _T_34[9:0]) begin
        image_2_268 <= io_pixelVal_in_2_6;
      end else if (10'h10c == _T_31[9:0]) begin
        image_2_268 <= io_pixelVal_in_2_5;
      end else if (10'h10c == _T_28[9:0]) begin
        image_2_268 <= io_pixelVal_in_2_4;
      end else if (10'h10c == _T_25[9:0]) begin
        image_2_268 <= io_pixelVal_in_2_3;
      end else if (10'h10c == _T_22[9:0]) begin
        image_2_268 <= io_pixelVal_in_2_2;
      end else if (10'h10c == _T_19[9:0]) begin
        image_2_268 <= io_pixelVal_in_2_1;
      end else if (10'h10c == _T_15[9:0]) begin
        image_2_268 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_269 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10d == _T_37[9:0]) begin
        image_2_269 <= io_pixelVal_in_2_7;
      end else if (10'h10d == _T_34[9:0]) begin
        image_2_269 <= io_pixelVal_in_2_6;
      end else if (10'h10d == _T_31[9:0]) begin
        image_2_269 <= io_pixelVal_in_2_5;
      end else if (10'h10d == _T_28[9:0]) begin
        image_2_269 <= io_pixelVal_in_2_4;
      end else if (10'h10d == _T_25[9:0]) begin
        image_2_269 <= io_pixelVal_in_2_3;
      end else if (10'h10d == _T_22[9:0]) begin
        image_2_269 <= io_pixelVal_in_2_2;
      end else if (10'h10d == _T_19[9:0]) begin
        image_2_269 <= io_pixelVal_in_2_1;
      end else if (10'h10d == _T_15[9:0]) begin
        image_2_269 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_270 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10e == _T_37[9:0]) begin
        image_2_270 <= io_pixelVal_in_2_7;
      end else if (10'h10e == _T_34[9:0]) begin
        image_2_270 <= io_pixelVal_in_2_6;
      end else if (10'h10e == _T_31[9:0]) begin
        image_2_270 <= io_pixelVal_in_2_5;
      end else if (10'h10e == _T_28[9:0]) begin
        image_2_270 <= io_pixelVal_in_2_4;
      end else if (10'h10e == _T_25[9:0]) begin
        image_2_270 <= io_pixelVal_in_2_3;
      end else if (10'h10e == _T_22[9:0]) begin
        image_2_270 <= io_pixelVal_in_2_2;
      end else if (10'h10e == _T_19[9:0]) begin
        image_2_270 <= io_pixelVal_in_2_1;
      end else if (10'h10e == _T_15[9:0]) begin
        image_2_270 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_271 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10f == _T_37[9:0]) begin
        image_2_271 <= io_pixelVal_in_2_7;
      end else if (10'h10f == _T_34[9:0]) begin
        image_2_271 <= io_pixelVal_in_2_6;
      end else if (10'h10f == _T_31[9:0]) begin
        image_2_271 <= io_pixelVal_in_2_5;
      end else if (10'h10f == _T_28[9:0]) begin
        image_2_271 <= io_pixelVal_in_2_4;
      end else if (10'h10f == _T_25[9:0]) begin
        image_2_271 <= io_pixelVal_in_2_3;
      end else if (10'h10f == _T_22[9:0]) begin
        image_2_271 <= io_pixelVal_in_2_2;
      end else if (10'h10f == _T_19[9:0]) begin
        image_2_271 <= io_pixelVal_in_2_1;
      end else if (10'h10f == _T_15[9:0]) begin
        image_2_271 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_272 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h110 == _T_37[9:0]) begin
        image_2_272 <= io_pixelVal_in_2_7;
      end else if (10'h110 == _T_34[9:0]) begin
        image_2_272 <= io_pixelVal_in_2_6;
      end else if (10'h110 == _T_31[9:0]) begin
        image_2_272 <= io_pixelVal_in_2_5;
      end else if (10'h110 == _T_28[9:0]) begin
        image_2_272 <= io_pixelVal_in_2_4;
      end else if (10'h110 == _T_25[9:0]) begin
        image_2_272 <= io_pixelVal_in_2_3;
      end else if (10'h110 == _T_22[9:0]) begin
        image_2_272 <= io_pixelVal_in_2_2;
      end else if (10'h110 == _T_19[9:0]) begin
        image_2_272 <= io_pixelVal_in_2_1;
      end else if (10'h110 == _T_15[9:0]) begin
        image_2_272 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_273 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h111 == _T_37[9:0]) begin
        image_2_273 <= io_pixelVal_in_2_7;
      end else if (10'h111 == _T_34[9:0]) begin
        image_2_273 <= io_pixelVal_in_2_6;
      end else if (10'h111 == _T_31[9:0]) begin
        image_2_273 <= io_pixelVal_in_2_5;
      end else if (10'h111 == _T_28[9:0]) begin
        image_2_273 <= io_pixelVal_in_2_4;
      end else if (10'h111 == _T_25[9:0]) begin
        image_2_273 <= io_pixelVal_in_2_3;
      end else if (10'h111 == _T_22[9:0]) begin
        image_2_273 <= io_pixelVal_in_2_2;
      end else if (10'h111 == _T_19[9:0]) begin
        image_2_273 <= io_pixelVal_in_2_1;
      end else if (10'h111 == _T_15[9:0]) begin
        image_2_273 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_274 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h112 == _T_37[9:0]) begin
        image_2_274 <= io_pixelVal_in_2_7;
      end else if (10'h112 == _T_34[9:0]) begin
        image_2_274 <= io_pixelVal_in_2_6;
      end else if (10'h112 == _T_31[9:0]) begin
        image_2_274 <= io_pixelVal_in_2_5;
      end else if (10'h112 == _T_28[9:0]) begin
        image_2_274 <= io_pixelVal_in_2_4;
      end else if (10'h112 == _T_25[9:0]) begin
        image_2_274 <= io_pixelVal_in_2_3;
      end else if (10'h112 == _T_22[9:0]) begin
        image_2_274 <= io_pixelVal_in_2_2;
      end else if (10'h112 == _T_19[9:0]) begin
        image_2_274 <= io_pixelVal_in_2_1;
      end else if (10'h112 == _T_15[9:0]) begin
        image_2_274 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_275 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h113 == _T_37[9:0]) begin
        image_2_275 <= io_pixelVal_in_2_7;
      end else if (10'h113 == _T_34[9:0]) begin
        image_2_275 <= io_pixelVal_in_2_6;
      end else if (10'h113 == _T_31[9:0]) begin
        image_2_275 <= io_pixelVal_in_2_5;
      end else if (10'h113 == _T_28[9:0]) begin
        image_2_275 <= io_pixelVal_in_2_4;
      end else if (10'h113 == _T_25[9:0]) begin
        image_2_275 <= io_pixelVal_in_2_3;
      end else if (10'h113 == _T_22[9:0]) begin
        image_2_275 <= io_pixelVal_in_2_2;
      end else if (10'h113 == _T_19[9:0]) begin
        image_2_275 <= io_pixelVal_in_2_1;
      end else if (10'h113 == _T_15[9:0]) begin
        image_2_275 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_276 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h114 == _T_37[9:0]) begin
        image_2_276 <= io_pixelVal_in_2_7;
      end else if (10'h114 == _T_34[9:0]) begin
        image_2_276 <= io_pixelVal_in_2_6;
      end else if (10'h114 == _T_31[9:0]) begin
        image_2_276 <= io_pixelVal_in_2_5;
      end else if (10'h114 == _T_28[9:0]) begin
        image_2_276 <= io_pixelVal_in_2_4;
      end else if (10'h114 == _T_25[9:0]) begin
        image_2_276 <= io_pixelVal_in_2_3;
      end else if (10'h114 == _T_22[9:0]) begin
        image_2_276 <= io_pixelVal_in_2_2;
      end else if (10'h114 == _T_19[9:0]) begin
        image_2_276 <= io_pixelVal_in_2_1;
      end else if (10'h114 == _T_15[9:0]) begin
        image_2_276 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_277 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h115 == _T_37[9:0]) begin
        image_2_277 <= io_pixelVal_in_2_7;
      end else if (10'h115 == _T_34[9:0]) begin
        image_2_277 <= io_pixelVal_in_2_6;
      end else if (10'h115 == _T_31[9:0]) begin
        image_2_277 <= io_pixelVal_in_2_5;
      end else if (10'h115 == _T_28[9:0]) begin
        image_2_277 <= io_pixelVal_in_2_4;
      end else if (10'h115 == _T_25[9:0]) begin
        image_2_277 <= io_pixelVal_in_2_3;
      end else if (10'h115 == _T_22[9:0]) begin
        image_2_277 <= io_pixelVal_in_2_2;
      end else if (10'h115 == _T_19[9:0]) begin
        image_2_277 <= io_pixelVal_in_2_1;
      end else if (10'h115 == _T_15[9:0]) begin
        image_2_277 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_278 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h116 == _T_37[9:0]) begin
        image_2_278 <= io_pixelVal_in_2_7;
      end else if (10'h116 == _T_34[9:0]) begin
        image_2_278 <= io_pixelVal_in_2_6;
      end else if (10'h116 == _T_31[9:0]) begin
        image_2_278 <= io_pixelVal_in_2_5;
      end else if (10'h116 == _T_28[9:0]) begin
        image_2_278 <= io_pixelVal_in_2_4;
      end else if (10'h116 == _T_25[9:0]) begin
        image_2_278 <= io_pixelVal_in_2_3;
      end else if (10'h116 == _T_22[9:0]) begin
        image_2_278 <= io_pixelVal_in_2_2;
      end else if (10'h116 == _T_19[9:0]) begin
        image_2_278 <= io_pixelVal_in_2_1;
      end else if (10'h116 == _T_15[9:0]) begin
        image_2_278 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_279 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h117 == _T_37[9:0]) begin
        image_2_279 <= io_pixelVal_in_2_7;
      end else if (10'h117 == _T_34[9:0]) begin
        image_2_279 <= io_pixelVal_in_2_6;
      end else if (10'h117 == _T_31[9:0]) begin
        image_2_279 <= io_pixelVal_in_2_5;
      end else if (10'h117 == _T_28[9:0]) begin
        image_2_279 <= io_pixelVal_in_2_4;
      end else if (10'h117 == _T_25[9:0]) begin
        image_2_279 <= io_pixelVal_in_2_3;
      end else if (10'h117 == _T_22[9:0]) begin
        image_2_279 <= io_pixelVal_in_2_2;
      end else if (10'h117 == _T_19[9:0]) begin
        image_2_279 <= io_pixelVal_in_2_1;
      end else if (10'h117 == _T_15[9:0]) begin
        image_2_279 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_280 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h118 == _T_37[9:0]) begin
        image_2_280 <= io_pixelVal_in_2_7;
      end else if (10'h118 == _T_34[9:0]) begin
        image_2_280 <= io_pixelVal_in_2_6;
      end else if (10'h118 == _T_31[9:0]) begin
        image_2_280 <= io_pixelVal_in_2_5;
      end else if (10'h118 == _T_28[9:0]) begin
        image_2_280 <= io_pixelVal_in_2_4;
      end else if (10'h118 == _T_25[9:0]) begin
        image_2_280 <= io_pixelVal_in_2_3;
      end else if (10'h118 == _T_22[9:0]) begin
        image_2_280 <= io_pixelVal_in_2_2;
      end else if (10'h118 == _T_19[9:0]) begin
        image_2_280 <= io_pixelVal_in_2_1;
      end else if (10'h118 == _T_15[9:0]) begin
        image_2_280 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_281 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h119 == _T_37[9:0]) begin
        image_2_281 <= io_pixelVal_in_2_7;
      end else if (10'h119 == _T_34[9:0]) begin
        image_2_281 <= io_pixelVal_in_2_6;
      end else if (10'h119 == _T_31[9:0]) begin
        image_2_281 <= io_pixelVal_in_2_5;
      end else if (10'h119 == _T_28[9:0]) begin
        image_2_281 <= io_pixelVal_in_2_4;
      end else if (10'h119 == _T_25[9:0]) begin
        image_2_281 <= io_pixelVal_in_2_3;
      end else if (10'h119 == _T_22[9:0]) begin
        image_2_281 <= io_pixelVal_in_2_2;
      end else if (10'h119 == _T_19[9:0]) begin
        image_2_281 <= io_pixelVal_in_2_1;
      end else if (10'h119 == _T_15[9:0]) begin
        image_2_281 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_282 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11a == _T_37[9:0]) begin
        image_2_282 <= io_pixelVal_in_2_7;
      end else if (10'h11a == _T_34[9:0]) begin
        image_2_282 <= io_pixelVal_in_2_6;
      end else if (10'h11a == _T_31[9:0]) begin
        image_2_282 <= io_pixelVal_in_2_5;
      end else if (10'h11a == _T_28[9:0]) begin
        image_2_282 <= io_pixelVal_in_2_4;
      end else if (10'h11a == _T_25[9:0]) begin
        image_2_282 <= io_pixelVal_in_2_3;
      end else if (10'h11a == _T_22[9:0]) begin
        image_2_282 <= io_pixelVal_in_2_2;
      end else if (10'h11a == _T_19[9:0]) begin
        image_2_282 <= io_pixelVal_in_2_1;
      end else if (10'h11a == _T_15[9:0]) begin
        image_2_282 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_283 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11b == _T_37[9:0]) begin
        image_2_283 <= io_pixelVal_in_2_7;
      end else if (10'h11b == _T_34[9:0]) begin
        image_2_283 <= io_pixelVal_in_2_6;
      end else if (10'h11b == _T_31[9:0]) begin
        image_2_283 <= io_pixelVal_in_2_5;
      end else if (10'h11b == _T_28[9:0]) begin
        image_2_283 <= io_pixelVal_in_2_4;
      end else if (10'h11b == _T_25[9:0]) begin
        image_2_283 <= io_pixelVal_in_2_3;
      end else if (10'h11b == _T_22[9:0]) begin
        image_2_283 <= io_pixelVal_in_2_2;
      end else if (10'h11b == _T_19[9:0]) begin
        image_2_283 <= io_pixelVal_in_2_1;
      end else if (10'h11b == _T_15[9:0]) begin
        image_2_283 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_284 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11c == _T_37[9:0]) begin
        image_2_284 <= io_pixelVal_in_2_7;
      end else if (10'h11c == _T_34[9:0]) begin
        image_2_284 <= io_pixelVal_in_2_6;
      end else if (10'h11c == _T_31[9:0]) begin
        image_2_284 <= io_pixelVal_in_2_5;
      end else if (10'h11c == _T_28[9:0]) begin
        image_2_284 <= io_pixelVal_in_2_4;
      end else if (10'h11c == _T_25[9:0]) begin
        image_2_284 <= io_pixelVal_in_2_3;
      end else if (10'h11c == _T_22[9:0]) begin
        image_2_284 <= io_pixelVal_in_2_2;
      end else if (10'h11c == _T_19[9:0]) begin
        image_2_284 <= io_pixelVal_in_2_1;
      end else if (10'h11c == _T_15[9:0]) begin
        image_2_284 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_285 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11d == _T_37[9:0]) begin
        image_2_285 <= io_pixelVal_in_2_7;
      end else if (10'h11d == _T_34[9:0]) begin
        image_2_285 <= io_pixelVal_in_2_6;
      end else if (10'h11d == _T_31[9:0]) begin
        image_2_285 <= io_pixelVal_in_2_5;
      end else if (10'h11d == _T_28[9:0]) begin
        image_2_285 <= io_pixelVal_in_2_4;
      end else if (10'h11d == _T_25[9:0]) begin
        image_2_285 <= io_pixelVal_in_2_3;
      end else if (10'h11d == _T_22[9:0]) begin
        image_2_285 <= io_pixelVal_in_2_2;
      end else if (10'h11d == _T_19[9:0]) begin
        image_2_285 <= io_pixelVal_in_2_1;
      end else if (10'h11d == _T_15[9:0]) begin
        image_2_285 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_286 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11e == _T_37[9:0]) begin
        image_2_286 <= io_pixelVal_in_2_7;
      end else if (10'h11e == _T_34[9:0]) begin
        image_2_286 <= io_pixelVal_in_2_6;
      end else if (10'h11e == _T_31[9:0]) begin
        image_2_286 <= io_pixelVal_in_2_5;
      end else if (10'h11e == _T_28[9:0]) begin
        image_2_286 <= io_pixelVal_in_2_4;
      end else if (10'h11e == _T_25[9:0]) begin
        image_2_286 <= io_pixelVal_in_2_3;
      end else if (10'h11e == _T_22[9:0]) begin
        image_2_286 <= io_pixelVal_in_2_2;
      end else if (10'h11e == _T_19[9:0]) begin
        image_2_286 <= io_pixelVal_in_2_1;
      end else if (10'h11e == _T_15[9:0]) begin
        image_2_286 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_287 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11f == _T_37[9:0]) begin
        image_2_287 <= io_pixelVal_in_2_7;
      end else if (10'h11f == _T_34[9:0]) begin
        image_2_287 <= io_pixelVal_in_2_6;
      end else if (10'h11f == _T_31[9:0]) begin
        image_2_287 <= io_pixelVal_in_2_5;
      end else if (10'h11f == _T_28[9:0]) begin
        image_2_287 <= io_pixelVal_in_2_4;
      end else if (10'h11f == _T_25[9:0]) begin
        image_2_287 <= io_pixelVal_in_2_3;
      end else if (10'h11f == _T_22[9:0]) begin
        image_2_287 <= io_pixelVal_in_2_2;
      end else if (10'h11f == _T_19[9:0]) begin
        image_2_287 <= io_pixelVal_in_2_1;
      end else if (10'h11f == _T_15[9:0]) begin
        image_2_287 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_288 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h120 == _T_37[9:0]) begin
        image_2_288 <= io_pixelVal_in_2_7;
      end else if (10'h120 == _T_34[9:0]) begin
        image_2_288 <= io_pixelVal_in_2_6;
      end else if (10'h120 == _T_31[9:0]) begin
        image_2_288 <= io_pixelVal_in_2_5;
      end else if (10'h120 == _T_28[9:0]) begin
        image_2_288 <= io_pixelVal_in_2_4;
      end else if (10'h120 == _T_25[9:0]) begin
        image_2_288 <= io_pixelVal_in_2_3;
      end else if (10'h120 == _T_22[9:0]) begin
        image_2_288 <= io_pixelVal_in_2_2;
      end else if (10'h120 == _T_19[9:0]) begin
        image_2_288 <= io_pixelVal_in_2_1;
      end else if (10'h120 == _T_15[9:0]) begin
        image_2_288 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_289 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h121 == _T_37[9:0]) begin
        image_2_289 <= io_pixelVal_in_2_7;
      end else if (10'h121 == _T_34[9:0]) begin
        image_2_289 <= io_pixelVal_in_2_6;
      end else if (10'h121 == _T_31[9:0]) begin
        image_2_289 <= io_pixelVal_in_2_5;
      end else if (10'h121 == _T_28[9:0]) begin
        image_2_289 <= io_pixelVal_in_2_4;
      end else if (10'h121 == _T_25[9:0]) begin
        image_2_289 <= io_pixelVal_in_2_3;
      end else if (10'h121 == _T_22[9:0]) begin
        image_2_289 <= io_pixelVal_in_2_2;
      end else if (10'h121 == _T_19[9:0]) begin
        image_2_289 <= io_pixelVal_in_2_1;
      end else if (10'h121 == _T_15[9:0]) begin
        image_2_289 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_290 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h122 == _T_37[9:0]) begin
        image_2_290 <= io_pixelVal_in_2_7;
      end else if (10'h122 == _T_34[9:0]) begin
        image_2_290 <= io_pixelVal_in_2_6;
      end else if (10'h122 == _T_31[9:0]) begin
        image_2_290 <= io_pixelVal_in_2_5;
      end else if (10'h122 == _T_28[9:0]) begin
        image_2_290 <= io_pixelVal_in_2_4;
      end else if (10'h122 == _T_25[9:0]) begin
        image_2_290 <= io_pixelVal_in_2_3;
      end else if (10'h122 == _T_22[9:0]) begin
        image_2_290 <= io_pixelVal_in_2_2;
      end else if (10'h122 == _T_19[9:0]) begin
        image_2_290 <= io_pixelVal_in_2_1;
      end else if (10'h122 == _T_15[9:0]) begin
        image_2_290 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_291 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h123 == _T_37[9:0]) begin
        image_2_291 <= io_pixelVal_in_2_7;
      end else if (10'h123 == _T_34[9:0]) begin
        image_2_291 <= io_pixelVal_in_2_6;
      end else if (10'h123 == _T_31[9:0]) begin
        image_2_291 <= io_pixelVal_in_2_5;
      end else if (10'h123 == _T_28[9:0]) begin
        image_2_291 <= io_pixelVal_in_2_4;
      end else if (10'h123 == _T_25[9:0]) begin
        image_2_291 <= io_pixelVal_in_2_3;
      end else if (10'h123 == _T_22[9:0]) begin
        image_2_291 <= io_pixelVal_in_2_2;
      end else if (10'h123 == _T_19[9:0]) begin
        image_2_291 <= io_pixelVal_in_2_1;
      end else if (10'h123 == _T_15[9:0]) begin
        image_2_291 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_292 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h124 == _T_37[9:0]) begin
        image_2_292 <= io_pixelVal_in_2_7;
      end else if (10'h124 == _T_34[9:0]) begin
        image_2_292 <= io_pixelVal_in_2_6;
      end else if (10'h124 == _T_31[9:0]) begin
        image_2_292 <= io_pixelVal_in_2_5;
      end else if (10'h124 == _T_28[9:0]) begin
        image_2_292 <= io_pixelVal_in_2_4;
      end else if (10'h124 == _T_25[9:0]) begin
        image_2_292 <= io_pixelVal_in_2_3;
      end else if (10'h124 == _T_22[9:0]) begin
        image_2_292 <= io_pixelVal_in_2_2;
      end else if (10'h124 == _T_19[9:0]) begin
        image_2_292 <= io_pixelVal_in_2_1;
      end else if (10'h124 == _T_15[9:0]) begin
        image_2_292 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_293 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h125 == _T_37[9:0]) begin
        image_2_293 <= io_pixelVal_in_2_7;
      end else if (10'h125 == _T_34[9:0]) begin
        image_2_293 <= io_pixelVal_in_2_6;
      end else if (10'h125 == _T_31[9:0]) begin
        image_2_293 <= io_pixelVal_in_2_5;
      end else if (10'h125 == _T_28[9:0]) begin
        image_2_293 <= io_pixelVal_in_2_4;
      end else if (10'h125 == _T_25[9:0]) begin
        image_2_293 <= io_pixelVal_in_2_3;
      end else if (10'h125 == _T_22[9:0]) begin
        image_2_293 <= io_pixelVal_in_2_2;
      end else if (10'h125 == _T_19[9:0]) begin
        image_2_293 <= io_pixelVal_in_2_1;
      end else if (10'h125 == _T_15[9:0]) begin
        image_2_293 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_294 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h126 == _T_37[9:0]) begin
        image_2_294 <= io_pixelVal_in_2_7;
      end else if (10'h126 == _T_34[9:0]) begin
        image_2_294 <= io_pixelVal_in_2_6;
      end else if (10'h126 == _T_31[9:0]) begin
        image_2_294 <= io_pixelVal_in_2_5;
      end else if (10'h126 == _T_28[9:0]) begin
        image_2_294 <= io_pixelVal_in_2_4;
      end else if (10'h126 == _T_25[9:0]) begin
        image_2_294 <= io_pixelVal_in_2_3;
      end else if (10'h126 == _T_22[9:0]) begin
        image_2_294 <= io_pixelVal_in_2_2;
      end else if (10'h126 == _T_19[9:0]) begin
        image_2_294 <= io_pixelVal_in_2_1;
      end else if (10'h126 == _T_15[9:0]) begin
        image_2_294 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_295 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h127 == _T_37[9:0]) begin
        image_2_295 <= io_pixelVal_in_2_7;
      end else if (10'h127 == _T_34[9:0]) begin
        image_2_295 <= io_pixelVal_in_2_6;
      end else if (10'h127 == _T_31[9:0]) begin
        image_2_295 <= io_pixelVal_in_2_5;
      end else if (10'h127 == _T_28[9:0]) begin
        image_2_295 <= io_pixelVal_in_2_4;
      end else if (10'h127 == _T_25[9:0]) begin
        image_2_295 <= io_pixelVal_in_2_3;
      end else if (10'h127 == _T_22[9:0]) begin
        image_2_295 <= io_pixelVal_in_2_2;
      end else if (10'h127 == _T_19[9:0]) begin
        image_2_295 <= io_pixelVal_in_2_1;
      end else if (10'h127 == _T_15[9:0]) begin
        image_2_295 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_296 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h128 == _T_37[9:0]) begin
        image_2_296 <= io_pixelVal_in_2_7;
      end else if (10'h128 == _T_34[9:0]) begin
        image_2_296 <= io_pixelVal_in_2_6;
      end else if (10'h128 == _T_31[9:0]) begin
        image_2_296 <= io_pixelVal_in_2_5;
      end else if (10'h128 == _T_28[9:0]) begin
        image_2_296 <= io_pixelVal_in_2_4;
      end else if (10'h128 == _T_25[9:0]) begin
        image_2_296 <= io_pixelVal_in_2_3;
      end else if (10'h128 == _T_22[9:0]) begin
        image_2_296 <= io_pixelVal_in_2_2;
      end else if (10'h128 == _T_19[9:0]) begin
        image_2_296 <= io_pixelVal_in_2_1;
      end else if (10'h128 == _T_15[9:0]) begin
        image_2_296 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_297 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h129 == _T_37[9:0]) begin
        image_2_297 <= io_pixelVal_in_2_7;
      end else if (10'h129 == _T_34[9:0]) begin
        image_2_297 <= io_pixelVal_in_2_6;
      end else if (10'h129 == _T_31[9:0]) begin
        image_2_297 <= io_pixelVal_in_2_5;
      end else if (10'h129 == _T_28[9:0]) begin
        image_2_297 <= io_pixelVal_in_2_4;
      end else if (10'h129 == _T_25[9:0]) begin
        image_2_297 <= io_pixelVal_in_2_3;
      end else if (10'h129 == _T_22[9:0]) begin
        image_2_297 <= io_pixelVal_in_2_2;
      end else if (10'h129 == _T_19[9:0]) begin
        image_2_297 <= io_pixelVal_in_2_1;
      end else if (10'h129 == _T_15[9:0]) begin
        image_2_297 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_298 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12a == _T_37[9:0]) begin
        image_2_298 <= io_pixelVal_in_2_7;
      end else if (10'h12a == _T_34[9:0]) begin
        image_2_298 <= io_pixelVal_in_2_6;
      end else if (10'h12a == _T_31[9:0]) begin
        image_2_298 <= io_pixelVal_in_2_5;
      end else if (10'h12a == _T_28[9:0]) begin
        image_2_298 <= io_pixelVal_in_2_4;
      end else if (10'h12a == _T_25[9:0]) begin
        image_2_298 <= io_pixelVal_in_2_3;
      end else if (10'h12a == _T_22[9:0]) begin
        image_2_298 <= io_pixelVal_in_2_2;
      end else if (10'h12a == _T_19[9:0]) begin
        image_2_298 <= io_pixelVal_in_2_1;
      end else if (10'h12a == _T_15[9:0]) begin
        image_2_298 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_299 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12b == _T_37[9:0]) begin
        image_2_299 <= io_pixelVal_in_2_7;
      end else if (10'h12b == _T_34[9:0]) begin
        image_2_299 <= io_pixelVal_in_2_6;
      end else if (10'h12b == _T_31[9:0]) begin
        image_2_299 <= io_pixelVal_in_2_5;
      end else if (10'h12b == _T_28[9:0]) begin
        image_2_299 <= io_pixelVal_in_2_4;
      end else if (10'h12b == _T_25[9:0]) begin
        image_2_299 <= io_pixelVal_in_2_3;
      end else if (10'h12b == _T_22[9:0]) begin
        image_2_299 <= io_pixelVal_in_2_2;
      end else if (10'h12b == _T_19[9:0]) begin
        image_2_299 <= io_pixelVal_in_2_1;
      end else if (10'h12b == _T_15[9:0]) begin
        image_2_299 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_300 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12c == _T_37[9:0]) begin
        image_2_300 <= io_pixelVal_in_2_7;
      end else if (10'h12c == _T_34[9:0]) begin
        image_2_300 <= io_pixelVal_in_2_6;
      end else if (10'h12c == _T_31[9:0]) begin
        image_2_300 <= io_pixelVal_in_2_5;
      end else if (10'h12c == _T_28[9:0]) begin
        image_2_300 <= io_pixelVal_in_2_4;
      end else if (10'h12c == _T_25[9:0]) begin
        image_2_300 <= io_pixelVal_in_2_3;
      end else if (10'h12c == _T_22[9:0]) begin
        image_2_300 <= io_pixelVal_in_2_2;
      end else if (10'h12c == _T_19[9:0]) begin
        image_2_300 <= io_pixelVal_in_2_1;
      end else if (10'h12c == _T_15[9:0]) begin
        image_2_300 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_301 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12d == _T_37[9:0]) begin
        image_2_301 <= io_pixelVal_in_2_7;
      end else if (10'h12d == _T_34[9:0]) begin
        image_2_301 <= io_pixelVal_in_2_6;
      end else if (10'h12d == _T_31[9:0]) begin
        image_2_301 <= io_pixelVal_in_2_5;
      end else if (10'h12d == _T_28[9:0]) begin
        image_2_301 <= io_pixelVal_in_2_4;
      end else if (10'h12d == _T_25[9:0]) begin
        image_2_301 <= io_pixelVal_in_2_3;
      end else if (10'h12d == _T_22[9:0]) begin
        image_2_301 <= io_pixelVal_in_2_2;
      end else if (10'h12d == _T_19[9:0]) begin
        image_2_301 <= io_pixelVal_in_2_1;
      end else if (10'h12d == _T_15[9:0]) begin
        image_2_301 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_302 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12e == _T_37[9:0]) begin
        image_2_302 <= io_pixelVal_in_2_7;
      end else if (10'h12e == _T_34[9:0]) begin
        image_2_302 <= io_pixelVal_in_2_6;
      end else if (10'h12e == _T_31[9:0]) begin
        image_2_302 <= io_pixelVal_in_2_5;
      end else if (10'h12e == _T_28[9:0]) begin
        image_2_302 <= io_pixelVal_in_2_4;
      end else if (10'h12e == _T_25[9:0]) begin
        image_2_302 <= io_pixelVal_in_2_3;
      end else if (10'h12e == _T_22[9:0]) begin
        image_2_302 <= io_pixelVal_in_2_2;
      end else if (10'h12e == _T_19[9:0]) begin
        image_2_302 <= io_pixelVal_in_2_1;
      end else if (10'h12e == _T_15[9:0]) begin
        image_2_302 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_303 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12f == _T_37[9:0]) begin
        image_2_303 <= io_pixelVal_in_2_7;
      end else if (10'h12f == _T_34[9:0]) begin
        image_2_303 <= io_pixelVal_in_2_6;
      end else if (10'h12f == _T_31[9:0]) begin
        image_2_303 <= io_pixelVal_in_2_5;
      end else if (10'h12f == _T_28[9:0]) begin
        image_2_303 <= io_pixelVal_in_2_4;
      end else if (10'h12f == _T_25[9:0]) begin
        image_2_303 <= io_pixelVal_in_2_3;
      end else if (10'h12f == _T_22[9:0]) begin
        image_2_303 <= io_pixelVal_in_2_2;
      end else if (10'h12f == _T_19[9:0]) begin
        image_2_303 <= io_pixelVal_in_2_1;
      end else if (10'h12f == _T_15[9:0]) begin
        image_2_303 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_304 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h130 == _T_37[9:0]) begin
        image_2_304 <= io_pixelVal_in_2_7;
      end else if (10'h130 == _T_34[9:0]) begin
        image_2_304 <= io_pixelVal_in_2_6;
      end else if (10'h130 == _T_31[9:0]) begin
        image_2_304 <= io_pixelVal_in_2_5;
      end else if (10'h130 == _T_28[9:0]) begin
        image_2_304 <= io_pixelVal_in_2_4;
      end else if (10'h130 == _T_25[9:0]) begin
        image_2_304 <= io_pixelVal_in_2_3;
      end else if (10'h130 == _T_22[9:0]) begin
        image_2_304 <= io_pixelVal_in_2_2;
      end else if (10'h130 == _T_19[9:0]) begin
        image_2_304 <= io_pixelVal_in_2_1;
      end else if (10'h130 == _T_15[9:0]) begin
        image_2_304 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_305 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h131 == _T_37[9:0]) begin
        image_2_305 <= io_pixelVal_in_2_7;
      end else if (10'h131 == _T_34[9:0]) begin
        image_2_305 <= io_pixelVal_in_2_6;
      end else if (10'h131 == _T_31[9:0]) begin
        image_2_305 <= io_pixelVal_in_2_5;
      end else if (10'h131 == _T_28[9:0]) begin
        image_2_305 <= io_pixelVal_in_2_4;
      end else if (10'h131 == _T_25[9:0]) begin
        image_2_305 <= io_pixelVal_in_2_3;
      end else if (10'h131 == _T_22[9:0]) begin
        image_2_305 <= io_pixelVal_in_2_2;
      end else if (10'h131 == _T_19[9:0]) begin
        image_2_305 <= io_pixelVal_in_2_1;
      end else if (10'h131 == _T_15[9:0]) begin
        image_2_305 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_306 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h132 == _T_37[9:0]) begin
        image_2_306 <= io_pixelVal_in_2_7;
      end else if (10'h132 == _T_34[9:0]) begin
        image_2_306 <= io_pixelVal_in_2_6;
      end else if (10'h132 == _T_31[9:0]) begin
        image_2_306 <= io_pixelVal_in_2_5;
      end else if (10'h132 == _T_28[9:0]) begin
        image_2_306 <= io_pixelVal_in_2_4;
      end else if (10'h132 == _T_25[9:0]) begin
        image_2_306 <= io_pixelVal_in_2_3;
      end else if (10'h132 == _T_22[9:0]) begin
        image_2_306 <= io_pixelVal_in_2_2;
      end else if (10'h132 == _T_19[9:0]) begin
        image_2_306 <= io_pixelVal_in_2_1;
      end else if (10'h132 == _T_15[9:0]) begin
        image_2_306 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_307 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h133 == _T_37[9:0]) begin
        image_2_307 <= io_pixelVal_in_2_7;
      end else if (10'h133 == _T_34[9:0]) begin
        image_2_307 <= io_pixelVal_in_2_6;
      end else if (10'h133 == _T_31[9:0]) begin
        image_2_307 <= io_pixelVal_in_2_5;
      end else if (10'h133 == _T_28[9:0]) begin
        image_2_307 <= io_pixelVal_in_2_4;
      end else if (10'h133 == _T_25[9:0]) begin
        image_2_307 <= io_pixelVal_in_2_3;
      end else if (10'h133 == _T_22[9:0]) begin
        image_2_307 <= io_pixelVal_in_2_2;
      end else if (10'h133 == _T_19[9:0]) begin
        image_2_307 <= io_pixelVal_in_2_1;
      end else if (10'h133 == _T_15[9:0]) begin
        image_2_307 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_308 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h134 == _T_37[9:0]) begin
        image_2_308 <= io_pixelVal_in_2_7;
      end else if (10'h134 == _T_34[9:0]) begin
        image_2_308 <= io_pixelVal_in_2_6;
      end else if (10'h134 == _T_31[9:0]) begin
        image_2_308 <= io_pixelVal_in_2_5;
      end else if (10'h134 == _T_28[9:0]) begin
        image_2_308 <= io_pixelVal_in_2_4;
      end else if (10'h134 == _T_25[9:0]) begin
        image_2_308 <= io_pixelVal_in_2_3;
      end else if (10'h134 == _T_22[9:0]) begin
        image_2_308 <= io_pixelVal_in_2_2;
      end else if (10'h134 == _T_19[9:0]) begin
        image_2_308 <= io_pixelVal_in_2_1;
      end else if (10'h134 == _T_15[9:0]) begin
        image_2_308 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_309 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h135 == _T_37[9:0]) begin
        image_2_309 <= io_pixelVal_in_2_7;
      end else if (10'h135 == _T_34[9:0]) begin
        image_2_309 <= io_pixelVal_in_2_6;
      end else if (10'h135 == _T_31[9:0]) begin
        image_2_309 <= io_pixelVal_in_2_5;
      end else if (10'h135 == _T_28[9:0]) begin
        image_2_309 <= io_pixelVal_in_2_4;
      end else if (10'h135 == _T_25[9:0]) begin
        image_2_309 <= io_pixelVal_in_2_3;
      end else if (10'h135 == _T_22[9:0]) begin
        image_2_309 <= io_pixelVal_in_2_2;
      end else if (10'h135 == _T_19[9:0]) begin
        image_2_309 <= io_pixelVal_in_2_1;
      end else if (10'h135 == _T_15[9:0]) begin
        image_2_309 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_310 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h136 == _T_37[9:0]) begin
        image_2_310 <= io_pixelVal_in_2_7;
      end else if (10'h136 == _T_34[9:0]) begin
        image_2_310 <= io_pixelVal_in_2_6;
      end else if (10'h136 == _T_31[9:0]) begin
        image_2_310 <= io_pixelVal_in_2_5;
      end else if (10'h136 == _T_28[9:0]) begin
        image_2_310 <= io_pixelVal_in_2_4;
      end else if (10'h136 == _T_25[9:0]) begin
        image_2_310 <= io_pixelVal_in_2_3;
      end else if (10'h136 == _T_22[9:0]) begin
        image_2_310 <= io_pixelVal_in_2_2;
      end else if (10'h136 == _T_19[9:0]) begin
        image_2_310 <= io_pixelVal_in_2_1;
      end else if (10'h136 == _T_15[9:0]) begin
        image_2_310 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_311 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h137 == _T_37[9:0]) begin
        image_2_311 <= io_pixelVal_in_2_7;
      end else if (10'h137 == _T_34[9:0]) begin
        image_2_311 <= io_pixelVal_in_2_6;
      end else if (10'h137 == _T_31[9:0]) begin
        image_2_311 <= io_pixelVal_in_2_5;
      end else if (10'h137 == _T_28[9:0]) begin
        image_2_311 <= io_pixelVal_in_2_4;
      end else if (10'h137 == _T_25[9:0]) begin
        image_2_311 <= io_pixelVal_in_2_3;
      end else if (10'h137 == _T_22[9:0]) begin
        image_2_311 <= io_pixelVal_in_2_2;
      end else if (10'h137 == _T_19[9:0]) begin
        image_2_311 <= io_pixelVal_in_2_1;
      end else if (10'h137 == _T_15[9:0]) begin
        image_2_311 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_312 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h138 == _T_37[9:0]) begin
        image_2_312 <= io_pixelVal_in_2_7;
      end else if (10'h138 == _T_34[9:0]) begin
        image_2_312 <= io_pixelVal_in_2_6;
      end else if (10'h138 == _T_31[9:0]) begin
        image_2_312 <= io_pixelVal_in_2_5;
      end else if (10'h138 == _T_28[9:0]) begin
        image_2_312 <= io_pixelVal_in_2_4;
      end else if (10'h138 == _T_25[9:0]) begin
        image_2_312 <= io_pixelVal_in_2_3;
      end else if (10'h138 == _T_22[9:0]) begin
        image_2_312 <= io_pixelVal_in_2_2;
      end else if (10'h138 == _T_19[9:0]) begin
        image_2_312 <= io_pixelVal_in_2_1;
      end else if (10'h138 == _T_15[9:0]) begin
        image_2_312 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_313 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h139 == _T_37[9:0]) begin
        image_2_313 <= io_pixelVal_in_2_7;
      end else if (10'h139 == _T_34[9:0]) begin
        image_2_313 <= io_pixelVal_in_2_6;
      end else if (10'h139 == _T_31[9:0]) begin
        image_2_313 <= io_pixelVal_in_2_5;
      end else if (10'h139 == _T_28[9:0]) begin
        image_2_313 <= io_pixelVal_in_2_4;
      end else if (10'h139 == _T_25[9:0]) begin
        image_2_313 <= io_pixelVal_in_2_3;
      end else if (10'h139 == _T_22[9:0]) begin
        image_2_313 <= io_pixelVal_in_2_2;
      end else if (10'h139 == _T_19[9:0]) begin
        image_2_313 <= io_pixelVal_in_2_1;
      end else if (10'h139 == _T_15[9:0]) begin
        image_2_313 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_314 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13a == _T_37[9:0]) begin
        image_2_314 <= io_pixelVal_in_2_7;
      end else if (10'h13a == _T_34[9:0]) begin
        image_2_314 <= io_pixelVal_in_2_6;
      end else if (10'h13a == _T_31[9:0]) begin
        image_2_314 <= io_pixelVal_in_2_5;
      end else if (10'h13a == _T_28[9:0]) begin
        image_2_314 <= io_pixelVal_in_2_4;
      end else if (10'h13a == _T_25[9:0]) begin
        image_2_314 <= io_pixelVal_in_2_3;
      end else if (10'h13a == _T_22[9:0]) begin
        image_2_314 <= io_pixelVal_in_2_2;
      end else if (10'h13a == _T_19[9:0]) begin
        image_2_314 <= io_pixelVal_in_2_1;
      end else if (10'h13a == _T_15[9:0]) begin
        image_2_314 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_315 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13b == _T_37[9:0]) begin
        image_2_315 <= io_pixelVal_in_2_7;
      end else if (10'h13b == _T_34[9:0]) begin
        image_2_315 <= io_pixelVal_in_2_6;
      end else if (10'h13b == _T_31[9:0]) begin
        image_2_315 <= io_pixelVal_in_2_5;
      end else if (10'h13b == _T_28[9:0]) begin
        image_2_315 <= io_pixelVal_in_2_4;
      end else if (10'h13b == _T_25[9:0]) begin
        image_2_315 <= io_pixelVal_in_2_3;
      end else if (10'h13b == _T_22[9:0]) begin
        image_2_315 <= io_pixelVal_in_2_2;
      end else if (10'h13b == _T_19[9:0]) begin
        image_2_315 <= io_pixelVal_in_2_1;
      end else if (10'h13b == _T_15[9:0]) begin
        image_2_315 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_316 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13c == _T_37[9:0]) begin
        image_2_316 <= io_pixelVal_in_2_7;
      end else if (10'h13c == _T_34[9:0]) begin
        image_2_316 <= io_pixelVal_in_2_6;
      end else if (10'h13c == _T_31[9:0]) begin
        image_2_316 <= io_pixelVal_in_2_5;
      end else if (10'h13c == _T_28[9:0]) begin
        image_2_316 <= io_pixelVal_in_2_4;
      end else if (10'h13c == _T_25[9:0]) begin
        image_2_316 <= io_pixelVal_in_2_3;
      end else if (10'h13c == _T_22[9:0]) begin
        image_2_316 <= io_pixelVal_in_2_2;
      end else if (10'h13c == _T_19[9:0]) begin
        image_2_316 <= io_pixelVal_in_2_1;
      end else if (10'h13c == _T_15[9:0]) begin
        image_2_316 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_317 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13d == _T_37[9:0]) begin
        image_2_317 <= io_pixelVal_in_2_7;
      end else if (10'h13d == _T_34[9:0]) begin
        image_2_317 <= io_pixelVal_in_2_6;
      end else if (10'h13d == _T_31[9:0]) begin
        image_2_317 <= io_pixelVal_in_2_5;
      end else if (10'h13d == _T_28[9:0]) begin
        image_2_317 <= io_pixelVal_in_2_4;
      end else if (10'h13d == _T_25[9:0]) begin
        image_2_317 <= io_pixelVal_in_2_3;
      end else if (10'h13d == _T_22[9:0]) begin
        image_2_317 <= io_pixelVal_in_2_2;
      end else if (10'h13d == _T_19[9:0]) begin
        image_2_317 <= io_pixelVal_in_2_1;
      end else if (10'h13d == _T_15[9:0]) begin
        image_2_317 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_318 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13e == _T_37[9:0]) begin
        image_2_318 <= io_pixelVal_in_2_7;
      end else if (10'h13e == _T_34[9:0]) begin
        image_2_318 <= io_pixelVal_in_2_6;
      end else if (10'h13e == _T_31[9:0]) begin
        image_2_318 <= io_pixelVal_in_2_5;
      end else if (10'h13e == _T_28[9:0]) begin
        image_2_318 <= io_pixelVal_in_2_4;
      end else if (10'h13e == _T_25[9:0]) begin
        image_2_318 <= io_pixelVal_in_2_3;
      end else if (10'h13e == _T_22[9:0]) begin
        image_2_318 <= io_pixelVal_in_2_2;
      end else if (10'h13e == _T_19[9:0]) begin
        image_2_318 <= io_pixelVal_in_2_1;
      end else if (10'h13e == _T_15[9:0]) begin
        image_2_318 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_319 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13f == _T_37[9:0]) begin
        image_2_319 <= io_pixelVal_in_2_7;
      end else if (10'h13f == _T_34[9:0]) begin
        image_2_319 <= io_pixelVal_in_2_6;
      end else if (10'h13f == _T_31[9:0]) begin
        image_2_319 <= io_pixelVal_in_2_5;
      end else if (10'h13f == _T_28[9:0]) begin
        image_2_319 <= io_pixelVal_in_2_4;
      end else if (10'h13f == _T_25[9:0]) begin
        image_2_319 <= io_pixelVal_in_2_3;
      end else if (10'h13f == _T_22[9:0]) begin
        image_2_319 <= io_pixelVal_in_2_2;
      end else if (10'h13f == _T_19[9:0]) begin
        image_2_319 <= io_pixelVal_in_2_1;
      end else if (10'h13f == _T_15[9:0]) begin
        image_2_319 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_320 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h140 == _T_37[9:0]) begin
        image_2_320 <= io_pixelVal_in_2_7;
      end else if (10'h140 == _T_34[9:0]) begin
        image_2_320 <= io_pixelVal_in_2_6;
      end else if (10'h140 == _T_31[9:0]) begin
        image_2_320 <= io_pixelVal_in_2_5;
      end else if (10'h140 == _T_28[9:0]) begin
        image_2_320 <= io_pixelVal_in_2_4;
      end else if (10'h140 == _T_25[9:0]) begin
        image_2_320 <= io_pixelVal_in_2_3;
      end else if (10'h140 == _T_22[9:0]) begin
        image_2_320 <= io_pixelVal_in_2_2;
      end else if (10'h140 == _T_19[9:0]) begin
        image_2_320 <= io_pixelVal_in_2_1;
      end else if (10'h140 == _T_15[9:0]) begin
        image_2_320 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_321 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h141 == _T_37[9:0]) begin
        image_2_321 <= io_pixelVal_in_2_7;
      end else if (10'h141 == _T_34[9:0]) begin
        image_2_321 <= io_pixelVal_in_2_6;
      end else if (10'h141 == _T_31[9:0]) begin
        image_2_321 <= io_pixelVal_in_2_5;
      end else if (10'h141 == _T_28[9:0]) begin
        image_2_321 <= io_pixelVal_in_2_4;
      end else if (10'h141 == _T_25[9:0]) begin
        image_2_321 <= io_pixelVal_in_2_3;
      end else if (10'h141 == _T_22[9:0]) begin
        image_2_321 <= io_pixelVal_in_2_2;
      end else if (10'h141 == _T_19[9:0]) begin
        image_2_321 <= io_pixelVal_in_2_1;
      end else if (10'h141 == _T_15[9:0]) begin
        image_2_321 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_322 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h142 == _T_37[9:0]) begin
        image_2_322 <= io_pixelVal_in_2_7;
      end else if (10'h142 == _T_34[9:0]) begin
        image_2_322 <= io_pixelVal_in_2_6;
      end else if (10'h142 == _T_31[9:0]) begin
        image_2_322 <= io_pixelVal_in_2_5;
      end else if (10'h142 == _T_28[9:0]) begin
        image_2_322 <= io_pixelVal_in_2_4;
      end else if (10'h142 == _T_25[9:0]) begin
        image_2_322 <= io_pixelVal_in_2_3;
      end else if (10'h142 == _T_22[9:0]) begin
        image_2_322 <= io_pixelVal_in_2_2;
      end else if (10'h142 == _T_19[9:0]) begin
        image_2_322 <= io_pixelVal_in_2_1;
      end else if (10'h142 == _T_15[9:0]) begin
        image_2_322 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_323 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h143 == _T_37[9:0]) begin
        image_2_323 <= io_pixelVal_in_2_7;
      end else if (10'h143 == _T_34[9:0]) begin
        image_2_323 <= io_pixelVal_in_2_6;
      end else if (10'h143 == _T_31[9:0]) begin
        image_2_323 <= io_pixelVal_in_2_5;
      end else if (10'h143 == _T_28[9:0]) begin
        image_2_323 <= io_pixelVal_in_2_4;
      end else if (10'h143 == _T_25[9:0]) begin
        image_2_323 <= io_pixelVal_in_2_3;
      end else if (10'h143 == _T_22[9:0]) begin
        image_2_323 <= io_pixelVal_in_2_2;
      end else if (10'h143 == _T_19[9:0]) begin
        image_2_323 <= io_pixelVal_in_2_1;
      end else if (10'h143 == _T_15[9:0]) begin
        image_2_323 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_324 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h144 == _T_37[9:0]) begin
        image_2_324 <= io_pixelVal_in_2_7;
      end else if (10'h144 == _T_34[9:0]) begin
        image_2_324 <= io_pixelVal_in_2_6;
      end else if (10'h144 == _T_31[9:0]) begin
        image_2_324 <= io_pixelVal_in_2_5;
      end else if (10'h144 == _T_28[9:0]) begin
        image_2_324 <= io_pixelVal_in_2_4;
      end else if (10'h144 == _T_25[9:0]) begin
        image_2_324 <= io_pixelVal_in_2_3;
      end else if (10'h144 == _T_22[9:0]) begin
        image_2_324 <= io_pixelVal_in_2_2;
      end else if (10'h144 == _T_19[9:0]) begin
        image_2_324 <= io_pixelVal_in_2_1;
      end else if (10'h144 == _T_15[9:0]) begin
        image_2_324 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_325 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h145 == _T_37[9:0]) begin
        image_2_325 <= io_pixelVal_in_2_7;
      end else if (10'h145 == _T_34[9:0]) begin
        image_2_325 <= io_pixelVal_in_2_6;
      end else if (10'h145 == _T_31[9:0]) begin
        image_2_325 <= io_pixelVal_in_2_5;
      end else if (10'h145 == _T_28[9:0]) begin
        image_2_325 <= io_pixelVal_in_2_4;
      end else if (10'h145 == _T_25[9:0]) begin
        image_2_325 <= io_pixelVal_in_2_3;
      end else if (10'h145 == _T_22[9:0]) begin
        image_2_325 <= io_pixelVal_in_2_2;
      end else if (10'h145 == _T_19[9:0]) begin
        image_2_325 <= io_pixelVal_in_2_1;
      end else if (10'h145 == _T_15[9:0]) begin
        image_2_325 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_326 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h146 == _T_37[9:0]) begin
        image_2_326 <= io_pixelVal_in_2_7;
      end else if (10'h146 == _T_34[9:0]) begin
        image_2_326 <= io_pixelVal_in_2_6;
      end else if (10'h146 == _T_31[9:0]) begin
        image_2_326 <= io_pixelVal_in_2_5;
      end else if (10'h146 == _T_28[9:0]) begin
        image_2_326 <= io_pixelVal_in_2_4;
      end else if (10'h146 == _T_25[9:0]) begin
        image_2_326 <= io_pixelVal_in_2_3;
      end else if (10'h146 == _T_22[9:0]) begin
        image_2_326 <= io_pixelVal_in_2_2;
      end else if (10'h146 == _T_19[9:0]) begin
        image_2_326 <= io_pixelVal_in_2_1;
      end else if (10'h146 == _T_15[9:0]) begin
        image_2_326 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_327 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h147 == _T_37[9:0]) begin
        image_2_327 <= io_pixelVal_in_2_7;
      end else if (10'h147 == _T_34[9:0]) begin
        image_2_327 <= io_pixelVal_in_2_6;
      end else if (10'h147 == _T_31[9:0]) begin
        image_2_327 <= io_pixelVal_in_2_5;
      end else if (10'h147 == _T_28[9:0]) begin
        image_2_327 <= io_pixelVal_in_2_4;
      end else if (10'h147 == _T_25[9:0]) begin
        image_2_327 <= io_pixelVal_in_2_3;
      end else if (10'h147 == _T_22[9:0]) begin
        image_2_327 <= io_pixelVal_in_2_2;
      end else if (10'h147 == _T_19[9:0]) begin
        image_2_327 <= io_pixelVal_in_2_1;
      end else if (10'h147 == _T_15[9:0]) begin
        image_2_327 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_328 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h148 == _T_37[9:0]) begin
        image_2_328 <= io_pixelVal_in_2_7;
      end else if (10'h148 == _T_34[9:0]) begin
        image_2_328 <= io_pixelVal_in_2_6;
      end else if (10'h148 == _T_31[9:0]) begin
        image_2_328 <= io_pixelVal_in_2_5;
      end else if (10'h148 == _T_28[9:0]) begin
        image_2_328 <= io_pixelVal_in_2_4;
      end else if (10'h148 == _T_25[9:0]) begin
        image_2_328 <= io_pixelVal_in_2_3;
      end else if (10'h148 == _T_22[9:0]) begin
        image_2_328 <= io_pixelVal_in_2_2;
      end else if (10'h148 == _T_19[9:0]) begin
        image_2_328 <= io_pixelVal_in_2_1;
      end else if (10'h148 == _T_15[9:0]) begin
        image_2_328 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_329 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h149 == _T_37[9:0]) begin
        image_2_329 <= io_pixelVal_in_2_7;
      end else if (10'h149 == _T_34[9:0]) begin
        image_2_329 <= io_pixelVal_in_2_6;
      end else if (10'h149 == _T_31[9:0]) begin
        image_2_329 <= io_pixelVal_in_2_5;
      end else if (10'h149 == _T_28[9:0]) begin
        image_2_329 <= io_pixelVal_in_2_4;
      end else if (10'h149 == _T_25[9:0]) begin
        image_2_329 <= io_pixelVal_in_2_3;
      end else if (10'h149 == _T_22[9:0]) begin
        image_2_329 <= io_pixelVal_in_2_2;
      end else if (10'h149 == _T_19[9:0]) begin
        image_2_329 <= io_pixelVal_in_2_1;
      end else if (10'h149 == _T_15[9:0]) begin
        image_2_329 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_330 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14a == _T_37[9:0]) begin
        image_2_330 <= io_pixelVal_in_2_7;
      end else if (10'h14a == _T_34[9:0]) begin
        image_2_330 <= io_pixelVal_in_2_6;
      end else if (10'h14a == _T_31[9:0]) begin
        image_2_330 <= io_pixelVal_in_2_5;
      end else if (10'h14a == _T_28[9:0]) begin
        image_2_330 <= io_pixelVal_in_2_4;
      end else if (10'h14a == _T_25[9:0]) begin
        image_2_330 <= io_pixelVal_in_2_3;
      end else if (10'h14a == _T_22[9:0]) begin
        image_2_330 <= io_pixelVal_in_2_2;
      end else if (10'h14a == _T_19[9:0]) begin
        image_2_330 <= io_pixelVal_in_2_1;
      end else if (10'h14a == _T_15[9:0]) begin
        image_2_330 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_331 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14b == _T_37[9:0]) begin
        image_2_331 <= io_pixelVal_in_2_7;
      end else if (10'h14b == _T_34[9:0]) begin
        image_2_331 <= io_pixelVal_in_2_6;
      end else if (10'h14b == _T_31[9:0]) begin
        image_2_331 <= io_pixelVal_in_2_5;
      end else if (10'h14b == _T_28[9:0]) begin
        image_2_331 <= io_pixelVal_in_2_4;
      end else if (10'h14b == _T_25[9:0]) begin
        image_2_331 <= io_pixelVal_in_2_3;
      end else if (10'h14b == _T_22[9:0]) begin
        image_2_331 <= io_pixelVal_in_2_2;
      end else if (10'h14b == _T_19[9:0]) begin
        image_2_331 <= io_pixelVal_in_2_1;
      end else if (10'h14b == _T_15[9:0]) begin
        image_2_331 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_332 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14c == _T_37[9:0]) begin
        image_2_332 <= io_pixelVal_in_2_7;
      end else if (10'h14c == _T_34[9:0]) begin
        image_2_332 <= io_pixelVal_in_2_6;
      end else if (10'h14c == _T_31[9:0]) begin
        image_2_332 <= io_pixelVal_in_2_5;
      end else if (10'h14c == _T_28[9:0]) begin
        image_2_332 <= io_pixelVal_in_2_4;
      end else if (10'h14c == _T_25[9:0]) begin
        image_2_332 <= io_pixelVal_in_2_3;
      end else if (10'h14c == _T_22[9:0]) begin
        image_2_332 <= io_pixelVal_in_2_2;
      end else if (10'h14c == _T_19[9:0]) begin
        image_2_332 <= io_pixelVal_in_2_1;
      end else if (10'h14c == _T_15[9:0]) begin
        image_2_332 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_333 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14d == _T_37[9:0]) begin
        image_2_333 <= io_pixelVal_in_2_7;
      end else if (10'h14d == _T_34[9:0]) begin
        image_2_333 <= io_pixelVal_in_2_6;
      end else if (10'h14d == _T_31[9:0]) begin
        image_2_333 <= io_pixelVal_in_2_5;
      end else if (10'h14d == _T_28[9:0]) begin
        image_2_333 <= io_pixelVal_in_2_4;
      end else if (10'h14d == _T_25[9:0]) begin
        image_2_333 <= io_pixelVal_in_2_3;
      end else if (10'h14d == _T_22[9:0]) begin
        image_2_333 <= io_pixelVal_in_2_2;
      end else if (10'h14d == _T_19[9:0]) begin
        image_2_333 <= io_pixelVal_in_2_1;
      end else if (10'h14d == _T_15[9:0]) begin
        image_2_333 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_334 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14e == _T_37[9:0]) begin
        image_2_334 <= io_pixelVal_in_2_7;
      end else if (10'h14e == _T_34[9:0]) begin
        image_2_334 <= io_pixelVal_in_2_6;
      end else if (10'h14e == _T_31[9:0]) begin
        image_2_334 <= io_pixelVal_in_2_5;
      end else if (10'h14e == _T_28[9:0]) begin
        image_2_334 <= io_pixelVal_in_2_4;
      end else if (10'h14e == _T_25[9:0]) begin
        image_2_334 <= io_pixelVal_in_2_3;
      end else if (10'h14e == _T_22[9:0]) begin
        image_2_334 <= io_pixelVal_in_2_2;
      end else if (10'h14e == _T_19[9:0]) begin
        image_2_334 <= io_pixelVal_in_2_1;
      end else if (10'h14e == _T_15[9:0]) begin
        image_2_334 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_335 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14f == _T_37[9:0]) begin
        image_2_335 <= io_pixelVal_in_2_7;
      end else if (10'h14f == _T_34[9:0]) begin
        image_2_335 <= io_pixelVal_in_2_6;
      end else if (10'h14f == _T_31[9:0]) begin
        image_2_335 <= io_pixelVal_in_2_5;
      end else if (10'h14f == _T_28[9:0]) begin
        image_2_335 <= io_pixelVal_in_2_4;
      end else if (10'h14f == _T_25[9:0]) begin
        image_2_335 <= io_pixelVal_in_2_3;
      end else if (10'h14f == _T_22[9:0]) begin
        image_2_335 <= io_pixelVal_in_2_2;
      end else if (10'h14f == _T_19[9:0]) begin
        image_2_335 <= io_pixelVal_in_2_1;
      end else if (10'h14f == _T_15[9:0]) begin
        image_2_335 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_336 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h150 == _T_37[9:0]) begin
        image_2_336 <= io_pixelVal_in_2_7;
      end else if (10'h150 == _T_34[9:0]) begin
        image_2_336 <= io_pixelVal_in_2_6;
      end else if (10'h150 == _T_31[9:0]) begin
        image_2_336 <= io_pixelVal_in_2_5;
      end else if (10'h150 == _T_28[9:0]) begin
        image_2_336 <= io_pixelVal_in_2_4;
      end else if (10'h150 == _T_25[9:0]) begin
        image_2_336 <= io_pixelVal_in_2_3;
      end else if (10'h150 == _T_22[9:0]) begin
        image_2_336 <= io_pixelVal_in_2_2;
      end else if (10'h150 == _T_19[9:0]) begin
        image_2_336 <= io_pixelVal_in_2_1;
      end else if (10'h150 == _T_15[9:0]) begin
        image_2_336 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_337 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h151 == _T_37[9:0]) begin
        image_2_337 <= io_pixelVal_in_2_7;
      end else if (10'h151 == _T_34[9:0]) begin
        image_2_337 <= io_pixelVal_in_2_6;
      end else if (10'h151 == _T_31[9:0]) begin
        image_2_337 <= io_pixelVal_in_2_5;
      end else if (10'h151 == _T_28[9:0]) begin
        image_2_337 <= io_pixelVal_in_2_4;
      end else if (10'h151 == _T_25[9:0]) begin
        image_2_337 <= io_pixelVal_in_2_3;
      end else if (10'h151 == _T_22[9:0]) begin
        image_2_337 <= io_pixelVal_in_2_2;
      end else if (10'h151 == _T_19[9:0]) begin
        image_2_337 <= io_pixelVal_in_2_1;
      end else if (10'h151 == _T_15[9:0]) begin
        image_2_337 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_338 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h152 == _T_37[9:0]) begin
        image_2_338 <= io_pixelVal_in_2_7;
      end else if (10'h152 == _T_34[9:0]) begin
        image_2_338 <= io_pixelVal_in_2_6;
      end else if (10'h152 == _T_31[9:0]) begin
        image_2_338 <= io_pixelVal_in_2_5;
      end else if (10'h152 == _T_28[9:0]) begin
        image_2_338 <= io_pixelVal_in_2_4;
      end else if (10'h152 == _T_25[9:0]) begin
        image_2_338 <= io_pixelVal_in_2_3;
      end else if (10'h152 == _T_22[9:0]) begin
        image_2_338 <= io_pixelVal_in_2_2;
      end else if (10'h152 == _T_19[9:0]) begin
        image_2_338 <= io_pixelVal_in_2_1;
      end else if (10'h152 == _T_15[9:0]) begin
        image_2_338 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_339 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h153 == _T_37[9:0]) begin
        image_2_339 <= io_pixelVal_in_2_7;
      end else if (10'h153 == _T_34[9:0]) begin
        image_2_339 <= io_pixelVal_in_2_6;
      end else if (10'h153 == _T_31[9:0]) begin
        image_2_339 <= io_pixelVal_in_2_5;
      end else if (10'h153 == _T_28[9:0]) begin
        image_2_339 <= io_pixelVal_in_2_4;
      end else if (10'h153 == _T_25[9:0]) begin
        image_2_339 <= io_pixelVal_in_2_3;
      end else if (10'h153 == _T_22[9:0]) begin
        image_2_339 <= io_pixelVal_in_2_2;
      end else if (10'h153 == _T_19[9:0]) begin
        image_2_339 <= io_pixelVal_in_2_1;
      end else if (10'h153 == _T_15[9:0]) begin
        image_2_339 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_340 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h154 == _T_37[9:0]) begin
        image_2_340 <= io_pixelVal_in_2_7;
      end else if (10'h154 == _T_34[9:0]) begin
        image_2_340 <= io_pixelVal_in_2_6;
      end else if (10'h154 == _T_31[9:0]) begin
        image_2_340 <= io_pixelVal_in_2_5;
      end else if (10'h154 == _T_28[9:0]) begin
        image_2_340 <= io_pixelVal_in_2_4;
      end else if (10'h154 == _T_25[9:0]) begin
        image_2_340 <= io_pixelVal_in_2_3;
      end else if (10'h154 == _T_22[9:0]) begin
        image_2_340 <= io_pixelVal_in_2_2;
      end else if (10'h154 == _T_19[9:0]) begin
        image_2_340 <= io_pixelVal_in_2_1;
      end else if (10'h154 == _T_15[9:0]) begin
        image_2_340 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_341 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h155 == _T_37[9:0]) begin
        image_2_341 <= io_pixelVal_in_2_7;
      end else if (10'h155 == _T_34[9:0]) begin
        image_2_341 <= io_pixelVal_in_2_6;
      end else if (10'h155 == _T_31[9:0]) begin
        image_2_341 <= io_pixelVal_in_2_5;
      end else if (10'h155 == _T_28[9:0]) begin
        image_2_341 <= io_pixelVal_in_2_4;
      end else if (10'h155 == _T_25[9:0]) begin
        image_2_341 <= io_pixelVal_in_2_3;
      end else if (10'h155 == _T_22[9:0]) begin
        image_2_341 <= io_pixelVal_in_2_2;
      end else if (10'h155 == _T_19[9:0]) begin
        image_2_341 <= io_pixelVal_in_2_1;
      end else if (10'h155 == _T_15[9:0]) begin
        image_2_341 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_342 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h156 == _T_37[9:0]) begin
        image_2_342 <= io_pixelVal_in_2_7;
      end else if (10'h156 == _T_34[9:0]) begin
        image_2_342 <= io_pixelVal_in_2_6;
      end else if (10'h156 == _T_31[9:0]) begin
        image_2_342 <= io_pixelVal_in_2_5;
      end else if (10'h156 == _T_28[9:0]) begin
        image_2_342 <= io_pixelVal_in_2_4;
      end else if (10'h156 == _T_25[9:0]) begin
        image_2_342 <= io_pixelVal_in_2_3;
      end else if (10'h156 == _T_22[9:0]) begin
        image_2_342 <= io_pixelVal_in_2_2;
      end else if (10'h156 == _T_19[9:0]) begin
        image_2_342 <= io_pixelVal_in_2_1;
      end else if (10'h156 == _T_15[9:0]) begin
        image_2_342 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_343 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h157 == _T_37[9:0]) begin
        image_2_343 <= io_pixelVal_in_2_7;
      end else if (10'h157 == _T_34[9:0]) begin
        image_2_343 <= io_pixelVal_in_2_6;
      end else if (10'h157 == _T_31[9:0]) begin
        image_2_343 <= io_pixelVal_in_2_5;
      end else if (10'h157 == _T_28[9:0]) begin
        image_2_343 <= io_pixelVal_in_2_4;
      end else if (10'h157 == _T_25[9:0]) begin
        image_2_343 <= io_pixelVal_in_2_3;
      end else if (10'h157 == _T_22[9:0]) begin
        image_2_343 <= io_pixelVal_in_2_2;
      end else if (10'h157 == _T_19[9:0]) begin
        image_2_343 <= io_pixelVal_in_2_1;
      end else if (10'h157 == _T_15[9:0]) begin
        image_2_343 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_344 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h158 == _T_37[9:0]) begin
        image_2_344 <= io_pixelVal_in_2_7;
      end else if (10'h158 == _T_34[9:0]) begin
        image_2_344 <= io_pixelVal_in_2_6;
      end else if (10'h158 == _T_31[9:0]) begin
        image_2_344 <= io_pixelVal_in_2_5;
      end else if (10'h158 == _T_28[9:0]) begin
        image_2_344 <= io_pixelVal_in_2_4;
      end else if (10'h158 == _T_25[9:0]) begin
        image_2_344 <= io_pixelVal_in_2_3;
      end else if (10'h158 == _T_22[9:0]) begin
        image_2_344 <= io_pixelVal_in_2_2;
      end else if (10'h158 == _T_19[9:0]) begin
        image_2_344 <= io_pixelVal_in_2_1;
      end else if (10'h158 == _T_15[9:0]) begin
        image_2_344 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_345 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h159 == _T_37[9:0]) begin
        image_2_345 <= io_pixelVal_in_2_7;
      end else if (10'h159 == _T_34[9:0]) begin
        image_2_345 <= io_pixelVal_in_2_6;
      end else if (10'h159 == _T_31[9:0]) begin
        image_2_345 <= io_pixelVal_in_2_5;
      end else if (10'h159 == _T_28[9:0]) begin
        image_2_345 <= io_pixelVal_in_2_4;
      end else if (10'h159 == _T_25[9:0]) begin
        image_2_345 <= io_pixelVal_in_2_3;
      end else if (10'h159 == _T_22[9:0]) begin
        image_2_345 <= io_pixelVal_in_2_2;
      end else if (10'h159 == _T_19[9:0]) begin
        image_2_345 <= io_pixelVal_in_2_1;
      end else if (10'h159 == _T_15[9:0]) begin
        image_2_345 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_346 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15a == _T_37[9:0]) begin
        image_2_346 <= io_pixelVal_in_2_7;
      end else if (10'h15a == _T_34[9:0]) begin
        image_2_346 <= io_pixelVal_in_2_6;
      end else if (10'h15a == _T_31[9:0]) begin
        image_2_346 <= io_pixelVal_in_2_5;
      end else if (10'h15a == _T_28[9:0]) begin
        image_2_346 <= io_pixelVal_in_2_4;
      end else if (10'h15a == _T_25[9:0]) begin
        image_2_346 <= io_pixelVal_in_2_3;
      end else if (10'h15a == _T_22[9:0]) begin
        image_2_346 <= io_pixelVal_in_2_2;
      end else if (10'h15a == _T_19[9:0]) begin
        image_2_346 <= io_pixelVal_in_2_1;
      end else if (10'h15a == _T_15[9:0]) begin
        image_2_346 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_347 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15b == _T_37[9:0]) begin
        image_2_347 <= io_pixelVal_in_2_7;
      end else if (10'h15b == _T_34[9:0]) begin
        image_2_347 <= io_pixelVal_in_2_6;
      end else if (10'h15b == _T_31[9:0]) begin
        image_2_347 <= io_pixelVal_in_2_5;
      end else if (10'h15b == _T_28[9:0]) begin
        image_2_347 <= io_pixelVal_in_2_4;
      end else if (10'h15b == _T_25[9:0]) begin
        image_2_347 <= io_pixelVal_in_2_3;
      end else if (10'h15b == _T_22[9:0]) begin
        image_2_347 <= io_pixelVal_in_2_2;
      end else if (10'h15b == _T_19[9:0]) begin
        image_2_347 <= io_pixelVal_in_2_1;
      end else if (10'h15b == _T_15[9:0]) begin
        image_2_347 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_348 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15c == _T_37[9:0]) begin
        image_2_348 <= io_pixelVal_in_2_7;
      end else if (10'h15c == _T_34[9:0]) begin
        image_2_348 <= io_pixelVal_in_2_6;
      end else if (10'h15c == _T_31[9:0]) begin
        image_2_348 <= io_pixelVal_in_2_5;
      end else if (10'h15c == _T_28[9:0]) begin
        image_2_348 <= io_pixelVal_in_2_4;
      end else if (10'h15c == _T_25[9:0]) begin
        image_2_348 <= io_pixelVal_in_2_3;
      end else if (10'h15c == _T_22[9:0]) begin
        image_2_348 <= io_pixelVal_in_2_2;
      end else if (10'h15c == _T_19[9:0]) begin
        image_2_348 <= io_pixelVal_in_2_1;
      end else if (10'h15c == _T_15[9:0]) begin
        image_2_348 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_349 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15d == _T_37[9:0]) begin
        image_2_349 <= io_pixelVal_in_2_7;
      end else if (10'h15d == _T_34[9:0]) begin
        image_2_349 <= io_pixelVal_in_2_6;
      end else if (10'h15d == _T_31[9:0]) begin
        image_2_349 <= io_pixelVal_in_2_5;
      end else if (10'h15d == _T_28[9:0]) begin
        image_2_349 <= io_pixelVal_in_2_4;
      end else if (10'h15d == _T_25[9:0]) begin
        image_2_349 <= io_pixelVal_in_2_3;
      end else if (10'h15d == _T_22[9:0]) begin
        image_2_349 <= io_pixelVal_in_2_2;
      end else if (10'h15d == _T_19[9:0]) begin
        image_2_349 <= io_pixelVal_in_2_1;
      end else if (10'h15d == _T_15[9:0]) begin
        image_2_349 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_350 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15e == _T_37[9:0]) begin
        image_2_350 <= io_pixelVal_in_2_7;
      end else if (10'h15e == _T_34[9:0]) begin
        image_2_350 <= io_pixelVal_in_2_6;
      end else if (10'h15e == _T_31[9:0]) begin
        image_2_350 <= io_pixelVal_in_2_5;
      end else if (10'h15e == _T_28[9:0]) begin
        image_2_350 <= io_pixelVal_in_2_4;
      end else if (10'h15e == _T_25[9:0]) begin
        image_2_350 <= io_pixelVal_in_2_3;
      end else if (10'h15e == _T_22[9:0]) begin
        image_2_350 <= io_pixelVal_in_2_2;
      end else if (10'h15e == _T_19[9:0]) begin
        image_2_350 <= io_pixelVal_in_2_1;
      end else if (10'h15e == _T_15[9:0]) begin
        image_2_350 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_351 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15f == _T_37[9:0]) begin
        image_2_351 <= io_pixelVal_in_2_7;
      end else if (10'h15f == _T_34[9:0]) begin
        image_2_351 <= io_pixelVal_in_2_6;
      end else if (10'h15f == _T_31[9:0]) begin
        image_2_351 <= io_pixelVal_in_2_5;
      end else if (10'h15f == _T_28[9:0]) begin
        image_2_351 <= io_pixelVal_in_2_4;
      end else if (10'h15f == _T_25[9:0]) begin
        image_2_351 <= io_pixelVal_in_2_3;
      end else if (10'h15f == _T_22[9:0]) begin
        image_2_351 <= io_pixelVal_in_2_2;
      end else if (10'h15f == _T_19[9:0]) begin
        image_2_351 <= io_pixelVal_in_2_1;
      end else if (10'h15f == _T_15[9:0]) begin
        image_2_351 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_352 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h160 == _T_37[9:0]) begin
        image_2_352 <= io_pixelVal_in_2_7;
      end else if (10'h160 == _T_34[9:0]) begin
        image_2_352 <= io_pixelVal_in_2_6;
      end else if (10'h160 == _T_31[9:0]) begin
        image_2_352 <= io_pixelVal_in_2_5;
      end else if (10'h160 == _T_28[9:0]) begin
        image_2_352 <= io_pixelVal_in_2_4;
      end else if (10'h160 == _T_25[9:0]) begin
        image_2_352 <= io_pixelVal_in_2_3;
      end else if (10'h160 == _T_22[9:0]) begin
        image_2_352 <= io_pixelVal_in_2_2;
      end else if (10'h160 == _T_19[9:0]) begin
        image_2_352 <= io_pixelVal_in_2_1;
      end else if (10'h160 == _T_15[9:0]) begin
        image_2_352 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_353 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h161 == _T_37[9:0]) begin
        image_2_353 <= io_pixelVal_in_2_7;
      end else if (10'h161 == _T_34[9:0]) begin
        image_2_353 <= io_pixelVal_in_2_6;
      end else if (10'h161 == _T_31[9:0]) begin
        image_2_353 <= io_pixelVal_in_2_5;
      end else if (10'h161 == _T_28[9:0]) begin
        image_2_353 <= io_pixelVal_in_2_4;
      end else if (10'h161 == _T_25[9:0]) begin
        image_2_353 <= io_pixelVal_in_2_3;
      end else if (10'h161 == _T_22[9:0]) begin
        image_2_353 <= io_pixelVal_in_2_2;
      end else if (10'h161 == _T_19[9:0]) begin
        image_2_353 <= io_pixelVal_in_2_1;
      end else if (10'h161 == _T_15[9:0]) begin
        image_2_353 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_354 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h162 == _T_37[9:0]) begin
        image_2_354 <= io_pixelVal_in_2_7;
      end else if (10'h162 == _T_34[9:0]) begin
        image_2_354 <= io_pixelVal_in_2_6;
      end else if (10'h162 == _T_31[9:0]) begin
        image_2_354 <= io_pixelVal_in_2_5;
      end else if (10'h162 == _T_28[9:0]) begin
        image_2_354 <= io_pixelVal_in_2_4;
      end else if (10'h162 == _T_25[9:0]) begin
        image_2_354 <= io_pixelVal_in_2_3;
      end else if (10'h162 == _T_22[9:0]) begin
        image_2_354 <= io_pixelVal_in_2_2;
      end else if (10'h162 == _T_19[9:0]) begin
        image_2_354 <= io_pixelVal_in_2_1;
      end else if (10'h162 == _T_15[9:0]) begin
        image_2_354 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_355 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h163 == _T_37[9:0]) begin
        image_2_355 <= io_pixelVal_in_2_7;
      end else if (10'h163 == _T_34[9:0]) begin
        image_2_355 <= io_pixelVal_in_2_6;
      end else if (10'h163 == _T_31[9:0]) begin
        image_2_355 <= io_pixelVal_in_2_5;
      end else if (10'h163 == _T_28[9:0]) begin
        image_2_355 <= io_pixelVal_in_2_4;
      end else if (10'h163 == _T_25[9:0]) begin
        image_2_355 <= io_pixelVal_in_2_3;
      end else if (10'h163 == _T_22[9:0]) begin
        image_2_355 <= io_pixelVal_in_2_2;
      end else if (10'h163 == _T_19[9:0]) begin
        image_2_355 <= io_pixelVal_in_2_1;
      end else if (10'h163 == _T_15[9:0]) begin
        image_2_355 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_356 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h164 == _T_37[9:0]) begin
        image_2_356 <= io_pixelVal_in_2_7;
      end else if (10'h164 == _T_34[9:0]) begin
        image_2_356 <= io_pixelVal_in_2_6;
      end else if (10'h164 == _T_31[9:0]) begin
        image_2_356 <= io_pixelVal_in_2_5;
      end else if (10'h164 == _T_28[9:0]) begin
        image_2_356 <= io_pixelVal_in_2_4;
      end else if (10'h164 == _T_25[9:0]) begin
        image_2_356 <= io_pixelVal_in_2_3;
      end else if (10'h164 == _T_22[9:0]) begin
        image_2_356 <= io_pixelVal_in_2_2;
      end else if (10'h164 == _T_19[9:0]) begin
        image_2_356 <= io_pixelVal_in_2_1;
      end else if (10'h164 == _T_15[9:0]) begin
        image_2_356 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_357 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h165 == _T_37[9:0]) begin
        image_2_357 <= io_pixelVal_in_2_7;
      end else if (10'h165 == _T_34[9:0]) begin
        image_2_357 <= io_pixelVal_in_2_6;
      end else if (10'h165 == _T_31[9:0]) begin
        image_2_357 <= io_pixelVal_in_2_5;
      end else if (10'h165 == _T_28[9:0]) begin
        image_2_357 <= io_pixelVal_in_2_4;
      end else if (10'h165 == _T_25[9:0]) begin
        image_2_357 <= io_pixelVal_in_2_3;
      end else if (10'h165 == _T_22[9:0]) begin
        image_2_357 <= io_pixelVal_in_2_2;
      end else if (10'h165 == _T_19[9:0]) begin
        image_2_357 <= io_pixelVal_in_2_1;
      end else if (10'h165 == _T_15[9:0]) begin
        image_2_357 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_358 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h166 == _T_37[9:0]) begin
        image_2_358 <= io_pixelVal_in_2_7;
      end else if (10'h166 == _T_34[9:0]) begin
        image_2_358 <= io_pixelVal_in_2_6;
      end else if (10'h166 == _T_31[9:0]) begin
        image_2_358 <= io_pixelVal_in_2_5;
      end else if (10'h166 == _T_28[9:0]) begin
        image_2_358 <= io_pixelVal_in_2_4;
      end else if (10'h166 == _T_25[9:0]) begin
        image_2_358 <= io_pixelVal_in_2_3;
      end else if (10'h166 == _T_22[9:0]) begin
        image_2_358 <= io_pixelVal_in_2_2;
      end else if (10'h166 == _T_19[9:0]) begin
        image_2_358 <= io_pixelVal_in_2_1;
      end else if (10'h166 == _T_15[9:0]) begin
        image_2_358 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_359 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h167 == _T_37[9:0]) begin
        image_2_359 <= io_pixelVal_in_2_7;
      end else if (10'h167 == _T_34[9:0]) begin
        image_2_359 <= io_pixelVal_in_2_6;
      end else if (10'h167 == _T_31[9:0]) begin
        image_2_359 <= io_pixelVal_in_2_5;
      end else if (10'h167 == _T_28[9:0]) begin
        image_2_359 <= io_pixelVal_in_2_4;
      end else if (10'h167 == _T_25[9:0]) begin
        image_2_359 <= io_pixelVal_in_2_3;
      end else if (10'h167 == _T_22[9:0]) begin
        image_2_359 <= io_pixelVal_in_2_2;
      end else if (10'h167 == _T_19[9:0]) begin
        image_2_359 <= io_pixelVal_in_2_1;
      end else if (10'h167 == _T_15[9:0]) begin
        image_2_359 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_360 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h168 == _T_37[9:0]) begin
        image_2_360 <= io_pixelVal_in_2_7;
      end else if (10'h168 == _T_34[9:0]) begin
        image_2_360 <= io_pixelVal_in_2_6;
      end else if (10'h168 == _T_31[9:0]) begin
        image_2_360 <= io_pixelVal_in_2_5;
      end else if (10'h168 == _T_28[9:0]) begin
        image_2_360 <= io_pixelVal_in_2_4;
      end else if (10'h168 == _T_25[9:0]) begin
        image_2_360 <= io_pixelVal_in_2_3;
      end else if (10'h168 == _T_22[9:0]) begin
        image_2_360 <= io_pixelVal_in_2_2;
      end else if (10'h168 == _T_19[9:0]) begin
        image_2_360 <= io_pixelVal_in_2_1;
      end else if (10'h168 == _T_15[9:0]) begin
        image_2_360 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_361 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h169 == _T_37[9:0]) begin
        image_2_361 <= io_pixelVal_in_2_7;
      end else if (10'h169 == _T_34[9:0]) begin
        image_2_361 <= io_pixelVal_in_2_6;
      end else if (10'h169 == _T_31[9:0]) begin
        image_2_361 <= io_pixelVal_in_2_5;
      end else if (10'h169 == _T_28[9:0]) begin
        image_2_361 <= io_pixelVal_in_2_4;
      end else if (10'h169 == _T_25[9:0]) begin
        image_2_361 <= io_pixelVal_in_2_3;
      end else if (10'h169 == _T_22[9:0]) begin
        image_2_361 <= io_pixelVal_in_2_2;
      end else if (10'h169 == _T_19[9:0]) begin
        image_2_361 <= io_pixelVal_in_2_1;
      end else if (10'h169 == _T_15[9:0]) begin
        image_2_361 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_362 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16a == _T_37[9:0]) begin
        image_2_362 <= io_pixelVal_in_2_7;
      end else if (10'h16a == _T_34[9:0]) begin
        image_2_362 <= io_pixelVal_in_2_6;
      end else if (10'h16a == _T_31[9:0]) begin
        image_2_362 <= io_pixelVal_in_2_5;
      end else if (10'h16a == _T_28[9:0]) begin
        image_2_362 <= io_pixelVal_in_2_4;
      end else if (10'h16a == _T_25[9:0]) begin
        image_2_362 <= io_pixelVal_in_2_3;
      end else if (10'h16a == _T_22[9:0]) begin
        image_2_362 <= io_pixelVal_in_2_2;
      end else if (10'h16a == _T_19[9:0]) begin
        image_2_362 <= io_pixelVal_in_2_1;
      end else if (10'h16a == _T_15[9:0]) begin
        image_2_362 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_363 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16b == _T_37[9:0]) begin
        image_2_363 <= io_pixelVal_in_2_7;
      end else if (10'h16b == _T_34[9:0]) begin
        image_2_363 <= io_pixelVal_in_2_6;
      end else if (10'h16b == _T_31[9:0]) begin
        image_2_363 <= io_pixelVal_in_2_5;
      end else if (10'h16b == _T_28[9:0]) begin
        image_2_363 <= io_pixelVal_in_2_4;
      end else if (10'h16b == _T_25[9:0]) begin
        image_2_363 <= io_pixelVal_in_2_3;
      end else if (10'h16b == _T_22[9:0]) begin
        image_2_363 <= io_pixelVal_in_2_2;
      end else if (10'h16b == _T_19[9:0]) begin
        image_2_363 <= io_pixelVal_in_2_1;
      end else if (10'h16b == _T_15[9:0]) begin
        image_2_363 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_364 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16c == _T_37[9:0]) begin
        image_2_364 <= io_pixelVal_in_2_7;
      end else if (10'h16c == _T_34[9:0]) begin
        image_2_364 <= io_pixelVal_in_2_6;
      end else if (10'h16c == _T_31[9:0]) begin
        image_2_364 <= io_pixelVal_in_2_5;
      end else if (10'h16c == _T_28[9:0]) begin
        image_2_364 <= io_pixelVal_in_2_4;
      end else if (10'h16c == _T_25[9:0]) begin
        image_2_364 <= io_pixelVal_in_2_3;
      end else if (10'h16c == _T_22[9:0]) begin
        image_2_364 <= io_pixelVal_in_2_2;
      end else if (10'h16c == _T_19[9:0]) begin
        image_2_364 <= io_pixelVal_in_2_1;
      end else if (10'h16c == _T_15[9:0]) begin
        image_2_364 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_365 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16d == _T_37[9:0]) begin
        image_2_365 <= io_pixelVal_in_2_7;
      end else if (10'h16d == _T_34[9:0]) begin
        image_2_365 <= io_pixelVal_in_2_6;
      end else if (10'h16d == _T_31[9:0]) begin
        image_2_365 <= io_pixelVal_in_2_5;
      end else if (10'h16d == _T_28[9:0]) begin
        image_2_365 <= io_pixelVal_in_2_4;
      end else if (10'h16d == _T_25[9:0]) begin
        image_2_365 <= io_pixelVal_in_2_3;
      end else if (10'h16d == _T_22[9:0]) begin
        image_2_365 <= io_pixelVal_in_2_2;
      end else if (10'h16d == _T_19[9:0]) begin
        image_2_365 <= io_pixelVal_in_2_1;
      end else if (10'h16d == _T_15[9:0]) begin
        image_2_365 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_366 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16e == _T_37[9:0]) begin
        image_2_366 <= io_pixelVal_in_2_7;
      end else if (10'h16e == _T_34[9:0]) begin
        image_2_366 <= io_pixelVal_in_2_6;
      end else if (10'h16e == _T_31[9:0]) begin
        image_2_366 <= io_pixelVal_in_2_5;
      end else if (10'h16e == _T_28[9:0]) begin
        image_2_366 <= io_pixelVal_in_2_4;
      end else if (10'h16e == _T_25[9:0]) begin
        image_2_366 <= io_pixelVal_in_2_3;
      end else if (10'h16e == _T_22[9:0]) begin
        image_2_366 <= io_pixelVal_in_2_2;
      end else if (10'h16e == _T_19[9:0]) begin
        image_2_366 <= io_pixelVal_in_2_1;
      end else if (10'h16e == _T_15[9:0]) begin
        image_2_366 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_367 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16f == _T_37[9:0]) begin
        image_2_367 <= io_pixelVal_in_2_7;
      end else if (10'h16f == _T_34[9:0]) begin
        image_2_367 <= io_pixelVal_in_2_6;
      end else if (10'h16f == _T_31[9:0]) begin
        image_2_367 <= io_pixelVal_in_2_5;
      end else if (10'h16f == _T_28[9:0]) begin
        image_2_367 <= io_pixelVal_in_2_4;
      end else if (10'h16f == _T_25[9:0]) begin
        image_2_367 <= io_pixelVal_in_2_3;
      end else if (10'h16f == _T_22[9:0]) begin
        image_2_367 <= io_pixelVal_in_2_2;
      end else if (10'h16f == _T_19[9:0]) begin
        image_2_367 <= io_pixelVal_in_2_1;
      end else if (10'h16f == _T_15[9:0]) begin
        image_2_367 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_368 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h170 == _T_37[9:0]) begin
        image_2_368 <= io_pixelVal_in_2_7;
      end else if (10'h170 == _T_34[9:0]) begin
        image_2_368 <= io_pixelVal_in_2_6;
      end else if (10'h170 == _T_31[9:0]) begin
        image_2_368 <= io_pixelVal_in_2_5;
      end else if (10'h170 == _T_28[9:0]) begin
        image_2_368 <= io_pixelVal_in_2_4;
      end else if (10'h170 == _T_25[9:0]) begin
        image_2_368 <= io_pixelVal_in_2_3;
      end else if (10'h170 == _T_22[9:0]) begin
        image_2_368 <= io_pixelVal_in_2_2;
      end else if (10'h170 == _T_19[9:0]) begin
        image_2_368 <= io_pixelVal_in_2_1;
      end else if (10'h170 == _T_15[9:0]) begin
        image_2_368 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_369 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h171 == _T_37[9:0]) begin
        image_2_369 <= io_pixelVal_in_2_7;
      end else if (10'h171 == _T_34[9:0]) begin
        image_2_369 <= io_pixelVal_in_2_6;
      end else if (10'h171 == _T_31[9:0]) begin
        image_2_369 <= io_pixelVal_in_2_5;
      end else if (10'h171 == _T_28[9:0]) begin
        image_2_369 <= io_pixelVal_in_2_4;
      end else if (10'h171 == _T_25[9:0]) begin
        image_2_369 <= io_pixelVal_in_2_3;
      end else if (10'h171 == _T_22[9:0]) begin
        image_2_369 <= io_pixelVal_in_2_2;
      end else if (10'h171 == _T_19[9:0]) begin
        image_2_369 <= io_pixelVal_in_2_1;
      end else if (10'h171 == _T_15[9:0]) begin
        image_2_369 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_370 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h172 == _T_37[9:0]) begin
        image_2_370 <= io_pixelVal_in_2_7;
      end else if (10'h172 == _T_34[9:0]) begin
        image_2_370 <= io_pixelVal_in_2_6;
      end else if (10'h172 == _T_31[9:0]) begin
        image_2_370 <= io_pixelVal_in_2_5;
      end else if (10'h172 == _T_28[9:0]) begin
        image_2_370 <= io_pixelVal_in_2_4;
      end else if (10'h172 == _T_25[9:0]) begin
        image_2_370 <= io_pixelVal_in_2_3;
      end else if (10'h172 == _T_22[9:0]) begin
        image_2_370 <= io_pixelVal_in_2_2;
      end else if (10'h172 == _T_19[9:0]) begin
        image_2_370 <= io_pixelVal_in_2_1;
      end else if (10'h172 == _T_15[9:0]) begin
        image_2_370 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_371 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h173 == _T_37[9:0]) begin
        image_2_371 <= io_pixelVal_in_2_7;
      end else if (10'h173 == _T_34[9:0]) begin
        image_2_371 <= io_pixelVal_in_2_6;
      end else if (10'h173 == _T_31[9:0]) begin
        image_2_371 <= io_pixelVal_in_2_5;
      end else if (10'h173 == _T_28[9:0]) begin
        image_2_371 <= io_pixelVal_in_2_4;
      end else if (10'h173 == _T_25[9:0]) begin
        image_2_371 <= io_pixelVal_in_2_3;
      end else if (10'h173 == _T_22[9:0]) begin
        image_2_371 <= io_pixelVal_in_2_2;
      end else if (10'h173 == _T_19[9:0]) begin
        image_2_371 <= io_pixelVal_in_2_1;
      end else if (10'h173 == _T_15[9:0]) begin
        image_2_371 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_372 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h174 == _T_37[9:0]) begin
        image_2_372 <= io_pixelVal_in_2_7;
      end else if (10'h174 == _T_34[9:0]) begin
        image_2_372 <= io_pixelVal_in_2_6;
      end else if (10'h174 == _T_31[9:0]) begin
        image_2_372 <= io_pixelVal_in_2_5;
      end else if (10'h174 == _T_28[9:0]) begin
        image_2_372 <= io_pixelVal_in_2_4;
      end else if (10'h174 == _T_25[9:0]) begin
        image_2_372 <= io_pixelVal_in_2_3;
      end else if (10'h174 == _T_22[9:0]) begin
        image_2_372 <= io_pixelVal_in_2_2;
      end else if (10'h174 == _T_19[9:0]) begin
        image_2_372 <= io_pixelVal_in_2_1;
      end else if (10'h174 == _T_15[9:0]) begin
        image_2_372 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_373 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h175 == _T_37[9:0]) begin
        image_2_373 <= io_pixelVal_in_2_7;
      end else if (10'h175 == _T_34[9:0]) begin
        image_2_373 <= io_pixelVal_in_2_6;
      end else if (10'h175 == _T_31[9:0]) begin
        image_2_373 <= io_pixelVal_in_2_5;
      end else if (10'h175 == _T_28[9:0]) begin
        image_2_373 <= io_pixelVal_in_2_4;
      end else if (10'h175 == _T_25[9:0]) begin
        image_2_373 <= io_pixelVal_in_2_3;
      end else if (10'h175 == _T_22[9:0]) begin
        image_2_373 <= io_pixelVal_in_2_2;
      end else if (10'h175 == _T_19[9:0]) begin
        image_2_373 <= io_pixelVal_in_2_1;
      end else if (10'h175 == _T_15[9:0]) begin
        image_2_373 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_374 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h176 == _T_37[9:0]) begin
        image_2_374 <= io_pixelVal_in_2_7;
      end else if (10'h176 == _T_34[9:0]) begin
        image_2_374 <= io_pixelVal_in_2_6;
      end else if (10'h176 == _T_31[9:0]) begin
        image_2_374 <= io_pixelVal_in_2_5;
      end else if (10'h176 == _T_28[9:0]) begin
        image_2_374 <= io_pixelVal_in_2_4;
      end else if (10'h176 == _T_25[9:0]) begin
        image_2_374 <= io_pixelVal_in_2_3;
      end else if (10'h176 == _T_22[9:0]) begin
        image_2_374 <= io_pixelVal_in_2_2;
      end else if (10'h176 == _T_19[9:0]) begin
        image_2_374 <= io_pixelVal_in_2_1;
      end else if (10'h176 == _T_15[9:0]) begin
        image_2_374 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_375 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h177 == _T_37[9:0]) begin
        image_2_375 <= io_pixelVal_in_2_7;
      end else if (10'h177 == _T_34[9:0]) begin
        image_2_375 <= io_pixelVal_in_2_6;
      end else if (10'h177 == _T_31[9:0]) begin
        image_2_375 <= io_pixelVal_in_2_5;
      end else if (10'h177 == _T_28[9:0]) begin
        image_2_375 <= io_pixelVal_in_2_4;
      end else if (10'h177 == _T_25[9:0]) begin
        image_2_375 <= io_pixelVal_in_2_3;
      end else if (10'h177 == _T_22[9:0]) begin
        image_2_375 <= io_pixelVal_in_2_2;
      end else if (10'h177 == _T_19[9:0]) begin
        image_2_375 <= io_pixelVal_in_2_1;
      end else if (10'h177 == _T_15[9:0]) begin
        image_2_375 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_376 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h178 == _T_37[9:0]) begin
        image_2_376 <= io_pixelVal_in_2_7;
      end else if (10'h178 == _T_34[9:0]) begin
        image_2_376 <= io_pixelVal_in_2_6;
      end else if (10'h178 == _T_31[9:0]) begin
        image_2_376 <= io_pixelVal_in_2_5;
      end else if (10'h178 == _T_28[9:0]) begin
        image_2_376 <= io_pixelVal_in_2_4;
      end else if (10'h178 == _T_25[9:0]) begin
        image_2_376 <= io_pixelVal_in_2_3;
      end else if (10'h178 == _T_22[9:0]) begin
        image_2_376 <= io_pixelVal_in_2_2;
      end else if (10'h178 == _T_19[9:0]) begin
        image_2_376 <= io_pixelVal_in_2_1;
      end else if (10'h178 == _T_15[9:0]) begin
        image_2_376 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_377 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h179 == _T_37[9:0]) begin
        image_2_377 <= io_pixelVal_in_2_7;
      end else if (10'h179 == _T_34[9:0]) begin
        image_2_377 <= io_pixelVal_in_2_6;
      end else if (10'h179 == _T_31[9:0]) begin
        image_2_377 <= io_pixelVal_in_2_5;
      end else if (10'h179 == _T_28[9:0]) begin
        image_2_377 <= io_pixelVal_in_2_4;
      end else if (10'h179 == _T_25[9:0]) begin
        image_2_377 <= io_pixelVal_in_2_3;
      end else if (10'h179 == _T_22[9:0]) begin
        image_2_377 <= io_pixelVal_in_2_2;
      end else if (10'h179 == _T_19[9:0]) begin
        image_2_377 <= io_pixelVal_in_2_1;
      end else if (10'h179 == _T_15[9:0]) begin
        image_2_377 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_378 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17a == _T_37[9:0]) begin
        image_2_378 <= io_pixelVal_in_2_7;
      end else if (10'h17a == _T_34[9:0]) begin
        image_2_378 <= io_pixelVal_in_2_6;
      end else if (10'h17a == _T_31[9:0]) begin
        image_2_378 <= io_pixelVal_in_2_5;
      end else if (10'h17a == _T_28[9:0]) begin
        image_2_378 <= io_pixelVal_in_2_4;
      end else if (10'h17a == _T_25[9:0]) begin
        image_2_378 <= io_pixelVal_in_2_3;
      end else if (10'h17a == _T_22[9:0]) begin
        image_2_378 <= io_pixelVal_in_2_2;
      end else if (10'h17a == _T_19[9:0]) begin
        image_2_378 <= io_pixelVal_in_2_1;
      end else if (10'h17a == _T_15[9:0]) begin
        image_2_378 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_379 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17b == _T_37[9:0]) begin
        image_2_379 <= io_pixelVal_in_2_7;
      end else if (10'h17b == _T_34[9:0]) begin
        image_2_379 <= io_pixelVal_in_2_6;
      end else if (10'h17b == _T_31[9:0]) begin
        image_2_379 <= io_pixelVal_in_2_5;
      end else if (10'h17b == _T_28[9:0]) begin
        image_2_379 <= io_pixelVal_in_2_4;
      end else if (10'h17b == _T_25[9:0]) begin
        image_2_379 <= io_pixelVal_in_2_3;
      end else if (10'h17b == _T_22[9:0]) begin
        image_2_379 <= io_pixelVal_in_2_2;
      end else if (10'h17b == _T_19[9:0]) begin
        image_2_379 <= io_pixelVal_in_2_1;
      end else if (10'h17b == _T_15[9:0]) begin
        image_2_379 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_380 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17c == _T_37[9:0]) begin
        image_2_380 <= io_pixelVal_in_2_7;
      end else if (10'h17c == _T_34[9:0]) begin
        image_2_380 <= io_pixelVal_in_2_6;
      end else if (10'h17c == _T_31[9:0]) begin
        image_2_380 <= io_pixelVal_in_2_5;
      end else if (10'h17c == _T_28[9:0]) begin
        image_2_380 <= io_pixelVal_in_2_4;
      end else if (10'h17c == _T_25[9:0]) begin
        image_2_380 <= io_pixelVal_in_2_3;
      end else if (10'h17c == _T_22[9:0]) begin
        image_2_380 <= io_pixelVal_in_2_2;
      end else if (10'h17c == _T_19[9:0]) begin
        image_2_380 <= io_pixelVal_in_2_1;
      end else if (10'h17c == _T_15[9:0]) begin
        image_2_380 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_381 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17d == _T_37[9:0]) begin
        image_2_381 <= io_pixelVal_in_2_7;
      end else if (10'h17d == _T_34[9:0]) begin
        image_2_381 <= io_pixelVal_in_2_6;
      end else if (10'h17d == _T_31[9:0]) begin
        image_2_381 <= io_pixelVal_in_2_5;
      end else if (10'h17d == _T_28[9:0]) begin
        image_2_381 <= io_pixelVal_in_2_4;
      end else if (10'h17d == _T_25[9:0]) begin
        image_2_381 <= io_pixelVal_in_2_3;
      end else if (10'h17d == _T_22[9:0]) begin
        image_2_381 <= io_pixelVal_in_2_2;
      end else if (10'h17d == _T_19[9:0]) begin
        image_2_381 <= io_pixelVal_in_2_1;
      end else if (10'h17d == _T_15[9:0]) begin
        image_2_381 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_382 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17e == _T_37[9:0]) begin
        image_2_382 <= io_pixelVal_in_2_7;
      end else if (10'h17e == _T_34[9:0]) begin
        image_2_382 <= io_pixelVal_in_2_6;
      end else if (10'h17e == _T_31[9:0]) begin
        image_2_382 <= io_pixelVal_in_2_5;
      end else if (10'h17e == _T_28[9:0]) begin
        image_2_382 <= io_pixelVal_in_2_4;
      end else if (10'h17e == _T_25[9:0]) begin
        image_2_382 <= io_pixelVal_in_2_3;
      end else if (10'h17e == _T_22[9:0]) begin
        image_2_382 <= io_pixelVal_in_2_2;
      end else if (10'h17e == _T_19[9:0]) begin
        image_2_382 <= io_pixelVal_in_2_1;
      end else if (10'h17e == _T_15[9:0]) begin
        image_2_382 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_383 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17f == _T_37[9:0]) begin
        image_2_383 <= io_pixelVal_in_2_7;
      end else if (10'h17f == _T_34[9:0]) begin
        image_2_383 <= io_pixelVal_in_2_6;
      end else if (10'h17f == _T_31[9:0]) begin
        image_2_383 <= io_pixelVal_in_2_5;
      end else if (10'h17f == _T_28[9:0]) begin
        image_2_383 <= io_pixelVal_in_2_4;
      end else if (10'h17f == _T_25[9:0]) begin
        image_2_383 <= io_pixelVal_in_2_3;
      end else if (10'h17f == _T_22[9:0]) begin
        image_2_383 <= io_pixelVal_in_2_2;
      end else if (10'h17f == _T_19[9:0]) begin
        image_2_383 <= io_pixelVal_in_2_1;
      end else if (10'h17f == _T_15[9:0]) begin
        image_2_383 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_384 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h180 == _T_37[9:0]) begin
        image_2_384 <= io_pixelVal_in_2_7;
      end else if (10'h180 == _T_34[9:0]) begin
        image_2_384 <= io_pixelVal_in_2_6;
      end else if (10'h180 == _T_31[9:0]) begin
        image_2_384 <= io_pixelVal_in_2_5;
      end else if (10'h180 == _T_28[9:0]) begin
        image_2_384 <= io_pixelVal_in_2_4;
      end else if (10'h180 == _T_25[9:0]) begin
        image_2_384 <= io_pixelVal_in_2_3;
      end else if (10'h180 == _T_22[9:0]) begin
        image_2_384 <= io_pixelVal_in_2_2;
      end else if (10'h180 == _T_19[9:0]) begin
        image_2_384 <= io_pixelVal_in_2_1;
      end else if (10'h180 == _T_15[9:0]) begin
        image_2_384 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_385 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h181 == _T_37[9:0]) begin
        image_2_385 <= io_pixelVal_in_2_7;
      end else if (10'h181 == _T_34[9:0]) begin
        image_2_385 <= io_pixelVal_in_2_6;
      end else if (10'h181 == _T_31[9:0]) begin
        image_2_385 <= io_pixelVal_in_2_5;
      end else if (10'h181 == _T_28[9:0]) begin
        image_2_385 <= io_pixelVal_in_2_4;
      end else if (10'h181 == _T_25[9:0]) begin
        image_2_385 <= io_pixelVal_in_2_3;
      end else if (10'h181 == _T_22[9:0]) begin
        image_2_385 <= io_pixelVal_in_2_2;
      end else if (10'h181 == _T_19[9:0]) begin
        image_2_385 <= io_pixelVal_in_2_1;
      end else if (10'h181 == _T_15[9:0]) begin
        image_2_385 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_386 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h182 == _T_37[9:0]) begin
        image_2_386 <= io_pixelVal_in_2_7;
      end else if (10'h182 == _T_34[9:0]) begin
        image_2_386 <= io_pixelVal_in_2_6;
      end else if (10'h182 == _T_31[9:0]) begin
        image_2_386 <= io_pixelVal_in_2_5;
      end else if (10'h182 == _T_28[9:0]) begin
        image_2_386 <= io_pixelVal_in_2_4;
      end else if (10'h182 == _T_25[9:0]) begin
        image_2_386 <= io_pixelVal_in_2_3;
      end else if (10'h182 == _T_22[9:0]) begin
        image_2_386 <= io_pixelVal_in_2_2;
      end else if (10'h182 == _T_19[9:0]) begin
        image_2_386 <= io_pixelVal_in_2_1;
      end else if (10'h182 == _T_15[9:0]) begin
        image_2_386 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_387 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h183 == _T_37[9:0]) begin
        image_2_387 <= io_pixelVal_in_2_7;
      end else if (10'h183 == _T_34[9:0]) begin
        image_2_387 <= io_pixelVal_in_2_6;
      end else if (10'h183 == _T_31[9:0]) begin
        image_2_387 <= io_pixelVal_in_2_5;
      end else if (10'h183 == _T_28[9:0]) begin
        image_2_387 <= io_pixelVal_in_2_4;
      end else if (10'h183 == _T_25[9:0]) begin
        image_2_387 <= io_pixelVal_in_2_3;
      end else if (10'h183 == _T_22[9:0]) begin
        image_2_387 <= io_pixelVal_in_2_2;
      end else if (10'h183 == _T_19[9:0]) begin
        image_2_387 <= io_pixelVal_in_2_1;
      end else if (10'h183 == _T_15[9:0]) begin
        image_2_387 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_388 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h184 == _T_37[9:0]) begin
        image_2_388 <= io_pixelVal_in_2_7;
      end else if (10'h184 == _T_34[9:0]) begin
        image_2_388 <= io_pixelVal_in_2_6;
      end else if (10'h184 == _T_31[9:0]) begin
        image_2_388 <= io_pixelVal_in_2_5;
      end else if (10'h184 == _T_28[9:0]) begin
        image_2_388 <= io_pixelVal_in_2_4;
      end else if (10'h184 == _T_25[9:0]) begin
        image_2_388 <= io_pixelVal_in_2_3;
      end else if (10'h184 == _T_22[9:0]) begin
        image_2_388 <= io_pixelVal_in_2_2;
      end else if (10'h184 == _T_19[9:0]) begin
        image_2_388 <= io_pixelVal_in_2_1;
      end else if (10'h184 == _T_15[9:0]) begin
        image_2_388 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_389 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h185 == _T_37[9:0]) begin
        image_2_389 <= io_pixelVal_in_2_7;
      end else if (10'h185 == _T_34[9:0]) begin
        image_2_389 <= io_pixelVal_in_2_6;
      end else if (10'h185 == _T_31[9:0]) begin
        image_2_389 <= io_pixelVal_in_2_5;
      end else if (10'h185 == _T_28[9:0]) begin
        image_2_389 <= io_pixelVal_in_2_4;
      end else if (10'h185 == _T_25[9:0]) begin
        image_2_389 <= io_pixelVal_in_2_3;
      end else if (10'h185 == _T_22[9:0]) begin
        image_2_389 <= io_pixelVal_in_2_2;
      end else if (10'h185 == _T_19[9:0]) begin
        image_2_389 <= io_pixelVal_in_2_1;
      end else if (10'h185 == _T_15[9:0]) begin
        image_2_389 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_390 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h186 == _T_37[9:0]) begin
        image_2_390 <= io_pixelVal_in_2_7;
      end else if (10'h186 == _T_34[9:0]) begin
        image_2_390 <= io_pixelVal_in_2_6;
      end else if (10'h186 == _T_31[9:0]) begin
        image_2_390 <= io_pixelVal_in_2_5;
      end else if (10'h186 == _T_28[9:0]) begin
        image_2_390 <= io_pixelVal_in_2_4;
      end else if (10'h186 == _T_25[9:0]) begin
        image_2_390 <= io_pixelVal_in_2_3;
      end else if (10'h186 == _T_22[9:0]) begin
        image_2_390 <= io_pixelVal_in_2_2;
      end else if (10'h186 == _T_19[9:0]) begin
        image_2_390 <= io_pixelVal_in_2_1;
      end else if (10'h186 == _T_15[9:0]) begin
        image_2_390 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_391 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h187 == _T_37[9:0]) begin
        image_2_391 <= io_pixelVal_in_2_7;
      end else if (10'h187 == _T_34[9:0]) begin
        image_2_391 <= io_pixelVal_in_2_6;
      end else if (10'h187 == _T_31[9:0]) begin
        image_2_391 <= io_pixelVal_in_2_5;
      end else if (10'h187 == _T_28[9:0]) begin
        image_2_391 <= io_pixelVal_in_2_4;
      end else if (10'h187 == _T_25[9:0]) begin
        image_2_391 <= io_pixelVal_in_2_3;
      end else if (10'h187 == _T_22[9:0]) begin
        image_2_391 <= io_pixelVal_in_2_2;
      end else if (10'h187 == _T_19[9:0]) begin
        image_2_391 <= io_pixelVal_in_2_1;
      end else if (10'h187 == _T_15[9:0]) begin
        image_2_391 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_392 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h188 == _T_37[9:0]) begin
        image_2_392 <= io_pixelVal_in_2_7;
      end else if (10'h188 == _T_34[9:0]) begin
        image_2_392 <= io_pixelVal_in_2_6;
      end else if (10'h188 == _T_31[9:0]) begin
        image_2_392 <= io_pixelVal_in_2_5;
      end else if (10'h188 == _T_28[9:0]) begin
        image_2_392 <= io_pixelVal_in_2_4;
      end else if (10'h188 == _T_25[9:0]) begin
        image_2_392 <= io_pixelVal_in_2_3;
      end else if (10'h188 == _T_22[9:0]) begin
        image_2_392 <= io_pixelVal_in_2_2;
      end else if (10'h188 == _T_19[9:0]) begin
        image_2_392 <= io_pixelVal_in_2_1;
      end else if (10'h188 == _T_15[9:0]) begin
        image_2_392 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_393 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h189 == _T_37[9:0]) begin
        image_2_393 <= io_pixelVal_in_2_7;
      end else if (10'h189 == _T_34[9:0]) begin
        image_2_393 <= io_pixelVal_in_2_6;
      end else if (10'h189 == _T_31[9:0]) begin
        image_2_393 <= io_pixelVal_in_2_5;
      end else if (10'h189 == _T_28[9:0]) begin
        image_2_393 <= io_pixelVal_in_2_4;
      end else if (10'h189 == _T_25[9:0]) begin
        image_2_393 <= io_pixelVal_in_2_3;
      end else if (10'h189 == _T_22[9:0]) begin
        image_2_393 <= io_pixelVal_in_2_2;
      end else if (10'h189 == _T_19[9:0]) begin
        image_2_393 <= io_pixelVal_in_2_1;
      end else if (10'h189 == _T_15[9:0]) begin
        image_2_393 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_394 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18a == _T_37[9:0]) begin
        image_2_394 <= io_pixelVal_in_2_7;
      end else if (10'h18a == _T_34[9:0]) begin
        image_2_394 <= io_pixelVal_in_2_6;
      end else if (10'h18a == _T_31[9:0]) begin
        image_2_394 <= io_pixelVal_in_2_5;
      end else if (10'h18a == _T_28[9:0]) begin
        image_2_394 <= io_pixelVal_in_2_4;
      end else if (10'h18a == _T_25[9:0]) begin
        image_2_394 <= io_pixelVal_in_2_3;
      end else if (10'h18a == _T_22[9:0]) begin
        image_2_394 <= io_pixelVal_in_2_2;
      end else if (10'h18a == _T_19[9:0]) begin
        image_2_394 <= io_pixelVal_in_2_1;
      end else if (10'h18a == _T_15[9:0]) begin
        image_2_394 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_395 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18b == _T_37[9:0]) begin
        image_2_395 <= io_pixelVal_in_2_7;
      end else if (10'h18b == _T_34[9:0]) begin
        image_2_395 <= io_pixelVal_in_2_6;
      end else if (10'h18b == _T_31[9:0]) begin
        image_2_395 <= io_pixelVal_in_2_5;
      end else if (10'h18b == _T_28[9:0]) begin
        image_2_395 <= io_pixelVal_in_2_4;
      end else if (10'h18b == _T_25[9:0]) begin
        image_2_395 <= io_pixelVal_in_2_3;
      end else if (10'h18b == _T_22[9:0]) begin
        image_2_395 <= io_pixelVal_in_2_2;
      end else if (10'h18b == _T_19[9:0]) begin
        image_2_395 <= io_pixelVal_in_2_1;
      end else if (10'h18b == _T_15[9:0]) begin
        image_2_395 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_396 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18c == _T_37[9:0]) begin
        image_2_396 <= io_pixelVal_in_2_7;
      end else if (10'h18c == _T_34[9:0]) begin
        image_2_396 <= io_pixelVal_in_2_6;
      end else if (10'h18c == _T_31[9:0]) begin
        image_2_396 <= io_pixelVal_in_2_5;
      end else if (10'h18c == _T_28[9:0]) begin
        image_2_396 <= io_pixelVal_in_2_4;
      end else if (10'h18c == _T_25[9:0]) begin
        image_2_396 <= io_pixelVal_in_2_3;
      end else if (10'h18c == _T_22[9:0]) begin
        image_2_396 <= io_pixelVal_in_2_2;
      end else if (10'h18c == _T_19[9:0]) begin
        image_2_396 <= io_pixelVal_in_2_1;
      end else if (10'h18c == _T_15[9:0]) begin
        image_2_396 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_397 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18d == _T_37[9:0]) begin
        image_2_397 <= io_pixelVal_in_2_7;
      end else if (10'h18d == _T_34[9:0]) begin
        image_2_397 <= io_pixelVal_in_2_6;
      end else if (10'h18d == _T_31[9:0]) begin
        image_2_397 <= io_pixelVal_in_2_5;
      end else if (10'h18d == _T_28[9:0]) begin
        image_2_397 <= io_pixelVal_in_2_4;
      end else if (10'h18d == _T_25[9:0]) begin
        image_2_397 <= io_pixelVal_in_2_3;
      end else if (10'h18d == _T_22[9:0]) begin
        image_2_397 <= io_pixelVal_in_2_2;
      end else if (10'h18d == _T_19[9:0]) begin
        image_2_397 <= io_pixelVal_in_2_1;
      end else if (10'h18d == _T_15[9:0]) begin
        image_2_397 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_398 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18e == _T_37[9:0]) begin
        image_2_398 <= io_pixelVal_in_2_7;
      end else if (10'h18e == _T_34[9:0]) begin
        image_2_398 <= io_pixelVal_in_2_6;
      end else if (10'h18e == _T_31[9:0]) begin
        image_2_398 <= io_pixelVal_in_2_5;
      end else if (10'h18e == _T_28[9:0]) begin
        image_2_398 <= io_pixelVal_in_2_4;
      end else if (10'h18e == _T_25[9:0]) begin
        image_2_398 <= io_pixelVal_in_2_3;
      end else if (10'h18e == _T_22[9:0]) begin
        image_2_398 <= io_pixelVal_in_2_2;
      end else if (10'h18e == _T_19[9:0]) begin
        image_2_398 <= io_pixelVal_in_2_1;
      end else if (10'h18e == _T_15[9:0]) begin
        image_2_398 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_399 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18f == _T_37[9:0]) begin
        image_2_399 <= io_pixelVal_in_2_7;
      end else if (10'h18f == _T_34[9:0]) begin
        image_2_399 <= io_pixelVal_in_2_6;
      end else if (10'h18f == _T_31[9:0]) begin
        image_2_399 <= io_pixelVal_in_2_5;
      end else if (10'h18f == _T_28[9:0]) begin
        image_2_399 <= io_pixelVal_in_2_4;
      end else if (10'h18f == _T_25[9:0]) begin
        image_2_399 <= io_pixelVal_in_2_3;
      end else if (10'h18f == _T_22[9:0]) begin
        image_2_399 <= io_pixelVal_in_2_2;
      end else if (10'h18f == _T_19[9:0]) begin
        image_2_399 <= io_pixelVal_in_2_1;
      end else if (10'h18f == _T_15[9:0]) begin
        image_2_399 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_400 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h190 == _T_37[9:0]) begin
        image_2_400 <= io_pixelVal_in_2_7;
      end else if (10'h190 == _T_34[9:0]) begin
        image_2_400 <= io_pixelVal_in_2_6;
      end else if (10'h190 == _T_31[9:0]) begin
        image_2_400 <= io_pixelVal_in_2_5;
      end else if (10'h190 == _T_28[9:0]) begin
        image_2_400 <= io_pixelVal_in_2_4;
      end else if (10'h190 == _T_25[9:0]) begin
        image_2_400 <= io_pixelVal_in_2_3;
      end else if (10'h190 == _T_22[9:0]) begin
        image_2_400 <= io_pixelVal_in_2_2;
      end else if (10'h190 == _T_19[9:0]) begin
        image_2_400 <= io_pixelVal_in_2_1;
      end else if (10'h190 == _T_15[9:0]) begin
        image_2_400 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_401 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h191 == _T_37[9:0]) begin
        image_2_401 <= io_pixelVal_in_2_7;
      end else if (10'h191 == _T_34[9:0]) begin
        image_2_401 <= io_pixelVal_in_2_6;
      end else if (10'h191 == _T_31[9:0]) begin
        image_2_401 <= io_pixelVal_in_2_5;
      end else if (10'h191 == _T_28[9:0]) begin
        image_2_401 <= io_pixelVal_in_2_4;
      end else if (10'h191 == _T_25[9:0]) begin
        image_2_401 <= io_pixelVal_in_2_3;
      end else if (10'h191 == _T_22[9:0]) begin
        image_2_401 <= io_pixelVal_in_2_2;
      end else if (10'h191 == _T_19[9:0]) begin
        image_2_401 <= io_pixelVal_in_2_1;
      end else if (10'h191 == _T_15[9:0]) begin
        image_2_401 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_402 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h192 == _T_37[9:0]) begin
        image_2_402 <= io_pixelVal_in_2_7;
      end else if (10'h192 == _T_34[9:0]) begin
        image_2_402 <= io_pixelVal_in_2_6;
      end else if (10'h192 == _T_31[9:0]) begin
        image_2_402 <= io_pixelVal_in_2_5;
      end else if (10'h192 == _T_28[9:0]) begin
        image_2_402 <= io_pixelVal_in_2_4;
      end else if (10'h192 == _T_25[9:0]) begin
        image_2_402 <= io_pixelVal_in_2_3;
      end else if (10'h192 == _T_22[9:0]) begin
        image_2_402 <= io_pixelVal_in_2_2;
      end else if (10'h192 == _T_19[9:0]) begin
        image_2_402 <= io_pixelVal_in_2_1;
      end else if (10'h192 == _T_15[9:0]) begin
        image_2_402 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_403 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h193 == _T_37[9:0]) begin
        image_2_403 <= io_pixelVal_in_2_7;
      end else if (10'h193 == _T_34[9:0]) begin
        image_2_403 <= io_pixelVal_in_2_6;
      end else if (10'h193 == _T_31[9:0]) begin
        image_2_403 <= io_pixelVal_in_2_5;
      end else if (10'h193 == _T_28[9:0]) begin
        image_2_403 <= io_pixelVal_in_2_4;
      end else if (10'h193 == _T_25[9:0]) begin
        image_2_403 <= io_pixelVal_in_2_3;
      end else if (10'h193 == _T_22[9:0]) begin
        image_2_403 <= io_pixelVal_in_2_2;
      end else if (10'h193 == _T_19[9:0]) begin
        image_2_403 <= io_pixelVal_in_2_1;
      end else if (10'h193 == _T_15[9:0]) begin
        image_2_403 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_404 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h194 == _T_37[9:0]) begin
        image_2_404 <= io_pixelVal_in_2_7;
      end else if (10'h194 == _T_34[9:0]) begin
        image_2_404 <= io_pixelVal_in_2_6;
      end else if (10'h194 == _T_31[9:0]) begin
        image_2_404 <= io_pixelVal_in_2_5;
      end else if (10'h194 == _T_28[9:0]) begin
        image_2_404 <= io_pixelVal_in_2_4;
      end else if (10'h194 == _T_25[9:0]) begin
        image_2_404 <= io_pixelVal_in_2_3;
      end else if (10'h194 == _T_22[9:0]) begin
        image_2_404 <= io_pixelVal_in_2_2;
      end else if (10'h194 == _T_19[9:0]) begin
        image_2_404 <= io_pixelVal_in_2_1;
      end else if (10'h194 == _T_15[9:0]) begin
        image_2_404 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_405 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h195 == _T_37[9:0]) begin
        image_2_405 <= io_pixelVal_in_2_7;
      end else if (10'h195 == _T_34[9:0]) begin
        image_2_405 <= io_pixelVal_in_2_6;
      end else if (10'h195 == _T_31[9:0]) begin
        image_2_405 <= io_pixelVal_in_2_5;
      end else if (10'h195 == _T_28[9:0]) begin
        image_2_405 <= io_pixelVal_in_2_4;
      end else if (10'h195 == _T_25[9:0]) begin
        image_2_405 <= io_pixelVal_in_2_3;
      end else if (10'h195 == _T_22[9:0]) begin
        image_2_405 <= io_pixelVal_in_2_2;
      end else if (10'h195 == _T_19[9:0]) begin
        image_2_405 <= io_pixelVal_in_2_1;
      end else if (10'h195 == _T_15[9:0]) begin
        image_2_405 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_406 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h196 == _T_37[9:0]) begin
        image_2_406 <= io_pixelVal_in_2_7;
      end else if (10'h196 == _T_34[9:0]) begin
        image_2_406 <= io_pixelVal_in_2_6;
      end else if (10'h196 == _T_31[9:0]) begin
        image_2_406 <= io_pixelVal_in_2_5;
      end else if (10'h196 == _T_28[9:0]) begin
        image_2_406 <= io_pixelVal_in_2_4;
      end else if (10'h196 == _T_25[9:0]) begin
        image_2_406 <= io_pixelVal_in_2_3;
      end else if (10'h196 == _T_22[9:0]) begin
        image_2_406 <= io_pixelVal_in_2_2;
      end else if (10'h196 == _T_19[9:0]) begin
        image_2_406 <= io_pixelVal_in_2_1;
      end else if (10'h196 == _T_15[9:0]) begin
        image_2_406 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_407 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h197 == _T_37[9:0]) begin
        image_2_407 <= io_pixelVal_in_2_7;
      end else if (10'h197 == _T_34[9:0]) begin
        image_2_407 <= io_pixelVal_in_2_6;
      end else if (10'h197 == _T_31[9:0]) begin
        image_2_407 <= io_pixelVal_in_2_5;
      end else if (10'h197 == _T_28[9:0]) begin
        image_2_407 <= io_pixelVal_in_2_4;
      end else if (10'h197 == _T_25[9:0]) begin
        image_2_407 <= io_pixelVal_in_2_3;
      end else if (10'h197 == _T_22[9:0]) begin
        image_2_407 <= io_pixelVal_in_2_2;
      end else if (10'h197 == _T_19[9:0]) begin
        image_2_407 <= io_pixelVal_in_2_1;
      end else if (10'h197 == _T_15[9:0]) begin
        image_2_407 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_408 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h198 == _T_37[9:0]) begin
        image_2_408 <= io_pixelVal_in_2_7;
      end else if (10'h198 == _T_34[9:0]) begin
        image_2_408 <= io_pixelVal_in_2_6;
      end else if (10'h198 == _T_31[9:0]) begin
        image_2_408 <= io_pixelVal_in_2_5;
      end else if (10'h198 == _T_28[9:0]) begin
        image_2_408 <= io_pixelVal_in_2_4;
      end else if (10'h198 == _T_25[9:0]) begin
        image_2_408 <= io_pixelVal_in_2_3;
      end else if (10'h198 == _T_22[9:0]) begin
        image_2_408 <= io_pixelVal_in_2_2;
      end else if (10'h198 == _T_19[9:0]) begin
        image_2_408 <= io_pixelVal_in_2_1;
      end else if (10'h198 == _T_15[9:0]) begin
        image_2_408 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_409 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h199 == _T_37[9:0]) begin
        image_2_409 <= io_pixelVal_in_2_7;
      end else if (10'h199 == _T_34[9:0]) begin
        image_2_409 <= io_pixelVal_in_2_6;
      end else if (10'h199 == _T_31[9:0]) begin
        image_2_409 <= io_pixelVal_in_2_5;
      end else if (10'h199 == _T_28[9:0]) begin
        image_2_409 <= io_pixelVal_in_2_4;
      end else if (10'h199 == _T_25[9:0]) begin
        image_2_409 <= io_pixelVal_in_2_3;
      end else if (10'h199 == _T_22[9:0]) begin
        image_2_409 <= io_pixelVal_in_2_2;
      end else if (10'h199 == _T_19[9:0]) begin
        image_2_409 <= io_pixelVal_in_2_1;
      end else if (10'h199 == _T_15[9:0]) begin
        image_2_409 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_410 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19a == _T_37[9:0]) begin
        image_2_410 <= io_pixelVal_in_2_7;
      end else if (10'h19a == _T_34[9:0]) begin
        image_2_410 <= io_pixelVal_in_2_6;
      end else if (10'h19a == _T_31[9:0]) begin
        image_2_410 <= io_pixelVal_in_2_5;
      end else if (10'h19a == _T_28[9:0]) begin
        image_2_410 <= io_pixelVal_in_2_4;
      end else if (10'h19a == _T_25[9:0]) begin
        image_2_410 <= io_pixelVal_in_2_3;
      end else if (10'h19a == _T_22[9:0]) begin
        image_2_410 <= io_pixelVal_in_2_2;
      end else if (10'h19a == _T_19[9:0]) begin
        image_2_410 <= io_pixelVal_in_2_1;
      end else if (10'h19a == _T_15[9:0]) begin
        image_2_410 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_411 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19b == _T_37[9:0]) begin
        image_2_411 <= io_pixelVal_in_2_7;
      end else if (10'h19b == _T_34[9:0]) begin
        image_2_411 <= io_pixelVal_in_2_6;
      end else if (10'h19b == _T_31[9:0]) begin
        image_2_411 <= io_pixelVal_in_2_5;
      end else if (10'h19b == _T_28[9:0]) begin
        image_2_411 <= io_pixelVal_in_2_4;
      end else if (10'h19b == _T_25[9:0]) begin
        image_2_411 <= io_pixelVal_in_2_3;
      end else if (10'h19b == _T_22[9:0]) begin
        image_2_411 <= io_pixelVal_in_2_2;
      end else if (10'h19b == _T_19[9:0]) begin
        image_2_411 <= io_pixelVal_in_2_1;
      end else if (10'h19b == _T_15[9:0]) begin
        image_2_411 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_412 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19c == _T_37[9:0]) begin
        image_2_412 <= io_pixelVal_in_2_7;
      end else if (10'h19c == _T_34[9:0]) begin
        image_2_412 <= io_pixelVal_in_2_6;
      end else if (10'h19c == _T_31[9:0]) begin
        image_2_412 <= io_pixelVal_in_2_5;
      end else if (10'h19c == _T_28[9:0]) begin
        image_2_412 <= io_pixelVal_in_2_4;
      end else if (10'h19c == _T_25[9:0]) begin
        image_2_412 <= io_pixelVal_in_2_3;
      end else if (10'h19c == _T_22[9:0]) begin
        image_2_412 <= io_pixelVal_in_2_2;
      end else if (10'h19c == _T_19[9:0]) begin
        image_2_412 <= io_pixelVal_in_2_1;
      end else if (10'h19c == _T_15[9:0]) begin
        image_2_412 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_413 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19d == _T_37[9:0]) begin
        image_2_413 <= io_pixelVal_in_2_7;
      end else if (10'h19d == _T_34[9:0]) begin
        image_2_413 <= io_pixelVal_in_2_6;
      end else if (10'h19d == _T_31[9:0]) begin
        image_2_413 <= io_pixelVal_in_2_5;
      end else if (10'h19d == _T_28[9:0]) begin
        image_2_413 <= io_pixelVal_in_2_4;
      end else if (10'h19d == _T_25[9:0]) begin
        image_2_413 <= io_pixelVal_in_2_3;
      end else if (10'h19d == _T_22[9:0]) begin
        image_2_413 <= io_pixelVal_in_2_2;
      end else if (10'h19d == _T_19[9:0]) begin
        image_2_413 <= io_pixelVal_in_2_1;
      end else if (10'h19d == _T_15[9:0]) begin
        image_2_413 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_414 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19e == _T_37[9:0]) begin
        image_2_414 <= io_pixelVal_in_2_7;
      end else if (10'h19e == _T_34[9:0]) begin
        image_2_414 <= io_pixelVal_in_2_6;
      end else if (10'h19e == _T_31[9:0]) begin
        image_2_414 <= io_pixelVal_in_2_5;
      end else if (10'h19e == _T_28[9:0]) begin
        image_2_414 <= io_pixelVal_in_2_4;
      end else if (10'h19e == _T_25[9:0]) begin
        image_2_414 <= io_pixelVal_in_2_3;
      end else if (10'h19e == _T_22[9:0]) begin
        image_2_414 <= io_pixelVal_in_2_2;
      end else if (10'h19e == _T_19[9:0]) begin
        image_2_414 <= io_pixelVal_in_2_1;
      end else if (10'h19e == _T_15[9:0]) begin
        image_2_414 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_415 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19f == _T_37[9:0]) begin
        image_2_415 <= io_pixelVal_in_2_7;
      end else if (10'h19f == _T_34[9:0]) begin
        image_2_415 <= io_pixelVal_in_2_6;
      end else if (10'h19f == _T_31[9:0]) begin
        image_2_415 <= io_pixelVal_in_2_5;
      end else if (10'h19f == _T_28[9:0]) begin
        image_2_415 <= io_pixelVal_in_2_4;
      end else if (10'h19f == _T_25[9:0]) begin
        image_2_415 <= io_pixelVal_in_2_3;
      end else if (10'h19f == _T_22[9:0]) begin
        image_2_415 <= io_pixelVal_in_2_2;
      end else if (10'h19f == _T_19[9:0]) begin
        image_2_415 <= io_pixelVal_in_2_1;
      end else if (10'h19f == _T_15[9:0]) begin
        image_2_415 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_416 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a0 == _T_37[9:0]) begin
        image_2_416 <= io_pixelVal_in_2_7;
      end else if (10'h1a0 == _T_34[9:0]) begin
        image_2_416 <= io_pixelVal_in_2_6;
      end else if (10'h1a0 == _T_31[9:0]) begin
        image_2_416 <= io_pixelVal_in_2_5;
      end else if (10'h1a0 == _T_28[9:0]) begin
        image_2_416 <= io_pixelVal_in_2_4;
      end else if (10'h1a0 == _T_25[9:0]) begin
        image_2_416 <= io_pixelVal_in_2_3;
      end else if (10'h1a0 == _T_22[9:0]) begin
        image_2_416 <= io_pixelVal_in_2_2;
      end else if (10'h1a0 == _T_19[9:0]) begin
        image_2_416 <= io_pixelVal_in_2_1;
      end else if (10'h1a0 == _T_15[9:0]) begin
        image_2_416 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_417 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a1 == _T_37[9:0]) begin
        image_2_417 <= io_pixelVal_in_2_7;
      end else if (10'h1a1 == _T_34[9:0]) begin
        image_2_417 <= io_pixelVal_in_2_6;
      end else if (10'h1a1 == _T_31[9:0]) begin
        image_2_417 <= io_pixelVal_in_2_5;
      end else if (10'h1a1 == _T_28[9:0]) begin
        image_2_417 <= io_pixelVal_in_2_4;
      end else if (10'h1a1 == _T_25[9:0]) begin
        image_2_417 <= io_pixelVal_in_2_3;
      end else if (10'h1a1 == _T_22[9:0]) begin
        image_2_417 <= io_pixelVal_in_2_2;
      end else if (10'h1a1 == _T_19[9:0]) begin
        image_2_417 <= io_pixelVal_in_2_1;
      end else if (10'h1a1 == _T_15[9:0]) begin
        image_2_417 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_418 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a2 == _T_37[9:0]) begin
        image_2_418 <= io_pixelVal_in_2_7;
      end else if (10'h1a2 == _T_34[9:0]) begin
        image_2_418 <= io_pixelVal_in_2_6;
      end else if (10'h1a2 == _T_31[9:0]) begin
        image_2_418 <= io_pixelVal_in_2_5;
      end else if (10'h1a2 == _T_28[9:0]) begin
        image_2_418 <= io_pixelVal_in_2_4;
      end else if (10'h1a2 == _T_25[9:0]) begin
        image_2_418 <= io_pixelVal_in_2_3;
      end else if (10'h1a2 == _T_22[9:0]) begin
        image_2_418 <= io_pixelVal_in_2_2;
      end else if (10'h1a2 == _T_19[9:0]) begin
        image_2_418 <= io_pixelVal_in_2_1;
      end else if (10'h1a2 == _T_15[9:0]) begin
        image_2_418 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_419 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a3 == _T_37[9:0]) begin
        image_2_419 <= io_pixelVal_in_2_7;
      end else if (10'h1a3 == _T_34[9:0]) begin
        image_2_419 <= io_pixelVal_in_2_6;
      end else if (10'h1a3 == _T_31[9:0]) begin
        image_2_419 <= io_pixelVal_in_2_5;
      end else if (10'h1a3 == _T_28[9:0]) begin
        image_2_419 <= io_pixelVal_in_2_4;
      end else if (10'h1a3 == _T_25[9:0]) begin
        image_2_419 <= io_pixelVal_in_2_3;
      end else if (10'h1a3 == _T_22[9:0]) begin
        image_2_419 <= io_pixelVal_in_2_2;
      end else if (10'h1a3 == _T_19[9:0]) begin
        image_2_419 <= io_pixelVal_in_2_1;
      end else if (10'h1a3 == _T_15[9:0]) begin
        image_2_419 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_420 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a4 == _T_37[9:0]) begin
        image_2_420 <= io_pixelVal_in_2_7;
      end else if (10'h1a4 == _T_34[9:0]) begin
        image_2_420 <= io_pixelVal_in_2_6;
      end else if (10'h1a4 == _T_31[9:0]) begin
        image_2_420 <= io_pixelVal_in_2_5;
      end else if (10'h1a4 == _T_28[9:0]) begin
        image_2_420 <= io_pixelVal_in_2_4;
      end else if (10'h1a4 == _T_25[9:0]) begin
        image_2_420 <= io_pixelVal_in_2_3;
      end else if (10'h1a4 == _T_22[9:0]) begin
        image_2_420 <= io_pixelVal_in_2_2;
      end else if (10'h1a4 == _T_19[9:0]) begin
        image_2_420 <= io_pixelVal_in_2_1;
      end else if (10'h1a4 == _T_15[9:0]) begin
        image_2_420 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_421 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a5 == _T_37[9:0]) begin
        image_2_421 <= io_pixelVal_in_2_7;
      end else if (10'h1a5 == _T_34[9:0]) begin
        image_2_421 <= io_pixelVal_in_2_6;
      end else if (10'h1a5 == _T_31[9:0]) begin
        image_2_421 <= io_pixelVal_in_2_5;
      end else if (10'h1a5 == _T_28[9:0]) begin
        image_2_421 <= io_pixelVal_in_2_4;
      end else if (10'h1a5 == _T_25[9:0]) begin
        image_2_421 <= io_pixelVal_in_2_3;
      end else if (10'h1a5 == _T_22[9:0]) begin
        image_2_421 <= io_pixelVal_in_2_2;
      end else if (10'h1a5 == _T_19[9:0]) begin
        image_2_421 <= io_pixelVal_in_2_1;
      end else if (10'h1a5 == _T_15[9:0]) begin
        image_2_421 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_422 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a6 == _T_37[9:0]) begin
        image_2_422 <= io_pixelVal_in_2_7;
      end else if (10'h1a6 == _T_34[9:0]) begin
        image_2_422 <= io_pixelVal_in_2_6;
      end else if (10'h1a6 == _T_31[9:0]) begin
        image_2_422 <= io_pixelVal_in_2_5;
      end else if (10'h1a6 == _T_28[9:0]) begin
        image_2_422 <= io_pixelVal_in_2_4;
      end else if (10'h1a6 == _T_25[9:0]) begin
        image_2_422 <= io_pixelVal_in_2_3;
      end else if (10'h1a6 == _T_22[9:0]) begin
        image_2_422 <= io_pixelVal_in_2_2;
      end else if (10'h1a6 == _T_19[9:0]) begin
        image_2_422 <= io_pixelVal_in_2_1;
      end else if (10'h1a6 == _T_15[9:0]) begin
        image_2_422 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_423 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a7 == _T_37[9:0]) begin
        image_2_423 <= io_pixelVal_in_2_7;
      end else if (10'h1a7 == _T_34[9:0]) begin
        image_2_423 <= io_pixelVal_in_2_6;
      end else if (10'h1a7 == _T_31[9:0]) begin
        image_2_423 <= io_pixelVal_in_2_5;
      end else if (10'h1a7 == _T_28[9:0]) begin
        image_2_423 <= io_pixelVal_in_2_4;
      end else if (10'h1a7 == _T_25[9:0]) begin
        image_2_423 <= io_pixelVal_in_2_3;
      end else if (10'h1a7 == _T_22[9:0]) begin
        image_2_423 <= io_pixelVal_in_2_2;
      end else if (10'h1a7 == _T_19[9:0]) begin
        image_2_423 <= io_pixelVal_in_2_1;
      end else if (10'h1a7 == _T_15[9:0]) begin
        image_2_423 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_424 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a8 == _T_37[9:0]) begin
        image_2_424 <= io_pixelVal_in_2_7;
      end else if (10'h1a8 == _T_34[9:0]) begin
        image_2_424 <= io_pixelVal_in_2_6;
      end else if (10'h1a8 == _T_31[9:0]) begin
        image_2_424 <= io_pixelVal_in_2_5;
      end else if (10'h1a8 == _T_28[9:0]) begin
        image_2_424 <= io_pixelVal_in_2_4;
      end else if (10'h1a8 == _T_25[9:0]) begin
        image_2_424 <= io_pixelVal_in_2_3;
      end else if (10'h1a8 == _T_22[9:0]) begin
        image_2_424 <= io_pixelVal_in_2_2;
      end else if (10'h1a8 == _T_19[9:0]) begin
        image_2_424 <= io_pixelVal_in_2_1;
      end else if (10'h1a8 == _T_15[9:0]) begin
        image_2_424 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_425 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a9 == _T_37[9:0]) begin
        image_2_425 <= io_pixelVal_in_2_7;
      end else if (10'h1a9 == _T_34[9:0]) begin
        image_2_425 <= io_pixelVal_in_2_6;
      end else if (10'h1a9 == _T_31[9:0]) begin
        image_2_425 <= io_pixelVal_in_2_5;
      end else if (10'h1a9 == _T_28[9:0]) begin
        image_2_425 <= io_pixelVal_in_2_4;
      end else if (10'h1a9 == _T_25[9:0]) begin
        image_2_425 <= io_pixelVal_in_2_3;
      end else if (10'h1a9 == _T_22[9:0]) begin
        image_2_425 <= io_pixelVal_in_2_2;
      end else if (10'h1a9 == _T_19[9:0]) begin
        image_2_425 <= io_pixelVal_in_2_1;
      end else if (10'h1a9 == _T_15[9:0]) begin
        image_2_425 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_426 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1aa == _T_37[9:0]) begin
        image_2_426 <= io_pixelVal_in_2_7;
      end else if (10'h1aa == _T_34[9:0]) begin
        image_2_426 <= io_pixelVal_in_2_6;
      end else if (10'h1aa == _T_31[9:0]) begin
        image_2_426 <= io_pixelVal_in_2_5;
      end else if (10'h1aa == _T_28[9:0]) begin
        image_2_426 <= io_pixelVal_in_2_4;
      end else if (10'h1aa == _T_25[9:0]) begin
        image_2_426 <= io_pixelVal_in_2_3;
      end else if (10'h1aa == _T_22[9:0]) begin
        image_2_426 <= io_pixelVal_in_2_2;
      end else if (10'h1aa == _T_19[9:0]) begin
        image_2_426 <= io_pixelVal_in_2_1;
      end else if (10'h1aa == _T_15[9:0]) begin
        image_2_426 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_427 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ab == _T_37[9:0]) begin
        image_2_427 <= io_pixelVal_in_2_7;
      end else if (10'h1ab == _T_34[9:0]) begin
        image_2_427 <= io_pixelVal_in_2_6;
      end else if (10'h1ab == _T_31[9:0]) begin
        image_2_427 <= io_pixelVal_in_2_5;
      end else if (10'h1ab == _T_28[9:0]) begin
        image_2_427 <= io_pixelVal_in_2_4;
      end else if (10'h1ab == _T_25[9:0]) begin
        image_2_427 <= io_pixelVal_in_2_3;
      end else if (10'h1ab == _T_22[9:0]) begin
        image_2_427 <= io_pixelVal_in_2_2;
      end else if (10'h1ab == _T_19[9:0]) begin
        image_2_427 <= io_pixelVal_in_2_1;
      end else if (10'h1ab == _T_15[9:0]) begin
        image_2_427 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_428 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ac == _T_37[9:0]) begin
        image_2_428 <= io_pixelVal_in_2_7;
      end else if (10'h1ac == _T_34[9:0]) begin
        image_2_428 <= io_pixelVal_in_2_6;
      end else if (10'h1ac == _T_31[9:0]) begin
        image_2_428 <= io_pixelVal_in_2_5;
      end else if (10'h1ac == _T_28[9:0]) begin
        image_2_428 <= io_pixelVal_in_2_4;
      end else if (10'h1ac == _T_25[9:0]) begin
        image_2_428 <= io_pixelVal_in_2_3;
      end else if (10'h1ac == _T_22[9:0]) begin
        image_2_428 <= io_pixelVal_in_2_2;
      end else if (10'h1ac == _T_19[9:0]) begin
        image_2_428 <= io_pixelVal_in_2_1;
      end else if (10'h1ac == _T_15[9:0]) begin
        image_2_428 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_429 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ad == _T_37[9:0]) begin
        image_2_429 <= io_pixelVal_in_2_7;
      end else if (10'h1ad == _T_34[9:0]) begin
        image_2_429 <= io_pixelVal_in_2_6;
      end else if (10'h1ad == _T_31[9:0]) begin
        image_2_429 <= io_pixelVal_in_2_5;
      end else if (10'h1ad == _T_28[9:0]) begin
        image_2_429 <= io_pixelVal_in_2_4;
      end else if (10'h1ad == _T_25[9:0]) begin
        image_2_429 <= io_pixelVal_in_2_3;
      end else if (10'h1ad == _T_22[9:0]) begin
        image_2_429 <= io_pixelVal_in_2_2;
      end else if (10'h1ad == _T_19[9:0]) begin
        image_2_429 <= io_pixelVal_in_2_1;
      end else if (10'h1ad == _T_15[9:0]) begin
        image_2_429 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_430 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ae == _T_37[9:0]) begin
        image_2_430 <= io_pixelVal_in_2_7;
      end else if (10'h1ae == _T_34[9:0]) begin
        image_2_430 <= io_pixelVal_in_2_6;
      end else if (10'h1ae == _T_31[9:0]) begin
        image_2_430 <= io_pixelVal_in_2_5;
      end else if (10'h1ae == _T_28[9:0]) begin
        image_2_430 <= io_pixelVal_in_2_4;
      end else if (10'h1ae == _T_25[9:0]) begin
        image_2_430 <= io_pixelVal_in_2_3;
      end else if (10'h1ae == _T_22[9:0]) begin
        image_2_430 <= io_pixelVal_in_2_2;
      end else if (10'h1ae == _T_19[9:0]) begin
        image_2_430 <= io_pixelVal_in_2_1;
      end else if (10'h1ae == _T_15[9:0]) begin
        image_2_430 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_431 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1af == _T_37[9:0]) begin
        image_2_431 <= io_pixelVal_in_2_7;
      end else if (10'h1af == _T_34[9:0]) begin
        image_2_431 <= io_pixelVal_in_2_6;
      end else if (10'h1af == _T_31[9:0]) begin
        image_2_431 <= io_pixelVal_in_2_5;
      end else if (10'h1af == _T_28[9:0]) begin
        image_2_431 <= io_pixelVal_in_2_4;
      end else if (10'h1af == _T_25[9:0]) begin
        image_2_431 <= io_pixelVal_in_2_3;
      end else if (10'h1af == _T_22[9:0]) begin
        image_2_431 <= io_pixelVal_in_2_2;
      end else if (10'h1af == _T_19[9:0]) begin
        image_2_431 <= io_pixelVal_in_2_1;
      end else if (10'h1af == _T_15[9:0]) begin
        image_2_431 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_432 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b0 == _T_37[9:0]) begin
        image_2_432 <= io_pixelVal_in_2_7;
      end else if (10'h1b0 == _T_34[9:0]) begin
        image_2_432 <= io_pixelVal_in_2_6;
      end else if (10'h1b0 == _T_31[9:0]) begin
        image_2_432 <= io_pixelVal_in_2_5;
      end else if (10'h1b0 == _T_28[9:0]) begin
        image_2_432 <= io_pixelVal_in_2_4;
      end else if (10'h1b0 == _T_25[9:0]) begin
        image_2_432 <= io_pixelVal_in_2_3;
      end else if (10'h1b0 == _T_22[9:0]) begin
        image_2_432 <= io_pixelVal_in_2_2;
      end else if (10'h1b0 == _T_19[9:0]) begin
        image_2_432 <= io_pixelVal_in_2_1;
      end else if (10'h1b0 == _T_15[9:0]) begin
        image_2_432 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_433 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b1 == _T_37[9:0]) begin
        image_2_433 <= io_pixelVal_in_2_7;
      end else if (10'h1b1 == _T_34[9:0]) begin
        image_2_433 <= io_pixelVal_in_2_6;
      end else if (10'h1b1 == _T_31[9:0]) begin
        image_2_433 <= io_pixelVal_in_2_5;
      end else if (10'h1b1 == _T_28[9:0]) begin
        image_2_433 <= io_pixelVal_in_2_4;
      end else if (10'h1b1 == _T_25[9:0]) begin
        image_2_433 <= io_pixelVal_in_2_3;
      end else if (10'h1b1 == _T_22[9:0]) begin
        image_2_433 <= io_pixelVal_in_2_2;
      end else if (10'h1b1 == _T_19[9:0]) begin
        image_2_433 <= io_pixelVal_in_2_1;
      end else if (10'h1b1 == _T_15[9:0]) begin
        image_2_433 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_434 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b2 == _T_37[9:0]) begin
        image_2_434 <= io_pixelVal_in_2_7;
      end else if (10'h1b2 == _T_34[9:0]) begin
        image_2_434 <= io_pixelVal_in_2_6;
      end else if (10'h1b2 == _T_31[9:0]) begin
        image_2_434 <= io_pixelVal_in_2_5;
      end else if (10'h1b2 == _T_28[9:0]) begin
        image_2_434 <= io_pixelVal_in_2_4;
      end else if (10'h1b2 == _T_25[9:0]) begin
        image_2_434 <= io_pixelVal_in_2_3;
      end else if (10'h1b2 == _T_22[9:0]) begin
        image_2_434 <= io_pixelVal_in_2_2;
      end else if (10'h1b2 == _T_19[9:0]) begin
        image_2_434 <= io_pixelVal_in_2_1;
      end else if (10'h1b2 == _T_15[9:0]) begin
        image_2_434 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_435 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b3 == _T_37[9:0]) begin
        image_2_435 <= io_pixelVal_in_2_7;
      end else if (10'h1b3 == _T_34[9:0]) begin
        image_2_435 <= io_pixelVal_in_2_6;
      end else if (10'h1b3 == _T_31[9:0]) begin
        image_2_435 <= io_pixelVal_in_2_5;
      end else if (10'h1b3 == _T_28[9:0]) begin
        image_2_435 <= io_pixelVal_in_2_4;
      end else if (10'h1b3 == _T_25[9:0]) begin
        image_2_435 <= io_pixelVal_in_2_3;
      end else if (10'h1b3 == _T_22[9:0]) begin
        image_2_435 <= io_pixelVal_in_2_2;
      end else if (10'h1b3 == _T_19[9:0]) begin
        image_2_435 <= io_pixelVal_in_2_1;
      end else if (10'h1b3 == _T_15[9:0]) begin
        image_2_435 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_436 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b4 == _T_37[9:0]) begin
        image_2_436 <= io_pixelVal_in_2_7;
      end else if (10'h1b4 == _T_34[9:0]) begin
        image_2_436 <= io_pixelVal_in_2_6;
      end else if (10'h1b4 == _T_31[9:0]) begin
        image_2_436 <= io_pixelVal_in_2_5;
      end else if (10'h1b4 == _T_28[9:0]) begin
        image_2_436 <= io_pixelVal_in_2_4;
      end else if (10'h1b4 == _T_25[9:0]) begin
        image_2_436 <= io_pixelVal_in_2_3;
      end else if (10'h1b4 == _T_22[9:0]) begin
        image_2_436 <= io_pixelVal_in_2_2;
      end else if (10'h1b4 == _T_19[9:0]) begin
        image_2_436 <= io_pixelVal_in_2_1;
      end else if (10'h1b4 == _T_15[9:0]) begin
        image_2_436 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_437 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b5 == _T_37[9:0]) begin
        image_2_437 <= io_pixelVal_in_2_7;
      end else if (10'h1b5 == _T_34[9:0]) begin
        image_2_437 <= io_pixelVal_in_2_6;
      end else if (10'h1b5 == _T_31[9:0]) begin
        image_2_437 <= io_pixelVal_in_2_5;
      end else if (10'h1b5 == _T_28[9:0]) begin
        image_2_437 <= io_pixelVal_in_2_4;
      end else if (10'h1b5 == _T_25[9:0]) begin
        image_2_437 <= io_pixelVal_in_2_3;
      end else if (10'h1b5 == _T_22[9:0]) begin
        image_2_437 <= io_pixelVal_in_2_2;
      end else if (10'h1b5 == _T_19[9:0]) begin
        image_2_437 <= io_pixelVal_in_2_1;
      end else if (10'h1b5 == _T_15[9:0]) begin
        image_2_437 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_438 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b6 == _T_37[9:0]) begin
        image_2_438 <= io_pixelVal_in_2_7;
      end else if (10'h1b6 == _T_34[9:0]) begin
        image_2_438 <= io_pixelVal_in_2_6;
      end else if (10'h1b6 == _T_31[9:0]) begin
        image_2_438 <= io_pixelVal_in_2_5;
      end else if (10'h1b6 == _T_28[9:0]) begin
        image_2_438 <= io_pixelVal_in_2_4;
      end else if (10'h1b6 == _T_25[9:0]) begin
        image_2_438 <= io_pixelVal_in_2_3;
      end else if (10'h1b6 == _T_22[9:0]) begin
        image_2_438 <= io_pixelVal_in_2_2;
      end else if (10'h1b6 == _T_19[9:0]) begin
        image_2_438 <= io_pixelVal_in_2_1;
      end else if (10'h1b6 == _T_15[9:0]) begin
        image_2_438 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_439 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b7 == _T_37[9:0]) begin
        image_2_439 <= io_pixelVal_in_2_7;
      end else if (10'h1b7 == _T_34[9:0]) begin
        image_2_439 <= io_pixelVal_in_2_6;
      end else if (10'h1b7 == _T_31[9:0]) begin
        image_2_439 <= io_pixelVal_in_2_5;
      end else if (10'h1b7 == _T_28[9:0]) begin
        image_2_439 <= io_pixelVal_in_2_4;
      end else if (10'h1b7 == _T_25[9:0]) begin
        image_2_439 <= io_pixelVal_in_2_3;
      end else if (10'h1b7 == _T_22[9:0]) begin
        image_2_439 <= io_pixelVal_in_2_2;
      end else if (10'h1b7 == _T_19[9:0]) begin
        image_2_439 <= io_pixelVal_in_2_1;
      end else if (10'h1b7 == _T_15[9:0]) begin
        image_2_439 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_440 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b8 == _T_37[9:0]) begin
        image_2_440 <= io_pixelVal_in_2_7;
      end else if (10'h1b8 == _T_34[9:0]) begin
        image_2_440 <= io_pixelVal_in_2_6;
      end else if (10'h1b8 == _T_31[9:0]) begin
        image_2_440 <= io_pixelVal_in_2_5;
      end else if (10'h1b8 == _T_28[9:0]) begin
        image_2_440 <= io_pixelVal_in_2_4;
      end else if (10'h1b8 == _T_25[9:0]) begin
        image_2_440 <= io_pixelVal_in_2_3;
      end else if (10'h1b8 == _T_22[9:0]) begin
        image_2_440 <= io_pixelVal_in_2_2;
      end else if (10'h1b8 == _T_19[9:0]) begin
        image_2_440 <= io_pixelVal_in_2_1;
      end else if (10'h1b8 == _T_15[9:0]) begin
        image_2_440 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_441 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b9 == _T_37[9:0]) begin
        image_2_441 <= io_pixelVal_in_2_7;
      end else if (10'h1b9 == _T_34[9:0]) begin
        image_2_441 <= io_pixelVal_in_2_6;
      end else if (10'h1b9 == _T_31[9:0]) begin
        image_2_441 <= io_pixelVal_in_2_5;
      end else if (10'h1b9 == _T_28[9:0]) begin
        image_2_441 <= io_pixelVal_in_2_4;
      end else if (10'h1b9 == _T_25[9:0]) begin
        image_2_441 <= io_pixelVal_in_2_3;
      end else if (10'h1b9 == _T_22[9:0]) begin
        image_2_441 <= io_pixelVal_in_2_2;
      end else if (10'h1b9 == _T_19[9:0]) begin
        image_2_441 <= io_pixelVal_in_2_1;
      end else if (10'h1b9 == _T_15[9:0]) begin
        image_2_441 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_442 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ba == _T_37[9:0]) begin
        image_2_442 <= io_pixelVal_in_2_7;
      end else if (10'h1ba == _T_34[9:0]) begin
        image_2_442 <= io_pixelVal_in_2_6;
      end else if (10'h1ba == _T_31[9:0]) begin
        image_2_442 <= io_pixelVal_in_2_5;
      end else if (10'h1ba == _T_28[9:0]) begin
        image_2_442 <= io_pixelVal_in_2_4;
      end else if (10'h1ba == _T_25[9:0]) begin
        image_2_442 <= io_pixelVal_in_2_3;
      end else if (10'h1ba == _T_22[9:0]) begin
        image_2_442 <= io_pixelVal_in_2_2;
      end else if (10'h1ba == _T_19[9:0]) begin
        image_2_442 <= io_pixelVal_in_2_1;
      end else if (10'h1ba == _T_15[9:0]) begin
        image_2_442 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_443 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1bb == _T_37[9:0]) begin
        image_2_443 <= io_pixelVal_in_2_7;
      end else if (10'h1bb == _T_34[9:0]) begin
        image_2_443 <= io_pixelVal_in_2_6;
      end else if (10'h1bb == _T_31[9:0]) begin
        image_2_443 <= io_pixelVal_in_2_5;
      end else if (10'h1bb == _T_28[9:0]) begin
        image_2_443 <= io_pixelVal_in_2_4;
      end else if (10'h1bb == _T_25[9:0]) begin
        image_2_443 <= io_pixelVal_in_2_3;
      end else if (10'h1bb == _T_22[9:0]) begin
        image_2_443 <= io_pixelVal_in_2_2;
      end else if (10'h1bb == _T_19[9:0]) begin
        image_2_443 <= io_pixelVal_in_2_1;
      end else if (10'h1bb == _T_15[9:0]) begin
        image_2_443 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_444 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1bc == _T_37[9:0]) begin
        image_2_444 <= io_pixelVal_in_2_7;
      end else if (10'h1bc == _T_34[9:0]) begin
        image_2_444 <= io_pixelVal_in_2_6;
      end else if (10'h1bc == _T_31[9:0]) begin
        image_2_444 <= io_pixelVal_in_2_5;
      end else if (10'h1bc == _T_28[9:0]) begin
        image_2_444 <= io_pixelVal_in_2_4;
      end else if (10'h1bc == _T_25[9:0]) begin
        image_2_444 <= io_pixelVal_in_2_3;
      end else if (10'h1bc == _T_22[9:0]) begin
        image_2_444 <= io_pixelVal_in_2_2;
      end else if (10'h1bc == _T_19[9:0]) begin
        image_2_444 <= io_pixelVal_in_2_1;
      end else if (10'h1bc == _T_15[9:0]) begin
        image_2_444 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_445 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1bd == _T_37[9:0]) begin
        image_2_445 <= io_pixelVal_in_2_7;
      end else if (10'h1bd == _T_34[9:0]) begin
        image_2_445 <= io_pixelVal_in_2_6;
      end else if (10'h1bd == _T_31[9:0]) begin
        image_2_445 <= io_pixelVal_in_2_5;
      end else if (10'h1bd == _T_28[9:0]) begin
        image_2_445 <= io_pixelVal_in_2_4;
      end else if (10'h1bd == _T_25[9:0]) begin
        image_2_445 <= io_pixelVal_in_2_3;
      end else if (10'h1bd == _T_22[9:0]) begin
        image_2_445 <= io_pixelVal_in_2_2;
      end else if (10'h1bd == _T_19[9:0]) begin
        image_2_445 <= io_pixelVal_in_2_1;
      end else if (10'h1bd == _T_15[9:0]) begin
        image_2_445 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_446 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1be == _T_37[9:0]) begin
        image_2_446 <= io_pixelVal_in_2_7;
      end else if (10'h1be == _T_34[9:0]) begin
        image_2_446 <= io_pixelVal_in_2_6;
      end else if (10'h1be == _T_31[9:0]) begin
        image_2_446 <= io_pixelVal_in_2_5;
      end else if (10'h1be == _T_28[9:0]) begin
        image_2_446 <= io_pixelVal_in_2_4;
      end else if (10'h1be == _T_25[9:0]) begin
        image_2_446 <= io_pixelVal_in_2_3;
      end else if (10'h1be == _T_22[9:0]) begin
        image_2_446 <= io_pixelVal_in_2_2;
      end else if (10'h1be == _T_19[9:0]) begin
        image_2_446 <= io_pixelVal_in_2_1;
      end else if (10'h1be == _T_15[9:0]) begin
        image_2_446 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_447 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1bf == _T_37[9:0]) begin
        image_2_447 <= io_pixelVal_in_2_7;
      end else if (10'h1bf == _T_34[9:0]) begin
        image_2_447 <= io_pixelVal_in_2_6;
      end else if (10'h1bf == _T_31[9:0]) begin
        image_2_447 <= io_pixelVal_in_2_5;
      end else if (10'h1bf == _T_28[9:0]) begin
        image_2_447 <= io_pixelVal_in_2_4;
      end else if (10'h1bf == _T_25[9:0]) begin
        image_2_447 <= io_pixelVal_in_2_3;
      end else if (10'h1bf == _T_22[9:0]) begin
        image_2_447 <= io_pixelVal_in_2_2;
      end else if (10'h1bf == _T_19[9:0]) begin
        image_2_447 <= io_pixelVal_in_2_1;
      end else if (10'h1bf == _T_15[9:0]) begin
        image_2_447 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_448 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c0 == _T_37[9:0]) begin
        image_2_448 <= io_pixelVal_in_2_7;
      end else if (10'h1c0 == _T_34[9:0]) begin
        image_2_448 <= io_pixelVal_in_2_6;
      end else if (10'h1c0 == _T_31[9:0]) begin
        image_2_448 <= io_pixelVal_in_2_5;
      end else if (10'h1c0 == _T_28[9:0]) begin
        image_2_448 <= io_pixelVal_in_2_4;
      end else if (10'h1c0 == _T_25[9:0]) begin
        image_2_448 <= io_pixelVal_in_2_3;
      end else if (10'h1c0 == _T_22[9:0]) begin
        image_2_448 <= io_pixelVal_in_2_2;
      end else if (10'h1c0 == _T_19[9:0]) begin
        image_2_448 <= io_pixelVal_in_2_1;
      end else if (10'h1c0 == _T_15[9:0]) begin
        image_2_448 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_449 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c1 == _T_37[9:0]) begin
        image_2_449 <= io_pixelVal_in_2_7;
      end else if (10'h1c1 == _T_34[9:0]) begin
        image_2_449 <= io_pixelVal_in_2_6;
      end else if (10'h1c1 == _T_31[9:0]) begin
        image_2_449 <= io_pixelVal_in_2_5;
      end else if (10'h1c1 == _T_28[9:0]) begin
        image_2_449 <= io_pixelVal_in_2_4;
      end else if (10'h1c1 == _T_25[9:0]) begin
        image_2_449 <= io_pixelVal_in_2_3;
      end else if (10'h1c1 == _T_22[9:0]) begin
        image_2_449 <= io_pixelVal_in_2_2;
      end else if (10'h1c1 == _T_19[9:0]) begin
        image_2_449 <= io_pixelVal_in_2_1;
      end else if (10'h1c1 == _T_15[9:0]) begin
        image_2_449 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_450 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c2 == _T_37[9:0]) begin
        image_2_450 <= io_pixelVal_in_2_7;
      end else if (10'h1c2 == _T_34[9:0]) begin
        image_2_450 <= io_pixelVal_in_2_6;
      end else if (10'h1c2 == _T_31[9:0]) begin
        image_2_450 <= io_pixelVal_in_2_5;
      end else if (10'h1c2 == _T_28[9:0]) begin
        image_2_450 <= io_pixelVal_in_2_4;
      end else if (10'h1c2 == _T_25[9:0]) begin
        image_2_450 <= io_pixelVal_in_2_3;
      end else if (10'h1c2 == _T_22[9:0]) begin
        image_2_450 <= io_pixelVal_in_2_2;
      end else if (10'h1c2 == _T_19[9:0]) begin
        image_2_450 <= io_pixelVal_in_2_1;
      end else if (10'h1c2 == _T_15[9:0]) begin
        image_2_450 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_451 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c3 == _T_37[9:0]) begin
        image_2_451 <= io_pixelVal_in_2_7;
      end else if (10'h1c3 == _T_34[9:0]) begin
        image_2_451 <= io_pixelVal_in_2_6;
      end else if (10'h1c3 == _T_31[9:0]) begin
        image_2_451 <= io_pixelVal_in_2_5;
      end else if (10'h1c3 == _T_28[9:0]) begin
        image_2_451 <= io_pixelVal_in_2_4;
      end else if (10'h1c3 == _T_25[9:0]) begin
        image_2_451 <= io_pixelVal_in_2_3;
      end else if (10'h1c3 == _T_22[9:0]) begin
        image_2_451 <= io_pixelVal_in_2_2;
      end else if (10'h1c3 == _T_19[9:0]) begin
        image_2_451 <= io_pixelVal_in_2_1;
      end else if (10'h1c3 == _T_15[9:0]) begin
        image_2_451 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_452 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c4 == _T_37[9:0]) begin
        image_2_452 <= io_pixelVal_in_2_7;
      end else if (10'h1c4 == _T_34[9:0]) begin
        image_2_452 <= io_pixelVal_in_2_6;
      end else if (10'h1c4 == _T_31[9:0]) begin
        image_2_452 <= io_pixelVal_in_2_5;
      end else if (10'h1c4 == _T_28[9:0]) begin
        image_2_452 <= io_pixelVal_in_2_4;
      end else if (10'h1c4 == _T_25[9:0]) begin
        image_2_452 <= io_pixelVal_in_2_3;
      end else if (10'h1c4 == _T_22[9:0]) begin
        image_2_452 <= io_pixelVal_in_2_2;
      end else if (10'h1c4 == _T_19[9:0]) begin
        image_2_452 <= io_pixelVal_in_2_1;
      end else if (10'h1c4 == _T_15[9:0]) begin
        image_2_452 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_453 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c5 == _T_37[9:0]) begin
        image_2_453 <= io_pixelVal_in_2_7;
      end else if (10'h1c5 == _T_34[9:0]) begin
        image_2_453 <= io_pixelVal_in_2_6;
      end else if (10'h1c5 == _T_31[9:0]) begin
        image_2_453 <= io_pixelVal_in_2_5;
      end else if (10'h1c5 == _T_28[9:0]) begin
        image_2_453 <= io_pixelVal_in_2_4;
      end else if (10'h1c5 == _T_25[9:0]) begin
        image_2_453 <= io_pixelVal_in_2_3;
      end else if (10'h1c5 == _T_22[9:0]) begin
        image_2_453 <= io_pixelVal_in_2_2;
      end else if (10'h1c5 == _T_19[9:0]) begin
        image_2_453 <= io_pixelVal_in_2_1;
      end else if (10'h1c5 == _T_15[9:0]) begin
        image_2_453 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_454 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c6 == _T_37[9:0]) begin
        image_2_454 <= io_pixelVal_in_2_7;
      end else if (10'h1c6 == _T_34[9:0]) begin
        image_2_454 <= io_pixelVal_in_2_6;
      end else if (10'h1c6 == _T_31[9:0]) begin
        image_2_454 <= io_pixelVal_in_2_5;
      end else if (10'h1c6 == _T_28[9:0]) begin
        image_2_454 <= io_pixelVal_in_2_4;
      end else if (10'h1c6 == _T_25[9:0]) begin
        image_2_454 <= io_pixelVal_in_2_3;
      end else if (10'h1c6 == _T_22[9:0]) begin
        image_2_454 <= io_pixelVal_in_2_2;
      end else if (10'h1c6 == _T_19[9:0]) begin
        image_2_454 <= io_pixelVal_in_2_1;
      end else if (10'h1c6 == _T_15[9:0]) begin
        image_2_454 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_455 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c7 == _T_37[9:0]) begin
        image_2_455 <= io_pixelVal_in_2_7;
      end else if (10'h1c7 == _T_34[9:0]) begin
        image_2_455 <= io_pixelVal_in_2_6;
      end else if (10'h1c7 == _T_31[9:0]) begin
        image_2_455 <= io_pixelVal_in_2_5;
      end else if (10'h1c7 == _T_28[9:0]) begin
        image_2_455 <= io_pixelVal_in_2_4;
      end else if (10'h1c7 == _T_25[9:0]) begin
        image_2_455 <= io_pixelVal_in_2_3;
      end else if (10'h1c7 == _T_22[9:0]) begin
        image_2_455 <= io_pixelVal_in_2_2;
      end else if (10'h1c7 == _T_19[9:0]) begin
        image_2_455 <= io_pixelVal_in_2_1;
      end else if (10'h1c7 == _T_15[9:0]) begin
        image_2_455 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_456 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c8 == _T_37[9:0]) begin
        image_2_456 <= io_pixelVal_in_2_7;
      end else if (10'h1c8 == _T_34[9:0]) begin
        image_2_456 <= io_pixelVal_in_2_6;
      end else if (10'h1c8 == _T_31[9:0]) begin
        image_2_456 <= io_pixelVal_in_2_5;
      end else if (10'h1c8 == _T_28[9:0]) begin
        image_2_456 <= io_pixelVal_in_2_4;
      end else if (10'h1c8 == _T_25[9:0]) begin
        image_2_456 <= io_pixelVal_in_2_3;
      end else if (10'h1c8 == _T_22[9:0]) begin
        image_2_456 <= io_pixelVal_in_2_2;
      end else if (10'h1c8 == _T_19[9:0]) begin
        image_2_456 <= io_pixelVal_in_2_1;
      end else if (10'h1c8 == _T_15[9:0]) begin
        image_2_456 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_457 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c9 == _T_37[9:0]) begin
        image_2_457 <= io_pixelVal_in_2_7;
      end else if (10'h1c9 == _T_34[9:0]) begin
        image_2_457 <= io_pixelVal_in_2_6;
      end else if (10'h1c9 == _T_31[9:0]) begin
        image_2_457 <= io_pixelVal_in_2_5;
      end else if (10'h1c9 == _T_28[9:0]) begin
        image_2_457 <= io_pixelVal_in_2_4;
      end else if (10'h1c9 == _T_25[9:0]) begin
        image_2_457 <= io_pixelVal_in_2_3;
      end else if (10'h1c9 == _T_22[9:0]) begin
        image_2_457 <= io_pixelVal_in_2_2;
      end else if (10'h1c9 == _T_19[9:0]) begin
        image_2_457 <= io_pixelVal_in_2_1;
      end else if (10'h1c9 == _T_15[9:0]) begin
        image_2_457 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_458 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ca == _T_37[9:0]) begin
        image_2_458 <= io_pixelVal_in_2_7;
      end else if (10'h1ca == _T_34[9:0]) begin
        image_2_458 <= io_pixelVal_in_2_6;
      end else if (10'h1ca == _T_31[9:0]) begin
        image_2_458 <= io_pixelVal_in_2_5;
      end else if (10'h1ca == _T_28[9:0]) begin
        image_2_458 <= io_pixelVal_in_2_4;
      end else if (10'h1ca == _T_25[9:0]) begin
        image_2_458 <= io_pixelVal_in_2_3;
      end else if (10'h1ca == _T_22[9:0]) begin
        image_2_458 <= io_pixelVal_in_2_2;
      end else if (10'h1ca == _T_19[9:0]) begin
        image_2_458 <= io_pixelVal_in_2_1;
      end else if (10'h1ca == _T_15[9:0]) begin
        image_2_458 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_459 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1cb == _T_37[9:0]) begin
        image_2_459 <= io_pixelVal_in_2_7;
      end else if (10'h1cb == _T_34[9:0]) begin
        image_2_459 <= io_pixelVal_in_2_6;
      end else if (10'h1cb == _T_31[9:0]) begin
        image_2_459 <= io_pixelVal_in_2_5;
      end else if (10'h1cb == _T_28[9:0]) begin
        image_2_459 <= io_pixelVal_in_2_4;
      end else if (10'h1cb == _T_25[9:0]) begin
        image_2_459 <= io_pixelVal_in_2_3;
      end else if (10'h1cb == _T_22[9:0]) begin
        image_2_459 <= io_pixelVal_in_2_2;
      end else if (10'h1cb == _T_19[9:0]) begin
        image_2_459 <= io_pixelVal_in_2_1;
      end else if (10'h1cb == _T_15[9:0]) begin
        image_2_459 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_460 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1cc == _T_37[9:0]) begin
        image_2_460 <= io_pixelVal_in_2_7;
      end else if (10'h1cc == _T_34[9:0]) begin
        image_2_460 <= io_pixelVal_in_2_6;
      end else if (10'h1cc == _T_31[9:0]) begin
        image_2_460 <= io_pixelVal_in_2_5;
      end else if (10'h1cc == _T_28[9:0]) begin
        image_2_460 <= io_pixelVal_in_2_4;
      end else if (10'h1cc == _T_25[9:0]) begin
        image_2_460 <= io_pixelVal_in_2_3;
      end else if (10'h1cc == _T_22[9:0]) begin
        image_2_460 <= io_pixelVal_in_2_2;
      end else if (10'h1cc == _T_19[9:0]) begin
        image_2_460 <= io_pixelVal_in_2_1;
      end else if (10'h1cc == _T_15[9:0]) begin
        image_2_460 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_461 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1cd == _T_37[9:0]) begin
        image_2_461 <= io_pixelVal_in_2_7;
      end else if (10'h1cd == _T_34[9:0]) begin
        image_2_461 <= io_pixelVal_in_2_6;
      end else if (10'h1cd == _T_31[9:0]) begin
        image_2_461 <= io_pixelVal_in_2_5;
      end else if (10'h1cd == _T_28[9:0]) begin
        image_2_461 <= io_pixelVal_in_2_4;
      end else if (10'h1cd == _T_25[9:0]) begin
        image_2_461 <= io_pixelVal_in_2_3;
      end else if (10'h1cd == _T_22[9:0]) begin
        image_2_461 <= io_pixelVal_in_2_2;
      end else if (10'h1cd == _T_19[9:0]) begin
        image_2_461 <= io_pixelVal_in_2_1;
      end else if (10'h1cd == _T_15[9:0]) begin
        image_2_461 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_462 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ce == _T_37[9:0]) begin
        image_2_462 <= io_pixelVal_in_2_7;
      end else if (10'h1ce == _T_34[9:0]) begin
        image_2_462 <= io_pixelVal_in_2_6;
      end else if (10'h1ce == _T_31[9:0]) begin
        image_2_462 <= io_pixelVal_in_2_5;
      end else if (10'h1ce == _T_28[9:0]) begin
        image_2_462 <= io_pixelVal_in_2_4;
      end else if (10'h1ce == _T_25[9:0]) begin
        image_2_462 <= io_pixelVal_in_2_3;
      end else if (10'h1ce == _T_22[9:0]) begin
        image_2_462 <= io_pixelVal_in_2_2;
      end else if (10'h1ce == _T_19[9:0]) begin
        image_2_462 <= io_pixelVal_in_2_1;
      end else if (10'h1ce == _T_15[9:0]) begin
        image_2_462 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_463 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1cf == _T_37[9:0]) begin
        image_2_463 <= io_pixelVal_in_2_7;
      end else if (10'h1cf == _T_34[9:0]) begin
        image_2_463 <= io_pixelVal_in_2_6;
      end else if (10'h1cf == _T_31[9:0]) begin
        image_2_463 <= io_pixelVal_in_2_5;
      end else if (10'h1cf == _T_28[9:0]) begin
        image_2_463 <= io_pixelVal_in_2_4;
      end else if (10'h1cf == _T_25[9:0]) begin
        image_2_463 <= io_pixelVal_in_2_3;
      end else if (10'h1cf == _T_22[9:0]) begin
        image_2_463 <= io_pixelVal_in_2_2;
      end else if (10'h1cf == _T_19[9:0]) begin
        image_2_463 <= io_pixelVal_in_2_1;
      end else if (10'h1cf == _T_15[9:0]) begin
        image_2_463 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_464 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d0 == _T_37[9:0]) begin
        image_2_464 <= io_pixelVal_in_2_7;
      end else if (10'h1d0 == _T_34[9:0]) begin
        image_2_464 <= io_pixelVal_in_2_6;
      end else if (10'h1d0 == _T_31[9:0]) begin
        image_2_464 <= io_pixelVal_in_2_5;
      end else if (10'h1d0 == _T_28[9:0]) begin
        image_2_464 <= io_pixelVal_in_2_4;
      end else if (10'h1d0 == _T_25[9:0]) begin
        image_2_464 <= io_pixelVal_in_2_3;
      end else if (10'h1d0 == _T_22[9:0]) begin
        image_2_464 <= io_pixelVal_in_2_2;
      end else if (10'h1d0 == _T_19[9:0]) begin
        image_2_464 <= io_pixelVal_in_2_1;
      end else if (10'h1d0 == _T_15[9:0]) begin
        image_2_464 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_465 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d1 == _T_37[9:0]) begin
        image_2_465 <= io_pixelVal_in_2_7;
      end else if (10'h1d1 == _T_34[9:0]) begin
        image_2_465 <= io_pixelVal_in_2_6;
      end else if (10'h1d1 == _T_31[9:0]) begin
        image_2_465 <= io_pixelVal_in_2_5;
      end else if (10'h1d1 == _T_28[9:0]) begin
        image_2_465 <= io_pixelVal_in_2_4;
      end else if (10'h1d1 == _T_25[9:0]) begin
        image_2_465 <= io_pixelVal_in_2_3;
      end else if (10'h1d1 == _T_22[9:0]) begin
        image_2_465 <= io_pixelVal_in_2_2;
      end else if (10'h1d1 == _T_19[9:0]) begin
        image_2_465 <= io_pixelVal_in_2_1;
      end else if (10'h1d1 == _T_15[9:0]) begin
        image_2_465 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_466 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d2 == _T_37[9:0]) begin
        image_2_466 <= io_pixelVal_in_2_7;
      end else if (10'h1d2 == _T_34[9:0]) begin
        image_2_466 <= io_pixelVal_in_2_6;
      end else if (10'h1d2 == _T_31[9:0]) begin
        image_2_466 <= io_pixelVal_in_2_5;
      end else if (10'h1d2 == _T_28[9:0]) begin
        image_2_466 <= io_pixelVal_in_2_4;
      end else if (10'h1d2 == _T_25[9:0]) begin
        image_2_466 <= io_pixelVal_in_2_3;
      end else if (10'h1d2 == _T_22[9:0]) begin
        image_2_466 <= io_pixelVal_in_2_2;
      end else if (10'h1d2 == _T_19[9:0]) begin
        image_2_466 <= io_pixelVal_in_2_1;
      end else if (10'h1d2 == _T_15[9:0]) begin
        image_2_466 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_467 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d3 == _T_37[9:0]) begin
        image_2_467 <= io_pixelVal_in_2_7;
      end else if (10'h1d3 == _T_34[9:0]) begin
        image_2_467 <= io_pixelVal_in_2_6;
      end else if (10'h1d3 == _T_31[9:0]) begin
        image_2_467 <= io_pixelVal_in_2_5;
      end else if (10'h1d3 == _T_28[9:0]) begin
        image_2_467 <= io_pixelVal_in_2_4;
      end else if (10'h1d3 == _T_25[9:0]) begin
        image_2_467 <= io_pixelVal_in_2_3;
      end else if (10'h1d3 == _T_22[9:0]) begin
        image_2_467 <= io_pixelVal_in_2_2;
      end else if (10'h1d3 == _T_19[9:0]) begin
        image_2_467 <= io_pixelVal_in_2_1;
      end else if (10'h1d3 == _T_15[9:0]) begin
        image_2_467 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_468 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d4 == _T_37[9:0]) begin
        image_2_468 <= io_pixelVal_in_2_7;
      end else if (10'h1d4 == _T_34[9:0]) begin
        image_2_468 <= io_pixelVal_in_2_6;
      end else if (10'h1d4 == _T_31[9:0]) begin
        image_2_468 <= io_pixelVal_in_2_5;
      end else if (10'h1d4 == _T_28[9:0]) begin
        image_2_468 <= io_pixelVal_in_2_4;
      end else if (10'h1d4 == _T_25[9:0]) begin
        image_2_468 <= io_pixelVal_in_2_3;
      end else if (10'h1d4 == _T_22[9:0]) begin
        image_2_468 <= io_pixelVal_in_2_2;
      end else if (10'h1d4 == _T_19[9:0]) begin
        image_2_468 <= io_pixelVal_in_2_1;
      end else if (10'h1d4 == _T_15[9:0]) begin
        image_2_468 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_469 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d5 == _T_37[9:0]) begin
        image_2_469 <= io_pixelVal_in_2_7;
      end else if (10'h1d5 == _T_34[9:0]) begin
        image_2_469 <= io_pixelVal_in_2_6;
      end else if (10'h1d5 == _T_31[9:0]) begin
        image_2_469 <= io_pixelVal_in_2_5;
      end else if (10'h1d5 == _T_28[9:0]) begin
        image_2_469 <= io_pixelVal_in_2_4;
      end else if (10'h1d5 == _T_25[9:0]) begin
        image_2_469 <= io_pixelVal_in_2_3;
      end else if (10'h1d5 == _T_22[9:0]) begin
        image_2_469 <= io_pixelVal_in_2_2;
      end else if (10'h1d5 == _T_19[9:0]) begin
        image_2_469 <= io_pixelVal_in_2_1;
      end else if (10'h1d5 == _T_15[9:0]) begin
        image_2_469 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_470 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d6 == _T_37[9:0]) begin
        image_2_470 <= io_pixelVal_in_2_7;
      end else if (10'h1d6 == _T_34[9:0]) begin
        image_2_470 <= io_pixelVal_in_2_6;
      end else if (10'h1d6 == _T_31[9:0]) begin
        image_2_470 <= io_pixelVal_in_2_5;
      end else if (10'h1d6 == _T_28[9:0]) begin
        image_2_470 <= io_pixelVal_in_2_4;
      end else if (10'h1d6 == _T_25[9:0]) begin
        image_2_470 <= io_pixelVal_in_2_3;
      end else if (10'h1d6 == _T_22[9:0]) begin
        image_2_470 <= io_pixelVal_in_2_2;
      end else if (10'h1d6 == _T_19[9:0]) begin
        image_2_470 <= io_pixelVal_in_2_1;
      end else if (10'h1d6 == _T_15[9:0]) begin
        image_2_470 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_471 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d7 == _T_37[9:0]) begin
        image_2_471 <= io_pixelVal_in_2_7;
      end else if (10'h1d7 == _T_34[9:0]) begin
        image_2_471 <= io_pixelVal_in_2_6;
      end else if (10'h1d7 == _T_31[9:0]) begin
        image_2_471 <= io_pixelVal_in_2_5;
      end else if (10'h1d7 == _T_28[9:0]) begin
        image_2_471 <= io_pixelVal_in_2_4;
      end else if (10'h1d7 == _T_25[9:0]) begin
        image_2_471 <= io_pixelVal_in_2_3;
      end else if (10'h1d7 == _T_22[9:0]) begin
        image_2_471 <= io_pixelVal_in_2_2;
      end else if (10'h1d7 == _T_19[9:0]) begin
        image_2_471 <= io_pixelVal_in_2_1;
      end else if (10'h1d7 == _T_15[9:0]) begin
        image_2_471 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_472 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d8 == _T_37[9:0]) begin
        image_2_472 <= io_pixelVal_in_2_7;
      end else if (10'h1d8 == _T_34[9:0]) begin
        image_2_472 <= io_pixelVal_in_2_6;
      end else if (10'h1d8 == _T_31[9:0]) begin
        image_2_472 <= io_pixelVal_in_2_5;
      end else if (10'h1d8 == _T_28[9:0]) begin
        image_2_472 <= io_pixelVal_in_2_4;
      end else if (10'h1d8 == _T_25[9:0]) begin
        image_2_472 <= io_pixelVal_in_2_3;
      end else if (10'h1d8 == _T_22[9:0]) begin
        image_2_472 <= io_pixelVal_in_2_2;
      end else if (10'h1d8 == _T_19[9:0]) begin
        image_2_472 <= io_pixelVal_in_2_1;
      end else if (10'h1d8 == _T_15[9:0]) begin
        image_2_472 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_473 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d9 == _T_37[9:0]) begin
        image_2_473 <= io_pixelVal_in_2_7;
      end else if (10'h1d9 == _T_34[9:0]) begin
        image_2_473 <= io_pixelVal_in_2_6;
      end else if (10'h1d9 == _T_31[9:0]) begin
        image_2_473 <= io_pixelVal_in_2_5;
      end else if (10'h1d9 == _T_28[9:0]) begin
        image_2_473 <= io_pixelVal_in_2_4;
      end else if (10'h1d9 == _T_25[9:0]) begin
        image_2_473 <= io_pixelVal_in_2_3;
      end else if (10'h1d9 == _T_22[9:0]) begin
        image_2_473 <= io_pixelVal_in_2_2;
      end else if (10'h1d9 == _T_19[9:0]) begin
        image_2_473 <= io_pixelVal_in_2_1;
      end else if (10'h1d9 == _T_15[9:0]) begin
        image_2_473 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_474 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1da == _T_37[9:0]) begin
        image_2_474 <= io_pixelVal_in_2_7;
      end else if (10'h1da == _T_34[9:0]) begin
        image_2_474 <= io_pixelVal_in_2_6;
      end else if (10'h1da == _T_31[9:0]) begin
        image_2_474 <= io_pixelVal_in_2_5;
      end else if (10'h1da == _T_28[9:0]) begin
        image_2_474 <= io_pixelVal_in_2_4;
      end else if (10'h1da == _T_25[9:0]) begin
        image_2_474 <= io_pixelVal_in_2_3;
      end else if (10'h1da == _T_22[9:0]) begin
        image_2_474 <= io_pixelVal_in_2_2;
      end else if (10'h1da == _T_19[9:0]) begin
        image_2_474 <= io_pixelVal_in_2_1;
      end else if (10'h1da == _T_15[9:0]) begin
        image_2_474 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_475 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1db == _T_37[9:0]) begin
        image_2_475 <= io_pixelVal_in_2_7;
      end else if (10'h1db == _T_34[9:0]) begin
        image_2_475 <= io_pixelVal_in_2_6;
      end else if (10'h1db == _T_31[9:0]) begin
        image_2_475 <= io_pixelVal_in_2_5;
      end else if (10'h1db == _T_28[9:0]) begin
        image_2_475 <= io_pixelVal_in_2_4;
      end else if (10'h1db == _T_25[9:0]) begin
        image_2_475 <= io_pixelVal_in_2_3;
      end else if (10'h1db == _T_22[9:0]) begin
        image_2_475 <= io_pixelVal_in_2_2;
      end else if (10'h1db == _T_19[9:0]) begin
        image_2_475 <= io_pixelVal_in_2_1;
      end else if (10'h1db == _T_15[9:0]) begin
        image_2_475 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_476 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1dc == _T_37[9:0]) begin
        image_2_476 <= io_pixelVal_in_2_7;
      end else if (10'h1dc == _T_34[9:0]) begin
        image_2_476 <= io_pixelVal_in_2_6;
      end else if (10'h1dc == _T_31[9:0]) begin
        image_2_476 <= io_pixelVal_in_2_5;
      end else if (10'h1dc == _T_28[9:0]) begin
        image_2_476 <= io_pixelVal_in_2_4;
      end else if (10'h1dc == _T_25[9:0]) begin
        image_2_476 <= io_pixelVal_in_2_3;
      end else if (10'h1dc == _T_22[9:0]) begin
        image_2_476 <= io_pixelVal_in_2_2;
      end else if (10'h1dc == _T_19[9:0]) begin
        image_2_476 <= io_pixelVal_in_2_1;
      end else if (10'h1dc == _T_15[9:0]) begin
        image_2_476 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_477 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1dd == _T_37[9:0]) begin
        image_2_477 <= io_pixelVal_in_2_7;
      end else if (10'h1dd == _T_34[9:0]) begin
        image_2_477 <= io_pixelVal_in_2_6;
      end else if (10'h1dd == _T_31[9:0]) begin
        image_2_477 <= io_pixelVal_in_2_5;
      end else if (10'h1dd == _T_28[9:0]) begin
        image_2_477 <= io_pixelVal_in_2_4;
      end else if (10'h1dd == _T_25[9:0]) begin
        image_2_477 <= io_pixelVal_in_2_3;
      end else if (10'h1dd == _T_22[9:0]) begin
        image_2_477 <= io_pixelVal_in_2_2;
      end else if (10'h1dd == _T_19[9:0]) begin
        image_2_477 <= io_pixelVal_in_2_1;
      end else if (10'h1dd == _T_15[9:0]) begin
        image_2_477 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_478 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1de == _T_37[9:0]) begin
        image_2_478 <= io_pixelVal_in_2_7;
      end else if (10'h1de == _T_34[9:0]) begin
        image_2_478 <= io_pixelVal_in_2_6;
      end else if (10'h1de == _T_31[9:0]) begin
        image_2_478 <= io_pixelVal_in_2_5;
      end else if (10'h1de == _T_28[9:0]) begin
        image_2_478 <= io_pixelVal_in_2_4;
      end else if (10'h1de == _T_25[9:0]) begin
        image_2_478 <= io_pixelVal_in_2_3;
      end else if (10'h1de == _T_22[9:0]) begin
        image_2_478 <= io_pixelVal_in_2_2;
      end else if (10'h1de == _T_19[9:0]) begin
        image_2_478 <= io_pixelVal_in_2_1;
      end else if (10'h1de == _T_15[9:0]) begin
        image_2_478 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_479 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1df == _T_37[9:0]) begin
        image_2_479 <= io_pixelVal_in_2_7;
      end else if (10'h1df == _T_34[9:0]) begin
        image_2_479 <= io_pixelVal_in_2_6;
      end else if (10'h1df == _T_31[9:0]) begin
        image_2_479 <= io_pixelVal_in_2_5;
      end else if (10'h1df == _T_28[9:0]) begin
        image_2_479 <= io_pixelVal_in_2_4;
      end else if (10'h1df == _T_25[9:0]) begin
        image_2_479 <= io_pixelVal_in_2_3;
      end else if (10'h1df == _T_22[9:0]) begin
        image_2_479 <= io_pixelVal_in_2_2;
      end else if (10'h1df == _T_19[9:0]) begin
        image_2_479 <= io_pixelVal_in_2_1;
      end else if (10'h1df == _T_15[9:0]) begin
        image_2_479 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_480 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e0 == _T_37[9:0]) begin
        image_2_480 <= io_pixelVal_in_2_7;
      end else if (10'h1e0 == _T_34[9:0]) begin
        image_2_480 <= io_pixelVal_in_2_6;
      end else if (10'h1e0 == _T_31[9:0]) begin
        image_2_480 <= io_pixelVal_in_2_5;
      end else if (10'h1e0 == _T_28[9:0]) begin
        image_2_480 <= io_pixelVal_in_2_4;
      end else if (10'h1e0 == _T_25[9:0]) begin
        image_2_480 <= io_pixelVal_in_2_3;
      end else if (10'h1e0 == _T_22[9:0]) begin
        image_2_480 <= io_pixelVal_in_2_2;
      end else if (10'h1e0 == _T_19[9:0]) begin
        image_2_480 <= io_pixelVal_in_2_1;
      end else if (10'h1e0 == _T_15[9:0]) begin
        image_2_480 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_481 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e1 == _T_37[9:0]) begin
        image_2_481 <= io_pixelVal_in_2_7;
      end else if (10'h1e1 == _T_34[9:0]) begin
        image_2_481 <= io_pixelVal_in_2_6;
      end else if (10'h1e1 == _T_31[9:0]) begin
        image_2_481 <= io_pixelVal_in_2_5;
      end else if (10'h1e1 == _T_28[9:0]) begin
        image_2_481 <= io_pixelVal_in_2_4;
      end else if (10'h1e1 == _T_25[9:0]) begin
        image_2_481 <= io_pixelVal_in_2_3;
      end else if (10'h1e1 == _T_22[9:0]) begin
        image_2_481 <= io_pixelVal_in_2_2;
      end else if (10'h1e1 == _T_19[9:0]) begin
        image_2_481 <= io_pixelVal_in_2_1;
      end else if (10'h1e1 == _T_15[9:0]) begin
        image_2_481 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_482 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e2 == _T_37[9:0]) begin
        image_2_482 <= io_pixelVal_in_2_7;
      end else if (10'h1e2 == _T_34[9:0]) begin
        image_2_482 <= io_pixelVal_in_2_6;
      end else if (10'h1e2 == _T_31[9:0]) begin
        image_2_482 <= io_pixelVal_in_2_5;
      end else if (10'h1e2 == _T_28[9:0]) begin
        image_2_482 <= io_pixelVal_in_2_4;
      end else if (10'h1e2 == _T_25[9:0]) begin
        image_2_482 <= io_pixelVal_in_2_3;
      end else if (10'h1e2 == _T_22[9:0]) begin
        image_2_482 <= io_pixelVal_in_2_2;
      end else if (10'h1e2 == _T_19[9:0]) begin
        image_2_482 <= io_pixelVal_in_2_1;
      end else if (10'h1e2 == _T_15[9:0]) begin
        image_2_482 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_483 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e3 == _T_37[9:0]) begin
        image_2_483 <= io_pixelVal_in_2_7;
      end else if (10'h1e3 == _T_34[9:0]) begin
        image_2_483 <= io_pixelVal_in_2_6;
      end else if (10'h1e3 == _T_31[9:0]) begin
        image_2_483 <= io_pixelVal_in_2_5;
      end else if (10'h1e3 == _T_28[9:0]) begin
        image_2_483 <= io_pixelVal_in_2_4;
      end else if (10'h1e3 == _T_25[9:0]) begin
        image_2_483 <= io_pixelVal_in_2_3;
      end else if (10'h1e3 == _T_22[9:0]) begin
        image_2_483 <= io_pixelVal_in_2_2;
      end else if (10'h1e3 == _T_19[9:0]) begin
        image_2_483 <= io_pixelVal_in_2_1;
      end else if (10'h1e3 == _T_15[9:0]) begin
        image_2_483 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_484 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e4 == _T_37[9:0]) begin
        image_2_484 <= io_pixelVal_in_2_7;
      end else if (10'h1e4 == _T_34[9:0]) begin
        image_2_484 <= io_pixelVal_in_2_6;
      end else if (10'h1e4 == _T_31[9:0]) begin
        image_2_484 <= io_pixelVal_in_2_5;
      end else if (10'h1e4 == _T_28[9:0]) begin
        image_2_484 <= io_pixelVal_in_2_4;
      end else if (10'h1e4 == _T_25[9:0]) begin
        image_2_484 <= io_pixelVal_in_2_3;
      end else if (10'h1e4 == _T_22[9:0]) begin
        image_2_484 <= io_pixelVal_in_2_2;
      end else if (10'h1e4 == _T_19[9:0]) begin
        image_2_484 <= io_pixelVal_in_2_1;
      end else if (10'h1e4 == _T_15[9:0]) begin
        image_2_484 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_485 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e5 == _T_37[9:0]) begin
        image_2_485 <= io_pixelVal_in_2_7;
      end else if (10'h1e5 == _T_34[9:0]) begin
        image_2_485 <= io_pixelVal_in_2_6;
      end else if (10'h1e5 == _T_31[9:0]) begin
        image_2_485 <= io_pixelVal_in_2_5;
      end else if (10'h1e5 == _T_28[9:0]) begin
        image_2_485 <= io_pixelVal_in_2_4;
      end else if (10'h1e5 == _T_25[9:0]) begin
        image_2_485 <= io_pixelVal_in_2_3;
      end else if (10'h1e5 == _T_22[9:0]) begin
        image_2_485 <= io_pixelVal_in_2_2;
      end else if (10'h1e5 == _T_19[9:0]) begin
        image_2_485 <= io_pixelVal_in_2_1;
      end else if (10'h1e5 == _T_15[9:0]) begin
        image_2_485 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_486 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e6 == _T_37[9:0]) begin
        image_2_486 <= io_pixelVal_in_2_7;
      end else if (10'h1e6 == _T_34[9:0]) begin
        image_2_486 <= io_pixelVal_in_2_6;
      end else if (10'h1e6 == _T_31[9:0]) begin
        image_2_486 <= io_pixelVal_in_2_5;
      end else if (10'h1e6 == _T_28[9:0]) begin
        image_2_486 <= io_pixelVal_in_2_4;
      end else if (10'h1e6 == _T_25[9:0]) begin
        image_2_486 <= io_pixelVal_in_2_3;
      end else if (10'h1e6 == _T_22[9:0]) begin
        image_2_486 <= io_pixelVal_in_2_2;
      end else if (10'h1e6 == _T_19[9:0]) begin
        image_2_486 <= io_pixelVal_in_2_1;
      end else if (10'h1e6 == _T_15[9:0]) begin
        image_2_486 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_487 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e7 == _T_37[9:0]) begin
        image_2_487 <= io_pixelVal_in_2_7;
      end else if (10'h1e7 == _T_34[9:0]) begin
        image_2_487 <= io_pixelVal_in_2_6;
      end else if (10'h1e7 == _T_31[9:0]) begin
        image_2_487 <= io_pixelVal_in_2_5;
      end else if (10'h1e7 == _T_28[9:0]) begin
        image_2_487 <= io_pixelVal_in_2_4;
      end else if (10'h1e7 == _T_25[9:0]) begin
        image_2_487 <= io_pixelVal_in_2_3;
      end else if (10'h1e7 == _T_22[9:0]) begin
        image_2_487 <= io_pixelVal_in_2_2;
      end else if (10'h1e7 == _T_19[9:0]) begin
        image_2_487 <= io_pixelVal_in_2_1;
      end else if (10'h1e7 == _T_15[9:0]) begin
        image_2_487 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_488 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e8 == _T_37[9:0]) begin
        image_2_488 <= io_pixelVal_in_2_7;
      end else if (10'h1e8 == _T_34[9:0]) begin
        image_2_488 <= io_pixelVal_in_2_6;
      end else if (10'h1e8 == _T_31[9:0]) begin
        image_2_488 <= io_pixelVal_in_2_5;
      end else if (10'h1e8 == _T_28[9:0]) begin
        image_2_488 <= io_pixelVal_in_2_4;
      end else if (10'h1e8 == _T_25[9:0]) begin
        image_2_488 <= io_pixelVal_in_2_3;
      end else if (10'h1e8 == _T_22[9:0]) begin
        image_2_488 <= io_pixelVal_in_2_2;
      end else if (10'h1e8 == _T_19[9:0]) begin
        image_2_488 <= io_pixelVal_in_2_1;
      end else if (10'h1e8 == _T_15[9:0]) begin
        image_2_488 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_489 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e9 == _T_37[9:0]) begin
        image_2_489 <= io_pixelVal_in_2_7;
      end else if (10'h1e9 == _T_34[9:0]) begin
        image_2_489 <= io_pixelVal_in_2_6;
      end else if (10'h1e9 == _T_31[9:0]) begin
        image_2_489 <= io_pixelVal_in_2_5;
      end else if (10'h1e9 == _T_28[9:0]) begin
        image_2_489 <= io_pixelVal_in_2_4;
      end else if (10'h1e9 == _T_25[9:0]) begin
        image_2_489 <= io_pixelVal_in_2_3;
      end else if (10'h1e9 == _T_22[9:0]) begin
        image_2_489 <= io_pixelVal_in_2_2;
      end else if (10'h1e9 == _T_19[9:0]) begin
        image_2_489 <= io_pixelVal_in_2_1;
      end else if (10'h1e9 == _T_15[9:0]) begin
        image_2_489 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_490 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ea == _T_37[9:0]) begin
        image_2_490 <= io_pixelVal_in_2_7;
      end else if (10'h1ea == _T_34[9:0]) begin
        image_2_490 <= io_pixelVal_in_2_6;
      end else if (10'h1ea == _T_31[9:0]) begin
        image_2_490 <= io_pixelVal_in_2_5;
      end else if (10'h1ea == _T_28[9:0]) begin
        image_2_490 <= io_pixelVal_in_2_4;
      end else if (10'h1ea == _T_25[9:0]) begin
        image_2_490 <= io_pixelVal_in_2_3;
      end else if (10'h1ea == _T_22[9:0]) begin
        image_2_490 <= io_pixelVal_in_2_2;
      end else if (10'h1ea == _T_19[9:0]) begin
        image_2_490 <= io_pixelVal_in_2_1;
      end else if (10'h1ea == _T_15[9:0]) begin
        image_2_490 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_491 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1eb == _T_37[9:0]) begin
        image_2_491 <= io_pixelVal_in_2_7;
      end else if (10'h1eb == _T_34[9:0]) begin
        image_2_491 <= io_pixelVal_in_2_6;
      end else if (10'h1eb == _T_31[9:0]) begin
        image_2_491 <= io_pixelVal_in_2_5;
      end else if (10'h1eb == _T_28[9:0]) begin
        image_2_491 <= io_pixelVal_in_2_4;
      end else if (10'h1eb == _T_25[9:0]) begin
        image_2_491 <= io_pixelVal_in_2_3;
      end else if (10'h1eb == _T_22[9:0]) begin
        image_2_491 <= io_pixelVal_in_2_2;
      end else if (10'h1eb == _T_19[9:0]) begin
        image_2_491 <= io_pixelVal_in_2_1;
      end else if (10'h1eb == _T_15[9:0]) begin
        image_2_491 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_492 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ec == _T_37[9:0]) begin
        image_2_492 <= io_pixelVal_in_2_7;
      end else if (10'h1ec == _T_34[9:0]) begin
        image_2_492 <= io_pixelVal_in_2_6;
      end else if (10'h1ec == _T_31[9:0]) begin
        image_2_492 <= io_pixelVal_in_2_5;
      end else if (10'h1ec == _T_28[9:0]) begin
        image_2_492 <= io_pixelVal_in_2_4;
      end else if (10'h1ec == _T_25[9:0]) begin
        image_2_492 <= io_pixelVal_in_2_3;
      end else if (10'h1ec == _T_22[9:0]) begin
        image_2_492 <= io_pixelVal_in_2_2;
      end else if (10'h1ec == _T_19[9:0]) begin
        image_2_492 <= io_pixelVal_in_2_1;
      end else if (10'h1ec == _T_15[9:0]) begin
        image_2_492 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_493 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ed == _T_37[9:0]) begin
        image_2_493 <= io_pixelVal_in_2_7;
      end else if (10'h1ed == _T_34[9:0]) begin
        image_2_493 <= io_pixelVal_in_2_6;
      end else if (10'h1ed == _T_31[9:0]) begin
        image_2_493 <= io_pixelVal_in_2_5;
      end else if (10'h1ed == _T_28[9:0]) begin
        image_2_493 <= io_pixelVal_in_2_4;
      end else if (10'h1ed == _T_25[9:0]) begin
        image_2_493 <= io_pixelVal_in_2_3;
      end else if (10'h1ed == _T_22[9:0]) begin
        image_2_493 <= io_pixelVal_in_2_2;
      end else if (10'h1ed == _T_19[9:0]) begin
        image_2_493 <= io_pixelVal_in_2_1;
      end else if (10'h1ed == _T_15[9:0]) begin
        image_2_493 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_494 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ee == _T_37[9:0]) begin
        image_2_494 <= io_pixelVal_in_2_7;
      end else if (10'h1ee == _T_34[9:0]) begin
        image_2_494 <= io_pixelVal_in_2_6;
      end else if (10'h1ee == _T_31[9:0]) begin
        image_2_494 <= io_pixelVal_in_2_5;
      end else if (10'h1ee == _T_28[9:0]) begin
        image_2_494 <= io_pixelVal_in_2_4;
      end else if (10'h1ee == _T_25[9:0]) begin
        image_2_494 <= io_pixelVal_in_2_3;
      end else if (10'h1ee == _T_22[9:0]) begin
        image_2_494 <= io_pixelVal_in_2_2;
      end else if (10'h1ee == _T_19[9:0]) begin
        image_2_494 <= io_pixelVal_in_2_1;
      end else if (10'h1ee == _T_15[9:0]) begin
        image_2_494 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_495 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ef == _T_37[9:0]) begin
        image_2_495 <= io_pixelVal_in_2_7;
      end else if (10'h1ef == _T_34[9:0]) begin
        image_2_495 <= io_pixelVal_in_2_6;
      end else if (10'h1ef == _T_31[9:0]) begin
        image_2_495 <= io_pixelVal_in_2_5;
      end else if (10'h1ef == _T_28[9:0]) begin
        image_2_495 <= io_pixelVal_in_2_4;
      end else if (10'h1ef == _T_25[9:0]) begin
        image_2_495 <= io_pixelVal_in_2_3;
      end else if (10'h1ef == _T_22[9:0]) begin
        image_2_495 <= io_pixelVal_in_2_2;
      end else if (10'h1ef == _T_19[9:0]) begin
        image_2_495 <= io_pixelVal_in_2_1;
      end else if (10'h1ef == _T_15[9:0]) begin
        image_2_495 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_496 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f0 == _T_37[9:0]) begin
        image_2_496 <= io_pixelVal_in_2_7;
      end else if (10'h1f0 == _T_34[9:0]) begin
        image_2_496 <= io_pixelVal_in_2_6;
      end else if (10'h1f0 == _T_31[9:0]) begin
        image_2_496 <= io_pixelVal_in_2_5;
      end else if (10'h1f0 == _T_28[9:0]) begin
        image_2_496 <= io_pixelVal_in_2_4;
      end else if (10'h1f0 == _T_25[9:0]) begin
        image_2_496 <= io_pixelVal_in_2_3;
      end else if (10'h1f0 == _T_22[9:0]) begin
        image_2_496 <= io_pixelVal_in_2_2;
      end else if (10'h1f0 == _T_19[9:0]) begin
        image_2_496 <= io_pixelVal_in_2_1;
      end else if (10'h1f0 == _T_15[9:0]) begin
        image_2_496 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_497 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f1 == _T_37[9:0]) begin
        image_2_497 <= io_pixelVal_in_2_7;
      end else if (10'h1f1 == _T_34[9:0]) begin
        image_2_497 <= io_pixelVal_in_2_6;
      end else if (10'h1f1 == _T_31[9:0]) begin
        image_2_497 <= io_pixelVal_in_2_5;
      end else if (10'h1f1 == _T_28[9:0]) begin
        image_2_497 <= io_pixelVal_in_2_4;
      end else if (10'h1f1 == _T_25[9:0]) begin
        image_2_497 <= io_pixelVal_in_2_3;
      end else if (10'h1f1 == _T_22[9:0]) begin
        image_2_497 <= io_pixelVal_in_2_2;
      end else if (10'h1f1 == _T_19[9:0]) begin
        image_2_497 <= io_pixelVal_in_2_1;
      end else if (10'h1f1 == _T_15[9:0]) begin
        image_2_497 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_498 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f2 == _T_37[9:0]) begin
        image_2_498 <= io_pixelVal_in_2_7;
      end else if (10'h1f2 == _T_34[9:0]) begin
        image_2_498 <= io_pixelVal_in_2_6;
      end else if (10'h1f2 == _T_31[9:0]) begin
        image_2_498 <= io_pixelVal_in_2_5;
      end else if (10'h1f2 == _T_28[9:0]) begin
        image_2_498 <= io_pixelVal_in_2_4;
      end else if (10'h1f2 == _T_25[9:0]) begin
        image_2_498 <= io_pixelVal_in_2_3;
      end else if (10'h1f2 == _T_22[9:0]) begin
        image_2_498 <= io_pixelVal_in_2_2;
      end else if (10'h1f2 == _T_19[9:0]) begin
        image_2_498 <= io_pixelVal_in_2_1;
      end else if (10'h1f2 == _T_15[9:0]) begin
        image_2_498 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_499 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f3 == _T_37[9:0]) begin
        image_2_499 <= io_pixelVal_in_2_7;
      end else if (10'h1f3 == _T_34[9:0]) begin
        image_2_499 <= io_pixelVal_in_2_6;
      end else if (10'h1f3 == _T_31[9:0]) begin
        image_2_499 <= io_pixelVal_in_2_5;
      end else if (10'h1f3 == _T_28[9:0]) begin
        image_2_499 <= io_pixelVal_in_2_4;
      end else if (10'h1f3 == _T_25[9:0]) begin
        image_2_499 <= io_pixelVal_in_2_3;
      end else if (10'h1f3 == _T_22[9:0]) begin
        image_2_499 <= io_pixelVal_in_2_2;
      end else if (10'h1f3 == _T_19[9:0]) begin
        image_2_499 <= io_pixelVal_in_2_1;
      end else if (10'h1f3 == _T_15[9:0]) begin
        image_2_499 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_500 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f4 == _T_37[9:0]) begin
        image_2_500 <= io_pixelVal_in_2_7;
      end else if (10'h1f4 == _T_34[9:0]) begin
        image_2_500 <= io_pixelVal_in_2_6;
      end else if (10'h1f4 == _T_31[9:0]) begin
        image_2_500 <= io_pixelVal_in_2_5;
      end else if (10'h1f4 == _T_28[9:0]) begin
        image_2_500 <= io_pixelVal_in_2_4;
      end else if (10'h1f4 == _T_25[9:0]) begin
        image_2_500 <= io_pixelVal_in_2_3;
      end else if (10'h1f4 == _T_22[9:0]) begin
        image_2_500 <= io_pixelVal_in_2_2;
      end else if (10'h1f4 == _T_19[9:0]) begin
        image_2_500 <= io_pixelVal_in_2_1;
      end else if (10'h1f4 == _T_15[9:0]) begin
        image_2_500 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_501 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f5 == _T_37[9:0]) begin
        image_2_501 <= io_pixelVal_in_2_7;
      end else if (10'h1f5 == _T_34[9:0]) begin
        image_2_501 <= io_pixelVal_in_2_6;
      end else if (10'h1f5 == _T_31[9:0]) begin
        image_2_501 <= io_pixelVal_in_2_5;
      end else if (10'h1f5 == _T_28[9:0]) begin
        image_2_501 <= io_pixelVal_in_2_4;
      end else if (10'h1f5 == _T_25[9:0]) begin
        image_2_501 <= io_pixelVal_in_2_3;
      end else if (10'h1f5 == _T_22[9:0]) begin
        image_2_501 <= io_pixelVal_in_2_2;
      end else if (10'h1f5 == _T_19[9:0]) begin
        image_2_501 <= io_pixelVal_in_2_1;
      end else if (10'h1f5 == _T_15[9:0]) begin
        image_2_501 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_502 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f6 == _T_37[9:0]) begin
        image_2_502 <= io_pixelVal_in_2_7;
      end else if (10'h1f6 == _T_34[9:0]) begin
        image_2_502 <= io_pixelVal_in_2_6;
      end else if (10'h1f6 == _T_31[9:0]) begin
        image_2_502 <= io_pixelVal_in_2_5;
      end else if (10'h1f6 == _T_28[9:0]) begin
        image_2_502 <= io_pixelVal_in_2_4;
      end else if (10'h1f6 == _T_25[9:0]) begin
        image_2_502 <= io_pixelVal_in_2_3;
      end else if (10'h1f6 == _T_22[9:0]) begin
        image_2_502 <= io_pixelVal_in_2_2;
      end else if (10'h1f6 == _T_19[9:0]) begin
        image_2_502 <= io_pixelVal_in_2_1;
      end else if (10'h1f6 == _T_15[9:0]) begin
        image_2_502 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_503 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f7 == _T_37[9:0]) begin
        image_2_503 <= io_pixelVal_in_2_7;
      end else if (10'h1f7 == _T_34[9:0]) begin
        image_2_503 <= io_pixelVal_in_2_6;
      end else if (10'h1f7 == _T_31[9:0]) begin
        image_2_503 <= io_pixelVal_in_2_5;
      end else if (10'h1f7 == _T_28[9:0]) begin
        image_2_503 <= io_pixelVal_in_2_4;
      end else if (10'h1f7 == _T_25[9:0]) begin
        image_2_503 <= io_pixelVal_in_2_3;
      end else if (10'h1f7 == _T_22[9:0]) begin
        image_2_503 <= io_pixelVal_in_2_2;
      end else if (10'h1f7 == _T_19[9:0]) begin
        image_2_503 <= io_pixelVal_in_2_1;
      end else if (10'h1f7 == _T_15[9:0]) begin
        image_2_503 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_504 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f8 == _T_37[9:0]) begin
        image_2_504 <= io_pixelVal_in_2_7;
      end else if (10'h1f8 == _T_34[9:0]) begin
        image_2_504 <= io_pixelVal_in_2_6;
      end else if (10'h1f8 == _T_31[9:0]) begin
        image_2_504 <= io_pixelVal_in_2_5;
      end else if (10'h1f8 == _T_28[9:0]) begin
        image_2_504 <= io_pixelVal_in_2_4;
      end else if (10'h1f8 == _T_25[9:0]) begin
        image_2_504 <= io_pixelVal_in_2_3;
      end else if (10'h1f8 == _T_22[9:0]) begin
        image_2_504 <= io_pixelVal_in_2_2;
      end else if (10'h1f8 == _T_19[9:0]) begin
        image_2_504 <= io_pixelVal_in_2_1;
      end else if (10'h1f8 == _T_15[9:0]) begin
        image_2_504 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_505 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f9 == _T_37[9:0]) begin
        image_2_505 <= io_pixelVal_in_2_7;
      end else if (10'h1f9 == _T_34[9:0]) begin
        image_2_505 <= io_pixelVal_in_2_6;
      end else if (10'h1f9 == _T_31[9:0]) begin
        image_2_505 <= io_pixelVal_in_2_5;
      end else if (10'h1f9 == _T_28[9:0]) begin
        image_2_505 <= io_pixelVal_in_2_4;
      end else if (10'h1f9 == _T_25[9:0]) begin
        image_2_505 <= io_pixelVal_in_2_3;
      end else if (10'h1f9 == _T_22[9:0]) begin
        image_2_505 <= io_pixelVal_in_2_2;
      end else if (10'h1f9 == _T_19[9:0]) begin
        image_2_505 <= io_pixelVal_in_2_1;
      end else if (10'h1f9 == _T_15[9:0]) begin
        image_2_505 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_506 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1fa == _T_37[9:0]) begin
        image_2_506 <= io_pixelVal_in_2_7;
      end else if (10'h1fa == _T_34[9:0]) begin
        image_2_506 <= io_pixelVal_in_2_6;
      end else if (10'h1fa == _T_31[9:0]) begin
        image_2_506 <= io_pixelVal_in_2_5;
      end else if (10'h1fa == _T_28[9:0]) begin
        image_2_506 <= io_pixelVal_in_2_4;
      end else if (10'h1fa == _T_25[9:0]) begin
        image_2_506 <= io_pixelVal_in_2_3;
      end else if (10'h1fa == _T_22[9:0]) begin
        image_2_506 <= io_pixelVal_in_2_2;
      end else if (10'h1fa == _T_19[9:0]) begin
        image_2_506 <= io_pixelVal_in_2_1;
      end else if (10'h1fa == _T_15[9:0]) begin
        image_2_506 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_507 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1fb == _T_37[9:0]) begin
        image_2_507 <= io_pixelVal_in_2_7;
      end else if (10'h1fb == _T_34[9:0]) begin
        image_2_507 <= io_pixelVal_in_2_6;
      end else if (10'h1fb == _T_31[9:0]) begin
        image_2_507 <= io_pixelVal_in_2_5;
      end else if (10'h1fb == _T_28[9:0]) begin
        image_2_507 <= io_pixelVal_in_2_4;
      end else if (10'h1fb == _T_25[9:0]) begin
        image_2_507 <= io_pixelVal_in_2_3;
      end else if (10'h1fb == _T_22[9:0]) begin
        image_2_507 <= io_pixelVal_in_2_2;
      end else if (10'h1fb == _T_19[9:0]) begin
        image_2_507 <= io_pixelVal_in_2_1;
      end else if (10'h1fb == _T_15[9:0]) begin
        image_2_507 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_508 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1fc == _T_37[9:0]) begin
        image_2_508 <= io_pixelVal_in_2_7;
      end else if (10'h1fc == _T_34[9:0]) begin
        image_2_508 <= io_pixelVal_in_2_6;
      end else if (10'h1fc == _T_31[9:0]) begin
        image_2_508 <= io_pixelVal_in_2_5;
      end else if (10'h1fc == _T_28[9:0]) begin
        image_2_508 <= io_pixelVal_in_2_4;
      end else if (10'h1fc == _T_25[9:0]) begin
        image_2_508 <= io_pixelVal_in_2_3;
      end else if (10'h1fc == _T_22[9:0]) begin
        image_2_508 <= io_pixelVal_in_2_2;
      end else if (10'h1fc == _T_19[9:0]) begin
        image_2_508 <= io_pixelVal_in_2_1;
      end else if (10'h1fc == _T_15[9:0]) begin
        image_2_508 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_509 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1fd == _T_37[9:0]) begin
        image_2_509 <= io_pixelVal_in_2_7;
      end else if (10'h1fd == _T_34[9:0]) begin
        image_2_509 <= io_pixelVal_in_2_6;
      end else if (10'h1fd == _T_31[9:0]) begin
        image_2_509 <= io_pixelVal_in_2_5;
      end else if (10'h1fd == _T_28[9:0]) begin
        image_2_509 <= io_pixelVal_in_2_4;
      end else if (10'h1fd == _T_25[9:0]) begin
        image_2_509 <= io_pixelVal_in_2_3;
      end else if (10'h1fd == _T_22[9:0]) begin
        image_2_509 <= io_pixelVal_in_2_2;
      end else if (10'h1fd == _T_19[9:0]) begin
        image_2_509 <= io_pixelVal_in_2_1;
      end else if (10'h1fd == _T_15[9:0]) begin
        image_2_509 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_510 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1fe == _T_37[9:0]) begin
        image_2_510 <= io_pixelVal_in_2_7;
      end else if (10'h1fe == _T_34[9:0]) begin
        image_2_510 <= io_pixelVal_in_2_6;
      end else if (10'h1fe == _T_31[9:0]) begin
        image_2_510 <= io_pixelVal_in_2_5;
      end else if (10'h1fe == _T_28[9:0]) begin
        image_2_510 <= io_pixelVal_in_2_4;
      end else if (10'h1fe == _T_25[9:0]) begin
        image_2_510 <= io_pixelVal_in_2_3;
      end else if (10'h1fe == _T_22[9:0]) begin
        image_2_510 <= io_pixelVal_in_2_2;
      end else if (10'h1fe == _T_19[9:0]) begin
        image_2_510 <= io_pixelVal_in_2_1;
      end else if (10'h1fe == _T_15[9:0]) begin
        image_2_510 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_511 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ff == _T_37[9:0]) begin
        image_2_511 <= io_pixelVal_in_2_7;
      end else if (10'h1ff == _T_34[9:0]) begin
        image_2_511 <= io_pixelVal_in_2_6;
      end else if (10'h1ff == _T_31[9:0]) begin
        image_2_511 <= io_pixelVal_in_2_5;
      end else if (10'h1ff == _T_28[9:0]) begin
        image_2_511 <= io_pixelVal_in_2_4;
      end else if (10'h1ff == _T_25[9:0]) begin
        image_2_511 <= io_pixelVal_in_2_3;
      end else if (10'h1ff == _T_22[9:0]) begin
        image_2_511 <= io_pixelVal_in_2_2;
      end else if (10'h1ff == _T_19[9:0]) begin
        image_2_511 <= io_pixelVal_in_2_1;
      end else if (10'h1ff == _T_15[9:0]) begin
        image_2_511 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_512 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h200 == _T_37[9:0]) begin
        image_2_512 <= io_pixelVal_in_2_7;
      end else if (10'h200 == _T_34[9:0]) begin
        image_2_512 <= io_pixelVal_in_2_6;
      end else if (10'h200 == _T_31[9:0]) begin
        image_2_512 <= io_pixelVal_in_2_5;
      end else if (10'h200 == _T_28[9:0]) begin
        image_2_512 <= io_pixelVal_in_2_4;
      end else if (10'h200 == _T_25[9:0]) begin
        image_2_512 <= io_pixelVal_in_2_3;
      end else if (10'h200 == _T_22[9:0]) begin
        image_2_512 <= io_pixelVal_in_2_2;
      end else if (10'h200 == _T_19[9:0]) begin
        image_2_512 <= io_pixelVal_in_2_1;
      end else if (10'h200 == _T_15[9:0]) begin
        image_2_512 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_513 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h201 == _T_37[9:0]) begin
        image_2_513 <= io_pixelVal_in_2_7;
      end else if (10'h201 == _T_34[9:0]) begin
        image_2_513 <= io_pixelVal_in_2_6;
      end else if (10'h201 == _T_31[9:0]) begin
        image_2_513 <= io_pixelVal_in_2_5;
      end else if (10'h201 == _T_28[9:0]) begin
        image_2_513 <= io_pixelVal_in_2_4;
      end else if (10'h201 == _T_25[9:0]) begin
        image_2_513 <= io_pixelVal_in_2_3;
      end else if (10'h201 == _T_22[9:0]) begin
        image_2_513 <= io_pixelVal_in_2_2;
      end else if (10'h201 == _T_19[9:0]) begin
        image_2_513 <= io_pixelVal_in_2_1;
      end else if (10'h201 == _T_15[9:0]) begin
        image_2_513 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_514 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h202 == _T_37[9:0]) begin
        image_2_514 <= io_pixelVal_in_2_7;
      end else if (10'h202 == _T_34[9:0]) begin
        image_2_514 <= io_pixelVal_in_2_6;
      end else if (10'h202 == _T_31[9:0]) begin
        image_2_514 <= io_pixelVal_in_2_5;
      end else if (10'h202 == _T_28[9:0]) begin
        image_2_514 <= io_pixelVal_in_2_4;
      end else if (10'h202 == _T_25[9:0]) begin
        image_2_514 <= io_pixelVal_in_2_3;
      end else if (10'h202 == _T_22[9:0]) begin
        image_2_514 <= io_pixelVal_in_2_2;
      end else if (10'h202 == _T_19[9:0]) begin
        image_2_514 <= io_pixelVal_in_2_1;
      end else if (10'h202 == _T_15[9:0]) begin
        image_2_514 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_515 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h203 == _T_37[9:0]) begin
        image_2_515 <= io_pixelVal_in_2_7;
      end else if (10'h203 == _T_34[9:0]) begin
        image_2_515 <= io_pixelVal_in_2_6;
      end else if (10'h203 == _T_31[9:0]) begin
        image_2_515 <= io_pixelVal_in_2_5;
      end else if (10'h203 == _T_28[9:0]) begin
        image_2_515 <= io_pixelVal_in_2_4;
      end else if (10'h203 == _T_25[9:0]) begin
        image_2_515 <= io_pixelVal_in_2_3;
      end else if (10'h203 == _T_22[9:0]) begin
        image_2_515 <= io_pixelVal_in_2_2;
      end else if (10'h203 == _T_19[9:0]) begin
        image_2_515 <= io_pixelVal_in_2_1;
      end else if (10'h203 == _T_15[9:0]) begin
        image_2_515 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_516 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h204 == _T_37[9:0]) begin
        image_2_516 <= io_pixelVal_in_2_7;
      end else if (10'h204 == _T_34[9:0]) begin
        image_2_516 <= io_pixelVal_in_2_6;
      end else if (10'h204 == _T_31[9:0]) begin
        image_2_516 <= io_pixelVal_in_2_5;
      end else if (10'h204 == _T_28[9:0]) begin
        image_2_516 <= io_pixelVal_in_2_4;
      end else if (10'h204 == _T_25[9:0]) begin
        image_2_516 <= io_pixelVal_in_2_3;
      end else if (10'h204 == _T_22[9:0]) begin
        image_2_516 <= io_pixelVal_in_2_2;
      end else if (10'h204 == _T_19[9:0]) begin
        image_2_516 <= io_pixelVal_in_2_1;
      end else if (10'h204 == _T_15[9:0]) begin
        image_2_516 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_517 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h205 == _T_37[9:0]) begin
        image_2_517 <= io_pixelVal_in_2_7;
      end else if (10'h205 == _T_34[9:0]) begin
        image_2_517 <= io_pixelVal_in_2_6;
      end else if (10'h205 == _T_31[9:0]) begin
        image_2_517 <= io_pixelVal_in_2_5;
      end else if (10'h205 == _T_28[9:0]) begin
        image_2_517 <= io_pixelVal_in_2_4;
      end else if (10'h205 == _T_25[9:0]) begin
        image_2_517 <= io_pixelVal_in_2_3;
      end else if (10'h205 == _T_22[9:0]) begin
        image_2_517 <= io_pixelVal_in_2_2;
      end else if (10'h205 == _T_19[9:0]) begin
        image_2_517 <= io_pixelVal_in_2_1;
      end else if (10'h205 == _T_15[9:0]) begin
        image_2_517 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_518 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h206 == _T_37[9:0]) begin
        image_2_518 <= io_pixelVal_in_2_7;
      end else if (10'h206 == _T_34[9:0]) begin
        image_2_518 <= io_pixelVal_in_2_6;
      end else if (10'h206 == _T_31[9:0]) begin
        image_2_518 <= io_pixelVal_in_2_5;
      end else if (10'h206 == _T_28[9:0]) begin
        image_2_518 <= io_pixelVal_in_2_4;
      end else if (10'h206 == _T_25[9:0]) begin
        image_2_518 <= io_pixelVal_in_2_3;
      end else if (10'h206 == _T_22[9:0]) begin
        image_2_518 <= io_pixelVal_in_2_2;
      end else if (10'h206 == _T_19[9:0]) begin
        image_2_518 <= io_pixelVal_in_2_1;
      end else if (10'h206 == _T_15[9:0]) begin
        image_2_518 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_519 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h207 == _T_37[9:0]) begin
        image_2_519 <= io_pixelVal_in_2_7;
      end else if (10'h207 == _T_34[9:0]) begin
        image_2_519 <= io_pixelVal_in_2_6;
      end else if (10'h207 == _T_31[9:0]) begin
        image_2_519 <= io_pixelVal_in_2_5;
      end else if (10'h207 == _T_28[9:0]) begin
        image_2_519 <= io_pixelVal_in_2_4;
      end else if (10'h207 == _T_25[9:0]) begin
        image_2_519 <= io_pixelVal_in_2_3;
      end else if (10'h207 == _T_22[9:0]) begin
        image_2_519 <= io_pixelVal_in_2_2;
      end else if (10'h207 == _T_19[9:0]) begin
        image_2_519 <= io_pixelVal_in_2_1;
      end else if (10'h207 == _T_15[9:0]) begin
        image_2_519 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_520 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h208 == _T_37[9:0]) begin
        image_2_520 <= io_pixelVal_in_2_7;
      end else if (10'h208 == _T_34[9:0]) begin
        image_2_520 <= io_pixelVal_in_2_6;
      end else if (10'h208 == _T_31[9:0]) begin
        image_2_520 <= io_pixelVal_in_2_5;
      end else if (10'h208 == _T_28[9:0]) begin
        image_2_520 <= io_pixelVal_in_2_4;
      end else if (10'h208 == _T_25[9:0]) begin
        image_2_520 <= io_pixelVal_in_2_3;
      end else if (10'h208 == _T_22[9:0]) begin
        image_2_520 <= io_pixelVal_in_2_2;
      end else if (10'h208 == _T_19[9:0]) begin
        image_2_520 <= io_pixelVal_in_2_1;
      end else if (10'h208 == _T_15[9:0]) begin
        image_2_520 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_521 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h209 == _T_37[9:0]) begin
        image_2_521 <= io_pixelVal_in_2_7;
      end else if (10'h209 == _T_34[9:0]) begin
        image_2_521 <= io_pixelVal_in_2_6;
      end else if (10'h209 == _T_31[9:0]) begin
        image_2_521 <= io_pixelVal_in_2_5;
      end else if (10'h209 == _T_28[9:0]) begin
        image_2_521 <= io_pixelVal_in_2_4;
      end else if (10'h209 == _T_25[9:0]) begin
        image_2_521 <= io_pixelVal_in_2_3;
      end else if (10'h209 == _T_22[9:0]) begin
        image_2_521 <= io_pixelVal_in_2_2;
      end else if (10'h209 == _T_19[9:0]) begin
        image_2_521 <= io_pixelVal_in_2_1;
      end else if (10'h209 == _T_15[9:0]) begin
        image_2_521 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_522 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20a == _T_37[9:0]) begin
        image_2_522 <= io_pixelVal_in_2_7;
      end else if (10'h20a == _T_34[9:0]) begin
        image_2_522 <= io_pixelVal_in_2_6;
      end else if (10'h20a == _T_31[9:0]) begin
        image_2_522 <= io_pixelVal_in_2_5;
      end else if (10'h20a == _T_28[9:0]) begin
        image_2_522 <= io_pixelVal_in_2_4;
      end else if (10'h20a == _T_25[9:0]) begin
        image_2_522 <= io_pixelVal_in_2_3;
      end else if (10'h20a == _T_22[9:0]) begin
        image_2_522 <= io_pixelVal_in_2_2;
      end else if (10'h20a == _T_19[9:0]) begin
        image_2_522 <= io_pixelVal_in_2_1;
      end else if (10'h20a == _T_15[9:0]) begin
        image_2_522 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_523 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20b == _T_37[9:0]) begin
        image_2_523 <= io_pixelVal_in_2_7;
      end else if (10'h20b == _T_34[9:0]) begin
        image_2_523 <= io_pixelVal_in_2_6;
      end else if (10'h20b == _T_31[9:0]) begin
        image_2_523 <= io_pixelVal_in_2_5;
      end else if (10'h20b == _T_28[9:0]) begin
        image_2_523 <= io_pixelVal_in_2_4;
      end else if (10'h20b == _T_25[9:0]) begin
        image_2_523 <= io_pixelVal_in_2_3;
      end else if (10'h20b == _T_22[9:0]) begin
        image_2_523 <= io_pixelVal_in_2_2;
      end else if (10'h20b == _T_19[9:0]) begin
        image_2_523 <= io_pixelVal_in_2_1;
      end else if (10'h20b == _T_15[9:0]) begin
        image_2_523 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_524 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20c == _T_37[9:0]) begin
        image_2_524 <= io_pixelVal_in_2_7;
      end else if (10'h20c == _T_34[9:0]) begin
        image_2_524 <= io_pixelVal_in_2_6;
      end else if (10'h20c == _T_31[9:0]) begin
        image_2_524 <= io_pixelVal_in_2_5;
      end else if (10'h20c == _T_28[9:0]) begin
        image_2_524 <= io_pixelVal_in_2_4;
      end else if (10'h20c == _T_25[9:0]) begin
        image_2_524 <= io_pixelVal_in_2_3;
      end else if (10'h20c == _T_22[9:0]) begin
        image_2_524 <= io_pixelVal_in_2_2;
      end else if (10'h20c == _T_19[9:0]) begin
        image_2_524 <= io_pixelVal_in_2_1;
      end else if (10'h20c == _T_15[9:0]) begin
        image_2_524 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_525 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20d == _T_37[9:0]) begin
        image_2_525 <= io_pixelVal_in_2_7;
      end else if (10'h20d == _T_34[9:0]) begin
        image_2_525 <= io_pixelVal_in_2_6;
      end else if (10'h20d == _T_31[9:0]) begin
        image_2_525 <= io_pixelVal_in_2_5;
      end else if (10'h20d == _T_28[9:0]) begin
        image_2_525 <= io_pixelVal_in_2_4;
      end else if (10'h20d == _T_25[9:0]) begin
        image_2_525 <= io_pixelVal_in_2_3;
      end else if (10'h20d == _T_22[9:0]) begin
        image_2_525 <= io_pixelVal_in_2_2;
      end else if (10'h20d == _T_19[9:0]) begin
        image_2_525 <= io_pixelVal_in_2_1;
      end else if (10'h20d == _T_15[9:0]) begin
        image_2_525 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_526 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20e == _T_37[9:0]) begin
        image_2_526 <= io_pixelVal_in_2_7;
      end else if (10'h20e == _T_34[9:0]) begin
        image_2_526 <= io_pixelVal_in_2_6;
      end else if (10'h20e == _T_31[9:0]) begin
        image_2_526 <= io_pixelVal_in_2_5;
      end else if (10'h20e == _T_28[9:0]) begin
        image_2_526 <= io_pixelVal_in_2_4;
      end else if (10'h20e == _T_25[9:0]) begin
        image_2_526 <= io_pixelVal_in_2_3;
      end else if (10'h20e == _T_22[9:0]) begin
        image_2_526 <= io_pixelVal_in_2_2;
      end else if (10'h20e == _T_19[9:0]) begin
        image_2_526 <= io_pixelVal_in_2_1;
      end else if (10'h20e == _T_15[9:0]) begin
        image_2_526 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_527 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20f == _T_37[9:0]) begin
        image_2_527 <= io_pixelVal_in_2_7;
      end else if (10'h20f == _T_34[9:0]) begin
        image_2_527 <= io_pixelVal_in_2_6;
      end else if (10'h20f == _T_31[9:0]) begin
        image_2_527 <= io_pixelVal_in_2_5;
      end else if (10'h20f == _T_28[9:0]) begin
        image_2_527 <= io_pixelVal_in_2_4;
      end else if (10'h20f == _T_25[9:0]) begin
        image_2_527 <= io_pixelVal_in_2_3;
      end else if (10'h20f == _T_22[9:0]) begin
        image_2_527 <= io_pixelVal_in_2_2;
      end else if (10'h20f == _T_19[9:0]) begin
        image_2_527 <= io_pixelVal_in_2_1;
      end else if (10'h20f == _T_15[9:0]) begin
        image_2_527 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_528 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h210 == _T_37[9:0]) begin
        image_2_528 <= io_pixelVal_in_2_7;
      end else if (10'h210 == _T_34[9:0]) begin
        image_2_528 <= io_pixelVal_in_2_6;
      end else if (10'h210 == _T_31[9:0]) begin
        image_2_528 <= io_pixelVal_in_2_5;
      end else if (10'h210 == _T_28[9:0]) begin
        image_2_528 <= io_pixelVal_in_2_4;
      end else if (10'h210 == _T_25[9:0]) begin
        image_2_528 <= io_pixelVal_in_2_3;
      end else if (10'h210 == _T_22[9:0]) begin
        image_2_528 <= io_pixelVal_in_2_2;
      end else if (10'h210 == _T_19[9:0]) begin
        image_2_528 <= io_pixelVal_in_2_1;
      end else if (10'h210 == _T_15[9:0]) begin
        image_2_528 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_529 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h211 == _T_37[9:0]) begin
        image_2_529 <= io_pixelVal_in_2_7;
      end else if (10'h211 == _T_34[9:0]) begin
        image_2_529 <= io_pixelVal_in_2_6;
      end else if (10'h211 == _T_31[9:0]) begin
        image_2_529 <= io_pixelVal_in_2_5;
      end else if (10'h211 == _T_28[9:0]) begin
        image_2_529 <= io_pixelVal_in_2_4;
      end else if (10'h211 == _T_25[9:0]) begin
        image_2_529 <= io_pixelVal_in_2_3;
      end else if (10'h211 == _T_22[9:0]) begin
        image_2_529 <= io_pixelVal_in_2_2;
      end else if (10'h211 == _T_19[9:0]) begin
        image_2_529 <= io_pixelVal_in_2_1;
      end else if (10'h211 == _T_15[9:0]) begin
        image_2_529 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_530 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h212 == _T_37[9:0]) begin
        image_2_530 <= io_pixelVal_in_2_7;
      end else if (10'h212 == _T_34[9:0]) begin
        image_2_530 <= io_pixelVal_in_2_6;
      end else if (10'h212 == _T_31[9:0]) begin
        image_2_530 <= io_pixelVal_in_2_5;
      end else if (10'h212 == _T_28[9:0]) begin
        image_2_530 <= io_pixelVal_in_2_4;
      end else if (10'h212 == _T_25[9:0]) begin
        image_2_530 <= io_pixelVal_in_2_3;
      end else if (10'h212 == _T_22[9:0]) begin
        image_2_530 <= io_pixelVal_in_2_2;
      end else if (10'h212 == _T_19[9:0]) begin
        image_2_530 <= io_pixelVal_in_2_1;
      end else if (10'h212 == _T_15[9:0]) begin
        image_2_530 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_531 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h213 == _T_37[9:0]) begin
        image_2_531 <= io_pixelVal_in_2_7;
      end else if (10'h213 == _T_34[9:0]) begin
        image_2_531 <= io_pixelVal_in_2_6;
      end else if (10'h213 == _T_31[9:0]) begin
        image_2_531 <= io_pixelVal_in_2_5;
      end else if (10'h213 == _T_28[9:0]) begin
        image_2_531 <= io_pixelVal_in_2_4;
      end else if (10'h213 == _T_25[9:0]) begin
        image_2_531 <= io_pixelVal_in_2_3;
      end else if (10'h213 == _T_22[9:0]) begin
        image_2_531 <= io_pixelVal_in_2_2;
      end else if (10'h213 == _T_19[9:0]) begin
        image_2_531 <= io_pixelVal_in_2_1;
      end else if (10'h213 == _T_15[9:0]) begin
        image_2_531 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_532 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h214 == _T_37[9:0]) begin
        image_2_532 <= io_pixelVal_in_2_7;
      end else if (10'h214 == _T_34[9:0]) begin
        image_2_532 <= io_pixelVal_in_2_6;
      end else if (10'h214 == _T_31[9:0]) begin
        image_2_532 <= io_pixelVal_in_2_5;
      end else if (10'h214 == _T_28[9:0]) begin
        image_2_532 <= io_pixelVal_in_2_4;
      end else if (10'h214 == _T_25[9:0]) begin
        image_2_532 <= io_pixelVal_in_2_3;
      end else if (10'h214 == _T_22[9:0]) begin
        image_2_532 <= io_pixelVal_in_2_2;
      end else if (10'h214 == _T_19[9:0]) begin
        image_2_532 <= io_pixelVal_in_2_1;
      end else if (10'h214 == _T_15[9:0]) begin
        image_2_532 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_533 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h215 == _T_37[9:0]) begin
        image_2_533 <= io_pixelVal_in_2_7;
      end else if (10'h215 == _T_34[9:0]) begin
        image_2_533 <= io_pixelVal_in_2_6;
      end else if (10'h215 == _T_31[9:0]) begin
        image_2_533 <= io_pixelVal_in_2_5;
      end else if (10'h215 == _T_28[9:0]) begin
        image_2_533 <= io_pixelVal_in_2_4;
      end else if (10'h215 == _T_25[9:0]) begin
        image_2_533 <= io_pixelVal_in_2_3;
      end else if (10'h215 == _T_22[9:0]) begin
        image_2_533 <= io_pixelVal_in_2_2;
      end else if (10'h215 == _T_19[9:0]) begin
        image_2_533 <= io_pixelVal_in_2_1;
      end else if (10'h215 == _T_15[9:0]) begin
        image_2_533 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_534 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h216 == _T_37[9:0]) begin
        image_2_534 <= io_pixelVal_in_2_7;
      end else if (10'h216 == _T_34[9:0]) begin
        image_2_534 <= io_pixelVal_in_2_6;
      end else if (10'h216 == _T_31[9:0]) begin
        image_2_534 <= io_pixelVal_in_2_5;
      end else if (10'h216 == _T_28[9:0]) begin
        image_2_534 <= io_pixelVal_in_2_4;
      end else if (10'h216 == _T_25[9:0]) begin
        image_2_534 <= io_pixelVal_in_2_3;
      end else if (10'h216 == _T_22[9:0]) begin
        image_2_534 <= io_pixelVal_in_2_2;
      end else if (10'h216 == _T_19[9:0]) begin
        image_2_534 <= io_pixelVal_in_2_1;
      end else if (10'h216 == _T_15[9:0]) begin
        image_2_534 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_535 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h217 == _T_37[9:0]) begin
        image_2_535 <= io_pixelVal_in_2_7;
      end else if (10'h217 == _T_34[9:0]) begin
        image_2_535 <= io_pixelVal_in_2_6;
      end else if (10'h217 == _T_31[9:0]) begin
        image_2_535 <= io_pixelVal_in_2_5;
      end else if (10'h217 == _T_28[9:0]) begin
        image_2_535 <= io_pixelVal_in_2_4;
      end else if (10'h217 == _T_25[9:0]) begin
        image_2_535 <= io_pixelVal_in_2_3;
      end else if (10'h217 == _T_22[9:0]) begin
        image_2_535 <= io_pixelVal_in_2_2;
      end else if (10'h217 == _T_19[9:0]) begin
        image_2_535 <= io_pixelVal_in_2_1;
      end else if (10'h217 == _T_15[9:0]) begin
        image_2_535 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_536 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h218 == _T_37[9:0]) begin
        image_2_536 <= io_pixelVal_in_2_7;
      end else if (10'h218 == _T_34[9:0]) begin
        image_2_536 <= io_pixelVal_in_2_6;
      end else if (10'h218 == _T_31[9:0]) begin
        image_2_536 <= io_pixelVal_in_2_5;
      end else if (10'h218 == _T_28[9:0]) begin
        image_2_536 <= io_pixelVal_in_2_4;
      end else if (10'h218 == _T_25[9:0]) begin
        image_2_536 <= io_pixelVal_in_2_3;
      end else if (10'h218 == _T_22[9:0]) begin
        image_2_536 <= io_pixelVal_in_2_2;
      end else if (10'h218 == _T_19[9:0]) begin
        image_2_536 <= io_pixelVal_in_2_1;
      end else if (10'h218 == _T_15[9:0]) begin
        image_2_536 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_537 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h219 == _T_37[9:0]) begin
        image_2_537 <= io_pixelVal_in_2_7;
      end else if (10'h219 == _T_34[9:0]) begin
        image_2_537 <= io_pixelVal_in_2_6;
      end else if (10'h219 == _T_31[9:0]) begin
        image_2_537 <= io_pixelVal_in_2_5;
      end else if (10'h219 == _T_28[9:0]) begin
        image_2_537 <= io_pixelVal_in_2_4;
      end else if (10'h219 == _T_25[9:0]) begin
        image_2_537 <= io_pixelVal_in_2_3;
      end else if (10'h219 == _T_22[9:0]) begin
        image_2_537 <= io_pixelVal_in_2_2;
      end else if (10'h219 == _T_19[9:0]) begin
        image_2_537 <= io_pixelVal_in_2_1;
      end else if (10'h219 == _T_15[9:0]) begin
        image_2_537 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_538 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21a == _T_37[9:0]) begin
        image_2_538 <= io_pixelVal_in_2_7;
      end else if (10'h21a == _T_34[9:0]) begin
        image_2_538 <= io_pixelVal_in_2_6;
      end else if (10'h21a == _T_31[9:0]) begin
        image_2_538 <= io_pixelVal_in_2_5;
      end else if (10'h21a == _T_28[9:0]) begin
        image_2_538 <= io_pixelVal_in_2_4;
      end else if (10'h21a == _T_25[9:0]) begin
        image_2_538 <= io_pixelVal_in_2_3;
      end else if (10'h21a == _T_22[9:0]) begin
        image_2_538 <= io_pixelVal_in_2_2;
      end else if (10'h21a == _T_19[9:0]) begin
        image_2_538 <= io_pixelVal_in_2_1;
      end else if (10'h21a == _T_15[9:0]) begin
        image_2_538 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_539 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21b == _T_37[9:0]) begin
        image_2_539 <= io_pixelVal_in_2_7;
      end else if (10'h21b == _T_34[9:0]) begin
        image_2_539 <= io_pixelVal_in_2_6;
      end else if (10'h21b == _T_31[9:0]) begin
        image_2_539 <= io_pixelVal_in_2_5;
      end else if (10'h21b == _T_28[9:0]) begin
        image_2_539 <= io_pixelVal_in_2_4;
      end else if (10'h21b == _T_25[9:0]) begin
        image_2_539 <= io_pixelVal_in_2_3;
      end else if (10'h21b == _T_22[9:0]) begin
        image_2_539 <= io_pixelVal_in_2_2;
      end else if (10'h21b == _T_19[9:0]) begin
        image_2_539 <= io_pixelVal_in_2_1;
      end else if (10'h21b == _T_15[9:0]) begin
        image_2_539 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_540 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21c == _T_37[9:0]) begin
        image_2_540 <= io_pixelVal_in_2_7;
      end else if (10'h21c == _T_34[9:0]) begin
        image_2_540 <= io_pixelVal_in_2_6;
      end else if (10'h21c == _T_31[9:0]) begin
        image_2_540 <= io_pixelVal_in_2_5;
      end else if (10'h21c == _T_28[9:0]) begin
        image_2_540 <= io_pixelVal_in_2_4;
      end else if (10'h21c == _T_25[9:0]) begin
        image_2_540 <= io_pixelVal_in_2_3;
      end else if (10'h21c == _T_22[9:0]) begin
        image_2_540 <= io_pixelVal_in_2_2;
      end else if (10'h21c == _T_19[9:0]) begin
        image_2_540 <= io_pixelVal_in_2_1;
      end else if (10'h21c == _T_15[9:0]) begin
        image_2_540 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_541 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21d == _T_37[9:0]) begin
        image_2_541 <= io_pixelVal_in_2_7;
      end else if (10'h21d == _T_34[9:0]) begin
        image_2_541 <= io_pixelVal_in_2_6;
      end else if (10'h21d == _T_31[9:0]) begin
        image_2_541 <= io_pixelVal_in_2_5;
      end else if (10'h21d == _T_28[9:0]) begin
        image_2_541 <= io_pixelVal_in_2_4;
      end else if (10'h21d == _T_25[9:0]) begin
        image_2_541 <= io_pixelVal_in_2_3;
      end else if (10'h21d == _T_22[9:0]) begin
        image_2_541 <= io_pixelVal_in_2_2;
      end else if (10'h21d == _T_19[9:0]) begin
        image_2_541 <= io_pixelVal_in_2_1;
      end else if (10'h21d == _T_15[9:0]) begin
        image_2_541 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_542 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21e == _T_37[9:0]) begin
        image_2_542 <= io_pixelVal_in_2_7;
      end else if (10'h21e == _T_34[9:0]) begin
        image_2_542 <= io_pixelVal_in_2_6;
      end else if (10'h21e == _T_31[9:0]) begin
        image_2_542 <= io_pixelVal_in_2_5;
      end else if (10'h21e == _T_28[9:0]) begin
        image_2_542 <= io_pixelVal_in_2_4;
      end else if (10'h21e == _T_25[9:0]) begin
        image_2_542 <= io_pixelVal_in_2_3;
      end else if (10'h21e == _T_22[9:0]) begin
        image_2_542 <= io_pixelVal_in_2_2;
      end else if (10'h21e == _T_19[9:0]) begin
        image_2_542 <= io_pixelVal_in_2_1;
      end else if (10'h21e == _T_15[9:0]) begin
        image_2_542 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_543 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21f == _T_37[9:0]) begin
        image_2_543 <= io_pixelVal_in_2_7;
      end else if (10'h21f == _T_34[9:0]) begin
        image_2_543 <= io_pixelVal_in_2_6;
      end else if (10'h21f == _T_31[9:0]) begin
        image_2_543 <= io_pixelVal_in_2_5;
      end else if (10'h21f == _T_28[9:0]) begin
        image_2_543 <= io_pixelVal_in_2_4;
      end else if (10'h21f == _T_25[9:0]) begin
        image_2_543 <= io_pixelVal_in_2_3;
      end else if (10'h21f == _T_22[9:0]) begin
        image_2_543 <= io_pixelVal_in_2_2;
      end else if (10'h21f == _T_19[9:0]) begin
        image_2_543 <= io_pixelVal_in_2_1;
      end else if (10'h21f == _T_15[9:0]) begin
        image_2_543 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_544 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h220 == _T_37[9:0]) begin
        image_2_544 <= io_pixelVal_in_2_7;
      end else if (10'h220 == _T_34[9:0]) begin
        image_2_544 <= io_pixelVal_in_2_6;
      end else if (10'h220 == _T_31[9:0]) begin
        image_2_544 <= io_pixelVal_in_2_5;
      end else if (10'h220 == _T_28[9:0]) begin
        image_2_544 <= io_pixelVal_in_2_4;
      end else if (10'h220 == _T_25[9:0]) begin
        image_2_544 <= io_pixelVal_in_2_3;
      end else if (10'h220 == _T_22[9:0]) begin
        image_2_544 <= io_pixelVal_in_2_2;
      end else if (10'h220 == _T_19[9:0]) begin
        image_2_544 <= io_pixelVal_in_2_1;
      end else if (10'h220 == _T_15[9:0]) begin
        image_2_544 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_545 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h221 == _T_37[9:0]) begin
        image_2_545 <= io_pixelVal_in_2_7;
      end else if (10'h221 == _T_34[9:0]) begin
        image_2_545 <= io_pixelVal_in_2_6;
      end else if (10'h221 == _T_31[9:0]) begin
        image_2_545 <= io_pixelVal_in_2_5;
      end else if (10'h221 == _T_28[9:0]) begin
        image_2_545 <= io_pixelVal_in_2_4;
      end else if (10'h221 == _T_25[9:0]) begin
        image_2_545 <= io_pixelVal_in_2_3;
      end else if (10'h221 == _T_22[9:0]) begin
        image_2_545 <= io_pixelVal_in_2_2;
      end else if (10'h221 == _T_19[9:0]) begin
        image_2_545 <= io_pixelVal_in_2_1;
      end else if (10'h221 == _T_15[9:0]) begin
        image_2_545 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_546 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h222 == _T_37[9:0]) begin
        image_2_546 <= io_pixelVal_in_2_7;
      end else if (10'h222 == _T_34[9:0]) begin
        image_2_546 <= io_pixelVal_in_2_6;
      end else if (10'h222 == _T_31[9:0]) begin
        image_2_546 <= io_pixelVal_in_2_5;
      end else if (10'h222 == _T_28[9:0]) begin
        image_2_546 <= io_pixelVal_in_2_4;
      end else if (10'h222 == _T_25[9:0]) begin
        image_2_546 <= io_pixelVal_in_2_3;
      end else if (10'h222 == _T_22[9:0]) begin
        image_2_546 <= io_pixelVal_in_2_2;
      end else if (10'h222 == _T_19[9:0]) begin
        image_2_546 <= io_pixelVal_in_2_1;
      end else if (10'h222 == _T_15[9:0]) begin
        image_2_546 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_547 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h223 == _T_37[9:0]) begin
        image_2_547 <= io_pixelVal_in_2_7;
      end else if (10'h223 == _T_34[9:0]) begin
        image_2_547 <= io_pixelVal_in_2_6;
      end else if (10'h223 == _T_31[9:0]) begin
        image_2_547 <= io_pixelVal_in_2_5;
      end else if (10'h223 == _T_28[9:0]) begin
        image_2_547 <= io_pixelVal_in_2_4;
      end else if (10'h223 == _T_25[9:0]) begin
        image_2_547 <= io_pixelVal_in_2_3;
      end else if (10'h223 == _T_22[9:0]) begin
        image_2_547 <= io_pixelVal_in_2_2;
      end else if (10'h223 == _T_19[9:0]) begin
        image_2_547 <= io_pixelVal_in_2_1;
      end else if (10'h223 == _T_15[9:0]) begin
        image_2_547 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_548 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h224 == _T_37[9:0]) begin
        image_2_548 <= io_pixelVal_in_2_7;
      end else if (10'h224 == _T_34[9:0]) begin
        image_2_548 <= io_pixelVal_in_2_6;
      end else if (10'h224 == _T_31[9:0]) begin
        image_2_548 <= io_pixelVal_in_2_5;
      end else if (10'h224 == _T_28[9:0]) begin
        image_2_548 <= io_pixelVal_in_2_4;
      end else if (10'h224 == _T_25[9:0]) begin
        image_2_548 <= io_pixelVal_in_2_3;
      end else if (10'h224 == _T_22[9:0]) begin
        image_2_548 <= io_pixelVal_in_2_2;
      end else if (10'h224 == _T_19[9:0]) begin
        image_2_548 <= io_pixelVal_in_2_1;
      end else if (10'h224 == _T_15[9:0]) begin
        image_2_548 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_549 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h225 == _T_37[9:0]) begin
        image_2_549 <= io_pixelVal_in_2_7;
      end else if (10'h225 == _T_34[9:0]) begin
        image_2_549 <= io_pixelVal_in_2_6;
      end else if (10'h225 == _T_31[9:0]) begin
        image_2_549 <= io_pixelVal_in_2_5;
      end else if (10'h225 == _T_28[9:0]) begin
        image_2_549 <= io_pixelVal_in_2_4;
      end else if (10'h225 == _T_25[9:0]) begin
        image_2_549 <= io_pixelVal_in_2_3;
      end else if (10'h225 == _T_22[9:0]) begin
        image_2_549 <= io_pixelVal_in_2_2;
      end else if (10'h225 == _T_19[9:0]) begin
        image_2_549 <= io_pixelVal_in_2_1;
      end else if (10'h225 == _T_15[9:0]) begin
        image_2_549 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_550 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h226 == _T_37[9:0]) begin
        image_2_550 <= io_pixelVal_in_2_7;
      end else if (10'h226 == _T_34[9:0]) begin
        image_2_550 <= io_pixelVal_in_2_6;
      end else if (10'h226 == _T_31[9:0]) begin
        image_2_550 <= io_pixelVal_in_2_5;
      end else if (10'h226 == _T_28[9:0]) begin
        image_2_550 <= io_pixelVal_in_2_4;
      end else if (10'h226 == _T_25[9:0]) begin
        image_2_550 <= io_pixelVal_in_2_3;
      end else if (10'h226 == _T_22[9:0]) begin
        image_2_550 <= io_pixelVal_in_2_2;
      end else if (10'h226 == _T_19[9:0]) begin
        image_2_550 <= io_pixelVal_in_2_1;
      end else if (10'h226 == _T_15[9:0]) begin
        image_2_550 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_551 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h227 == _T_37[9:0]) begin
        image_2_551 <= io_pixelVal_in_2_7;
      end else if (10'h227 == _T_34[9:0]) begin
        image_2_551 <= io_pixelVal_in_2_6;
      end else if (10'h227 == _T_31[9:0]) begin
        image_2_551 <= io_pixelVal_in_2_5;
      end else if (10'h227 == _T_28[9:0]) begin
        image_2_551 <= io_pixelVal_in_2_4;
      end else if (10'h227 == _T_25[9:0]) begin
        image_2_551 <= io_pixelVal_in_2_3;
      end else if (10'h227 == _T_22[9:0]) begin
        image_2_551 <= io_pixelVal_in_2_2;
      end else if (10'h227 == _T_19[9:0]) begin
        image_2_551 <= io_pixelVal_in_2_1;
      end else if (10'h227 == _T_15[9:0]) begin
        image_2_551 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_552 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h228 == _T_37[9:0]) begin
        image_2_552 <= io_pixelVal_in_2_7;
      end else if (10'h228 == _T_34[9:0]) begin
        image_2_552 <= io_pixelVal_in_2_6;
      end else if (10'h228 == _T_31[9:0]) begin
        image_2_552 <= io_pixelVal_in_2_5;
      end else if (10'h228 == _T_28[9:0]) begin
        image_2_552 <= io_pixelVal_in_2_4;
      end else if (10'h228 == _T_25[9:0]) begin
        image_2_552 <= io_pixelVal_in_2_3;
      end else if (10'h228 == _T_22[9:0]) begin
        image_2_552 <= io_pixelVal_in_2_2;
      end else if (10'h228 == _T_19[9:0]) begin
        image_2_552 <= io_pixelVal_in_2_1;
      end else if (10'h228 == _T_15[9:0]) begin
        image_2_552 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_553 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h229 == _T_37[9:0]) begin
        image_2_553 <= io_pixelVal_in_2_7;
      end else if (10'h229 == _T_34[9:0]) begin
        image_2_553 <= io_pixelVal_in_2_6;
      end else if (10'h229 == _T_31[9:0]) begin
        image_2_553 <= io_pixelVal_in_2_5;
      end else if (10'h229 == _T_28[9:0]) begin
        image_2_553 <= io_pixelVal_in_2_4;
      end else if (10'h229 == _T_25[9:0]) begin
        image_2_553 <= io_pixelVal_in_2_3;
      end else if (10'h229 == _T_22[9:0]) begin
        image_2_553 <= io_pixelVal_in_2_2;
      end else if (10'h229 == _T_19[9:0]) begin
        image_2_553 <= io_pixelVal_in_2_1;
      end else if (10'h229 == _T_15[9:0]) begin
        image_2_553 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_554 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22a == _T_37[9:0]) begin
        image_2_554 <= io_pixelVal_in_2_7;
      end else if (10'h22a == _T_34[9:0]) begin
        image_2_554 <= io_pixelVal_in_2_6;
      end else if (10'h22a == _T_31[9:0]) begin
        image_2_554 <= io_pixelVal_in_2_5;
      end else if (10'h22a == _T_28[9:0]) begin
        image_2_554 <= io_pixelVal_in_2_4;
      end else if (10'h22a == _T_25[9:0]) begin
        image_2_554 <= io_pixelVal_in_2_3;
      end else if (10'h22a == _T_22[9:0]) begin
        image_2_554 <= io_pixelVal_in_2_2;
      end else if (10'h22a == _T_19[9:0]) begin
        image_2_554 <= io_pixelVal_in_2_1;
      end else if (10'h22a == _T_15[9:0]) begin
        image_2_554 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_555 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22b == _T_37[9:0]) begin
        image_2_555 <= io_pixelVal_in_2_7;
      end else if (10'h22b == _T_34[9:0]) begin
        image_2_555 <= io_pixelVal_in_2_6;
      end else if (10'h22b == _T_31[9:0]) begin
        image_2_555 <= io_pixelVal_in_2_5;
      end else if (10'h22b == _T_28[9:0]) begin
        image_2_555 <= io_pixelVal_in_2_4;
      end else if (10'h22b == _T_25[9:0]) begin
        image_2_555 <= io_pixelVal_in_2_3;
      end else if (10'h22b == _T_22[9:0]) begin
        image_2_555 <= io_pixelVal_in_2_2;
      end else if (10'h22b == _T_19[9:0]) begin
        image_2_555 <= io_pixelVal_in_2_1;
      end else if (10'h22b == _T_15[9:0]) begin
        image_2_555 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_556 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22c == _T_37[9:0]) begin
        image_2_556 <= io_pixelVal_in_2_7;
      end else if (10'h22c == _T_34[9:0]) begin
        image_2_556 <= io_pixelVal_in_2_6;
      end else if (10'h22c == _T_31[9:0]) begin
        image_2_556 <= io_pixelVal_in_2_5;
      end else if (10'h22c == _T_28[9:0]) begin
        image_2_556 <= io_pixelVal_in_2_4;
      end else if (10'h22c == _T_25[9:0]) begin
        image_2_556 <= io_pixelVal_in_2_3;
      end else if (10'h22c == _T_22[9:0]) begin
        image_2_556 <= io_pixelVal_in_2_2;
      end else if (10'h22c == _T_19[9:0]) begin
        image_2_556 <= io_pixelVal_in_2_1;
      end else if (10'h22c == _T_15[9:0]) begin
        image_2_556 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_557 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22d == _T_37[9:0]) begin
        image_2_557 <= io_pixelVal_in_2_7;
      end else if (10'h22d == _T_34[9:0]) begin
        image_2_557 <= io_pixelVal_in_2_6;
      end else if (10'h22d == _T_31[9:0]) begin
        image_2_557 <= io_pixelVal_in_2_5;
      end else if (10'h22d == _T_28[9:0]) begin
        image_2_557 <= io_pixelVal_in_2_4;
      end else if (10'h22d == _T_25[9:0]) begin
        image_2_557 <= io_pixelVal_in_2_3;
      end else if (10'h22d == _T_22[9:0]) begin
        image_2_557 <= io_pixelVal_in_2_2;
      end else if (10'h22d == _T_19[9:0]) begin
        image_2_557 <= io_pixelVal_in_2_1;
      end else if (10'h22d == _T_15[9:0]) begin
        image_2_557 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_558 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22e == _T_37[9:0]) begin
        image_2_558 <= io_pixelVal_in_2_7;
      end else if (10'h22e == _T_34[9:0]) begin
        image_2_558 <= io_pixelVal_in_2_6;
      end else if (10'h22e == _T_31[9:0]) begin
        image_2_558 <= io_pixelVal_in_2_5;
      end else if (10'h22e == _T_28[9:0]) begin
        image_2_558 <= io_pixelVal_in_2_4;
      end else if (10'h22e == _T_25[9:0]) begin
        image_2_558 <= io_pixelVal_in_2_3;
      end else if (10'h22e == _T_22[9:0]) begin
        image_2_558 <= io_pixelVal_in_2_2;
      end else if (10'h22e == _T_19[9:0]) begin
        image_2_558 <= io_pixelVal_in_2_1;
      end else if (10'h22e == _T_15[9:0]) begin
        image_2_558 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_559 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22f == _T_37[9:0]) begin
        image_2_559 <= io_pixelVal_in_2_7;
      end else if (10'h22f == _T_34[9:0]) begin
        image_2_559 <= io_pixelVal_in_2_6;
      end else if (10'h22f == _T_31[9:0]) begin
        image_2_559 <= io_pixelVal_in_2_5;
      end else if (10'h22f == _T_28[9:0]) begin
        image_2_559 <= io_pixelVal_in_2_4;
      end else if (10'h22f == _T_25[9:0]) begin
        image_2_559 <= io_pixelVal_in_2_3;
      end else if (10'h22f == _T_22[9:0]) begin
        image_2_559 <= io_pixelVal_in_2_2;
      end else if (10'h22f == _T_19[9:0]) begin
        image_2_559 <= io_pixelVal_in_2_1;
      end else if (10'h22f == _T_15[9:0]) begin
        image_2_559 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_560 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h230 == _T_37[9:0]) begin
        image_2_560 <= io_pixelVal_in_2_7;
      end else if (10'h230 == _T_34[9:0]) begin
        image_2_560 <= io_pixelVal_in_2_6;
      end else if (10'h230 == _T_31[9:0]) begin
        image_2_560 <= io_pixelVal_in_2_5;
      end else if (10'h230 == _T_28[9:0]) begin
        image_2_560 <= io_pixelVal_in_2_4;
      end else if (10'h230 == _T_25[9:0]) begin
        image_2_560 <= io_pixelVal_in_2_3;
      end else if (10'h230 == _T_22[9:0]) begin
        image_2_560 <= io_pixelVal_in_2_2;
      end else if (10'h230 == _T_19[9:0]) begin
        image_2_560 <= io_pixelVal_in_2_1;
      end else if (10'h230 == _T_15[9:0]) begin
        image_2_560 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_561 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h231 == _T_37[9:0]) begin
        image_2_561 <= io_pixelVal_in_2_7;
      end else if (10'h231 == _T_34[9:0]) begin
        image_2_561 <= io_pixelVal_in_2_6;
      end else if (10'h231 == _T_31[9:0]) begin
        image_2_561 <= io_pixelVal_in_2_5;
      end else if (10'h231 == _T_28[9:0]) begin
        image_2_561 <= io_pixelVal_in_2_4;
      end else if (10'h231 == _T_25[9:0]) begin
        image_2_561 <= io_pixelVal_in_2_3;
      end else if (10'h231 == _T_22[9:0]) begin
        image_2_561 <= io_pixelVal_in_2_2;
      end else if (10'h231 == _T_19[9:0]) begin
        image_2_561 <= io_pixelVal_in_2_1;
      end else if (10'h231 == _T_15[9:0]) begin
        image_2_561 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_562 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h232 == _T_37[9:0]) begin
        image_2_562 <= io_pixelVal_in_2_7;
      end else if (10'h232 == _T_34[9:0]) begin
        image_2_562 <= io_pixelVal_in_2_6;
      end else if (10'h232 == _T_31[9:0]) begin
        image_2_562 <= io_pixelVal_in_2_5;
      end else if (10'h232 == _T_28[9:0]) begin
        image_2_562 <= io_pixelVal_in_2_4;
      end else if (10'h232 == _T_25[9:0]) begin
        image_2_562 <= io_pixelVal_in_2_3;
      end else if (10'h232 == _T_22[9:0]) begin
        image_2_562 <= io_pixelVal_in_2_2;
      end else if (10'h232 == _T_19[9:0]) begin
        image_2_562 <= io_pixelVal_in_2_1;
      end else if (10'h232 == _T_15[9:0]) begin
        image_2_562 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_563 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h233 == _T_37[9:0]) begin
        image_2_563 <= io_pixelVal_in_2_7;
      end else if (10'h233 == _T_34[9:0]) begin
        image_2_563 <= io_pixelVal_in_2_6;
      end else if (10'h233 == _T_31[9:0]) begin
        image_2_563 <= io_pixelVal_in_2_5;
      end else if (10'h233 == _T_28[9:0]) begin
        image_2_563 <= io_pixelVal_in_2_4;
      end else if (10'h233 == _T_25[9:0]) begin
        image_2_563 <= io_pixelVal_in_2_3;
      end else if (10'h233 == _T_22[9:0]) begin
        image_2_563 <= io_pixelVal_in_2_2;
      end else if (10'h233 == _T_19[9:0]) begin
        image_2_563 <= io_pixelVal_in_2_1;
      end else if (10'h233 == _T_15[9:0]) begin
        image_2_563 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_564 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h234 == _T_37[9:0]) begin
        image_2_564 <= io_pixelVal_in_2_7;
      end else if (10'h234 == _T_34[9:0]) begin
        image_2_564 <= io_pixelVal_in_2_6;
      end else if (10'h234 == _T_31[9:0]) begin
        image_2_564 <= io_pixelVal_in_2_5;
      end else if (10'h234 == _T_28[9:0]) begin
        image_2_564 <= io_pixelVal_in_2_4;
      end else if (10'h234 == _T_25[9:0]) begin
        image_2_564 <= io_pixelVal_in_2_3;
      end else if (10'h234 == _T_22[9:0]) begin
        image_2_564 <= io_pixelVal_in_2_2;
      end else if (10'h234 == _T_19[9:0]) begin
        image_2_564 <= io_pixelVal_in_2_1;
      end else if (10'h234 == _T_15[9:0]) begin
        image_2_564 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_565 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h235 == _T_37[9:0]) begin
        image_2_565 <= io_pixelVal_in_2_7;
      end else if (10'h235 == _T_34[9:0]) begin
        image_2_565 <= io_pixelVal_in_2_6;
      end else if (10'h235 == _T_31[9:0]) begin
        image_2_565 <= io_pixelVal_in_2_5;
      end else if (10'h235 == _T_28[9:0]) begin
        image_2_565 <= io_pixelVal_in_2_4;
      end else if (10'h235 == _T_25[9:0]) begin
        image_2_565 <= io_pixelVal_in_2_3;
      end else if (10'h235 == _T_22[9:0]) begin
        image_2_565 <= io_pixelVal_in_2_2;
      end else if (10'h235 == _T_19[9:0]) begin
        image_2_565 <= io_pixelVal_in_2_1;
      end else if (10'h235 == _T_15[9:0]) begin
        image_2_565 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_566 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h236 == _T_37[9:0]) begin
        image_2_566 <= io_pixelVal_in_2_7;
      end else if (10'h236 == _T_34[9:0]) begin
        image_2_566 <= io_pixelVal_in_2_6;
      end else if (10'h236 == _T_31[9:0]) begin
        image_2_566 <= io_pixelVal_in_2_5;
      end else if (10'h236 == _T_28[9:0]) begin
        image_2_566 <= io_pixelVal_in_2_4;
      end else if (10'h236 == _T_25[9:0]) begin
        image_2_566 <= io_pixelVal_in_2_3;
      end else if (10'h236 == _T_22[9:0]) begin
        image_2_566 <= io_pixelVal_in_2_2;
      end else if (10'h236 == _T_19[9:0]) begin
        image_2_566 <= io_pixelVal_in_2_1;
      end else if (10'h236 == _T_15[9:0]) begin
        image_2_566 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_567 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h237 == _T_37[9:0]) begin
        image_2_567 <= io_pixelVal_in_2_7;
      end else if (10'h237 == _T_34[9:0]) begin
        image_2_567 <= io_pixelVal_in_2_6;
      end else if (10'h237 == _T_31[9:0]) begin
        image_2_567 <= io_pixelVal_in_2_5;
      end else if (10'h237 == _T_28[9:0]) begin
        image_2_567 <= io_pixelVal_in_2_4;
      end else if (10'h237 == _T_25[9:0]) begin
        image_2_567 <= io_pixelVal_in_2_3;
      end else if (10'h237 == _T_22[9:0]) begin
        image_2_567 <= io_pixelVal_in_2_2;
      end else if (10'h237 == _T_19[9:0]) begin
        image_2_567 <= io_pixelVal_in_2_1;
      end else if (10'h237 == _T_15[9:0]) begin
        image_2_567 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_568 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h238 == _T_37[9:0]) begin
        image_2_568 <= io_pixelVal_in_2_7;
      end else if (10'h238 == _T_34[9:0]) begin
        image_2_568 <= io_pixelVal_in_2_6;
      end else if (10'h238 == _T_31[9:0]) begin
        image_2_568 <= io_pixelVal_in_2_5;
      end else if (10'h238 == _T_28[9:0]) begin
        image_2_568 <= io_pixelVal_in_2_4;
      end else if (10'h238 == _T_25[9:0]) begin
        image_2_568 <= io_pixelVal_in_2_3;
      end else if (10'h238 == _T_22[9:0]) begin
        image_2_568 <= io_pixelVal_in_2_2;
      end else if (10'h238 == _T_19[9:0]) begin
        image_2_568 <= io_pixelVal_in_2_1;
      end else if (10'h238 == _T_15[9:0]) begin
        image_2_568 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_569 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h239 == _T_37[9:0]) begin
        image_2_569 <= io_pixelVal_in_2_7;
      end else if (10'h239 == _T_34[9:0]) begin
        image_2_569 <= io_pixelVal_in_2_6;
      end else if (10'h239 == _T_31[9:0]) begin
        image_2_569 <= io_pixelVal_in_2_5;
      end else if (10'h239 == _T_28[9:0]) begin
        image_2_569 <= io_pixelVal_in_2_4;
      end else if (10'h239 == _T_25[9:0]) begin
        image_2_569 <= io_pixelVal_in_2_3;
      end else if (10'h239 == _T_22[9:0]) begin
        image_2_569 <= io_pixelVal_in_2_2;
      end else if (10'h239 == _T_19[9:0]) begin
        image_2_569 <= io_pixelVal_in_2_1;
      end else if (10'h239 == _T_15[9:0]) begin
        image_2_569 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_570 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23a == _T_37[9:0]) begin
        image_2_570 <= io_pixelVal_in_2_7;
      end else if (10'h23a == _T_34[9:0]) begin
        image_2_570 <= io_pixelVal_in_2_6;
      end else if (10'h23a == _T_31[9:0]) begin
        image_2_570 <= io_pixelVal_in_2_5;
      end else if (10'h23a == _T_28[9:0]) begin
        image_2_570 <= io_pixelVal_in_2_4;
      end else if (10'h23a == _T_25[9:0]) begin
        image_2_570 <= io_pixelVal_in_2_3;
      end else if (10'h23a == _T_22[9:0]) begin
        image_2_570 <= io_pixelVal_in_2_2;
      end else if (10'h23a == _T_19[9:0]) begin
        image_2_570 <= io_pixelVal_in_2_1;
      end else if (10'h23a == _T_15[9:0]) begin
        image_2_570 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_571 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23b == _T_37[9:0]) begin
        image_2_571 <= io_pixelVal_in_2_7;
      end else if (10'h23b == _T_34[9:0]) begin
        image_2_571 <= io_pixelVal_in_2_6;
      end else if (10'h23b == _T_31[9:0]) begin
        image_2_571 <= io_pixelVal_in_2_5;
      end else if (10'h23b == _T_28[9:0]) begin
        image_2_571 <= io_pixelVal_in_2_4;
      end else if (10'h23b == _T_25[9:0]) begin
        image_2_571 <= io_pixelVal_in_2_3;
      end else if (10'h23b == _T_22[9:0]) begin
        image_2_571 <= io_pixelVal_in_2_2;
      end else if (10'h23b == _T_19[9:0]) begin
        image_2_571 <= io_pixelVal_in_2_1;
      end else if (10'h23b == _T_15[9:0]) begin
        image_2_571 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_572 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23c == _T_37[9:0]) begin
        image_2_572 <= io_pixelVal_in_2_7;
      end else if (10'h23c == _T_34[9:0]) begin
        image_2_572 <= io_pixelVal_in_2_6;
      end else if (10'h23c == _T_31[9:0]) begin
        image_2_572 <= io_pixelVal_in_2_5;
      end else if (10'h23c == _T_28[9:0]) begin
        image_2_572 <= io_pixelVal_in_2_4;
      end else if (10'h23c == _T_25[9:0]) begin
        image_2_572 <= io_pixelVal_in_2_3;
      end else if (10'h23c == _T_22[9:0]) begin
        image_2_572 <= io_pixelVal_in_2_2;
      end else if (10'h23c == _T_19[9:0]) begin
        image_2_572 <= io_pixelVal_in_2_1;
      end else if (10'h23c == _T_15[9:0]) begin
        image_2_572 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_573 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23d == _T_37[9:0]) begin
        image_2_573 <= io_pixelVal_in_2_7;
      end else if (10'h23d == _T_34[9:0]) begin
        image_2_573 <= io_pixelVal_in_2_6;
      end else if (10'h23d == _T_31[9:0]) begin
        image_2_573 <= io_pixelVal_in_2_5;
      end else if (10'h23d == _T_28[9:0]) begin
        image_2_573 <= io_pixelVal_in_2_4;
      end else if (10'h23d == _T_25[9:0]) begin
        image_2_573 <= io_pixelVal_in_2_3;
      end else if (10'h23d == _T_22[9:0]) begin
        image_2_573 <= io_pixelVal_in_2_2;
      end else if (10'h23d == _T_19[9:0]) begin
        image_2_573 <= io_pixelVal_in_2_1;
      end else if (10'h23d == _T_15[9:0]) begin
        image_2_573 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_574 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23e == _T_37[9:0]) begin
        image_2_574 <= io_pixelVal_in_2_7;
      end else if (10'h23e == _T_34[9:0]) begin
        image_2_574 <= io_pixelVal_in_2_6;
      end else if (10'h23e == _T_31[9:0]) begin
        image_2_574 <= io_pixelVal_in_2_5;
      end else if (10'h23e == _T_28[9:0]) begin
        image_2_574 <= io_pixelVal_in_2_4;
      end else if (10'h23e == _T_25[9:0]) begin
        image_2_574 <= io_pixelVal_in_2_3;
      end else if (10'h23e == _T_22[9:0]) begin
        image_2_574 <= io_pixelVal_in_2_2;
      end else if (10'h23e == _T_19[9:0]) begin
        image_2_574 <= io_pixelVal_in_2_1;
      end else if (10'h23e == _T_15[9:0]) begin
        image_2_574 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_575 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23f == _T_37[9:0]) begin
        image_2_575 <= io_pixelVal_in_2_7;
      end else if (10'h23f == _T_34[9:0]) begin
        image_2_575 <= io_pixelVal_in_2_6;
      end else if (10'h23f == _T_31[9:0]) begin
        image_2_575 <= io_pixelVal_in_2_5;
      end else if (10'h23f == _T_28[9:0]) begin
        image_2_575 <= io_pixelVal_in_2_4;
      end else if (10'h23f == _T_25[9:0]) begin
        image_2_575 <= io_pixelVal_in_2_3;
      end else if (10'h23f == _T_22[9:0]) begin
        image_2_575 <= io_pixelVal_in_2_2;
      end else if (10'h23f == _T_19[9:0]) begin
        image_2_575 <= io_pixelVal_in_2_1;
      end else if (10'h23f == _T_15[9:0]) begin
        image_2_575 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      pixelIndex <= 32'h0;
    end else if (io_valid_in) begin
      if (_T_90) begin
        pixelIndex <= 32'h0;
      end else begin
        pixelIndex <= _T_88;
      end
    end
  end
endmodule
module ImageProcessing(
  input         clock,
  input         reset,
  input  [5:0]  io_SPI_filterIndex,
  input         io_SPI_invert,
  input         io_SPI_distort,
  input  [10:0] io_rowIndex,
  input  [10:0] io_colIndex,
  output [3:0]  io_pixelVal_out_0,
  output [3:0]  io_pixelVal_out_1,
  output [3:0]  io_pixelVal_out_2
);
  wire  filter_clock; // @[ImageProcessing.scala 23:22]
  wire  filter_reset; // @[ImageProcessing.scala 23:22]
  wire [5:0] filter_io_SPI_filterIndex; // @[ImageProcessing.scala 23:22]
  wire  filter_io_SPI_distort; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_0; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_1; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_2; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_3; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_4; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_5; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_6; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_7; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_0; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_1; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_2; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_3; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_4; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_5; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_6; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_7; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_0; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_1; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_2; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_3; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_4; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_5; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_6; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_7; // @[ImageProcessing.scala 23:22]
  wire  filter_io_valid_out; // @[ImageProcessing.scala 23:22]
  wire  videoBuffer_clock; // @[ImageProcessing.scala 24:27]
  wire  videoBuffer_reset; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_0; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_1; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_2; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_3; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_4; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_5; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_6; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_7; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_0; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_1; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_2; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_3; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_4; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_5; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_6; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_7; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_0; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_1; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_2; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_3; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_4; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_5; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_6; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_7; // @[ImageProcessing.scala 24:27]
  wire  videoBuffer_io_valid_in; // @[ImageProcessing.scala 24:27]
  wire [10:0] videoBuffer_io_rowIndex; // @[ImageProcessing.scala 24:27]
  wire [10:0] videoBuffer_io_colIndex; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_out_0; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_out_1; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_out_2; // @[ImageProcessing.scala 24:27]
  Filter filter ( // @[ImageProcessing.scala 23:22]
    .clock(filter_clock),
    .reset(filter_reset),
    .io_SPI_filterIndex(filter_io_SPI_filterIndex),
    .io_SPI_distort(filter_io_SPI_distort),
    .io_pixelVal_out_0_0(filter_io_pixelVal_out_0_0),
    .io_pixelVal_out_0_1(filter_io_pixelVal_out_0_1),
    .io_pixelVal_out_0_2(filter_io_pixelVal_out_0_2),
    .io_pixelVal_out_0_3(filter_io_pixelVal_out_0_3),
    .io_pixelVal_out_0_4(filter_io_pixelVal_out_0_4),
    .io_pixelVal_out_0_5(filter_io_pixelVal_out_0_5),
    .io_pixelVal_out_0_6(filter_io_pixelVal_out_0_6),
    .io_pixelVal_out_0_7(filter_io_pixelVal_out_0_7),
    .io_pixelVal_out_1_0(filter_io_pixelVal_out_1_0),
    .io_pixelVal_out_1_1(filter_io_pixelVal_out_1_1),
    .io_pixelVal_out_1_2(filter_io_pixelVal_out_1_2),
    .io_pixelVal_out_1_3(filter_io_pixelVal_out_1_3),
    .io_pixelVal_out_1_4(filter_io_pixelVal_out_1_4),
    .io_pixelVal_out_1_5(filter_io_pixelVal_out_1_5),
    .io_pixelVal_out_1_6(filter_io_pixelVal_out_1_6),
    .io_pixelVal_out_1_7(filter_io_pixelVal_out_1_7),
    .io_pixelVal_out_2_0(filter_io_pixelVal_out_2_0),
    .io_pixelVal_out_2_1(filter_io_pixelVal_out_2_1),
    .io_pixelVal_out_2_2(filter_io_pixelVal_out_2_2),
    .io_pixelVal_out_2_3(filter_io_pixelVal_out_2_3),
    .io_pixelVal_out_2_4(filter_io_pixelVal_out_2_4),
    .io_pixelVal_out_2_5(filter_io_pixelVal_out_2_5),
    .io_pixelVal_out_2_6(filter_io_pixelVal_out_2_6),
    .io_pixelVal_out_2_7(filter_io_pixelVal_out_2_7),
    .io_valid_out(filter_io_valid_out)
  );
  VideoBuffer videoBuffer ( // @[ImageProcessing.scala 24:27]
    .clock(videoBuffer_clock),
    .reset(videoBuffer_reset),
    .io_pixelVal_in_0_0(videoBuffer_io_pixelVal_in_0_0),
    .io_pixelVal_in_0_1(videoBuffer_io_pixelVal_in_0_1),
    .io_pixelVal_in_0_2(videoBuffer_io_pixelVal_in_0_2),
    .io_pixelVal_in_0_3(videoBuffer_io_pixelVal_in_0_3),
    .io_pixelVal_in_0_4(videoBuffer_io_pixelVal_in_0_4),
    .io_pixelVal_in_0_5(videoBuffer_io_pixelVal_in_0_5),
    .io_pixelVal_in_0_6(videoBuffer_io_pixelVal_in_0_6),
    .io_pixelVal_in_0_7(videoBuffer_io_pixelVal_in_0_7),
    .io_pixelVal_in_1_0(videoBuffer_io_pixelVal_in_1_0),
    .io_pixelVal_in_1_1(videoBuffer_io_pixelVal_in_1_1),
    .io_pixelVal_in_1_2(videoBuffer_io_pixelVal_in_1_2),
    .io_pixelVal_in_1_3(videoBuffer_io_pixelVal_in_1_3),
    .io_pixelVal_in_1_4(videoBuffer_io_pixelVal_in_1_4),
    .io_pixelVal_in_1_5(videoBuffer_io_pixelVal_in_1_5),
    .io_pixelVal_in_1_6(videoBuffer_io_pixelVal_in_1_6),
    .io_pixelVal_in_1_7(videoBuffer_io_pixelVal_in_1_7),
    .io_pixelVal_in_2_0(videoBuffer_io_pixelVal_in_2_0),
    .io_pixelVal_in_2_1(videoBuffer_io_pixelVal_in_2_1),
    .io_pixelVal_in_2_2(videoBuffer_io_pixelVal_in_2_2),
    .io_pixelVal_in_2_3(videoBuffer_io_pixelVal_in_2_3),
    .io_pixelVal_in_2_4(videoBuffer_io_pixelVal_in_2_4),
    .io_pixelVal_in_2_5(videoBuffer_io_pixelVal_in_2_5),
    .io_pixelVal_in_2_6(videoBuffer_io_pixelVal_in_2_6),
    .io_pixelVal_in_2_7(videoBuffer_io_pixelVal_in_2_7),
    .io_valid_in(videoBuffer_io_valid_in),
    .io_rowIndex(videoBuffer_io_rowIndex),
    .io_colIndex(videoBuffer_io_colIndex),
    .io_pixelVal_out_0(videoBuffer_io_pixelVal_out_0),
    .io_pixelVal_out_1(videoBuffer_io_pixelVal_out_1),
    .io_pixelVal_out_2(videoBuffer_io_pixelVal_out_2)
  );
  assign io_pixelVal_out_0 = videoBuffer_io_pixelVal_out_0; // @[ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25]
  assign io_pixelVal_out_1 = videoBuffer_io_pixelVal_out_1; // @[ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25]
  assign io_pixelVal_out_2 = videoBuffer_io_pixelVal_out_2; // @[ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25]
  assign filter_clock = clock;
  assign filter_reset = reset;
  assign filter_io_SPI_filterIndex = io_SPI_filterIndex; // @[ImageProcessing.scala 29:29]
  assign filter_io_SPI_distort = io_SPI_distort; // @[ImageProcessing.scala 31:29]
  assign videoBuffer_clock = clock;
  assign videoBuffer_reset = reset;
  assign videoBuffer_io_pixelVal_in_0_0 = filter_io_pixelVal_out_0_0; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_1 = filter_io_pixelVal_out_0_1; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_2 = filter_io_pixelVal_out_0_2; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_3 = filter_io_pixelVal_out_0_3; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_4 = filter_io_pixelVal_out_0_4; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_5 = filter_io_pixelVal_out_0_5; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_6 = filter_io_pixelVal_out_0_6; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_7 = filter_io_pixelVal_out_0_7; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_0 = filter_io_pixelVal_out_1_0; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_1 = filter_io_pixelVal_out_1_1; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_2 = filter_io_pixelVal_out_1_2; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_3 = filter_io_pixelVal_out_1_3; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_4 = filter_io_pixelVal_out_1_4; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_5 = filter_io_pixelVal_out_1_5; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_6 = filter_io_pixelVal_out_1_6; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_7 = filter_io_pixelVal_out_1_7; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_0 = filter_io_pixelVal_out_2_0; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_1 = filter_io_pixelVal_out_2_1; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_2 = filter_io_pixelVal_out_2_2; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_3 = filter_io_pixelVal_out_2_3; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_4 = filter_io_pixelVal_out_2_4; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_5 = filter_io_pixelVal_out_2_5; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_6 = filter_io_pixelVal_out_2_6; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_7 = filter_io_pixelVal_out_2_7; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_valid_in = filter_io_valid_out; // @[ImageProcessing.scala 39:27]
  assign videoBuffer_io_rowIndex = io_rowIndex; // @[ImageProcessing.scala 26:27]
  assign videoBuffer_io_colIndex = io_colIndex; // @[ImageProcessing.scala 27:27]
endmodule
