module DotProd(
  input        clock,
  input        reset,
  input  [7:0] io_dataInA,
  input  [7:0] io_dataInB,
  output [8:0] io_dataOut,
  output       io_outputValid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] countVal; // @[Counter.scala 29:33]
  wire  countReset = countVal == 4'h8; // @[Counter.scala 38:24]
  wire [3:0] _T_2 = countVal + 4'h1; // @[Counter.scala 39:22]
  reg [8:0] accumulator; // @[DotProd.scala 19:28]
  wire [15:0] product = $signed(io_dataInA) * $signed(io_dataInB); // @[DotProd.scala 20:35]
  wire [15:0] _GEN_5 = {{7{accumulator[8]}},accumulator}; // @[DotProd.scala 21:30]
  wire [15:0] _T_6 = $signed(_GEN_5) + $signed(product); // @[DotProd.scala 21:30]
  wire [15:0] _GEN_4 = countReset ? $signed(16'sh0) : $signed(_T_6); // @[DotProd.scala 25:20]
  assign io_dataOut = _T_6[8:0]; // @[DotProd.scala 23:14]
  assign io_outputValid = countVal == 4'h8; // @[DotProd.scala 26:20 DotProd.scala 29:20]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  countVal = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  accumulator = _RAND_1[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      countVal <= 4'h0;
    end else if (countReset) begin
      countVal <= 4'h0;
    end else begin
      countVal <= _T_2;
    end
    if (reset) begin
      accumulator <= 9'sh0;
    end else begin
      accumulator <= _GEN_4[8:0];
    end
  end
endmodule
module KernelConvolution(
  input        clock,
  input        reset,
  input  [4:0] io_kernelVal_in,
  input  [3:0] io_pixelVal_in_0,
  input  [3:0] io_pixelVal_in_1,
  input  [3:0] io_pixelVal_in_2,
  input  [3:0] io_pixelVal_in_3,
  input  [3:0] io_pixelVal_in_4,
  input  [3:0] io_pixelVal_in_5,
  input  [3:0] io_pixelVal_in_6,
  output [8:0] io_pixelVal_out_0,
  output [8:0] io_pixelVal_out_1,
  output [8:0] io_pixelVal_out_2,
  output [8:0] io_pixelVal_out_3,
  output [8:0] io_pixelVal_out_4,
  output [8:0] io_pixelVal_out_5,
  output [8:0] io_pixelVal_out_6,
  output       io_valid_out
);
  wire  DotProd_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_1_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_1_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_1_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_1_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_1_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_1_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_2_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_2_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_2_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_2_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_2_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_2_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_3_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_3_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_3_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_3_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_3_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_3_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_4_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_4_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_4_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_4_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_4_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_4_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_5_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_5_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_5_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_5_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_5_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_5_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_6_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_6_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_6_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_6_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_6_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_6_io_outputValid; // @[KernelConvolution.scala 21:58]
  DotProd DotProd ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_clock),
    .reset(DotProd_reset),
    .io_dataInA(DotProd_io_dataInA),
    .io_dataInB(DotProd_io_dataInB),
    .io_dataOut(DotProd_io_dataOut),
    .io_outputValid(DotProd_io_outputValid)
  );
  DotProd DotProd_1 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_1_clock),
    .reset(DotProd_1_reset),
    .io_dataInA(DotProd_1_io_dataInA),
    .io_dataInB(DotProd_1_io_dataInB),
    .io_dataOut(DotProd_1_io_dataOut),
    .io_outputValid(DotProd_1_io_outputValid)
  );
  DotProd DotProd_2 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_2_clock),
    .reset(DotProd_2_reset),
    .io_dataInA(DotProd_2_io_dataInA),
    .io_dataInB(DotProd_2_io_dataInB),
    .io_dataOut(DotProd_2_io_dataOut),
    .io_outputValid(DotProd_2_io_outputValid)
  );
  DotProd DotProd_3 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_3_clock),
    .reset(DotProd_3_reset),
    .io_dataInA(DotProd_3_io_dataInA),
    .io_dataInB(DotProd_3_io_dataInB),
    .io_dataOut(DotProd_3_io_dataOut),
    .io_outputValid(DotProd_3_io_outputValid)
  );
  DotProd DotProd_4 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_4_clock),
    .reset(DotProd_4_reset),
    .io_dataInA(DotProd_4_io_dataInA),
    .io_dataInB(DotProd_4_io_dataInB),
    .io_dataOut(DotProd_4_io_dataOut),
    .io_outputValid(DotProd_4_io_outputValid)
  );
  DotProd DotProd_5 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_5_clock),
    .reset(DotProd_5_reset),
    .io_dataInA(DotProd_5_io_dataInA),
    .io_dataInB(DotProd_5_io_dataInB),
    .io_dataOut(DotProd_5_io_dataOut),
    .io_outputValid(DotProd_5_io_outputValid)
  );
  DotProd DotProd_6 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_6_clock),
    .reset(DotProd_6_reset),
    .io_dataInA(DotProd_6_io_dataInA),
    .io_dataInB(DotProd_6_io_dataInB),
    .io_dataOut(DotProd_6_io_dataOut),
    .io_outputValid(DotProd_6_io_outputValid)
  );
  assign io_pixelVal_out_0 = DotProd_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_1 = DotProd_1_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_2 = DotProd_2_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_3 = DotProd_3_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_4 = DotProd_4_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_5 = DotProd_5_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_6 = DotProd_6_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_valid_out = DotProd_io_outputValid; // @[KernelConvolution.scala 35:30]
  assign DotProd_clock = clock;
  assign DotProd_reset = reset;
  assign DotProd_io_dataInA = {{4'd0}, io_pixelVal_in_0}; // @[KernelConvolution.scala 21:32]
  assign DotProd_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_1_clock = clock;
  assign DotProd_1_reset = reset;
  assign DotProd_1_io_dataInA = {{4'd0}, io_pixelVal_in_1}; // @[KernelConvolution.scala 21:32]
  assign DotProd_1_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_2_clock = clock;
  assign DotProd_2_reset = reset;
  assign DotProd_2_io_dataInA = {{4'd0}, io_pixelVal_in_2}; // @[KernelConvolution.scala 21:32]
  assign DotProd_2_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_3_clock = clock;
  assign DotProd_3_reset = reset;
  assign DotProd_3_io_dataInA = {{4'd0}, io_pixelVal_in_3}; // @[KernelConvolution.scala 21:32]
  assign DotProd_3_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_4_clock = clock;
  assign DotProd_4_reset = reset;
  assign DotProd_4_io_dataInA = {{4'd0}, io_pixelVal_in_4}; // @[KernelConvolution.scala 21:32]
  assign DotProd_4_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_5_clock = clock;
  assign DotProd_5_reset = reset;
  assign DotProd_5_io_dataInA = {{4'd0}, io_pixelVal_in_5}; // @[KernelConvolution.scala 21:32]
  assign DotProd_5_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_6_clock = clock;
  assign DotProd_6_reset = reset;
  assign DotProd_6_io_dataInA = {{4'd0}, io_pixelVal_in_6}; // @[KernelConvolution.scala 21:32]
  assign DotProd_6_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
endmodule
module Filter(
  input        clock,
  input        reset,
  input  [5:0] io_SPI_filterIndex,
  input        io_SPI_invert,
  input        io_SPI_distort,
  output [3:0] io_pixelVal_out_0_0,
  output [3:0] io_pixelVal_out_0_1,
  output [3:0] io_pixelVal_out_0_2,
  output [3:0] io_pixelVal_out_0_3,
  output [3:0] io_pixelVal_out_0_4,
  output [3:0] io_pixelVal_out_0_5,
  output [3:0] io_pixelVal_out_0_6,
  output [3:0] io_pixelVal_out_1_0,
  output [3:0] io_pixelVal_out_1_1,
  output [3:0] io_pixelVal_out_1_2,
  output [3:0] io_pixelVal_out_1_3,
  output [3:0] io_pixelVal_out_1_4,
  output [3:0] io_pixelVal_out_1_5,
  output [3:0] io_pixelVal_out_1_6,
  output [3:0] io_pixelVal_out_2_0,
  output [3:0] io_pixelVal_out_2_1,
  output [3:0] io_pixelVal_out_2_2,
  output [3:0] io_pixelVal_out_2_3,
  output [3:0] io_pixelVal_out_2_4,
  output [3:0] io_pixelVal_out_2_5,
  output [3:0] io_pixelVal_out_2_6,
  output       io_valid_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
`endif // RANDOMIZE_REG_INIT
  wire  KernelConvolution_clock; // @[Filter.scala 186:36]
  wire  KernelConvolution_reset; // @[Filter.scala 186:36]
  wire [4:0] KernelConvolution_io_kernelVal_in; // @[Filter.scala 186:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_0; // @[Filter.scala 186:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_1; // @[Filter.scala 186:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_2; // @[Filter.scala 186:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_3; // @[Filter.scala 186:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_4; // @[Filter.scala 186:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_5; // @[Filter.scala 186:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_6; // @[Filter.scala 186:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_0; // @[Filter.scala 186:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_1; // @[Filter.scala 186:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_2; // @[Filter.scala 186:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_3; // @[Filter.scala 186:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_4; // @[Filter.scala 186:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_5; // @[Filter.scala 186:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_6; // @[Filter.scala 186:36]
  wire  KernelConvolution_io_valid_out; // @[Filter.scala 186:36]
  wire  KernelConvolution_1_clock; // @[Filter.scala 187:36]
  wire  KernelConvolution_1_reset; // @[Filter.scala 187:36]
  wire [4:0] KernelConvolution_1_io_kernelVal_in; // @[Filter.scala 187:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_0; // @[Filter.scala 187:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_1; // @[Filter.scala 187:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_2; // @[Filter.scala 187:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_3; // @[Filter.scala 187:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_4; // @[Filter.scala 187:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_5; // @[Filter.scala 187:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_6; // @[Filter.scala 187:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_0; // @[Filter.scala 187:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_1; // @[Filter.scala 187:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_2; // @[Filter.scala 187:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_3; // @[Filter.scala 187:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_4; // @[Filter.scala 187:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_5; // @[Filter.scala 187:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_6; // @[Filter.scala 187:36]
  wire  KernelConvolution_1_io_valid_out; // @[Filter.scala 187:36]
  wire  KernelConvolution_2_clock; // @[Filter.scala 188:36]
  wire  KernelConvolution_2_reset; // @[Filter.scala 188:36]
  wire [4:0] KernelConvolution_2_io_kernelVal_in; // @[Filter.scala 188:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_0; // @[Filter.scala 188:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_1; // @[Filter.scala 188:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_2; // @[Filter.scala 188:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_3; // @[Filter.scala 188:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_4; // @[Filter.scala 188:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_5; // @[Filter.scala 188:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_6; // @[Filter.scala 188:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_0; // @[Filter.scala 188:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_1; // @[Filter.scala 188:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_2; // @[Filter.scala 188:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_3; // @[Filter.scala 188:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_4; // @[Filter.scala 188:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_5; // @[Filter.scala 188:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_6; // @[Filter.scala 188:36]
  wire  KernelConvolution_2_io_valid_out; // @[Filter.scala 188:36]
  reg [3:0] kernelCounter; // @[Counter.scala 29:33]
  wire  kernelCountReset = kernelCounter == 4'h8; // @[Counter.scala 38:24]
  wire [3:0] _T_14 = kernelCounter + 4'h1; // @[Counter.scala 39:22]
  wire  _GEN_10910 = 3'h0 == io_SPI_filterIndex[2:0]; // @[Filter.scala 194:41]
  wire  _GEN_10911 = 4'h4 == kernelCounter; // @[Filter.scala 194:41]
  wire [4:0] _GEN_7 = _GEN_10910 & _GEN_10911 ? $signed(5'sh1) : $signed(5'sh0); // @[Filter.scala 194:41]
  wire  _GEN_10913 = 4'h5 == kernelCounter; // @[Filter.scala 194:41]
  wire [4:0] _GEN_8 = _GEN_10910 & _GEN_10913 ? $signed(5'sh0) : $signed(_GEN_7); // @[Filter.scala 194:41]
  wire  _GEN_10915 = 4'h6 == kernelCounter; // @[Filter.scala 194:41]
  wire [4:0] _GEN_9 = _GEN_10910 & _GEN_10915 ? $signed(5'sh0) : $signed(_GEN_8); // @[Filter.scala 194:41]
  wire  _GEN_10917 = 4'h7 == kernelCounter; // @[Filter.scala 194:41]
  wire [4:0] _GEN_10 = _GEN_10910 & _GEN_10917 ? $signed(5'sh0) : $signed(_GEN_9); // @[Filter.scala 194:41]
  wire  _GEN_10919 = 4'h8 == kernelCounter; // @[Filter.scala 194:41]
  wire [4:0] _GEN_11 = _GEN_10910 & _GEN_10919 ? $signed(5'sh0) : $signed(_GEN_10); // @[Filter.scala 194:41]
  wire  _GEN_10920 = 3'h1 == io_SPI_filterIndex[2:0]; // @[Filter.scala 194:41]
  wire  _GEN_10921 = 4'h0 == kernelCounter; // @[Filter.scala 194:41]
  wire [4:0] _GEN_12 = _GEN_10920 & _GEN_10921 ? $signed(5'sh1) : $signed(_GEN_11); // @[Filter.scala 194:41]
  wire  _GEN_10923 = 4'h1 == kernelCounter; // @[Filter.scala 194:41]
  wire [4:0] _GEN_13 = _GEN_10920 & _GEN_10923 ? $signed(5'sh1) : $signed(_GEN_12); // @[Filter.scala 194:41]
  wire  _GEN_10925 = 4'h2 == kernelCounter; // @[Filter.scala 194:41]
  wire [4:0] _GEN_14 = _GEN_10920 & _GEN_10925 ? $signed(5'sh1) : $signed(_GEN_13); // @[Filter.scala 194:41]
  wire  _GEN_10927 = 4'h3 == kernelCounter; // @[Filter.scala 194:41]
  wire [4:0] _GEN_15 = _GEN_10920 & _GEN_10927 ? $signed(5'sh1) : $signed(_GEN_14); // @[Filter.scala 194:41]
  wire [4:0] _GEN_16 = _GEN_10920 & _GEN_10911 ? $signed(5'sh1) : $signed(_GEN_15); // @[Filter.scala 194:41]
  wire [4:0] _GEN_17 = _GEN_10920 & _GEN_10913 ? $signed(5'sh1) : $signed(_GEN_16); // @[Filter.scala 194:41]
  wire [4:0] _GEN_18 = _GEN_10920 & _GEN_10915 ? $signed(5'sh1) : $signed(_GEN_17); // @[Filter.scala 194:41]
  wire [4:0] _GEN_19 = _GEN_10920 & _GEN_10917 ? $signed(5'sh1) : $signed(_GEN_18); // @[Filter.scala 194:41]
  wire [4:0] _GEN_20 = _GEN_10920 & _GEN_10919 ? $signed(5'sh1) : $signed(_GEN_19); // @[Filter.scala 194:41]
  wire  _GEN_10938 = 3'h2 == io_SPI_filterIndex[2:0]; // @[Filter.scala 194:41]
  wire [4:0] _GEN_21 = _GEN_10938 & _GEN_10921 ? $signed(5'sh1) : $signed(_GEN_20); // @[Filter.scala 194:41]
  wire [4:0] _GEN_22 = _GEN_10938 & _GEN_10923 ? $signed(5'sh2) : $signed(_GEN_21); // @[Filter.scala 194:41]
  wire [4:0] _GEN_23 = _GEN_10938 & _GEN_10925 ? $signed(5'sh1) : $signed(_GEN_22); // @[Filter.scala 194:41]
  wire [4:0] _GEN_24 = _GEN_10938 & _GEN_10927 ? $signed(5'sh2) : $signed(_GEN_23); // @[Filter.scala 194:41]
  wire [4:0] _GEN_25 = _GEN_10938 & _GEN_10911 ? $signed(5'sh4) : $signed(_GEN_24); // @[Filter.scala 194:41]
  wire [4:0] _GEN_26 = _GEN_10938 & _GEN_10913 ? $signed(5'sh2) : $signed(_GEN_25); // @[Filter.scala 194:41]
  wire [4:0] _GEN_27 = _GEN_10938 & _GEN_10915 ? $signed(5'sh1) : $signed(_GEN_26); // @[Filter.scala 194:41]
  wire [4:0] _GEN_28 = _GEN_10938 & _GEN_10917 ? $signed(5'sh2) : $signed(_GEN_27); // @[Filter.scala 194:41]
  wire [4:0] _GEN_29 = _GEN_10938 & _GEN_10919 ? $signed(5'sh1) : $signed(_GEN_28); // @[Filter.scala 194:41]
  wire  _GEN_10956 = 3'h3 == io_SPI_filterIndex[2:0]; // @[Filter.scala 194:41]
  wire [4:0] _GEN_30 = _GEN_10956 & _GEN_10921 ? $signed(5'sh0) : $signed(_GEN_29); // @[Filter.scala 194:41]
  wire [4:0] _GEN_31 = _GEN_10956 & _GEN_10923 ? $signed(-5'sh1) : $signed(_GEN_30); // @[Filter.scala 194:41]
  wire [4:0] _GEN_32 = _GEN_10956 & _GEN_10925 ? $signed(5'sh0) : $signed(_GEN_31); // @[Filter.scala 194:41]
  wire [4:0] _GEN_33 = _GEN_10956 & _GEN_10927 ? $signed(-5'sh1) : $signed(_GEN_32); // @[Filter.scala 194:41]
  wire [4:0] _GEN_34 = _GEN_10956 & _GEN_10911 ? $signed(5'sh4) : $signed(_GEN_33); // @[Filter.scala 194:41]
  wire [4:0] _GEN_35 = _GEN_10956 & _GEN_10913 ? $signed(-5'sh1) : $signed(_GEN_34); // @[Filter.scala 194:41]
  wire [4:0] _GEN_36 = _GEN_10956 & _GEN_10915 ? $signed(5'sh0) : $signed(_GEN_35); // @[Filter.scala 194:41]
  wire [4:0] _GEN_37 = _GEN_10956 & _GEN_10917 ? $signed(-5'sh1) : $signed(_GEN_36); // @[Filter.scala 194:41]
  wire [4:0] _GEN_38 = _GEN_10956 & _GEN_10919 ? $signed(5'sh0) : $signed(_GEN_37); // @[Filter.scala 194:41]
  wire  _GEN_10974 = 3'h4 == io_SPI_filterIndex[2:0]; // @[Filter.scala 194:41]
  wire [4:0] _GEN_39 = _GEN_10974 & _GEN_10921 ? $signed(-5'sh1) : $signed(_GEN_38); // @[Filter.scala 194:41]
  wire [4:0] _GEN_40 = _GEN_10974 & _GEN_10923 ? $signed(-5'sh1) : $signed(_GEN_39); // @[Filter.scala 194:41]
  wire [4:0] _GEN_41 = _GEN_10974 & _GEN_10925 ? $signed(-5'sh1) : $signed(_GEN_40); // @[Filter.scala 194:41]
  wire [4:0] _GEN_42 = _GEN_10974 & _GEN_10927 ? $signed(-5'sh1) : $signed(_GEN_41); // @[Filter.scala 194:41]
  wire [4:0] _GEN_43 = _GEN_10974 & _GEN_10911 ? $signed(5'sh8) : $signed(_GEN_42); // @[Filter.scala 194:41]
  wire [4:0] _GEN_44 = _GEN_10974 & _GEN_10913 ? $signed(-5'sh1) : $signed(_GEN_43); // @[Filter.scala 194:41]
  wire [4:0] _GEN_45 = _GEN_10974 & _GEN_10915 ? $signed(-5'sh1) : $signed(_GEN_44); // @[Filter.scala 194:41]
  wire [4:0] _GEN_46 = _GEN_10974 & _GEN_10917 ? $signed(-5'sh1) : $signed(_GEN_45); // @[Filter.scala 194:41]
  wire [4:0] _GEN_47 = _GEN_10974 & _GEN_10919 ? $signed(-5'sh1) : $signed(_GEN_46); // @[Filter.scala 194:41]
  wire  _GEN_10992 = 3'h5 == io_SPI_filterIndex[2:0]; // @[Filter.scala 194:41]
  wire [4:0] _GEN_48 = _GEN_10992 & _GEN_10921 ? $signed(5'sh0) : $signed(_GEN_47); // @[Filter.scala 194:41]
  wire [4:0] _GEN_49 = _GEN_10992 & _GEN_10923 ? $signed(-5'sh1) : $signed(_GEN_48); // @[Filter.scala 194:41]
  wire [4:0] _GEN_50 = _GEN_10992 & _GEN_10925 ? $signed(5'sh0) : $signed(_GEN_49); // @[Filter.scala 194:41]
  wire [4:0] _GEN_51 = _GEN_10992 & _GEN_10927 ? $signed(-5'sh1) : $signed(_GEN_50); // @[Filter.scala 194:41]
  wire [4:0] _GEN_52 = _GEN_10992 & _GEN_10911 ? $signed(5'sh5) : $signed(_GEN_51); // @[Filter.scala 194:41]
  wire [4:0] _GEN_53 = _GEN_10992 & _GEN_10913 ? $signed(-5'sh1) : $signed(_GEN_52); // @[Filter.scala 194:41]
  wire [4:0] _GEN_54 = _GEN_10992 & _GEN_10915 ? $signed(5'sh0) : $signed(_GEN_53); // @[Filter.scala 194:41]
  wire [4:0] _GEN_55 = _GEN_10992 & _GEN_10917 ? $signed(-5'sh1) : $signed(_GEN_54); // @[Filter.scala 194:41]
  reg [1:0] imageCounterX; // @[Counter.scala 29:33]
  wire  imageCounterXReset = imageCounterX == 2'h2; // @[Counter.scala 38:24]
  wire [1:0] _T_20 = imageCounterX + 2'h1; // @[Counter.scala 39:22]
  reg [1:0] imageCounterY; // @[Counter.scala 29:33]
  wire  _T_21 = imageCounterY == 2'h2; // @[Counter.scala 38:24]
  wire [1:0] _T_23 = imageCounterY + 2'h1; // @[Counter.scala 39:22]
  reg [31:0] pixelIndex; // @[Filter.scala 199:31]
  wire [32:0] _T_24 = {{1'd0}, pixelIndex}; // @[Filter.scala 202:31]
  wire [31:0] _GEN_0 = _T_24[31:0] % 32'h15; // @[Filter.scala 202:38]
  wire [4:0] _T_26 = _GEN_0[4:0]; // @[Filter.scala 202:38]
  wire [4:0] _GEN_11210 = {{3'd0}, imageCounterX}; // @[Filter.scala 202:53]
  wire [4:0] _T_28 = _T_26 + _GEN_11210; // @[Filter.scala 202:53]
  wire [4:0] _T_30 = _T_28 - 5'h1; // @[Filter.scala 202:69]
  wire [31:0] _T_33 = _T_24[31:0] / 32'h15; // @[Filter.scala 203:38]
  wire [31:0] _GEN_11211 = {{30'd0}, imageCounterY}; // @[Filter.scala 203:53]
  wire [31:0] _T_35 = _T_33 + _GEN_11211; // @[Filter.scala 203:53]
  wire [31:0] _T_37 = _T_35 - 32'h1; // @[Filter.scala 203:69]
  wire [36:0] _T_38 = _T_37 * 32'h15; // @[Filter.scala 204:42]
  wire [36:0] _GEN_11212 = {{32'd0}, _T_30}; // @[Filter.scala 204:57]
  wire [36:0] _T_40 = _T_38 + _GEN_11212; // @[Filter.scala 204:57]
  wire [3:0] _GEN_179 = 8'h8 == _T_40[7:0] ? 4'h1 : 4'h0; // @[Filter.scala 204:62]
  wire [3:0] _GEN_180 = 8'h9 == _T_40[7:0] ? 4'h2 : _GEN_179; // @[Filter.scala 204:62]
  wire [3:0] _GEN_181 = 8'ha == _T_40[7:0] ? 4'h2 : _GEN_180; // @[Filter.scala 204:62]
  wire [3:0] _GEN_182 = 8'hb == _T_40[7:0] ? 4'h2 : _GEN_181; // @[Filter.scala 204:62]
  wire [3:0] _GEN_183 = 8'hc == _T_40[7:0] ? 4'h1 : _GEN_182; // @[Filter.scala 204:62]
  wire [3:0] _GEN_184 = 8'hd == _T_40[7:0] ? 4'h0 : _GEN_183; // @[Filter.scala 204:62]
  wire [3:0] _GEN_185 = 8'he == _T_40[7:0] ? 4'h0 : _GEN_184; // @[Filter.scala 204:62]
  wire [3:0] _GEN_186 = 8'hf == _T_40[7:0] ? 4'h0 : _GEN_185; // @[Filter.scala 204:62]
  wire [3:0] _GEN_187 = 8'h10 == _T_40[7:0] ? 4'h0 : _GEN_186; // @[Filter.scala 204:62]
  wire [3:0] _GEN_188 = 8'h11 == _T_40[7:0] ? 4'h0 : _GEN_187; // @[Filter.scala 204:62]
  wire [3:0] _GEN_189 = 8'h12 == _T_40[7:0] ? 4'h0 : _GEN_188; // @[Filter.scala 204:62]
  wire [3:0] _GEN_190 = 8'h13 == _T_40[7:0] ? 4'h0 : _GEN_189; // @[Filter.scala 204:62]
  wire [3:0] _GEN_191 = 8'h14 == _T_40[7:0] ? 4'h0 : _GEN_190; // @[Filter.scala 204:62]
  wire [3:0] _GEN_192 = 8'h15 == _T_40[7:0] ? 4'h0 : _GEN_191; // @[Filter.scala 204:62]
  wire [3:0] _GEN_193 = 8'h16 == _T_40[7:0] ? 4'h0 : _GEN_192; // @[Filter.scala 204:62]
  wire [3:0] _GEN_194 = 8'h17 == _T_40[7:0] ? 4'h0 : _GEN_193; // @[Filter.scala 204:62]
  wire [3:0] _GEN_195 = 8'h18 == _T_40[7:0] ? 4'h0 : _GEN_194; // @[Filter.scala 204:62]
  wire [3:0] _GEN_196 = 8'h19 == _T_40[7:0] ? 4'h0 : _GEN_195; // @[Filter.scala 204:62]
  wire [3:0] _GEN_197 = 8'h1a == _T_40[7:0] ? 4'h0 : _GEN_196; // @[Filter.scala 204:62]
  wire [3:0] _GEN_198 = 8'h1b == _T_40[7:0] ? 4'h0 : _GEN_197; // @[Filter.scala 204:62]
  wire [3:0] _GEN_199 = 8'h1c == _T_40[7:0] ? 4'h2 : _GEN_198; // @[Filter.scala 204:62]
  wire [3:0] _GEN_200 = 8'h1d == _T_40[7:0] ? 4'h1 : _GEN_199; // @[Filter.scala 204:62]
  wire [3:0] _GEN_201 = 8'h1e == _T_40[7:0] ? 4'h0 : _GEN_200; // @[Filter.scala 204:62]
  wire [3:0] _GEN_202 = 8'h1f == _T_40[7:0] ? 4'h0 : _GEN_201; // @[Filter.scala 204:62]
  wire [3:0] _GEN_203 = 8'h20 == _T_40[7:0] ? 4'h0 : _GEN_202; // @[Filter.scala 204:62]
  wire [3:0] _GEN_204 = 8'h21 == _T_40[7:0] ? 4'h1 : _GEN_203; // @[Filter.scala 204:62]
  wire [3:0] _GEN_205 = 8'h22 == _T_40[7:0] ? 4'h2 : _GEN_204; // @[Filter.scala 204:62]
  wire [3:0] _GEN_206 = 8'h23 == _T_40[7:0] ? 4'h0 : _GEN_205; // @[Filter.scala 204:62]
  wire [3:0] _GEN_207 = 8'h24 == _T_40[7:0] ? 4'h0 : _GEN_206; // @[Filter.scala 204:62]
  wire [3:0] _GEN_208 = 8'h25 == _T_40[7:0] ? 4'h0 : _GEN_207; // @[Filter.scala 204:62]
  wire [3:0] _GEN_209 = 8'h26 == _T_40[7:0] ? 4'h0 : _GEN_208; // @[Filter.scala 204:62]
  wire [3:0] _GEN_210 = 8'h27 == _T_40[7:0] ? 4'h0 : _GEN_209; // @[Filter.scala 204:62]
  wire [3:0] _GEN_211 = 8'h28 == _T_40[7:0] ? 4'h0 : _GEN_210; // @[Filter.scala 204:62]
  wire [3:0] _GEN_212 = 8'h29 == _T_40[7:0] ? 4'h0 : _GEN_211; // @[Filter.scala 204:62]
  wire [3:0] _GEN_213 = 8'h2a == _T_40[7:0] ? 4'h0 : _GEN_212; // @[Filter.scala 204:62]
  wire [3:0] _GEN_214 = 8'h2b == _T_40[7:0] ? 4'h0 : _GEN_213; // @[Filter.scala 204:62]
  wire [3:0] _GEN_215 = 8'h2c == _T_40[7:0] ? 4'h0 : _GEN_214; // @[Filter.scala 204:62]
  wire [3:0] _GEN_216 = 8'h2d == _T_40[7:0] ? 4'h0 : _GEN_215; // @[Filter.scala 204:62]
  wire [3:0] _GEN_217 = 8'h2e == _T_40[7:0] ? 4'h0 : _GEN_216; // @[Filter.scala 204:62]
  wire [3:0] _GEN_218 = 8'h2f == _T_40[7:0] ? 4'h0 : _GEN_217; // @[Filter.scala 204:62]
  wire [3:0] _GEN_219 = 8'h30 == _T_40[7:0] ? 4'h2 : _GEN_218; // @[Filter.scala 204:62]
  wire [3:0] _GEN_220 = 8'h31 == _T_40[7:0] ? 4'h2 : _GEN_219; // @[Filter.scala 204:62]
  wire [3:0] _GEN_221 = 8'h32 == _T_40[7:0] ? 4'h0 : _GEN_220; // @[Filter.scala 204:62]
  wire [3:0] _GEN_222 = 8'h33 == _T_40[7:0] ? 4'h0 : _GEN_221; // @[Filter.scala 204:62]
  wire [3:0] _GEN_223 = 8'h34 == _T_40[7:0] ? 4'h0 : _GEN_222; // @[Filter.scala 204:62]
  wire [3:0] _GEN_224 = 8'h35 == _T_40[7:0] ? 4'h0 : _GEN_223; // @[Filter.scala 204:62]
  wire [3:0] _GEN_225 = 8'h36 == _T_40[7:0] ? 4'h0 : _GEN_224; // @[Filter.scala 204:62]
  wire [3:0] _GEN_226 = 8'h37 == _T_40[7:0] ? 4'h0 : _GEN_225; // @[Filter.scala 204:62]
  wire [3:0] _GEN_227 = 8'h38 == _T_40[7:0] ? 4'h2 : _GEN_226; // @[Filter.scala 204:62]
  wire [3:0] _GEN_228 = 8'h39 == _T_40[7:0] ? 4'h0 : _GEN_227; // @[Filter.scala 204:62]
  wire [3:0] _GEN_229 = 8'h3a == _T_40[7:0] ? 4'h0 : _GEN_228; // @[Filter.scala 204:62]
  wire [3:0] _GEN_230 = 8'h3b == _T_40[7:0] ? 4'h0 : _GEN_229; // @[Filter.scala 204:62]
  wire [3:0] _GEN_231 = 8'h3c == _T_40[7:0] ? 4'h0 : _GEN_230; // @[Filter.scala 204:62]
  wire [3:0] _GEN_232 = 8'h3d == _T_40[7:0] ? 4'h0 : _GEN_231; // @[Filter.scala 204:62]
  wire [3:0] _GEN_233 = 8'h3e == _T_40[7:0] ? 4'h0 : _GEN_232; // @[Filter.scala 204:62]
  wire [3:0] _GEN_234 = 8'h3f == _T_40[7:0] ? 4'h0 : _GEN_233; // @[Filter.scala 204:62]
  wire [3:0] _GEN_235 = 8'h40 == _T_40[7:0] ? 4'h0 : _GEN_234; // @[Filter.scala 204:62]
  wire [3:0] _GEN_236 = 8'h41 == _T_40[7:0] ? 4'h0 : _GEN_235; // @[Filter.scala 204:62]
  wire [3:0] _GEN_237 = 8'h42 == _T_40[7:0] ? 4'h0 : _GEN_236; // @[Filter.scala 204:62]
  wire [3:0] _GEN_238 = 8'h43 == _T_40[7:0] ? 4'h0 : _GEN_237; // @[Filter.scala 204:62]
  wire [3:0] _GEN_239 = 8'h44 == _T_40[7:0] ? 4'h1 : _GEN_238; // @[Filter.scala 204:62]
  wire [3:0] _GEN_240 = 8'h45 == _T_40[7:0] ? 4'h3 : _GEN_239; // @[Filter.scala 204:62]
  wire [3:0] _GEN_241 = 8'h46 == _T_40[7:0] ? 4'h7 : _GEN_240; // @[Filter.scala 204:62]
  wire [3:0] _GEN_242 = 8'h47 == _T_40[7:0] ? 4'h0 : _GEN_241; // @[Filter.scala 204:62]
  wire [3:0] _GEN_243 = 8'h48 == _T_40[7:0] ? 4'h0 : _GEN_242; // @[Filter.scala 204:62]
  wire [3:0] _GEN_244 = 8'h49 == _T_40[7:0] ? 4'h0 : _GEN_243; // @[Filter.scala 204:62]
  wire [3:0] _GEN_245 = 8'h4a == _T_40[7:0] ? 4'h0 : _GEN_244; // @[Filter.scala 204:62]
  wire [3:0] _GEN_246 = 8'h4b == _T_40[7:0] ? 4'h0 : _GEN_245; // @[Filter.scala 204:62]
  wire [3:0] _GEN_247 = 8'h4c == _T_40[7:0] ? 4'h0 : _GEN_246; // @[Filter.scala 204:62]
  wire [3:0] _GEN_248 = 8'h4d == _T_40[7:0] ? 4'h0 : _GEN_247; // @[Filter.scala 204:62]
  wire [3:0] _GEN_249 = 8'h4e == _T_40[7:0] ? 4'h2 : _GEN_248; // @[Filter.scala 204:62]
  wire [3:0] _GEN_250 = 8'h4f == _T_40[7:0] ? 4'h0 : _GEN_249; // @[Filter.scala 204:62]
  wire [3:0] _GEN_251 = 8'h50 == _T_40[7:0] ? 4'h0 : _GEN_250; // @[Filter.scala 204:62]
  wire [3:0] _GEN_252 = 8'h51 == _T_40[7:0] ? 4'h0 : _GEN_251; // @[Filter.scala 204:62]
  wire [3:0] _GEN_253 = 8'h52 == _T_40[7:0] ? 4'h0 : _GEN_252; // @[Filter.scala 204:62]
  wire [3:0] _GEN_254 = 8'h53 == _T_40[7:0] ? 4'h0 : _GEN_253; // @[Filter.scala 204:62]
  wire [3:0] _GEN_255 = 8'h54 == _T_40[7:0] ? 4'h0 : _GEN_254; // @[Filter.scala 204:62]
  wire [3:0] _GEN_256 = 8'h55 == _T_40[7:0] ? 4'h0 : _GEN_255; // @[Filter.scala 204:62]
  wire [3:0] _GEN_257 = 8'h56 == _T_40[7:0] ? 4'h0 : _GEN_256; // @[Filter.scala 204:62]
  wire [3:0] _GEN_258 = 8'h57 == _T_40[7:0] ? 4'h0 : _GEN_257; // @[Filter.scala 204:62]
  wire [3:0] _GEN_259 = 8'h58 == _T_40[7:0] ? 4'h0 : _GEN_258; // @[Filter.scala 204:62]
  wire [3:0] _GEN_260 = 8'h59 == _T_40[7:0] ? 4'h2 : _GEN_259; // @[Filter.scala 204:62]
  wire [3:0] _GEN_261 = 8'h5a == _T_40[7:0] ? 4'h2 : _GEN_260; // @[Filter.scala 204:62]
  wire [3:0] _GEN_262 = 8'h5b == _T_40[7:0] ? 4'h0 : _GEN_261; // @[Filter.scala 204:62]
  wire [3:0] _GEN_263 = 8'h5c == _T_40[7:0] ? 4'h0 : _GEN_262; // @[Filter.scala 204:62]
  wire [3:0] _GEN_264 = 8'h5d == _T_40[7:0] ? 4'h0 : _GEN_263; // @[Filter.scala 204:62]
  wire [3:0] _GEN_265 = 8'h5e == _T_40[7:0] ? 4'h4 : _GEN_264; // @[Filter.scala 204:62]
  wire [3:0] _GEN_266 = 8'h5f == _T_40[7:0] ? 4'h0 : _GEN_265; // @[Filter.scala 204:62]
  wire [3:0] _GEN_267 = 8'h60 == _T_40[7:0] ? 4'h0 : _GEN_266; // @[Filter.scala 204:62]
  wire [3:0] _GEN_268 = 8'h61 == _T_40[7:0] ? 4'h0 : _GEN_267; // @[Filter.scala 204:62]
  wire [3:0] _GEN_269 = 8'h62 == _T_40[7:0] ? 4'h0 : _GEN_268; // @[Filter.scala 204:62]
  wire [3:0] _GEN_270 = 8'h63 == _T_40[7:0] ? 4'h2 : _GEN_269; // @[Filter.scala 204:62]
  wire [3:0] _GEN_271 = 8'h64 == _T_40[7:0] ? 4'h0 : _GEN_270; // @[Filter.scala 204:62]
  wire [3:0] _GEN_272 = 8'h65 == _T_40[7:0] ? 4'h0 : _GEN_271; // @[Filter.scala 204:62]
  wire [3:0] _GEN_273 = 8'h66 == _T_40[7:0] ? 4'h0 : _GEN_272; // @[Filter.scala 204:62]
  wire [3:0] _GEN_274 = 8'h67 == _T_40[7:0] ? 4'h0 : _GEN_273; // @[Filter.scala 204:62]
  wire [3:0] _GEN_275 = 8'h68 == _T_40[7:0] ? 4'h0 : _GEN_274; // @[Filter.scala 204:62]
  wire [3:0] _GEN_276 = 8'h69 == _T_40[7:0] ? 4'h0 : _GEN_275; // @[Filter.scala 204:62]
  wire [3:0] _GEN_277 = 8'h6a == _T_40[7:0] ? 4'h0 : _GEN_276; // @[Filter.scala 204:62]
  wire [3:0] _GEN_278 = 8'h6b == _T_40[7:0] ? 4'h0 : _GEN_277; // @[Filter.scala 204:62]
  wire [3:0] _GEN_279 = 8'h6c == _T_40[7:0] ? 4'h0 : _GEN_278; // @[Filter.scala 204:62]
  wire [3:0] _GEN_280 = 8'h6d == _T_40[7:0] ? 4'h0 : _GEN_279; // @[Filter.scala 204:62]
  wire [3:0] _GEN_281 = 8'h6e == _T_40[7:0] ? 4'h2 : _GEN_280; // @[Filter.scala 204:62]
  wire [3:0] _GEN_282 = 8'h6f == _T_40[7:0] ? 4'h0 : _GEN_281; // @[Filter.scala 204:62]
  wire [3:0] _GEN_283 = 8'h70 == _T_40[7:0] ? 4'h0 : _GEN_282; // @[Filter.scala 204:62]
  wire [3:0] _GEN_284 = 8'h71 == _T_40[7:0] ? 4'h0 : _GEN_283; // @[Filter.scala 204:62]
  wire [3:0] _GEN_285 = 8'h72 == _T_40[7:0] ? 4'h2 : _GEN_284; // @[Filter.scala 204:62]
  wire [3:0] _GEN_286 = 8'h73 == _T_40[7:0] ? 4'h9 : _GEN_285; // @[Filter.scala 204:62]
  wire [3:0] _GEN_287 = 8'h74 == _T_40[7:0] ? 4'h2 : _GEN_286; // @[Filter.scala 204:62]
  wire [3:0] _GEN_288 = 8'h75 == _T_40[7:0] ? 4'h0 : _GEN_287; // @[Filter.scala 204:62]
  wire [3:0] _GEN_289 = 8'h76 == _T_40[7:0] ? 4'h0 : _GEN_288; // @[Filter.scala 204:62]
  wire [3:0] _GEN_290 = 8'h77 == _T_40[7:0] ? 4'h0 : _GEN_289; // @[Filter.scala 204:62]
  wire [3:0] _GEN_291 = 8'h78 == _T_40[7:0] ? 4'h1 : _GEN_290; // @[Filter.scala 204:62]
  wire [3:0] _GEN_292 = 8'h79 == _T_40[7:0] ? 4'h1 : _GEN_291; // @[Filter.scala 204:62]
  wire [3:0] _GEN_293 = 8'h7a == _T_40[7:0] ? 4'h0 : _GEN_292; // @[Filter.scala 204:62]
  wire [3:0] _GEN_294 = 8'h7b == _T_40[7:0] ? 4'h0 : _GEN_293; // @[Filter.scala 204:62]
  wire [3:0] _GEN_295 = 8'h7c == _T_40[7:0] ? 4'h0 : _GEN_294; // @[Filter.scala 204:62]
  wire [3:0] _GEN_296 = 8'h7d == _T_40[7:0] ? 4'h0 : _GEN_295; // @[Filter.scala 204:62]
  wire [3:0] _GEN_297 = 8'h7e == _T_40[7:0] ? 4'h0 : _GEN_296; // @[Filter.scala 204:62]
  wire [3:0] _GEN_298 = 8'h7f == _T_40[7:0] ? 4'h0 : _GEN_297; // @[Filter.scala 204:62]
  wire [3:0] _GEN_299 = 8'h80 == _T_40[7:0] ? 4'h0 : _GEN_298; // @[Filter.scala 204:62]
  wire [3:0] _GEN_300 = 8'h81 == _T_40[7:0] ? 4'h0 : _GEN_299; // @[Filter.scala 204:62]
  wire [3:0] _GEN_301 = 8'h82 == _T_40[7:0] ? 4'h2 : _GEN_300; // @[Filter.scala 204:62]
  wire [3:0] _GEN_302 = 8'h83 == _T_40[7:0] ? 4'h0 : _GEN_301; // @[Filter.scala 204:62]
  wire [3:0] _GEN_303 = 8'h84 == _T_40[7:0] ? 4'h0 : _GEN_302; // @[Filter.scala 204:62]
  wire [3:0] _GEN_304 = 8'h85 == _T_40[7:0] ? 4'h0 : _GEN_303; // @[Filter.scala 204:62]
  wire [3:0] _GEN_305 = 8'h86 == _T_40[7:0] ? 4'h7 : _GEN_304; // @[Filter.scala 204:62]
  wire [3:0] _GEN_306 = 8'h87 == _T_40[7:0] ? 4'h2 : _GEN_305; // @[Filter.scala 204:62]
  wire [3:0] _GEN_307 = 8'h88 == _T_40[7:0] ? 4'h0 : _GEN_306; // @[Filter.scala 204:62]
  wire [3:0] _GEN_308 = 8'h89 == _T_40[7:0] ? 4'h2 : _GEN_307; // @[Filter.scala 204:62]
  wire [3:0] _GEN_309 = 8'h8a == _T_40[7:0] ? 4'h7 : _GEN_308; // @[Filter.scala 204:62]
  wire [3:0] _GEN_310 = 8'h8b == _T_40[7:0] ? 4'h0 : _GEN_309; // @[Filter.scala 204:62]
  wire [3:0] _GEN_311 = 8'h8c == _T_40[7:0] ? 4'h0 : _GEN_310; // @[Filter.scala 204:62]
  wire [3:0] _GEN_312 = 8'h8d == _T_40[7:0] ? 4'h0 : _GEN_311; // @[Filter.scala 204:62]
  wire [3:0] _GEN_313 = 8'h8e == _T_40[7:0] ? 4'h2 : _GEN_312; // @[Filter.scala 204:62]
  wire [3:0] _GEN_314 = 8'h8f == _T_40[7:0] ? 4'h0 : _GEN_313; // @[Filter.scala 204:62]
  wire [3:0] _GEN_315 = 8'h90 == _T_40[7:0] ? 4'h0 : _GEN_314; // @[Filter.scala 204:62]
  wire [3:0] _GEN_316 = 8'h91 == _T_40[7:0] ? 4'h0 : _GEN_315; // @[Filter.scala 204:62]
  wire [3:0] _GEN_317 = 8'h92 == _T_40[7:0] ? 4'h0 : _GEN_316; // @[Filter.scala 204:62]
  wire [3:0] _GEN_318 = 8'h93 == _T_40[7:0] ? 4'h0 : _GEN_317; // @[Filter.scala 204:62]
  wire [3:0] _GEN_319 = 8'h94 == _T_40[7:0] ? 4'h0 : _GEN_318; // @[Filter.scala 204:62]
  wire [3:0] _GEN_320 = 8'h95 == _T_40[7:0] ? 4'h0 : _GEN_319; // @[Filter.scala 204:62]
  wire [3:0] _GEN_321 = 8'h96 == _T_40[7:0] ? 4'h0 : _GEN_320; // @[Filter.scala 204:62]
  wire [3:0] _GEN_322 = 8'h97 == _T_40[7:0] ? 4'h2 : _GEN_321; // @[Filter.scala 204:62]
  wire [3:0] _GEN_323 = 8'h98 == _T_40[7:0] ? 4'h2 : _GEN_322; // @[Filter.scala 204:62]
  wire [3:0] _GEN_324 = 8'h99 == _T_40[7:0] ? 4'h1 : _GEN_323; // @[Filter.scala 204:62]
  wire [3:0] _GEN_325 = 8'h9a == _T_40[7:0] ? 4'h0 : _GEN_324; // @[Filter.scala 204:62]
  wire [3:0] _GEN_326 = 8'h9b == _T_40[7:0] ? 4'h7 : _GEN_325; // @[Filter.scala 204:62]
  wire [3:0] _GEN_327 = 8'h9c == _T_40[7:0] ? 4'h7 : _GEN_326; // @[Filter.scala 204:62]
  wire [3:0] _GEN_328 = 8'h9d == _T_40[7:0] ? 4'h0 : _GEN_327; // @[Filter.scala 204:62]
  wire [3:0] _GEN_329 = 8'h9e == _T_40[7:0] ? 4'h7 : _GEN_328; // @[Filter.scala 204:62]
  wire [3:0] _GEN_330 = 8'h9f == _T_40[7:0] ? 4'h7 : _GEN_329; // @[Filter.scala 204:62]
  wire [3:0] _GEN_331 = 8'ha0 == _T_40[7:0] ? 4'h0 : _GEN_330; // @[Filter.scala 204:62]
  wire [3:0] _GEN_332 = 8'ha1 == _T_40[7:0] ? 4'h1 : _GEN_331; // @[Filter.scala 204:62]
  wire [3:0] _GEN_333 = 8'ha2 == _T_40[7:0] ? 4'h2 : _GEN_332; // @[Filter.scala 204:62]
  wire [3:0] _GEN_334 = 8'ha3 == _T_40[7:0] ? 4'h2 : _GEN_333; // @[Filter.scala 204:62]
  wire [3:0] _GEN_335 = 8'ha4 == _T_40[7:0] ? 4'h0 : _GEN_334; // @[Filter.scala 204:62]
  wire [3:0] _GEN_336 = 8'ha5 == _T_40[7:0] ? 4'h0 : _GEN_335; // @[Filter.scala 204:62]
  wire [3:0] _GEN_337 = 8'ha6 == _T_40[7:0] ? 4'h0 : _GEN_336; // @[Filter.scala 204:62]
  wire [3:0] _GEN_338 = 8'ha7 == _T_40[7:0] ? 4'h0 : _GEN_337; // @[Filter.scala 204:62]
  wire [3:0] _GEN_339 = 8'ha8 == _T_40[7:0] ? 4'h0 : _GEN_338; // @[Filter.scala 204:62]
  wire [3:0] _GEN_340 = 8'ha9 == _T_40[7:0] ? 4'h0 : _GEN_339; // @[Filter.scala 204:62]
  wire [3:0] _GEN_341 = 8'haa == _T_40[7:0] ? 4'h0 : _GEN_340; // @[Filter.scala 204:62]
  wire [3:0] _GEN_342 = 8'hab == _T_40[7:0] ? 4'h0 : _GEN_341; // @[Filter.scala 204:62]
  wire [3:0] _GEN_343 = 8'hac == _T_40[7:0] ? 4'h2 : _GEN_342; // @[Filter.scala 204:62]
  wire [3:0] _GEN_344 = 8'had == _T_40[7:0] ? 4'h0 : _GEN_343; // @[Filter.scala 204:62]
  wire [3:0] _GEN_345 = 8'hae == _T_40[7:0] ? 4'h1 : _GEN_344; // @[Filter.scala 204:62]
  wire [3:0] _GEN_346 = 8'haf == _T_40[7:0] ? 4'h3 : _GEN_345; // @[Filter.scala 204:62]
  wire [3:0] _GEN_347 = 8'hb0 == _T_40[7:0] ? 4'h1 : _GEN_346; // @[Filter.scala 204:62]
  wire [3:0] _GEN_348 = 8'hb1 == _T_40[7:0] ? 4'h0 : _GEN_347; // @[Filter.scala 204:62]
  wire [3:0] _GEN_349 = 8'hb2 == _T_40[7:0] ? 4'h0 : _GEN_348; // @[Filter.scala 204:62]
  wire [3:0] _GEN_350 = 8'hb3 == _T_40[7:0] ? 4'h0 : _GEN_349; // @[Filter.scala 204:62]
  wire [3:0] _GEN_351 = 8'hb4 == _T_40[7:0] ? 4'h1 : _GEN_350; // @[Filter.scala 204:62]
  wire [3:0] _GEN_352 = 8'hb5 == _T_40[7:0] ? 4'h3 : _GEN_351; // @[Filter.scala 204:62]
  wire [3:0] _GEN_353 = 8'hb6 == _T_40[7:0] ? 4'h1 : _GEN_352; // @[Filter.scala 204:62]
  wire [3:0] _GEN_354 = 8'hb7 == _T_40[7:0] ? 4'h0 : _GEN_353; // @[Filter.scala 204:62]
  wire [3:0] _GEN_355 = 8'hb8 == _T_40[7:0] ? 4'h2 : _GEN_354; // @[Filter.scala 204:62]
  wire [3:0] _GEN_356 = 8'hb9 == _T_40[7:0] ? 4'h0 : _GEN_355; // @[Filter.scala 204:62]
  wire [3:0] _GEN_357 = 8'hba == _T_40[7:0] ? 4'h0 : _GEN_356; // @[Filter.scala 204:62]
  wire [3:0] _GEN_358 = 8'hbb == _T_40[7:0] ? 4'h0 : _GEN_357; // @[Filter.scala 204:62]
  wire [3:0] _GEN_359 = 8'hbc == _T_40[7:0] ? 4'h0 : _GEN_358; // @[Filter.scala 204:62]
  wire [3:0] _GEN_360 = 8'hbd == _T_40[7:0] ? 4'h0 : _GEN_359; // @[Filter.scala 204:62]
  wire [3:0] _GEN_361 = 8'hbe == _T_40[7:0] ? 4'h0 : _GEN_360; // @[Filter.scala 204:62]
  wire [3:0] _GEN_362 = 8'hbf == _T_40[7:0] ? 4'h0 : _GEN_361; // @[Filter.scala 204:62]
  wire [3:0] _GEN_363 = 8'hc0 == _T_40[7:0] ? 4'h0 : _GEN_362; // @[Filter.scala 204:62]
  wire [3:0] _GEN_364 = 8'hc1 == _T_40[7:0] ? 4'h0 : _GEN_363; // @[Filter.scala 204:62]
  wire [3:0] _GEN_365 = 8'hc2 == _T_40[7:0] ? 4'h3 : _GEN_364; // @[Filter.scala 204:62]
  wire [3:0] _GEN_366 = 8'hc3 == _T_40[7:0] ? 4'h0 : _GEN_365; // @[Filter.scala 204:62]
  wire [3:0] _GEN_367 = 8'hc4 == _T_40[7:0] ? 4'h0 : _GEN_366; // @[Filter.scala 204:62]
  wire [3:0] _GEN_368 = 8'hc5 == _T_40[7:0] ? 4'h2 : _GEN_367; // @[Filter.scala 204:62]
  wire [3:0] _GEN_369 = 8'hc6 == _T_40[7:0] ? 4'h3 : _GEN_368; // @[Filter.scala 204:62]
  wire [3:0] _GEN_370 = 8'hc7 == _T_40[7:0] ? 4'h2 : _GEN_369; // @[Filter.scala 204:62]
  wire [3:0] _GEN_371 = 8'hc8 == _T_40[7:0] ? 4'h3 : _GEN_370; // @[Filter.scala 204:62]
  wire [3:0] _GEN_372 = 8'hc9 == _T_40[7:0] ? 4'h2 : _GEN_371; // @[Filter.scala 204:62]
  wire [3:0] _GEN_373 = 8'hca == _T_40[7:0] ? 4'h0 : _GEN_372; // @[Filter.scala 204:62]
  wire [3:0] _GEN_374 = 8'hcb == _T_40[7:0] ? 4'h0 : _GEN_373; // @[Filter.scala 204:62]
  wire [3:0] _GEN_375 = 8'hcc == _T_40[7:0] ? 4'h3 : _GEN_374; // @[Filter.scala 204:62]
  wire [3:0] _GEN_376 = 8'hcd == _T_40[7:0] ? 4'h0 : _GEN_375; // @[Filter.scala 204:62]
  wire [3:0] _GEN_377 = 8'hce == _T_40[7:0] ? 4'h0 : _GEN_376; // @[Filter.scala 204:62]
  wire [3:0] _GEN_378 = 8'hcf == _T_40[7:0] ? 4'h0 : _GEN_377; // @[Filter.scala 204:62]
  wire [3:0] _GEN_379 = 8'hd0 == _T_40[7:0] ? 4'h0 : _GEN_378; // @[Filter.scala 204:62]
  wire [3:0] _GEN_380 = 8'hd1 == _T_40[7:0] ? 4'h0 : _GEN_379; // @[Filter.scala 204:62]
  wire [3:0] _GEN_381 = 8'hd2 == _T_40[7:0] ? 4'h0 : _GEN_380; // @[Filter.scala 204:62]
  wire [3:0] _GEN_382 = 8'hd3 == _T_40[7:0] ? 4'h0 : _GEN_381; // @[Filter.scala 204:62]
  wire [3:0] _GEN_383 = 8'hd4 == _T_40[7:0] ? 4'h0 : _GEN_382; // @[Filter.scala 204:62]
  wire [3:0] _GEN_384 = 8'hd5 == _T_40[7:0] ? 4'h0 : _GEN_383; // @[Filter.scala 204:62]
  wire [3:0] _GEN_385 = 8'hd6 == _T_40[7:0] ? 4'h0 : _GEN_384; // @[Filter.scala 204:62]
  wire [3:0] _GEN_386 = 8'hd7 == _T_40[7:0] ? 4'h2 : _GEN_385; // @[Filter.scala 204:62]
  wire [3:0] _GEN_387 = 8'hd8 == _T_40[7:0] ? 4'h2 : _GEN_386; // @[Filter.scala 204:62]
  wire [3:0] _GEN_388 = 8'hd9 == _T_40[7:0] ? 4'h0 : _GEN_387; // @[Filter.scala 204:62]
  wire [3:0] _GEN_389 = 8'hda == _T_40[7:0] ? 4'h7 : _GEN_388; // @[Filter.scala 204:62]
  wire [3:0] _GEN_390 = 8'hdb == _T_40[7:0] ? 4'h1 : _GEN_389; // @[Filter.scala 204:62]
  wire [3:0] _GEN_391 = 8'hdc == _T_40[7:0] ? 4'h4 : _GEN_390; // @[Filter.scala 204:62]
  wire [3:0] _GEN_392 = 8'hdd == _T_40[7:0] ? 4'h1 : _GEN_391; // @[Filter.scala 204:62]
  wire [3:0] _GEN_393 = 8'hde == _T_40[7:0] ? 4'h7 : _GEN_392; // @[Filter.scala 204:62]
  wire [3:0] _GEN_394 = 8'hdf == _T_40[7:0] ? 4'h0 : _GEN_393; // @[Filter.scala 204:62]
  wire [3:0] _GEN_395 = 8'he0 == _T_40[7:0] ? 4'h2 : _GEN_394; // @[Filter.scala 204:62]
  wire [3:0] _GEN_396 = 8'he1 == _T_40[7:0] ? 4'h2 : _GEN_395; // @[Filter.scala 204:62]
  wire [3:0] _GEN_397 = 8'he2 == _T_40[7:0] ? 4'h0 : _GEN_396; // @[Filter.scala 204:62]
  wire [3:0] _GEN_398 = 8'he3 == _T_40[7:0] ? 4'h0 : _GEN_397; // @[Filter.scala 204:62]
  wire [3:0] _GEN_399 = 8'he4 == _T_40[7:0] ? 4'h0 : _GEN_398; // @[Filter.scala 204:62]
  wire [3:0] _GEN_400 = 8'he5 == _T_40[7:0] ? 4'h0 : _GEN_399; // @[Filter.scala 204:62]
  wire [3:0] _GEN_401 = 8'he6 == _T_40[7:0] ? 4'h0 : _GEN_400; // @[Filter.scala 204:62]
  wire [3:0] _GEN_402 = 8'he7 == _T_40[7:0] ? 4'h0 : _GEN_401; // @[Filter.scala 204:62]
  wire [3:0] _GEN_403 = 8'he8 == _T_40[7:0] ? 4'h0 : _GEN_402; // @[Filter.scala 204:62]
  wire [3:0] _GEN_404 = 8'he9 == _T_40[7:0] ? 4'h0 : _GEN_403; // @[Filter.scala 204:62]
  wire [3:0] _GEN_405 = 8'hea == _T_40[7:0] ? 4'h0 : _GEN_404; // @[Filter.scala 204:62]
  wire [3:0] _GEN_406 = 8'heb == _T_40[7:0] ? 4'h0 : _GEN_405; // @[Filter.scala 204:62]
  wire [3:0] _GEN_407 = 8'hec == _T_40[7:0] ? 4'h0 : _GEN_406; // @[Filter.scala 204:62]
  wire [3:0] _GEN_408 = 8'hed == _T_40[7:0] ? 4'h0 : _GEN_407; // @[Filter.scala 204:62]
  wire [3:0] _GEN_409 = 8'hee == _T_40[7:0] ? 4'h0 : _GEN_408; // @[Filter.scala 204:62]
  wire [3:0] _GEN_410 = 8'hef == _T_40[7:0] ? 4'h0 : _GEN_409; // @[Filter.scala 204:62]
  wire [3:0] _GEN_411 = 8'hf0 == _T_40[7:0] ? 4'h0 : _GEN_410; // @[Filter.scala 204:62]
  wire [3:0] _GEN_412 = 8'hf1 == _T_40[7:0] ? 4'h0 : _GEN_411; // @[Filter.scala 204:62]
  wire [3:0] _GEN_413 = 8'hf2 == _T_40[7:0] ? 4'h0 : _GEN_412; // @[Filter.scala 204:62]
  wire [3:0] _GEN_414 = 8'hf3 == _T_40[7:0] ? 4'h0 : _GEN_413; // @[Filter.scala 204:62]
  wire [3:0] _GEN_415 = 8'hf4 == _T_40[7:0] ? 4'h0 : _GEN_414; // @[Filter.scala 204:62]
  wire [3:0] _GEN_416 = 8'hf5 == _T_40[7:0] ? 4'h0 : _GEN_415; // @[Filter.scala 204:62]
  wire [3:0] _GEN_417 = 8'hf6 == _T_40[7:0] ? 4'h0 : _GEN_416; // @[Filter.scala 204:62]
  wire [3:0] _GEN_418 = 8'hf7 == _T_40[7:0] ? 4'h0 : _GEN_417; // @[Filter.scala 204:62]
  wire [3:0] _GEN_419 = 8'hf8 == _T_40[7:0] ? 4'h0 : _GEN_418; // @[Filter.scala 204:62]
  wire [3:0] _GEN_420 = 8'hf9 == _T_40[7:0] ? 4'h0 : _GEN_419; // @[Filter.scala 204:62]
  wire [3:0] _GEN_421 = 8'hfa == _T_40[7:0] ? 4'h0 : _GEN_420; // @[Filter.scala 204:62]
  wire [3:0] _GEN_422 = 8'hfb == _T_40[7:0] ? 4'h0 : _GEN_421; // @[Filter.scala 204:62]
  wire [4:0] _GEN_11213 = {{1'd0}, _GEN_422}; // @[Filter.scala 204:62]
  wire [8:0] _T_42 = _GEN_11213 * 5'h14; // @[Filter.scala 204:62]
  wire [3:0] _GEN_472 = 8'h31 == _T_40[7:0] ? 4'h3 : _GEN_219; // @[Filter.scala 204:102]
  wire [3:0] _GEN_473 = 8'h32 == _T_40[7:0] ? 4'h3 : _GEN_472; // @[Filter.scala 204:102]
  wire [3:0] _GEN_474 = 8'h33 == _T_40[7:0] ? 4'h6 : _GEN_473; // @[Filter.scala 204:102]
  wire [3:0] _GEN_475 = 8'h34 == _T_40[7:0] ? 4'h6 : _GEN_474; // @[Filter.scala 204:102]
  wire [3:0] _GEN_476 = 8'h35 == _T_40[7:0] ? 4'h0 : _GEN_475; // @[Filter.scala 204:102]
  wire [3:0] _GEN_477 = 8'h36 == _T_40[7:0] ? 4'h0 : _GEN_476; // @[Filter.scala 204:102]
  wire [3:0] _GEN_478 = 8'h37 == _T_40[7:0] ? 4'h0 : _GEN_477; // @[Filter.scala 204:102]
  wire [3:0] _GEN_479 = 8'h38 == _T_40[7:0] ? 4'h2 : _GEN_478; // @[Filter.scala 204:102]
  wire [3:0] _GEN_480 = 8'h39 == _T_40[7:0] ? 4'h0 : _GEN_479; // @[Filter.scala 204:102]
  wire [3:0] _GEN_481 = 8'h3a == _T_40[7:0] ? 4'h0 : _GEN_480; // @[Filter.scala 204:102]
  wire [3:0] _GEN_482 = 8'h3b == _T_40[7:0] ? 4'h0 : _GEN_481; // @[Filter.scala 204:102]
  wire [3:0] _GEN_483 = 8'h3c == _T_40[7:0] ? 4'h0 : _GEN_482; // @[Filter.scala 204:102]
  wire [3:0] _GEN_484 = 8'h3d == _T_40[7:0] ? 4'h0 : _GEN_483; // @[Filter.scala 204:102]
  wire [3:0] _GEN_485 = 8'h3e == _T_40[7:0] ? 4'h0 : _GEN_484; // @[Filter.scala 204:102]
  wire [3:0] _GEN_486 = 8'h3f == _T_40[7:0] ? 4'h0 : _GEN_485; // @[Filter.scala 204:102]
  wire [3:0] _GEN_487 = 8'h40 == _T_40[7:0] ? 4'h0 : _GEN_486; // @[Filter.scala 204:102]
  wire [3:0] _GEN_488 = 8'h41 == _T_40[7:0] ? 4'h0 : _GEN_487; // @[Filter.scala 204:102]
  wire [3:0] _GEN_489 = 8'h42 == _T_40[7:0] ? 4'h0 : _GEN_488; // @[Filter.scala 204:102]
  wire [3:0] _GEN_490 = 8'h43 == _T_40[7:0] ? 4'h0 : _GEN_489; // @[Filter.scala 204:102]
  wire [3:0] _GEN_491 = 8'h44 == _T_40[7:0] ? 4'h1 : _GEN_490; // @[Filter.scala 204:102]
  wire [3:0] _GEN_492 = 8'h45 == _T_40[7:0] ? 4'h4 : _GEN_491; // @[Filter.scala 204:102]
  wire [3:0] _GEN_493 = 8'h46 == _T_40[7:0] ? 4'hb : _GEN_492; // @[Filter.scala 204:102]
  wire [3:0] _GEN_494 = 8'h47 == _T_40[7:0] ? 4'h0 : _GEN_493; // @[Filter.scala 204:102]
  wire [3:0] _GEN_495 = 8'h48 == _T_40[7:0] ? 4'h0 : _GEN_494; // @[Filter.scala 204:102]
  wire [3:0] _GEN_496 = 8'h49 == _T_40[7:0] ? 4'h0 : _GEN_495; // @[Filter.scala 204:102]
  wire [3:0] _GEN_497 = 8'h4a == _T_40[7:0] ? 4'h6 : _GEN_496; // @[Filter.scala 204:102]
  wire [3:0] _GEN_498 = 8'h4b == _T_40[7:0] ? 4'h0 : _GEN_497; // @[Filter.scala 204:102]
  wire [3:0] _GEN_499 = 8'h4c == _T_40[7:0] ? 4'h3 : _GEN_498; // @[Filter.scala 204:102]
  wire [3:0] _GEN_500 = 8'h4d == _T_40[7:0] ? 4'h3 : _GEN_499; // @[Filter.scala 204:102]
  wire [3:0] _GEN_501 = 8'h4e == _T_40[7:0] ? 4'h2 : _GEN_500; // @[Filter.scala 204:102]
  wire [3:0] _GEN_502 = 8'h4f == _T_40[7:0] ? 4'h0 : _GEN_501; // @[Filter.scala 204:102]
  wire [3:0] _GEN_503 = 8'h50 == _T_40[7:0] ? 4'h0 : _GEN_502; // @[Filter.scala 204:102]
  wire [3:0] _GEN_504 = 8'h51 == _T_40[7:0] ? 4'h0 : _GEN_503; // @[Filter.scala 204:102]
  wire [3:0] _GEN_505 = 8'h52 == _T_40[7:0] ? 4'h0 : _GEN_504; // @[Filter.scala 204:102]
  wire [3:0] _GEN_506 = 8'h53 == _T_40[7:0] ? 4'h0 : _GEN_505; // @[Filter.scala 204:102]
  wire [3:0] _GEN_507 = 8'h54 == _T_40[7:0] ? 4'h0 : _GEN_506; // @[Filter.scala 204:102]
  wire [3:0] _GEN_508 = 8'h55 == _T_40[7:0] ? 4'h0 : _GEN_507; // @[Filter.scala 204:102]
  wire [3:0] _GEN_509 = 8'h56 == _T_40[7:0] ? 4'h0 : _GEN_508; // @[Filter.scala 204:102]
  wire [3:0] _GEN_510 = 8'h57 == _T_40[7:0] ? 4'h0 : _GEN_509; // @[Filter.scala 204:102]
  wire [3:0] _GEN_511 = 8'h58 == _T_40[7:0] ? 4'h0 : _GEN_510; // @[Filter.scala 204:102]
  wire [3:0] _GEN_512 = 8'h59 == _T_40[7:0] ? 4'h2 : _GEN_511; // @[Filter.scala 204:102]
  wire [3:0] _GEN_513 = 8'h5a == _T_40[7:0] ? 4'h3 : _GEN_512; // @[Filter.scala 204:102]
  wire [3:0] _GEN_514 = 8'h5b == _T_40[7:0] ? 4'h0 : _GEN_513; // @[Filter.scala 204:102]
  wire [3:0] _GEN_515 = 8'h5c == _T_40[7:0] ? 4'h0 : _GEN_514; // @[Filter.scala 204:102]
  wire [3:0] _GEN_516 = 8'h5d == _T_40[7:0] ? 4'h3 : _GEN_515; // @[Filter.scala 204:102]
  wire [3:0] _GEN_517 = 8'h5e == _T_40[7:0] ? 4'hd : _GEN_516; // @[Filter.scala 204:102]
  wire [3:0] _GEN_518 = 8'h5f == _T_40[7:0] ? 4'h3 : _GEN_517; // @[Filter.scala 204:102]
  wire [3:0] _GEN_519 = 8'h60 == _T_40[7:0] ? 4'h0 : _GEN_518; // @[Filter.scala 204:102]
  wire [3:0] _GEN_520 = 8'h61 == _T_40[7:0] ? 4'h6 : _GEN_519; // @[Filter.scala 204:102]
  wire [3:0] _GEN_521 = 8'h62 == _T_40[7:0] ? 4'h0 : _GEN_520; // @[Filter.scala 204:102]
  wire [3:0] _GEN_522 = 8'h63 == _T_40[7:0] ? 4'h2 : _GEN_521; // @[Filter.scala 204:102]
  wire [3:0] _GEN_523 = 8'h64 == _T_40[7:0] ? 4'h0 : _GEN_522; // @[Filter.scala 204:102]
  wire [3:0] _GEN_524 = 8'h65 == _T_40[7:0] ? 4'h0 : _GEN_523; // @[Filter.scala 204:102]
  wire [3:0] _GEN_525 = 8'h66 == _T_40[7:0] ? 4'h0 : _GEN_524; // @[Filter.scala 204:102]
  wire [3:0] _GEN_526 = 8'h67 == _T_40[7:0] ? 4'h0 : _GEN_525; // @[Filter.scala 204:102]
  wire [3:0] _GEN_527 = 8'h68 == _T_40[7:0] ? 4'h0 : _GEN_526; // @[Filter.scala 204:102]
  wire [3:0] _GEN_528 = 8'h69 == _T_40[7:0] ? 4'h0 : _GEN_527; // @[Filter.scala 204:102]
  wire [3:0] _GEN_529 = 8'h6a == _T_40[7:0] ? 4'h0 : _GEN_528; // @[Filter.scala 204:102]
  wire [3:0] _GEN_530 = 8'h6b == _T_40[7:0] ? 4'h0 : _GEN_529; // @[Filter.scala 204:102]
  wire [3:0] _GEN_531 = 8'h6c == _T_40[7:0] ? 4'h0 : _GEN_530; // @[Filter.scala 204:102]
  wire [3:0] _GEN_532 = 8'h6d == _T_40[7:0] ? 4'h0 : _GEN_531; // @[Filter.scala 204:102]
  wire [3:0] _GEN_533 = 8'h6e == _T_40[7:0] ? 4'h2 : _GEN_532; // @[Filter.scala 204:102]
  wire [3:0] _GEN_534 = 8'h6f == _T_40[7:0] ? 4'h0 : _GEN_533; // @[Filter.scala 204:102]
  wire [3:0] _GEN_535 = 8'h70 == _T_40[7:0] ? 4'h0 : _GEN_534; // @[Filter.scala 204:102]
  wire [3:0] _GEN_536 = 8'h71 == _T_40[7:0] ? 4'h0 : _GEN_535; // @[Filter.scala 204:102]
  wire [3:0] _GEN_537 = 8'h72 == _T_40[7:0] ? 4'h6 : _GEN_536; // @[Filter.scala 204:102]
  wire [3:0] _GEN_538 = 8'h73 == _T_40[7:0] ? 4'he : _GEN_537; // @[Filter.scala 204:102]
  wire [3:0] _GEN_539 = 8'h74 == _T_40[7:0] ? 4'h6 : _GEN_538; // @[Filter.scala 204:102]
  wire [3:0] _GEN_540 = 8'h75 == _T_40[7:0] ? 4'h0 : _GEN_539; // @[Filter.scala 204:102]
  wire [3:0] _GEN_541 = 8'h76 == _T_40[7:0] ? 4'h6 : _GEN_540; // @[Filter.scala 204:102]
  wire [3:0] _GEN_542 = 8'h77 == _T_40[7:0] ? 4'h3 : _GEN_541; // @[Filter.scala 204:102]
  wire [3:0] _GEN_543 = 8'h78 == _T_40[7:0] ? 4'h4 : _GEN_542; // @[Filter.scala 204:102]
  wire [3:0] _GEN_544 = 8'h79 == _T_40[7:0] ? 4'h1 : _GEN_543; // @[Filter.scala 204:102]
  wire [3:0] _GEN_545 = 8'h7a == _T_40[7:0] ? 4'h0 : _GEN_544; // @[Filter.scala 204:102]
  wire [3:0] _GEN_546 = 8'h7b == _T_40[7:0] ? 4'h0 : _GEN_545; // @[Filter.scala 204:102]
  wire [3:0] _GEN_547 = 8'h7c == _T_40[7:0] ? 4'h0 : _GEN_546; // @[Filter.scala 204:102]
  wire [3:0] _GEN_548 = 8'h7d == _T_40[7:0] ? 4'h0 : _GEN_547; // @[Filter.scala 204:102]
  wire [3:0] _GEN_549 = 8'h7e == _T_40[7:0] ? 4'h0 : _GEN_548; // @[Filter.scala 204:102]
  wire [3:0] _GEN_550 = 8'h7f == _T_40[7:0] ? 4'h0 : _GEN_549; // @[Filter.scala 204:102]
  wire [3:0] _GEN_551 = 8'h80 == _T_40[7:0] ? 4'h0 : _GEN_550; // @[Filter.scala 204:102]
  wire [3:0] _GEN_552 = 8'h81 == _T_40[7:0] ? 4'h0 : _GEN_551; // @[Filter.scala 204:102]
  wire [3:0] _GEN_553 = 8'h82 == _T_40[7:0] ? 4'h2 : _GEN_552; // @[Filter.scala 204:102]
  wire [3:0] _GEN_554 = 8'h83 == _T_40[7:0] ? 4'h3 : _GEN_553; // @[Filter.scala 204:102]
  wire [3:0] _GEN_555 = 8'h84 == _T_40[7:0] ? 4'h6 : _GEN_554; // @[Filter.scala 204:102]
  wire [3:0] _GEN_556 = 8'h85 == _T_40[7:0] ? 4'h6 : _GEN_555; // @[Filter.scala 204:102]
  wire [3:0] _GEN_557 = 8'h86 == _T_40[7:0] ? 4'he : _GEN_556; // @[Filter.scala 204:102]
  wire [3:0] _GEN_558 = 8'h87 == _T_40[7:0] ? 4'ha : _GEN_557; // @[Filter.scala 204:102]
  wire [3:0] _GEN_559 = 8'h88 == _T_40[7:0] ? 4'h6 : _GEN_558; // @[Filter.scala 204:102]
  wire [3:0] _GEN_560 = 8'h89 == _T_40[7:0] ? 4'ha : _GEN_559; // @[Filter.scala 204:102]
  wire [3:0] _GEN_561 = 8'h8a == _T_40[7:0] ? 4'he : _GEN_560; // @[Filter.scala 204:102]
  wire [3:0] _GEN_562 = 8'h8b == _T_40[7:0] ? 4'h3 : _GEN_561; // @[Filter.scala 204:102]
  wire [3:0] _GEN_563 = 8'h8c == _T_40[7:0] ? 4'h3 : _GEN_562; // @[Filter.scala 204:102]
  wire [3:0] _GEN_564 = 8'h8d == _T_40[7:0] ? 4'h0 : _GEN_563; // @[Filter.scala 204:102]
  wire [3:0] _GEN_565 = 8'h8e == _T_40[7:0] ? 4'h2 : _GEN_564; // @[Filter.scala 204:102]
  wire [3:0] _GEN_566 = 8'h8f == _T_40[7:0] ? 4'h0 : _GEN_565; // @[Filter.scala 204:102]
  wire [3:0] _GEN_567 = 8'h90 == _T_40[7:0] ? 4'h0 : _GEN_566; // @[Filter.scala 204:102]
  wire [3:0] _GEN_568 = 8'h91 == _T_40[7:0] ? 4'h0 : _GEN_567; // @[Filter.scala 204:102]
  wire [3:0] _GEN_569 = 8'h92 == _T_40[7:0] ? 4'h0 : _GEN_568; // @[Filter.scala 204:102]
  wire [3:0] _GEN_570 = 8'h93 == _T_40[7:0] ? 4'h0 : _GEN_569; // @[Filter.scala 204:102]
  wire [3:0] _GEN_571 = 8'h94 == _T_40[7:0] ? 4'h0 : _GEN_570; // @[Filter.scala 204:102]
  wire [3:0] _GEN_572 = 8'h95 == _T_40[7:0] ? 4'h0 : _GEN_571; // @[Filter.scala 204:102]
  wire [3:0] _GEN_573 = 8'h96 == _T_40[7:0] ? 4'h0 : _GEN_572; // @[Filter.scala 204:102]
  wire [3:0] _GEN_574 = 8'h97 == _T_40[7:0] ? 4'h2 : _GEN_573; // @[Filter.scala 204:102]
  wire [3:0] _GEN_575 = 8'h98 == _T_40[7:0] ? 4'h2 : _GEN_574; // @[Filter.scala 204:102]
  wire [3:0] _GEN_576 = 8'h99 == _T_40[7:0] ? 4'h1 : _GEN_575; // @[Filter.scala 204:102]
  wire [3:0] _GEN_577 = 8'h9a == _T_40[7:0] ? 4'h3 : _GEN_576; // @[Filter.scala 204:102]
  wire [3:0] _GEN_578 = 8'h9b == _T_40[7:0] ? 4'he : _GEN_577; // @[Filter.scala 204:102]
  wire [3:0] _GEN_579 = 8'h9c == _T_40[7:0] ? 4'he : _GEN_578; // @[Filter.scala 204:102]
  wire [3:0] _GEN_580 = 8'h9d == _T_40[7:0] ? 4'h0 : _GEN_579; // @[Filter.scala 204:102]
  wire [3:0] _GEN_581 = 8'h9e == _T_40[7:0] ? 4'he : _GEN_580; // @[Filter.scala 204:102]
  wire [3:0] _GEN_582 = 8'h9f == _T_40[7:0] ? 4'he : _GEN_581; // @[Filter.scala 204:102]
  wire [3:0] _GEN_583 = 8'ha0 == _T_40[7:0] ? 4'h3 : _GEN_582; // @[Filter.scala 204:102]
  wire [3:0] _GEN_584 = 8'ha1 == _T_40[7:0] ? 4'h1 : _GEN_583; // @[Filter.scala 204:102]
  wire [3:0] _GEN_585 = 8'ha2 == _T_40[7:0] ? 4'h2 : _GEN_584; // @[Filter.scala 204:102]
  wire [3:0] _GEN_586 = 8'ha3 == _T_40[7:0] ? 4'h2 : _GEN_585; // @[Filter.scala 204:102]
  wire [3:0] _GEN_587 = 8'ha4 == _T_40[7:0] ? 4'h0 : _GEN_586; // @[Filter.scala 204:102]
  wire [3:0] _GEN_588 = 8'ha5 == _T_40[7:0] ? 4'h0 : _GEN_587; // @[Filter.scala 204:102]
  wire [3:0] _GEN_589 = 8'ha6 == _T_40[7:0] ? 4'h0 : _GEN_588; // @[Filter.scala 204:102]
  wire [3:0] _GEN_590 = 8'ha7 == _T_40[7:0] ? 4'h0 : _GEN_589; // @[Filter.scala 204:102]
  wire [3:0] _GEN_591 = 8'ha8 == _T_40[7:0] ? 4'h0 : _GEN_590; // @[Filter.scala 204:102]
  wire [3:0] _GEN_592 = 8'ha9 == _T_40[7:0] ? 4'h0 : _GEN_591; // @[Filter.scala 204:102]
  wire [3:0] _GEN_593 = 8'haa == _T_40[7:0] ? 4'h0 : _GEN_592; // @[Filter.scala 204:102]
  wire [3:0] _GEN_594 = 8'hab == _T_40[7:0] ? 4'h0 : _GEN_593; // @[Filter.scala 204:102]
  wire [3:0] _GEN_595 = 8'hac == _T_40[7:0] ? 4'h2 : _GEN_594; // @[Filter.scala 204:102]
  wire [3:0] _GEN_596 = 8'had == _T_40[7:0] ? 4'h3 : _GEN_595; // @[Filter.scala 204:102]
  wire [3:0] _GEN_597 = 8'hae == _T_40[7:0] ? 4'h4 : _GEN_596; // @[Filter.scala 204:102]
  wire [3:0] _GEN_598 = 8'haf == _T_40[7:0] ? 4'h3 : _GEN_597; // @[Filter.scala 204:102]
  wire [3:0] _GEN_599 = 8'hb0 == _T_40[7:0] ? 4'h4 : _GEN_598; // @[Filter.scala 204:102]
  wire [3:0] _GEN_600 = 8'hb1 == _T_40[7:0] ? 4'h3 : _GEN_599; // @[Filter.scala 204:102]
  wire [3:0] _GEN_601 = 8'hb2 == _T_40[7:0] ? 4'h0 : _GEN_600; // @[Filter.scala 204:102]
  wire [3:0] _GEN_602 = 8'hb3 == _T_40[7:0] ? 4'h3 : _GEN_601; // @[Filter.scala 204:102]
  wire [3:0] _GEN_603 = 8'hb4 == _T_40[7:0] ? 4'h4 : _GEN_602; // @[Filter.scala 204:102]
  wire [3:0] _GEN_604 = 8'hb5 == _T_40[7:0] ? 4'h3 : _GEN_603; // @[Filter.scala 204:102]
  wire [3:0] _GEN_605 = 8'hb6 == _T_40[7:0] ? 4'h4 : _GEN_604; // @[Filter.scala 204:102]
  wire [3:0] _GEN_606 = 8'hb7 == _T_40[7:0] ? 4'h3 : _GEN_605; // @[Filter.scala 204:102]
  wire [3:0] _GEN_607 = 8'hb8 == _T_40[7:0] ? 4'h2 : _GEN_606; // @[Filter.scala 204:102]
  wire [3:0] _GEN_608 = 8'hb9 == _T_40[7:0] ? 4'h0 : _GEN_607; // @[Filter.scala 204:102]
  wire [3:0] _GEN_609 = 8'hba == _T_40[7:0] ? 4'h0 : _GEN_608; // @[Filter.scala 204:102]
  wire [3:0] _GEN_610 = 8'hbb == _T_40[7:0] ? 4'h0 : _GEN_609; // @[Filter.scala 204:102]
  wire [3:0] _GEN_611 = 8'hbc == _T_40[7:0] ? 4'h0 : _GEN_610; // @[Filter.scala 204:102]
  wire [3:0] _GEN_612 = 8'hbd == _T_40[7:0] ? 4'h0 : _GEN_611; // @[Filter.scala 204:102]
  wire [3:0] _GEN_613 = 8'hbe == _T_40[7:0] ? 4'h0 : _GEN_612; // @[Filter.scala 204:102]
  wire [3:0] _GEN_614 = 8'hbf == _T_40[7:0] ? 4'h0 : _GEN_613; // @[Filter.scala 204:102]
  wire [3:0] _GEN_615 = 8'hc0 == _T_40[7:0] ? 4'h0 : _GEN_614; // @[Filter.scala 204:102]
  wire [3:0] _GEN_616 = 8'hc1 == _T_40[7:0] ? 4'h0 : _GEN_615; // @[Filter.scala 204:102]
  wire [3:0] _GEN_617 = 8'hc2 == _T_40[7:0] ? 4'h8 : _GEN_616; // @[Filter.scala 204:102]
  wire [3:0] _GEN_618 = 8'hc3 == _T_40[7:0] ? 4'hc : _GEN_617; // @[Filter.scala 204:102]
  wire [3:0] _GEN_619 = 8'hc4 == _T_40[7:0] ? 4'h0 : _GEN_618; // @[Filter.scala 204:102]
  wire [3:0] _GEN_620 = 8'hc5 == _T_40[7:0] ? 4'h2 : _GEN_619; // @[Filter.scala 204:102]
  wire [3:0] _GEN_621 = 8'hc6 == _T_40[7:0] ? 4'h3 : _GEN_620; // @[Filter.scala 204:102]
  wire [3:0] _GEN_622 = 8'hc7 == _T_40[7:0] ? 4'h2 : _GEN_621; // @[Filter.scala 204:102]
  wire [3:0] _GEN_623 = 8'hc8 == _T_40[7:0] ? 4'h3 : _GEN_622; // @[Filter.scala 204:102]
  wire [3:0] _GEN_624 = 8'hc9 == _T_40[7:0] ? 4'h2 : _GEN_623; // @[Filter.scala 204:102]
  wire [3:0] _GEN_625 = 8'hca == _T_40[7:0] ? 4'h0 : _GEN_624; // @[Filter.scala 204:102]
  wire [3:0] _GEN_626 = 8'hcb == _T_40[7:0] ? 4'hc : _GEN_625; // @[Filter.scala 204:102]
  wire [3:0] _GEN_627 = 8'hcc == _T_40[7:0] ? 4'h8 : _GEN_626; // @[Filter.scala 204:102]
  wire [3:0] _GEN_628 = 8'hcd == _T_40[7:0] ? 4'h0 : _GEN_627; // @[Filter.scala 204:102]
  wire [3:0] _GEN_629 = 8'hce == _T_40[7:0] ? 4'h0 : _GEN_628; // @[Filter.scala 204:102]
  wire [3:0] _GEN_630 = 8'hcf == _T_40[7:0] ? 4'h0 : _GEN_629; // @[Filter.scala 204:102]
  wire [3:0] _GEN_631 = 8'hd0 == _T_40[7:0] ? 4'h0 : _GEN_630; // @[Filter.scala 204:102]
  wire [3:0] _GEN_632 = 8'hd1 == _T_40[7:0] ? 4'h0 : _GEN_631; // @[Filter.scala 204:102]
  wire [3:0] _GEN_633 = 8'hd2 == _T_40[7:0] ? 4'h0 : _GEN_632; // @[Filter.scala 204:102]
  wire [3:0] _GEN_634 = 8'hd3 == _T_40[7:0] ? 4'h0 : _GEN_633; // @[Filter.scala 204:102]
  wire [3:0] _GEN_635 = 8'hd4 == _T_40[7:0] ? 4'h0 : _GEN_634; // @[Filter.scala 204:102]
  wire [3:0] _GEN_636 = 8'hd5 == _T_40[7:0] ? 4'h0 : _GEN_635; // @[Filter.scala 204:102]
  wire [3:0] _GEN_637 = 8'hd6 == _T_40[7:0] ? 4'h0 : _GEN_636; // @[Filter.scala 204:102]
  wire [3:0] _GEN_638 = 8'hd7 == _T_40[7:0] ? 4'h3 : _GEN_637; // @[Filter.scala 204:102]
  wire [3:0] _GEN_639 = 8'hd8 == _T_40[7:0] ? 4'h6 : _GEN_638; // @[Filter.scala 204:102]
  wire [3:0] _GEN_640 = 8'hd9 == _T_40[7:0] ? 4'h0 : _GEN_639; // @[Filter.scala 204:102]
  wire [3:0] _GEN_641 = 8'hda == _T_40[7:0] ? 4'hb : _GEN_640; // @[Filter.scala 204:102]
  wire [3:0] _GEN_642 = 8'hdb == _T_40[7:0] ? 4'h1 : _GEN_641; // @[Filter.scala 204:102]
  wire [3:0] _GEN_643 = 8'hdc == _T_40[7:0] ? 4'h4 : _GEN_642; // @[Filter.scala 204:102]
  wire [3:0] _GEN_644 = 8'hdd == _T_40[7:0] ? 4'h1 : _GEN_643; // @[Filter.scala 204:102]
  wire [3:0] _GEN_645 = 8'hde == _T_40[7:0] ? 4'hb : _GEN_644; // @[Filter.scala 204:102]
  wire [3:0] _GEN_646 = 8'hdf == _T_40[7:0] ? 4'h0 : _GEN_645; // @[Filter.scala 204:102]
  wire [3:0] _GEN_647 = 8'he0 == _T_40[7:0] ? 4'h6 : _GEN_646; // @[Filter.scala 204:102]
  wire [3:0] _GEN_648 = 8'he1 == _T_40[7:0] ? 4'h3 : _GEN_647; // @[Filter.scala 204:102]
  wire [3:0] _GEN_649 = 8'he2 == _T_40[7:0] ? 4'h0 : _GEN_648; // @[Filter.scala 204:102]
  wire [3:0] _GEN_650 = 8'he3 == _T_40[7:0] ? 4'h0 : _GEN_649; // @[Filter.scala 204:102]
  wire [3:0] _GEN_651 = 8'he4 == _T_40[7:0] ? 4'h0 : _GEN_650; // @[Filter.scala 204:102]
  wire [3:0] _GEN_652 = 8'he5 == _T_40[7:0] ? 4'h0 : _GEN_651; // @[Filter.scala 204:102]
  wire [3:0] _GEN_653 = 8'he6 == _T_40[7:0] ? 4'h0 : _GEN_652; // @[Filter.scala 204:102]
  wire [3:0] _GEN_654 = 8'he7 == _T_40[7:0] ? 4'h0 : _GEN_653; // @[Filter.scala 204:102]
  wire [3:0] _GEN_655 = 8'he8 == _T_40[7:0] ? 4'h0 : _GEN_654; // @[Filter.scala 204:102]
  wire [3:0] _GEN_656 = 8'he9 == _T_40[7:0] ? 4'h0 : _GEN_655; // @[Filter.scala 204:102]
  wire [3:0] _GEN_657 = 8'hea == _T_40[7:0] ? 4'h0 : _GEN_656; // @[Filter.scala 204:102]
  wire [3:0] _GEN_658 = 8'heb == _T_40[7:0] ? 4'h0 : _GEN_657; // @[Filter.scala 204:102]
  wire [3:0] _GEN_659 = 8'hec == _T_40[7:0] ? 4'h0 : _GEN_658; // @[Filter.scala 204:102]
  wire [3:0] _GEN_660 = 8'hed == _T_40[7:0] ? 4'h0 : _GEN_659; // @[Filter.scala 204:102]
  wire [3:0] _GEN_661 = 8'hee == _T_40[7:0] ? 4'h0 : _GEN_660; // @[Filter.scala 204:102]
  wire [3:0] _GEN_662 = 8'hef == _T_40[7:0] ? 4'h0 : _GEN_661; // @[Filter.scala 204:102]
  wire [3:0] _GEN_663 = 8'hf0 == _T_40[7:0] ? 4'h0 : _GEN_662; // @[Filter.scala 204:102]
  wire [3:0] _GEN_664 = 8'hf1 == _T_40[7:0] ? 4'h0 : _GEN_663; // @[Filter.scala 204:102]
  wire [3:0] _GEN_665 = 8'hf2 == _T_40[7:0] ? 4'h0 : _GEN_664; // @[Filter.scala 204:102]
  wire [3:0] _GEN_666 = 8'hf3 == _T_40[7:0] ? 4'h0 : _GEN_665; // @[Filter.scala 204:102]
  wire [3:0] _GEN_667 = 8'hf4 == _T_40[7:0] ? 4'h0 : _GEN_666; // @[Filter.scala 204:102]
  wire [3:0] _GEN_668 = 8'hf5 == _T_40[7:0] ? 4'h0 : _GEN_667; // @[Filter.scala 204:102]
  wire [3:0] _GEN_669 = 8'hf6 == _T_40[7:0] ? 4'h0 : _GEN_668; // @[Filter.scala 204:102]
  wire [3:0] _GEN_670 = 8'hf7 == _T_40[7:0] ? 4'h0 : _GEN_669; // @[Filter.scala 204:102]
  wire [3:0] _GEN_671 = 8'hf8 == _T_40[7:0] ? 4'h0 : _GEN_670; // @[Filter.scala 204:102]
  wire [3:0] _GEN_672 = 8'hf9 == _T_40[7:0] ? 4'h0 : _GEN_671; // @[Filter.scala 204:102]
  wire [3:0] _GEN_673 = 8'hfa == _T_40[7:0] ? 4'h0 : _GEN_672; // @[Filter.scala 204:102]
  wire [3:0] _GEN_674 = 8'hfb == _T_40[7:0] ? 4'h0 : _GEN_673; // @[Filter.scala 204:102]
  wire [6:0] _GEN_11215 = {{3'd0}, _GEN_674}; // @[Filter.scala 204:102]
  wire [10:0] _T_47 = _GEN_11215 * 7'h46; // @[Filter.scala 204:102]
  wire [10:0] _GEN_11216 = {{2'd0}, _T_42}; // @[Filter.scala 204:69]
  wire [10:0] _T_49 = _GEN_11216 + _T_47; // @[Filter.scala 204:69]
  wire [3:0] _GEN_683 = 8'h8 == _T_40[7:0] ? 4'h3 : 4'h0; // @[Filter.scala 204:142]
  wire [3:0] _GEN_684 = 8'h9 == _T_40[7:0] ? 4'h6 : _GEN_683; // @[Filter.scala 204:142]
  wire [3:0] _GEN_685 = 8'ha == _T_40[7:0] ? 4'h6 : _GEN_684; // @[Filter.scala 204:142]
  wire [3:0] _GEN_686 = 8'hb == _T_40[7:0] ? 4'h6 : _GEN_685; // @[Filter.scala 204:142]
  wire [3:0] _GEN_687 = 8'hc == _T_40[7:0] ? 4'h3 : _GEN_686; // @[Filter.scala 204:142]
  wire [3:0] _GEN_688 = 8'hd == _T_40[7:0] ? 4'h0 : _GEN_687; // @[Filter.scala 204:142]
  wire [3:0] _GEN_689 = 8'he == _T_40[7:0] ? 4'h0 : _GEN_688; // @[Filter.scala 204:142]
  wire [3:0] _GEN_690 = 8'hf == _T_40[7:0] ? 4'h0 : _GEN_689; // @[Filter.scala 204:142]
  wire [3:0] _GEN_691 = 8'h10 == _T_40[7:0] ? 4'h0 : _GEN_690; // @[Filter.scala 204:142]
  wire [3:0] _GEN_692 = 8'h11 == _T_40[7:0] ? 4'h0 : _GEN_691; // @[Filter.scala 204:142]
  wire [3:0] _GEN_693 = 8'h12 == _T_40[7:0] ? 4'h0 : _GEN_692; // @[Filter.scala 204:142]
  wire [3:0] _GEN_694 = 8'h13 == _T_40[7:0] ? 4'h0 : _GEN_693; // @[Filter.scala 204:142]
  wire [3:0] _GEN_695 = 8'h14 == _T_40[7:0] ? 4'h0 : _GEN_694; // @[Filter.scala 204:142]
  wire [3:0] _GEN_696 = 8'h15 == _T_40[7:0] ? 4'h0 : _GEN_695; // @[Filter.scala 204:142]
  wire [3:0] _GEN_697 = 8'h16 == _T_40[7:0] ? 4'h0 : _GEN_696; // @[Filter.scala 204:142]
  wire [3:0] _GEN_698 = 8'h17 == _T_40[7:0] ? 4'h0 : _GEN_697; // @[Filter.scala 204:142]
  wire [3:0] _GEN_699 = 8'h18 == _T_40[7:0] ? 4'h0 : _GEN_698; // @[Filter.scala 204:142]
  wire [3:0] _GEN_700 = 8'h19 == _T_40[7:0] ? 4'h0 : _GEN_699; // @[Filter.scala 204:142]
  wire [3:0] _GEN_701 = 8'h1a == _T_40[7:0] ? 4'h0 : _GEN_700; // @[Filter.scala 204:142]
  wire [3:0] _GEN_702 = 8'h1b == _T_40[7:0] ? 4'h0 : _GEN_701; // @[Filter.scala 204:142]
  wire [3:0] _GEN_703 = 8'h1c == _T_40[7:0] ? 4'h6 : _GEN_702; // @[Filter.scala 204:142]
  wire [3:0] _GEN_704 = 8'h1d == _T_40[7:0] ? 4'h3 : _GEN_703; // @[Filter.scala 204:142]
  wire [3:0] _GEN_705 = 8'h1e == _T_40[7:0] ? 4'h0 : _GEN_704; // @[Filter.scala 204:142]
  wire [3:0] _GEN_706 = 8'h1f == _T_40[7:0] ? 4'h0 : _GEN_705; // @[Filter.scala 204:142]
  wire [3:0] _GEN_707 = 8'h20 == _T_40[7:0] ? 4'h0 : _GEN_706; // @[Filter.scala 204:142]
  wire [3:0] _GEN_708 = 8'h21 == _T_40[7:0] ? 4'h3 : _GEN_707; // @[Filter.scala 204:142]
  wire [3:0] _GEN_709 = 8'h22 == _T_40[7:0] ? 4'h6 : _GEN_708; // @[Filter.scala 204:142]
  wire [3:0] _GEN_710 = 8'h23 == _T_40[7:0] ? 4'h0 : _GEN_709; // @[Filter.scala 204:142]
  wire [3:0] _GEN_711 = 8'h24 == _T_40[7:0] ? 4'h0 : _GEN_710; // @[Filter.scala 204:142]
  wire [3:0] _GEN_712 = 8'h25 == _T_40[7:0] ? 4'h0 : _GEN_711; // @[Filter.scala 204:142]
  wire [3:0] _GEN_713 = 8'h26 == _T_40[7:0] ? 4'h0 : _GEN_712; // @[Filter.scala 204:142]
  wire [3:0] _GEN_714 = 8'h27 == _T_40[7:0] ? 4'h0 : _GEN_713; // @[Filter.scala 204:142]
  wire [3:0] _GEN_715 = 8'h28 == _T_40[7:0] ? 4'h0 : _GEN_714; // @[Filter.scala 204:142]
  wire [3:0] _GEN_716 = 8'h29 == _T_40[7:0] ? 4'h0 : _GEN_715; // @[Filter.scala 204:142]
  wire [3:0] _GEN_717 = 8'h2a == _T_40[7:0] ? 4'h0 : _GEN_716; // @[Filter.scala 204:142]
  wire [3:0] _GEN_718 = 8'h2b == _T_40[7:0] ? 4'h0 : _GEN_717; // @[Filter.scala 204:142]
  wire [3:0] _GEN_719 = 8'h2c == _T_40[7:0] ? 4'h0 : _GEN_718; // @[Filter.scala 204:142]
  wire [3:0] _GEN_720 = 8'h2d == _T_40[7:0] ? 4'h0 : _GEN_719; // @[Filter.scala 204:142]
  wire [3:0] _GEN_721 = 8'h2e == _T_40[7:0] ? 4'h0 : _GEN_720; // @[Filter.scala 204:142]
  wire [3:0] _GEN_722 = 8'h2f == _T_40[7:0] ? 4'h0 : _GEN_721; // @[Filter.scala 204:142]
  wire [3:0] _GEN_723 = 8'h30 == _T_40[7:0] ? 4'h6 : _GEN_722; // @[Filter.scala 204:142]
  wire [3:0] _GEN_724 = 8'h31 == _T_40[7:0] ? 4'h3 : _GEN_723; // @[Filter.scala 204:142]
  wire [3:0] _GEN_725 = 8'h32 == _T_40[7:0] ? 4'h0 : _GEN_724; // @[Filter.scala 204:142]
  wire [3:0] _GEN_726 = 8'h33 == _T_40[7:0] ? 4'h1 : _GEN_725; // @[Filter.scala 204:142]
  wire [3:0] _GEN_727 = 8'h34 == _T_40[7:0] ? 4'h1 : _GEN_726; // @[Filter.scala 204:142]
  wire [3:0] _GEN_728 = 8'h35 == _T_40[7:0] ? 4'h0 : _GEN_727; // @[Filter.scala 204:142]
  wire [3:0] _GEN_729 = 8'h36 == _T_40[7:0] ? 4'h0 : _GEN_728; // @[Filter.scala 204:142]
  wire [3:0] _GEN_730 = 8'h37 == _T_40[7:0] ? 4'h0 : _GEN_729; // @[Filter.scala 204:142]
  wire [3:0] _GEN_731 = 8'h38 == _T_40[7:0] ? 4'h6 : _GEN_730; // @[Filter.scala 204:142]
  wire [3:0] _GEN_732 = 8'h39 == _T_40[7:0] ? 4'h0 : _GEN_731; // @[Filter.scala 204:142]
  wire [3:0] _GEN_733 = 8'h3a == _T_40[7:0] ? 4'h0 : _GEN_732; // @[Filter.scala 204:142]
  wire [3:0] _GEN_734 = 8'h3b == _T_40[7:0] ? 4'h0 : _GEN_733; // @[Filter.scala 204:142]
  wire [3:0] _GEN_735 = 8'h3c == _T_40[7:0] ? 4'h0 : _GEN_734; // @[Filter.scala 204:142]
  wire [3:0] _GEN_736 = 8'h3d == _T_40[7:0] ? 4'h0 : _GEN_735; // @[Filter.scala 204:142]
  wire [3:0] _GEN_737 = 8'h3e == _T_40[7:0] ? 4'h0 : _GEN_736; // @[Filter.scala 204:142]
  wire [3:0] _GEN_738 = 8'h3f == _T_40[7:0] ? 4'h0 : _GEN_737; // @[Filter.scala 204:142]
  wire [3:0] _GEN_739 = 8'h40 == _T_40[7:0] ? 4'h0 : _GEN_738; // @[Filter.scala 204:142]
  wire [3:0] _GEN_740 = 8'h41 == _T_40[7:0] ? 4'h0 : _GEN_739; // @[Filter.scala 204:142]
  wire [3:0] _GEN_741 = 8'h42 == _T_40[7:0] ? 4'h0 : _GEN_740; // @[Filter.scala 204:142]
  wire [3:0] _GEN_742 = 8'h43 == _T_40[7:0] ? 4'h0 : _GEN_741; // @[Filter.scala 204:142]
  wire [3:0] _GEN_743 = 8'h44 == _T_40[7:0] ? 4'h3 : _GEN_742; // @[Filter.scala 204:142]
  wire [3:0] _GEN_744 = 8'h45 == _T_40[7:0] ? 4'h6 : _GEN_743; // @[Filter.scala 204:142]
  wire [3:0] _GEN_745 = 8'h46 == _T_40[7:0] ? 4'h9 : _GEN_744; // @[Filter.scala 204:142]
  wire [3:0] _GEN_746 = 8'h47 == _T_40[7:0] ? 4'h0 : _GEN_745; // @[Filter.scala 204:142]
  wire [3:0] _GEN_747 = 8'h48 == _T_40[7:0] ? 4'h0 : _GEN_746; // @[Filter.scala 204:142]
  wire [3:0] _GEN_748 = 8'h49 == _T_40[7:0] ? 4'h0 : _GEN_747; // @[Filter.scala 204:142]
  wire [3:0] _GEN_749 = 8'h4a == _T_40[7:0] ? 4'h1 : _GEN_748; // @[Filter.scala 204:142]
  wire [3:0] _GEN_750 = 8'h4b == _T_40[7:0] ? 4'h0 : _GEN_749; // @[Filter.scala 204:142]
  wire [3:0] _GEN_751 = 8'h4c == _T_40[7:0] ? 4'h0 : _GEN_750; // @[Filter.scala 204:142]
  wire [3:0] _GEN_752 = 8'h4d == _T_40[7:0] ? 4'h0 : _GEN_751; // @[Filter.scala 204:142]
  wire [3:0] _GEN_753 = 8'h4e == _T_40[7:0] ? 4'h6 : _GEN_752; // @[Filter.scala 204:142]
  wire [3:0] _GEN_754 = 8'h4f == _T_40[7:0] ? 4'h0 : _GEN_753; // @[Filter.scala 204:142]
  wire [3:0] _GEN_755 = 8'h50 == _T_40[7:0] ? 4'h0 : _GEN_754; // @[Filter.scala 204:142]
  wire [3:0] _GEN_756 = 8'h51 == _T_40[7:0] ? 4'h0 : _GEN_755; // @[Filter.scala 204:142]
  wire [3:0] _GEN_757 = 8'h52 == _T_40[7:0] ? 4'h0 : _GEN_756; // @[Filter.scala 204:142]
  wire [3:0] _GEN_758 = 8'h53 == _T_40[7:0] ? 4'h0 : _GEN_757; // @[Filter.scala 204:142]
  wire [3:0] _GEN_759 = 8'h54 == _T_40[7:0] ? 4'h0 : _GEN_758; // @[Filter.scala 204:142]
  wire [3:0] _GEN_760 = 8'h55 == _T_40[7:0] ? 4'h0 : _GEN_759; // @[Filter.scala 204:142]
  wire [3:0] _GEN_761 = 8'h56 == _T_40[7:0] ? 4'h0 : _GEN_760; // @[Filter.scala 204:142]
  wire [3:0] _GEN_762 = 8'h57 == _T_40[7:0] ? 4'h0 : _GEN_761; // @[Filter.scala 204:142]
  wire [3:0] _GEN_763 = 8'h58 == _T_40[7:0] ? 4'h0 : _GEN_762; // @[Filter.scala 204:142]
  wire [3:0] _GEN_764 = 8'h59 == _T_40[7:0] ? 4'h6 : _GEN_763; // @[Filter.scala 204:142]
  wire [3:0] _GEN_765 = 8'h5a == _T_40[7:0] ? 4'h3 : _GEN_764; // @[Filter.scala 204:142]
  wire [3:0] _GEN_766 = 8'h5b == _T_40[7:0] ? 4'h0 : _GEN_765; // @[Filter.scala 204:142]
  wire [3:0] _GEN_767 = 8'h5c == _T_40[7:0] ? 4'h0 : _GEN_766; // @[Filter.scala 204:142]
  wire [3:0] _GEN_768 = 8'h5d == _T_40[7:0] ? 4'h0 : _GEN_767; // @[Filter.scala 204:142]
  wire [3:0] _GEN_769 = 8'h5e == _T_40[7:0] ? 4'h7 : _GEN_768; // @[Filter.scala 204:142]
  wire [3:0] _GEN_770 = 8'h5f == _T_40[7:0] ? 4'h0 : _GEN_769; // @[Filter.scala 204:142]
  wire [3:0] _GEN_771 = 8'h60 == _T_40[7:0] ? 4'h0 : _GEN_770; // @[Filter.scala 204:142]
  wire [3:0] _GEN_772 = 8'h61 == _T_40[7:0] ? 4'h1 : _GEN_771; // @[Filter.scala 204:142]
  wire [3:0] _GEN_773 = 8'h62 == _T_40[7:0] ? 4'h0 : _GEN_772; // @[Filter.scala 204:142]
  wire [3:0] _GEN_774 = 8'h63 == _T_40[7:0] ? 4'h6 : _GEN_773; // @[Filter.scala 204:142]
  wire [3:0] _GEN_775 = 8'h64 == _T_40[7:0] ? 4'h0 : _GEN_774; // @[Filter.scala 204:142]
  wire [3:0] _GEN_776 = 8'h65 == _T_40[7:0] ? 4'h0 : _GEN_775; // @[Filter.scala 204:142]
  wire [3:0] _GEN_777 = 8'h66 == _T_40[7:0] ? 4'h0 : _GEN_776; // @[Filter.scala 204:142]
  wire [3:0] _GEN_778 = 8'h67 == _T_40[7:0] ? 4'h0 : _GEN_777; // @[Filter.scala 204:142]
  wire [3:0] _GEN_779 = 8'h68 == _T_40[7:0] ? 4'h0 : _GEN_778; // @[Filter.scala 204:142]
  wire [3:0] _GEN_780 = 8'h69 == _T_40[7:0] ? 4'h0 : _GEN_779; // @[Filter.scala 204:142]
  wire [3:0] _GEN_781 = 8'h6a == _T_40[7:0] ? 4'h0 : _GEN_780; // @[Filter.scala 204:142]
  wire [3:0] _GEN_782 = 8'h6b == _T_40[7:0] ? 4'h0 : _GEN_781; // @[Filter.scala 204:142]
  wire [3:0] _GEN_783 = 8'h6c == _T_40[7:0] ? 4'h0 : _GEN_782; // @[Filter.scala 204:142]
  wire [3:0] _GEN_784 = 8'h6d == _T_40[7:0] ? 4'h0 : _GEN_783; // @[Filter.scala 204:142]
  wire [3:0] _GEN_785 = 8'h6e == _T_40[7:0] ? 4'h6 : _GEN_784; // @[Filter.scala 204:142]
  wire [3:0] _GEN_786 = 8'h6f == _T_40[7:0] ? 4'h0 : _GEN_785; // @[Filter.scala 204:142]
  wire [3:0] _GEN_787 = 8'h70 == _T_40[7:0] ? 4'h0 : _GEN_786; // @[Filter.scala 204:142]
  wire [3:0] _GEN_788 = 8'h71 == _T_40[7:0] ? 4'h0 : _GEN_787; // @[Filter.scala 204:142]
  wire [3:0] _GEN_789 = 8'h72 == _T_40[7:0] ? 4'h3 : _GEN_788; // @[Filter.scala 204:142]
  wire [3:0] _GEN_790 = 8'h73 == _T_40[7:0] ? 4'hc : _GEN_789; // @[Filter.scala 204:142]
  wire [3:0] _GEN_791 = 8'h74 == _T_40[7:0] ? 4'h3 : _GEN_790; // @[Filter.scala 204:142]
  wire [3:0] _GEN_792 = 8'h75 == _T_40[7:0] ? 4'h0 : _GEN_791; // @[Filter.scala 204:142]
  wire [3:0] _GEN_793 = 8'h76 == _T_40[7:0] ? 4'h1 : _GEN_792; // @[Filter.scala 204:142]
  wire [3:0] _GEN_794 = 8'h77 == _T_40[7:0] ? 4'h0 : _GEN_793; // @[Filter.scala 204:142]
  wire [3:0] _GEN_795 = 8'h78 == _T_40[7:0] ? 4'h3 : _GEN_794; // @[Filter.scala 204:142]
  wire [3:0] _GEN_796 = 8'h79 == _T_40[7:0] ? 4'h3 : _GEN_795; // @[Filter.scala 204:142]
  wire [3:0] _GEN_797 = 8'h7a == _T_40[7:0] ? 4'h0 : _GEN_796; // @[Filter.scala 204:142]
  wire [3:0] _GEN_798 = 8'h7b == _T_40[7:0] ? 4'h0 : _GEN_797; // @[Filter.scala 204:142]
  wire [3:0] _GEN_799 = 8'h7c == _T_40[7:0] ? 4'h0 : _GEN_798; // @[Filter.scala 204:142]
  wire [3:0] _GEN_800 = 8'h7d == _T_40[7:0] ? 4'h0 : _GEN_799; // @[Filter.scala 204:142]
  wire [3:0] _GEN_801 = 8'h7e == _T_40[7:0] ? 4'h0 : _GEN_800; // @[Filter.scala 204:142]
  wire [3:0] _GEN_802 = 8'h7f == _T_40[7:0] ? 4'h0 : _GEN_801; // @[Filter.scala 204:142]
  wire [3:0] _GEN_803 = 8'h80 == _T_40[7:0] ? 4'h0 : _GEN_802; // @[Filter.scala 204:142]
  wire [3:0] _GEN_804 = 8'h81 == _T_40[7:0] ? 4'h0 : _GEN_803; // @[Filter.scala 204:142]
  wire [3:0] _GEN_805 = 8'h82 == _T_40[7:0] ? 4'h6 : _GEN_804; // @[Filter.scala 204:142]
  wire [3:0] _GEN_806 = 8'h83 == _T_40[7:0] ? 4'h0 : _GEN_805; // @[Filter.scala 204:142]
  wire [3:0] _GEN_807 = 8'h84 == _T_40[7:0] ? 4'h1 : _GEN_806; // @[Filter.scala 204:142]
  wire [3:0] _GEN_808 = 8'h85 == _T_40[7:0] ? 4'h1 : _GEN_807; // @[Filter.scala 204:142]
  wire [3:0] _GEN_809 = 8'h86 == _T_40[7:0] ? 4'ha : _GEN_808; // @[Filter.scala 204:142]
  wire [3:0] _GEN_810 = 8'h87 == _T_40[7:0] ? 4'h4 : _GEN_809; // @[Filter.scala 204:142]
  wire [3:0] _GEN_811 = 8'h88 == _T_40[7:0] ? 4'h1 : _GEN_810; // @[Filter.scala 204:142]
  wire [3:0] _GEN_812 = 8'h89 == _T_40[7:0] ? 4'h4 : _GEN_811; // @[Filter.scala 204:142]
  wire [3:0] _GEN_813 = 8'h8a == _T_40[7:0] ? 4'ha : _GEN_812; // @[Filter.scala 204:142]
  wire [3:0] _GEN_814 = 8'h8b == _T_40[7:0] ? 4'h0 : _GEN_813; // @[Filter.scala 204:142]
  wire [3:0] _GEN_815 = 8'h8c == _T_40[7:0] ? 4'h0 : _GEN_814; // @[Filter.scala 204:142]
  wire [3:0] _GEN_816 = 8'h8d == _T_40[7:0] ? 4'h0 : _GEN_815; // @[Filter.scala 204:142]
  wire [3:0] _GEN_817 = 8'h8e == _T_40[7:0] ? 4'h6 : _GEN_816; // @[Filter.scala 204:142]
  wire [3:0] _GEN_818 = 8'h8f == _T_40[7:0] ? 4'h0 : _GEN_817; // @[Filter.scala 204:142]
  wire [3:0] _GEN_819 = 8'h90 == _T_40[7:0] ? 4'h0 : _GEN_818; // @[Filter.scala 204:142]
  wire [3:0] _GEN_820 = 8'h91 == _T_40[7:0] ? 4'h0 : _GEN_819; // @[Filter.scala 204:142]
  wire [3:0] _GEN_821 = 8'h92 == _T_40[7:0] ? 4'h0 : _GEN_820; // @[Filter.scala 204:142]
  wire [3:0] _GEN_822 = 8'h93 == _T_40[7:0] ? 4'h0 : _GEN_821; // @[Filter.scala 204:142]
  wire [3:0] _GEN_823 = 8'h94 == _T_40[7:0] ? 4'h0 : _GEN_822; // @[Filter.scala 204:142]
  wire [3:0] _GEN_824 = 8'h95 == _T_40[7:0] ? 4'h0 : _GEN_823; // @[Filter.scala 204:142]
  wire [3:0] _GEN_825 = 8'h96 == _T_40[7:0] ? 4'h0 : _GEN_824; // @[Filter.scala 204:142]
  wire [3:0] _GEN_826 = 8'h97 == _T_40[7:0] ? 4'h6 : _GEN_825; // @[Filter.scala 204:142]
  wire [3:0] _GEN_827 = 8'h98 == _T_40[7:0] ? 4'h6 : _GEN_826; // @[Filter.scala 204:142]
  wire [3:0] _GEN_828 = 8'h99 == _T_40[7:0] ? 4'h3 : _GEN_827; // @[Filter.scala 204:142]
  wire [3:0] _GEN_829 = 8'h9a == _T_40[7:0] ? 4'h0 : _GEN_828; // @[Filter.scala 204:142]
  wire [3:0] _GEN_830 = 8'h9b == _T_40[7:0] ? 4'ha : _GEN_829; // @[Filter.scala 204:142]
  wire [3:0] _GEN_831 = 8'h9c == _T_40[7:0] ? 4'ha : _GEN_830; // @[Filter.scala 204:142]
  wire [3:0] _GEN_832 = 8'h9d == _T_40[7:0] ? 4'h0 : _GEN_831; // @[Filter.scala 204:142]
  wire [3:0] _GEN_833 = 8'h9e == _T_40[7:0] ? 4'ha : _GEN_832; // @[Filter.scala 204:142]
  wire [3:0] _GEN_834 = 8'h9f == _T_40[7:0] ? 4'ha : _GEN_833; // @[Filter.scala 204:142]
  wire [3:0] _GEN_835 = 8'ha0 == _T_40[7:0] ? 4'h0 : _GEN_834; // @[Filter.scala 204:142]
  wire [3:0] _GEN_836 = 8'ha1 == _T_40[7:0] ? 4'h3 : _GEN_835; // @[Filter.scala 204:142]
  wire [3:0] _GEN_837 = 8'ha2 == _T_40[7:0] ? 4'h6 : _GEN_836; // @[Filter.scala 204:142]
  wire [3:0] _GEN_838 = 8'ha3 == _T_40[7:0] ? 4'h6 : _GEN_837; // @[Filter.scala 204:142]
  wire [3:0] _GEN_839 = 8'ha4 == _T_40[7:0] ? 4'h0 : _GEN_838; // @[Filter.scala 204:142]
  wire [3:0] _GEN_840 = 8'ha5 == _T_40[7:0] ? 4'h0 : _GEN_839; // @[Filter.scala 204:142]
  wire [3:0] _GEN_841 = 8'ha6 == _T_40[7:0] ? 4'h0 : _GEN_840; // @[Filter.scala 204:142]
  wire [3:0] _GEN_842 = 8'ha7 == _T_40[7:0] ? 4'h0 : _GEN_841; // @[Filter.scala 204:142]
  wire [3:0] _GEN_843 = 8'ha8 == _T_40[7:0] ? 4'h0 : _GEN_842; // @[Filter.scala 204:142]
  wire [3:0] _GEN_844 = 8'ha9 == _T_40[7:0] ? 4'h0 : _GEN_843; // @[Filter.scala 204:142]
  wire [3:0] _GEN_845 = 8'haa == _T_40[7:0] ? 4'h0 : _GEN_844; // @[Filter.scala 204:142]
  wire [3:0] _GEN_846 = 8'hab == _T_40[7:0] ? 4'h0 : _GEN_845; // @[Filter.scala 204:142]
  wire [3:0] _GEN_847 = 8'hac == _T_40[7:0] ? 4'h6 : _GEN_846; // @[Filter.scala 204:142]
  wire [3:0] _GEN_848 = 8'had == _T_40[7:0] ? 4'h0 : _GEN_847; // @[Filter.scala 204:142]
  wire [3:0] _GEN_849 = 8'hae == _T_40[7:0] ? 4'h3 : _GEN_848; // @[Filter.scala 204:142]
  wire [3:0] _GEN_850 = 8'haf == _T_40[7:0] ? 4'h9 : _GEN_849; // @[Filter.scala 204:142]
  wire [3:0] _GEN_851 = 8'hb0 == _T_40[7:0] ? 4'h3 : _GEN_850; // @[Filter.scala 204:142]
  wire [3:0] _GEN_852 = 8'hb1 == _T_40[7:0] ? 4'h0 : _GEN_851; // @[Filter.scala 204:142]
  wire [3:0] _GEN_853 = 8'hb2 == _T_40[7:0] ? 4'h0 : _GEN_852; // @[Filter.scala 204:142]
  wire [3:0] _GEN_854 = 8'hb3 == _T_40[7:0] ? 4'h0 : _GEN_853; // @[Filter.scala 204:142]
  wire [3:0] _GEN_855 = 8'hb4 == _T_40[7:0] ? 4'h3 : _GEN_854; // @[Filter.scala 204:142]
  wire [3:0] _GEN_856 = 8'hb5 == _T_40[7:0] ? 4'h9 : _GEN_855; // @[Filter.scala 204:142]
  wire [3:0] _GEN_857 = 8'hb6 == _T_40[7:0] ? 4'h3 : _GEN_856; // @[Filter.scala 204:142]
  wire [3:0] _GEN_858 = 8'hb7 == _T_40[7:0] ? 4'h0 : _GEN_857; // @[Filter.scala 204:142]
  wire [3:0] _GEN_859 = 8'hb8 == _T_40[7:0] ? 4'h6 : _GEN_858; // @[Filter.scala 204:142]
  wire [3:0] _GEN_860 = 8'hb9 == _T_40[7:0] ? 4'h0 : _GEN_859; // @[Filter.scala 204:142]
  wire [3:0] _GEN_861 = 8'hba == _T_40[7:0] ? 4'h0 : _GEN_860; // @[Filter.scala 204:142]
  wire [3:0] _GEN_862 = 8'hbb == _T_40[7:0] ? 4'h0 : _GEN_861; // @[Filter.scala 204:142]
  wire [3:0] _GEN_863 = 8'hbc == _T_40[7:0] ? 4'h0 : _GEN_862; // @[Filter.scala 204:142]
  wire [3:0] _GEN_864 = 8'hbd == _T_40[7:0] ? 4'h0 : _GEN_863; // @[Filter.scala 204:142]
  wire [3:0] _GEN_865 = 8'hbe == _T_40[7:0] ? 4'h0 : _GEN_864; // @[Filter.scala 204:142]
  wire [3:0] _GEN_866 = 8'hbf == _T_40[7:0] ? 4'h0 : _GEN_865; // @[Filter.scala 204:142]
  wire [3:0] _GEN_867 = 8'hc0 == _T_40[7:0] ? 4'h0 : _GEN_866; // @[Filter.scala 204:142]
  wire [3:0] _GEN_868 = 8'hc1 == _T_40[7:0] ? 4'h0 : _GEN_867; // @[Filter.scala 204:142]
  wire [3:0] _GEN_869 = 8'hc2 == _T_40[7:0] ? 4'h7 : _GEN_868; // @[Filter.scala 204:142]
  wire [3:0] _GEN_870 = 8'hc3 == _T_40[7:0] ? 4'h2 : _GEN_869; // @[Filter.scala 204:142]
  wire [3:0] _GEN_871 = 8'hc4 == _T_40[7:0] ? 4'h0 : _GEN_870; // @[Filter.scala 204:142]
  wire [3:0] _GEN_872 = 8'hc5 == _T_40[7:0] ? 4'h6 : _GEN_871; // @[Filter.scala 204:142]
  wire [3:0] _GEN_873 = 8'hc6 == _T_40[7:0] ? 4'h9 : _GEN_872; // @[Filter.scala 204:142]
  wire [3:0] _GEN_874 = 8'hc7 == _T_40[7:0] ? 4'h6 : _GEN_873; // @[Filter.scala 204:142]
  wire [3:0] _GEN_875 = 8'hc8 == _T_40[7:0] ? 4'h9 : _GEN_874; // @[Filter.scala 204:142]
  wire [3:0] _GEN_876 = 8'hc9 == _T_40[7:0] ? 4'h6 : _GEN_875; // @[Filter.scala 204:142]
  wire [3:0] _GEN_877 = 8'hca == _T_40[7:0] ? 4'h0 : _GEN_876; // @[Filter.scala 204:142]
  wire [3:0] _GEN_878 = 8'hcb == _T_40[7:0] ? 4'h2 : _GEN_877; // @[Filter.scala 204:142]
  wire [3:0] _GEN_879 = 8'hcc == _T_40[7:0] ? 4'h7 : _GEN_878; // @[Filter.scala 204:142]
  wire [3:0] _GEN_880 = 8'hcd == _T_40[7:0] ? 4'h0 : _GEN_879; // @[Filter.scala 204:142]
  wire [3:0] _GEN_881 = 8'hce == _T_40[7:0] ? 4'h0 : _GEN_880; // @[Filter.scala 204:142]
  wire [3:0] _GEN_882 = 8'hcf == _T_40[7:0] ? 4'h0 : _GEN_881; // @[Filter.scala 204:142]
  wire [3:0] _GEN_883 = 8'hd0 == _T_40[7:0] ? 4'h0 : _GEN_882; // @[Filter.scala 204:142]
  wire [3:0] _GEN_884 = 8'hd1 == _T_40[7:0] ? 4'h0 : _GEN_883; // @[Filter.scala 204:142]
  wire [3:0] _GEN_885 = 8'hd2 == _T_40[7:0] ? 4'h0 : _GEN_884; // @[Filter.scala 204:142]
  wire [3:0] _GEN_886 = 8'hd3 == _T_40[7:0] ? 4'h0 : _GEN_885; // @[Filter.scala 204:142]
  wire [3:0] _GEN_887 = 8'hd4 == _T_40[7:0] ? 4'h0 : _GEN_886; // @[Filter.scala 204:142]
  wire [3:0] _GEN_888 = 8'hd5 == _T_40[7:0] ? 4'h0 : _GEN_887; // @[Filter.scala 204:142]
  wire [3:0] _GEN_889 = 8'hd6 == _T_40[7:0] ? 4'h0 : _GEN_888; // @[Filter.scala 204:142]
  wire [3:0] _GEN_890 = 8'hd7 == _T_40[7:0] ? 4'h3 : _GEN_889; // @[Filter.scala 204:142]
  wire [3:0] _GEN_891 = 8'hd8 == _T_40[7:0] ? 4'h3 : _GEN_890; // @[Filter.scala 204:142]
  wire [3:0] _GEN_892 = 8'hd9 == _T_40[7:0] ? 4'h0 : _GEN_891; // @[Filter.scala 204:142]
  wire [3:0] _GEN_893 = 8'hda == _T_40[7:0] ? 4'h9 : _GEN_892; // @[Filter.scala 204:142]
  wire [3:0] _GEN_894 = 8'hdb == _T_40[7:0] ? 4'h3 : _GEN_893; // @[Filter.scala 204:142]
  wire [3:0] _GEN_895 = 8'hdc == _T_40[7:0] ? 4'hc : _GEN_894; // @[Filter.scala 204:142]
  wire [3:0] _GEN_896 = 8'hdd == _T_40[7:0] ? 4'h3 : _GEN_895; // @[Filter.scala 204:142]
  wire [3:0] _GEN_897 = 8'hde == _T_40[7:0] ? 4'h9 : _GEN_896; // @[Filter.scala 204:142]
  wire [3:0] _GEN_898 = 8'hdf == _T_40[7:0] ? 4'h0 : _GEN_897; // @[Filter.scala 204:142]
  wire [3:0] _GEN_899 = 8'he0 == _T_40[7:0] ? 4'h3 : _GEN_898; // @[Filter.scala 204:142]
  wire [3:0] _GEN_900 = 8'he1 == _T_40[7:0] ? 4'h3 : _GEN_899; // @[Filter.scala 204:142]
  wire [3:0] _GEN_901 = 8'he2 == _T_40[7:0] ? 4'h0 : _GEN_900; // @[Filter.scala 204:142]
  wire [3:0] _GEN_902 = 8'he3 == _T_40[7:0] ? 4'h0 : _GEN_901; // @[Filter.scala 204:142]
  wire [3:0] _GEN_903 = 8'he4 == _T_40[7:0] ? 4'h0 : _GEN_902; // @[Filter.scala 204:142]
  wire [3:0] _GEN_904 = 8'he5 == _T_40[7:0] ? 4'h0 : _GEN_903; // @[Filter.scala 204:142]
  wire [3:0] _GEN_905 = 8'he6 == _T_40[7:0] ? 4'h0 : _GEN_904; // @[Filter.scala 204:142]
  wire [3:0] _GEN_906 = 8'he7 == _T_40[7:0] ? 4'h0 : _GEN_905; // @[Filter.scala 204:142]
  wire [3:0] _GEN_907 = 8'he8 == _T_40[7:0] ? 4'h0 : _GEN_906; // @[Filter.scala 204:142]
  wire [3:0] _GEN_908 = 8'he9 == _T_40[7:0] ? 4'h0 : _GEN_907; // @[Filter.scala 204:142]
  wire [3:0] _GEN_909 = 8'hea == _T_40[7:0] ? 4'h0 : _GEN_908; // @[Filter.scala 204:142]
  wire [3:0] _GEN_910 = 8'heb == _T_40[7:0] ? 4'h0 : _GEN_909; // @[Filter.scala 204:142]
  wire [3:0] _GEN_911 = 8'hec == _T_40[7:0] ? 4'h0 : _GEN_910; // @[Filter.scala 204:142]
  wire [3:0] _GEN_912 = 8'hed == _T_40[7:0] ? 4'h0 : _GEN_911; // @[Filter.scala 204:142]
  wire [3:0] _GEN_913 = 8'hee == _T_40[7:0] ? 4'h0 : _GEN_912; // @[Filter.scala 204:142]
  wire [3:0] _GEN_914 = 8'hef == _T_40[7:0] ? 4'h0 : _GEN_913; // @[Filter.scala 204:142]
  wire [3:0] _GEN_915 = 8'hf0 == _T_40[7:0] ? 4'h0 : _GEN_914; // @[Filter.scala 204:142]
  wire [3:0] _GEN_916 = 8'hf1 == _T_40[7:0] ? 4'h0 : _GEN_915; // @[Filter.scala 204:142]
  wire [3:0] _GEN_917 = 8'hf2 == _T_40[7:0] ? 4'h0 : _GEN_916; // @[Filter.scala 204:142]
  wire [3:0] _GEN_918 = 8'hf3 == _T_40[7:0] ? 4'h0 : _GEN_917; // @[Filter.scala 204:142]
  wire [3:0] _GEN_919 = 8'hf4 == _T_40[7:0] ? 4'h0 : _GEN_918; // @[Filter.scala 204:142]
  wire [3:0] _GEN_920 = 8'hf5 == _T_40[7:0] ? 4'h0 : _GEN_919; // @[Filter.scala 204:142]
  wire [3:0] _GEN_921 = 8'hf6 == _T_40[7:0] ? 4'h0 : _GEN_920; // @[Filter.scala 204:142]
  wire [3:0] _GEN_922 = 8'hf7 == _T_40[7:0] ? 4'h0 : _GEN_921; // @[Filter.scala 204:142]
  wire [3:0] _GEN_923 = 8'hf8 == _T_40[7:0] ? 4'h0 : _GEN_922; // @[Filter.scala 204:142]
  wire [3:0] _GEN_924 = 8'hf9 == _T_40[7:0] ? 4'h0 : _GEN_923; // @[Filter.scala 204:142]
  wire [3:0] _GEN_925 = 8'hfa == _T_40[7:0] ? 4'h0 : _GEN_924; // @[Filter.scala 204:142]
  wire [3:0] _GEN_926 = 8'hfb == _T_40[7:0] ? 4'h0 : _GEN_925; // @[Filter.scala 204:142]
  wire [7:0] _T_54 = _GEN_926 * 4'ha; // @[Filter.scala 204:142]
  wire [10:0] _GEN_11218 = {{3'd0}, _T_54}; // @[Filter.scala 204:109]
  wire [10:0] _T_56 = _T_49 + _GEN_11218; // @[Filter.scala 204:109]
  wire [10:0] _T_57 = _T_56 / 11'h64; // @[Filter.scala 204:150]
  wire  _T_59 = _T_30 >= 5'h15; // @[Filter.scala 207:31]
  wire  _T_63 = _T_37 >= 32'hc; // @[Filter.scala 207:63]
  wire  _T_64 = _T_59 | _T_63; // @[Filter.scala 207:58]
  wire [10:0] _GEN_1179 = io_SPI_distort ? _T_57 : {{7'd0}, _GEN_422}; // @[Filter.scala 209:35]
  wire [10:0] _GEN_1180 = _T_64 ? 11'h0 : _GEN_1179; // @[Filter.scala 207:80]
  wire [10:0] _GEN_1433 = io_SPI_distort ? _T_57 : {{7'd0}, _GEN_674}; // @[Filter.scala 209:35]
  wire [10:0] _GEN_1434 = _T_64 ? 11'h0 : _GEN_1433; // @[Filter.scala 207:80]
  wire [10:0] _GEN_1687 = io_SPI_distort ? _T_57 : {{7'd0}, _GEN_926}; // @[Filter.scala 209:35]
  wire [10:0] _GEN_1688 = _T_64 ? 11'h0 : _GEN_1687; // @[Filter.scala 207:80]
  wire [31:0] _T_92 = pixelIndex + 32'h1; // @[Filter.scala 202:31]
  wire [31:0] _GEN_1 = _T_92 % 32'h15; // @[Filter.scala 202:38]
  wire [4:0] _T_93 = _GEN_1[4:0]; // @[Filter.scala 202:38]
  wire [4:0] _T_95 = _T_93 + _GEN_11210; // @[Filter.scala 202:53]
  wire [4:0] _T_97 = _T_95 - 5'h1; // @[Filter.scala 202:69]
  wire [31:0] _T_100 = _T_92 / 32'h15; // @[Filter.scala 203:38]
  wire [31:0] _T_102 = _T_100 + _GEN_11211; // @[Filter.scala 203:53]
  wire [31:0] _T_104 = _T_102 - 32'h1; // @[Filter.scala 203:69]
  wire [36:0] _T_105 = _T_104 * 32'h15; // @[Filter.scala 204:42]
  wire [36:0] _GEN_11224 = {{32'd0}, _T_97}; // @[Filter.scala 204:57]
  wire [36:0] _T_107 = _T_105 + _GEN_11224; // @[Filter.scala 204:57]
  wire [3:0] _GEN_1697 = 8'h8 == _T_107[7:0] ? 4'h1 : 4'h0; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1698 = 8'h9 == _T_107[7:0] ? 4'h2 : _GEN_1697; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1699 = 8'ha == _T_107[7:0] ? 4'h2 : _GEN_1698; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1700 = 8'hb == _T_107[7:0] ? 4'h2 : _GEN_1699; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1701 = 8'hc == _T_107[7:0] ? 4'h1 : _GEN_1700; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1702 = 8'hd == _T_107[7:0] ? 4'h0 : _GEN_1701; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1703 = 8'he == _T_107[7:0] ? 4'h0 : _GEN_1702; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1704 = 8'hf == _T_107[7:0] ? 4'h0 : _GEN_1703; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1705 = 8'h10 == _T_107[7:0] ? 4'h0 : _GEN_1704; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1706 = 8'h11 == _T_107[7:0] ? 4'h0 : _GEN_1705; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1707 = 8'h12 == _T_107[7:0] ? 4'h0 : _GEN_1706; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1708 = 8'h13 == _T_107[7:0] ? 4'h0 : _GEN_1707; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1709 = 8'h14 == _T_107[7:0] ? 4'h0 : _GEN_1708; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1710 = 8'h15 == _T_107[7:0] ? 4'h0 : _GEN_1709; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1711 = 8'h16 == _T_107[7:0] ? 4'h0 : _GEN_1710; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1712 = 8'h17 == _T_107[7:0] ? 4'h0 : _GEN_1711; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1713 = 8'h18 == _T_107[7:0] ? 4'h0 : _GEN_1712; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1714 = 8'h19 == _T_107[7:0] ? 4'h0 : _GEN_1713; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1715 = 8'h1a == _T_107[7:0] ? 4'h0 : _GEN_1714; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1716 = 8'h1b == _T_107[7:0] ? 4'h0 : _GEN_1715; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1717 = 8'h1c == _T_107[7:0] ? 4'h2 : _GEN_1716; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1718 = 8'h1d == _T_107[7:0] ? 4'h1 : _GEN_1717; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1719 = 8'h1e == _T_107[7:0] ? 4'h0 : _GEN_1718; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1720 = 8'h1f == _T_107[7:0] ? 4'h0 : _GEN_1719; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1721 = 8'h20 == _T_107[7:0] ? 4'h0 : _GEN_1720; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1722 = 8'h21 == _T_107[7:0] ? 4'h1 : _GEN_1721; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1723 = 8'h22 == _T_107[7:0] ? 4'h2 : _GEN_1722; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1724 = 8'h23 == _T_107[7:0] ? 4'h0 : _GEN_1723; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1725 = 8'h24 == _T_107[7:0] ? 4'h0 : _GEN_1724; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1726 = 8'h25 == _T_107[7:0] ? 4'h0 : _GEN_1725; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1727 = 8'h26 == _T_107[7:0] ? 4'h0 : _GEN_1726; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1728 = 8'h27 == _T_107[7:0] ? 4'h0 : _GEN_1727; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1729 = 8'h28 == _T_107[7:0] ? 4'h0 : _GEN_1728; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1730 = 8'h29 == _T_107[7:0] ? 4'h0 : _GEN_1729; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1731 = 8'h2a == _T_107[7:0] ? 4'h0 : _GEN_1730; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1732 = 8'h2b == _T_107[7:0] ? 4'h0 : _GEN_1731; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1733 = 8'h2c == _T_107[7:0] ? 4'h0 : _GEN_1732; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1734 = 8'h2d == _T_107[7:0] ? 4'h0 : _GEN_1733; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1735 = 8'h2e == _T_107[7:0] ? 4'h0 : _GEN_1734; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1736 = 8'h2f == _T_107[7:0] ? 4'h0 : _GEN_1735; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1737 = 8'h30 == _T_107[7:0] ? 4'h2 : _GEN_1736; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1738 = 8'h31 == _T_107[7:0] ? 4'h2 : _GEN_1737; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1739 = 8'h32 == _T_107[7:0] ? 4'h0 : _GEN_1738; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1740 = 8'h33 == _T_107[7:0] ? 4'h0 : _GEN_1739; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1741 = 8'h34 == _T_107[7:0] ? 4'h0 : _GEN_1740; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1742 = 8'h35 == _T_107[7:0] ? 4'h0 : _GEN_1741; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1743 = 8'h36 == _T_107[7:0] ? 4'h0 : _GEN_1742; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1744 = 8'h37 == _T_107[7:0] ? 4'h0 : _GEN_1743; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1745 = 8'h38 == _T_107[7:0] ? 4'h2 : _GEN_1744; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1746 = 8'h39 == _T_107[7:0] ? 4'h0 : _GEN_1745; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1747 = 8'h3a == _T_107[7:0] ? 4'h0 : _GEN_1746; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1748 = 8'h3b == _T_107[7:0] ? 4'h0 : _GEN_1747; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1749 = 8'h3c == _T_107[7:0] ? 4'h0 : _GEN_1748; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1750 = 8'h3d == _T_107[7:0] ? 4'h0 : _GEN_1749; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1751 = 8'h3e == _T_107[7:0] ? 4'h0 : _GEN_1750; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1752 = 8'h3f == _T_107[7:0] ? 4'h0 : _GEN_1751; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1753 = 8'h40 == _T_107[7:0] ? 4'h0 : _GEN_1752; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1754 = 8'h41 == _T_107[7:0] ? 4'h0 : _GEN_1753; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1755 = 8'h42 == _T_107[7:0] ? 4'h0 : _GEN_1754; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1756 = 8'h43 == _T_107[7:0] ? 4'h0 : _GEN_1755; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1757 = 8'h44 == _T_107[7:0] ? 4'h1 : _GEN_1756; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1758 = 8'h45 == _T_107[7:0] ? 4'h3 : _GEN_1757; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1759 = 8'h46 == _T_107[7:0] ? 4'h7 : _GEN_1758; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1760 = 8'h47 == _T_107[7:0] ? 4'h0 : _GEN_1759; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1761 = 8'h48 == _T_107[7:0] ? 4'h0 : _GEN_1760; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1762 = 8'h49 == _T_107[7:0] ? 4'h0 : _GEN_1761; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1763 = 8'h4a == _T_107[7:0] ? 4'h0 : _GEN_1762; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1764 = 8'h4b == _T_107[7:0] ? 4'h0 : _GEN_1763; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1765 = 8'h4c == _T_107[7:0] ? 4'h0 : _GEN_1764; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1766 = 8'h4d == _T_107[7:0] ? 4'h0 : _GEN_1765; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1767 = 8'h4e == _T_107[7:0] ? 4'h2 : _GEN_1766; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1768 = 8'h4f == _T_107[7:0] ? 4'h0 : _GEN_1767; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1769 = 8'h50 == _T_107[7:0] ? 4'h0 : _GEN_1768; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1770 = 8'h51 == _T_107[7:0] ? 4'h0 : _GEN_1769; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1771 = 8'h52 == _T_107[7:0] ? 4'h0 : _GEN_1770; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1772 = 8'h53 == _T_107[7:0] ? 4'h0 : _GEN_1771; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1773 = 8'h54 == _T_107[7:0] ? 4'h0 : _GEN_1772; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1774 = 8'h55 == _T_107[7:0] ? 4'h0 : _GEN_1773; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1775 = 8'h56 == _T_107[7:0] ? 4'h0 : _GEN_1774; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1776 = 8'h57 == _T_107[7:0] ? 4'h0 : _GEN_1775; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1777 = 8'h58 == _T_107[7:0] ? 4'h0 : _GEN_1776; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1778 = 8'h59 == _T_107[7:0] ? 4'h2 : _GEN_1777; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1779 = 8'h5a == _T_107[7:0] ? 4'h2 : _GEN_1778; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1780 = 8'h5b == _T_107[7:0] ? 4'h0 : _GEN_1779; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1781 = 8'h5c == _T_107[7:0] ? 4'h0 : _GEN_1780; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1782 = 8'h5d == _T_107[7:0] ? 4'h0 : _GEN_1781; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1783 = 8'h5e == _T_107[7:0] ? 4'h4 : _GEN_1782; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1784 = 8'h5f == _T_107[7:0] ? 4'h0 : _GEN_1783; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1785 = 8'h60 == _T_107[7:0] ? 4'h0 : _GEN_1784; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1786 = 8'h61 == _T_107[7:0] ? 4'h0 : _GEN_1785; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1787 = 8'h62 == _T_107[7:0] ? 4'h0 : _GEN_1786; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1788 = 8'h63 == _T_107[7:0] ? 4'h2 : _GEN_1787; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1789 = 8'h64 == _T_107[7:0] ? 4'h0 : _GEN_1788; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1790 = 8'h65 == _T_107[7:0] ? 4'h0 : _GEN_1789; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1791 = 8'h66 == _T_107[7:0] ? 4'h0 : _GEN_1790; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1792 = 8'h67 == _T_107[7:0] ? 4'h0 : _GEN_1791; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1793 = 8'h68 == _T_107[7:0] ? 4'h0 : _GEN_1792; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1794 = 8'h69 == _T_107[7:0] ? 4'h0 : _GEN_1793; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1795 = 8'h6a == _T_107[7:0] ? 4'h0 : _GEN_1794; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1796 = 8'h6b == _T_107[7:0] ? 4'h0 : _GEN_1795; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1797 = 8'h6c == _T_107[7:0] ? 4'h0 : _GEN_1796; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1798 = 8'h6d == _T_107[7:0] ? 4'h0 : _GEN_1797; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1799 = 8'h6e == _T_107[7:0] ? 4'h2 : _GEN_1798; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1800 = 8'h6f == _T_107[7:0] ? 4'h0 : _GEN_1799; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1801 = 8'h70 == _T_107[7:0] ? 4'h0 : _GEN_1800; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1802 = 8'h71 == _T_107[7:0] ? 4'h0 : _GEN_1801; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1803 = 8'h72 == _T_107[7:0] ? 4'h2 : _GEN_1802; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1804 = 8'h73 == _T_107[7:0] ? 4'h9 : _GEN_1803; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1805 = 8'h74 == _T_107[7:0] ? 4'h2 : _GEN_1804; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1806 = 8'h75 == _T_107[7:0] ? 4'h0 : _GEN_1805; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1807 = 8'h76 == _T_107[7:0] ? 4'h0 : _GEN_1806; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1808 = 8'h77 == _T_107[7:0] ? 4'h0 : _GEN_1807; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1809 = 8'h78 == _T_107[7:0] ? 4'h1 : _GEN_1808; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1810 = 8'h79 == _T_107[7:0] ? 4'h1 : _GEN_1809; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1811 = 8'h7a == _T_107[7:0] ? 4'h0 : _GEN_1810; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1812 = 8'h7b == _T_107[7:0] ? 4'h0 : _GEN_1811; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1813 = 8'h7c == _T_107[7:0] ? 4'h0 : _GEN_1812; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1814 = 8'h7d == _T_107[7:0] ? 4'h0 : _GEN_1813; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1815 = 8'h7e == _T_107[7:0] ? 4'h0 : _GEN_1814; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1816 = 8'h7f == _T_107[7:0] ? 4'h0 : _GEN_1815; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1817 = 8'h80 == _T_107[7:0] ? 4'h0 : _GEN_1816; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1818 = 8'h81 == _T_107[7:0] ? 4'h0 : _GEN_1817; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1819 = 8'h82 == _T_107[7:0] ? 4'h2 : _GEN_1818; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1820 = 8'h83 == _T_107[7:0] ? 4'h0 : _GEN_1819; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1821 = 8'h84 == _T_107[7:0] ? 4'h0 : _GEN_1820; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1822 = 8'h85 == _T_107[7:0] ? 4'h0 : _GEN_1821; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1823 = 8'h86 == _T_107[7:0] ? 4'h7 : _GEN_1822; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1824 = 8'h87 == _T_107[7:0] ? 4'h2 : _GEN_1823; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1825 = 8'h88 == _T_107[7:0] ? 4'h0 : _GEN_1824; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1826 = 8'h89 == _T_107[7:0] ? 4'h2 : _GEN_1825; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1827 = 8'h8a == _T_107[7:0] ? 4'h7 : _GEN_1826; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1828 = 8'h8b == _T_107[7:0] ? 4'h0 : _GEN_1827; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1829 = 8'h8c == _T_107[7:0] ? 4'h0 : _GEN_1828; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1830 = 8'h8d == _T_107[7:0] ? 4'h0 : _GEN_1829; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1831 = 8'h8e == _T_107[7:0] ? 4'h2 : _GEN_1830; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1832 = 8'h8f == _T_107[7:0] ? 4'h0 : _GEN_1831; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1833 = 8'h90 == _T_107[7:0] ? 4'h0 : _GEN_1832; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1834 = 8'h91 == _T_107[7:0] ? 4'h0 : _GEN_1833; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1835 = 8'h92 == _T_107[7:0] ? 4'h0 : _GEN_1834; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1836 = 8'h93 == _T_107[7:0] ? 4'h0 : _GEN_1835; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1837 = 8'h94 == _T_107[7:0] ? 4'h0 : _GEN_1836; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1838 = 8'h95 == _T_107[7:0] ? 4'h0 : _GEN_1837; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1839 = 8'h96 == _T_107[7:0] ? 4'h0 : _GEN_1838; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1840 = 8'h97 == _T_107[7:0] ? 4'h2 : _GEN_1839; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1841 = 8'h98 == _T_107[7:0] ? 4'h2 : _GEN_1840; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1842 = 8'h99 == _T_107[7:0] ? 4'h1 : _GEN_1841; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1843 = 8'h9a == _T_107[7:0] ? 4'h0 : _GEN_1842; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1844 = 8'h9b == _T_107[7:0] ? 4'h7 : _GEN_1843; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1845 = 8'h9c == _T_107[7:0] ? 4'h7 : _GEN_1844; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1846 = 8'h9d == _T_107[7:0] ? 4'h0 : _GEN_1845; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1847 = 8'h9e == _T_107[7:0] ? 4'h7 : _GEN_1846; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1848 = 8'h9f == _T_107[7:0] ? 4'h7 : _GEN_1847; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1849 = 8'ha0 == _T_107[7:0] ? 4'h0 : _GEN_1848; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1850 = 8'ha1 == _T_107[7:0] ? 4'h1 : _GEN_1849; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1851 = 8'ha2 == _T_107[7:0] ? 4'h2 : _GEN_1850; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1852 = 8'ha3 == _T_107[7:0] ? 4'h2 : _GEN_1851; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1853 = 8'ha4 == _T_107[7:0] ? 4'h0 : _GEN_1852; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1854 = 8'ha5 == _T_107[7:0] ? 4'h0 : _GEN_1853; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1855 = 8'ha6 == _T_107[7:0] ? 4'h0 : _GEN_1854; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1856 = 8'ha7 == _T_107[7:0] ? 4'h0 : _GEN_1855; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1857 = 8'ha8 == _T_107[7:0] ? 4'h0 : _GEN_1856; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1858 = 8'ha9 == _T_107[7:0] ? 4'h0 : _GEN_1857; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1859 = 8'haa == _T_107[7:0] ? 4'h0 : _GEN_1858; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1860 = 8'hab == _T_107[7:0] ? 4'h0 : _GEN_1859; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1861 = 8'hac == _T_107[7:0] ? 4'h2 : _GEN_1860; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1862 = 8'had == _T_107[7:0] ? 4'h0 : _GEN_1861; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1863 = 8'hae == _T_107[7:0] ? 4'h1 : _GEN_1862; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1864 = 8'haf == _T_107[7:0] ? 4'h3 : _GEN_1863; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1865 = 8'hb0 == _T_107[7:0] ? 4'h1 : _GEN_1864; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1866 = 8'hb1 == _T_107[7:0] ? 4'h0 : _GEN_1865; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1867 = 8'hb2 == _T_107[7:0] ? 4'h0 : _GEN_1866; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1868 = 8'hb3 == _T_107[7:0] ? 4'h0 : _GEN_1867; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1869 = 8'hb4 == _T_107[7:0] ? 4'h1 : _GEN_1868; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1870 = 8'hb5 == _T_107[7:0] ? 4'h3 : _GEN_1869; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1871 = 8'hb6 == _T_107[7:0] ? 4'h1 : _GEN_1870; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1872 = 8'hb7 == _T_107[7:0] ? 4'h0 : _GEN_1871; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1873 = 8'hb8 == _T_107[7:0] ? 4'h2 : _GEN_1872; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1874 = 8'hb9 == _T_107[7:0] ? 4'h0 : _GEN_1873; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1875 = 8'hba == _T_107[7:0] ? 4'h0 : _GEN_1874; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1876 = 8'hbb == _T_107[7:0] ? 4'h0 : _GEN_1875; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1877 = 8'hbc == _T_107[7:0] ? 4'h0 : _GEN_1876; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1878 = 8'hbd == _T_107[7:0] ? 4'h0 : _GEN_1877; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1879 = 8'hbe == _T_107[7:0] ? 4'h0 : _GEN_1878; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1880 = 8'hbf == _T_107[7:0] ? 4'h0 : _GEN_1879; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1881 = 8'hc0 == _T_107[7:0] ? 4'h0 : _GEN_1880; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1882 = 8'hc1 == _T_107[7:0] ? 4'h0 : _GEN_1881; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1883 = 8'hc2 == _T_107[7:0] ? 4'h3 : _GEN_1882; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1884 = 8'hc3 == _T_107[7:0] ? 4'h0 : _GEN_1883; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1885 = 8'hc4 == _T_107[7:0] ? 4'h0 : _GEN_1884; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1886 = 8'hc5 == _T_107[7:0] ? 4'h2 : _GEN_1885; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1887 = 8'hc6 == _T_107[7:0] ? 4'h3 : _GEN_1886; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1888 = 8'hc7 == _T_107[7:0] ? 4'h2 : _GEN_1887; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1889 = 8'hc8 == _T_107[7:0] ? 4'h3 : _GEN_1888; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1890 = 8'hc9 == _T_107[7:0] ? 4'h2 : _GEN_1889; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1891 = 8'hca == _T_107[7:0] ? 4'h0 : _GEN_1890; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1892 = 8'hcb == _T_107[7:0] ? 4'h0 : _GEN_1891; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1893 = 8'hcc == _T_107[7:0] ? 4'h3 : _GEN_1892; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1894 = 8'hcd == _T_107[7:0] ? 4'h0 : _GEN_1893; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1895 = 8'hce == _T_107[7:0] ? 4'h0 : _GEN_1894; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1896 = 8'hcf == _T_107[7:0] ? 4'h0 : _GEN_1895; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1897 = 8'hd0 == _T_107[7:0] ? 4'h0 : _GEN_1896; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1898 = 8'hd1 == _T_107[7:0] ? 4'h0 : _GEN_1897; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1899 = 8'hd2 == _T_107[7:0] ? 4'h0 : _GEN_1898; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1900 = 8'hd3 == _T_107[7:0] ? 4'h0 : _GEN_1899; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1901 = 8'hd4 == _T_107[7:0] ? 4'h0 : _GEN_1900; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1902 = 8'hd5 == _T_107[7:0] ? 4'h0 : _GEN_1901; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1903 = 8'hd6 == _T_107[7:0] ? 4'h0 : _GEN_1902; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1904 = 8'hd7 == _T_107[7:0] ? 4'h2 : _GEN_1903; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1905 = 8'hd8 == _T_107[7:0] ? 4'h2 : _GEN_1904; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1906 = 8'hd9 == _T_107[7:0] ? 4'h0 : _GEN_1905; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1907 = 8'hda == _T_107[7:0] ? 4'h7 : _GEN_1906; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1908 = 8'hdb == _T_107[7:0] ? 4'h1 : _GEN_1907; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1909 = 8'hdc == _T_107[7:0] ? 4'h4 : _GEN_1908; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1910 = 8'hdd == _T_107[7:0] ? 4'h1 : _GEN_1909; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1911 = 8'hde == _T_107[7:0] ? 4'h7 : _GEN_1910; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1912 = 8'hdf == _T_107[7:0] ? 4'h0 : _GEN_1911; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1913 = 8'he0 == _T_107[7:0] ? 4'h2 : _GEN_1912; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1914 = 8'he1 == _T_107[7:0] ? 4'h2 : _GEN_1913; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1915 = 8'he2 == _T_107[7:0] ? 4'h0 : _GEN_1914; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1916 = 8'he3 == _T_107[7:0] ? 4'h0 : _GEN_1915; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1917 = 8'he4 == _T_107[7:0] ? 4'h0 : _GEN_1916; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1918 = 8'he5 == _T_107[7:0] ? 4'h0 : _GEN_1917; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1919 = 8'he6 == _T_107[7:0] ? 4'h0 : _GEN_1918; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1920 = 8'he7 == _T_107[7:0] ? 4'h0 : _GEN_1919; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1921 = 8'he8 == _T_107[7:0] ? 4'h0 : _GEN_1920; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1922 = 8'he9 == _T_107[7:0] ? 4'h0 : _GEN_1921; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1923 = 8'hea == _T_107[7:0] ? 4'h0 : _GEN_1922; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1924 = 8'heb == _T_107[7:0] ? 4'h0 : _GEN_1923; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1925 = 8'hec == _T_107[7:0] ? 4'h0 : _GEN_1924; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1926 = 8'hed == _T_107[7:0] ? 4'h0 : _GEN_1925; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1927 = 8'hee == _T_107[7:0] ? 4'h0 : _GEN_1926; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1928 = 8'hef == _T_107[7:0] ? 4'h0 : _GEN_1927; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1929 = 8'hf0 == _T_107[7:0] ? 4'h0 : _GEN_1928; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1930 = 8'hf1 == _T_107[7:0] ? 4'h0 : _GEN_1929; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1931 = 8'hf2 == _T_107[7:0] ? 4'h0 : _GEN_1930; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1932 = 8'hf3 == _T_107[7:0] ? 4'h0 : _GEN_1931; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1933 = 8'hf4 == _T_107[7:0] ? 4'h0 : _GEN_1932; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1934 = 8'hf5 == _T_107[7:0] ? 4'h0 : _GEN_1933; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1935 = 8'hf6 == _T_107[7:0] ? 4'h0 : _GEN_1934; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1936 = 8'hf7 == _T_107[7:0] ? 4'h0 : _GEN_1935; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1937 = 8'hf8 == _T_107[7:0] ? 4'h0 : _GEN_1936; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1938 = 8'hf9 == _T_107[7:0] ? 4'h0 : _GEN_1937; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1939 = 8'hfa == _T_107[7:0] ? 4'h0 : _GEN_1938; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1940 = 8'hfb == _T_107[7:0] ? 4'h0 : _GEN_1939; // @[Filter.scala 204:62]
  wire [4:0] _GEN_11225 = {{1'd0}, _GEN_1940}; // @[Filter.scala 204:62]
  wire [8:0] _T_109 = _GEN_11225 * 5'h14; // @[Filter.scala 204:62]
  wire [3:0] _GEN_1990 = 8'h31 == _T_107[7:0] ? 4'h3 : _GEN_1737; // @[Filter.scala 204:102]
  wire [3:0] _GEN_1991 = 8'h32 == _T_107[7:0] ? 4'h3 : _GEN_1990; // @[Filter.scala 204:102]
  wire [3:0] _GEN_1992 = 8'h33 == _T_107[7:0] ? 4'h6 : _GEN_1991; // @[Filter.scala 204:102]
  wire [3:0] _GEN_1993 = 8'h34 == _T_107[7:0] ? 4'h6 : _GEN_1992; // @[Filter.scala 204:102]
  wire [3:0] _GEN_1994 = 8'h35 == _T_107[7:0] ? 4'h0 : _GEN_1993; // @[Filter.scala 204:102]
  wire [3:0] _GEN_1995 = 8'h36 == _T_107[7:0] ? 4'h0 : _GEN_1994; // @[Filter.scala 204:102]
  wire [3:0] _GEN_1996 = 8'h37 == _T_107[7:0] ? 4'h0 : _GEN_1995; // @[Filter.scala 204:102]
  wire [3:0] _GEN_1997 = 8'h38 == _T_107[7:0] ? 4'h2 : _GEN_1996; // @[Filter.scala 204:102]
  wire [3:0] _GEN_1998 = 8'h39 == _T_107[7:0] ? 4'h0 : _GEN_1997; // @[Filter.scala 204:102]
  wire [3:0] _GEN_1999 = 8'h3a == _T_107[7:0] ? 4'h0 : _GEN_1998; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2000 = 8'h3b == _T_107[7:0] ? 4'h0 : _GEN_1999; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2001 = 8'h3c == _T_107[7:0] ? 4'h0 : _GEN_2000; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2002 = 8'h3d == _T_107[7:0] ? 4'h0 : _GEN_2001; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2003 = 8'h3e == _T_107[7:0] ? 4'h0 : _GEN_2002; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2004 = 8'h3f == _T_107[7:0] ? 4'h0 : _GEN_2003; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2005 = 8'h40 == _T_107[7:0] ? 4'h0 : _GEN_2004; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2006 = 8'h41 == _T_107[7:0] ? 4'h0 : _GEN_2005; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2007 = 8'h42 == _T_107[7:0] ? 4'h0 : _GEN_2006; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2008 = 8'h43 == _T_107[7:0] ? 4'h0 : _GEN_2007; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2009 = 8'h44 == _T_107[7:0] ? 4'h1 : _GEN_2008; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2010 = 8'h45 == _T_107[7:0] ? 4'h4 : _GEN_2009; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2011 = 8'h46 == _T_107[7:0] ? 4'hb : _GEN_2010; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2012 = 8'h47 == _T_107[7:0] ? 4'h0 : _GEN_2011; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2013 = 8'h48 == _T_107[7:0] ? 4'h0 : _GEN_2012; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2014 = 8'h49 == _T_107[7:0] ? 4'h0 : _GEN_2013; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2015 = 8'h4a == _T_107[7:0] ? 4'h6 : _GEN_2014; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2016 = 8'h4b == _T_107[7:0] ? 4'h0 : _GEN_2015; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2017 = 8'h4c == _T_107[7:0] ? 4'h3 : _GEN_2016; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2018 = 8'h4d == _T_107[7:0] ? 4'h3 : _GEN_2017; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2019 = 8'h4e == _T_107[7:0] ? 4'h2 : _GEN_2018; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2020 = 8'h4f == _T_107[7:0] ? 4'h0 : _GEN_2019; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2021 = 8'h50 == _T_107[7:0] ? 4'h0 : _GEN_2020; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2022 = 8'h51 == _T_107[7:0] ? 4'h0 : _GEN_2021; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2023 = 8'h52 == _T_107[7:0] ? 4'h0 : _GEN_2022; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2024 = 8'h53 == _T_107[7:0] ? 4'h0 : _GEN_2023; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2025 = 8'h54 == _T_107[7:0] ? 4'h0 : _GEN_2024; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2026 = 8'h55 == _T_107[7:0] ? 4'h0 : _GEN_2025; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2027 = 8'h56 == _T_107[7:0] ? 4'h0 : _GEN_2026; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2028 = 8'h57 == _T_107[7:0] ? 4'h0 : _GEN_2027; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2029 = 8'h58 == _T_107[7:0] ? 4'h0 : _GEN_2028; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2030 = 8'h59 == _T_107[7:0] ? 4'h2 : _GEN_2029; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2031 = 8'h5a == _T_107[7:0] ? 4'h3 : _GEN_2030; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2032 = 8'h5b == _T_107[7:0] ? 4'h0 : _GEN_2031; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2033 = 8'h5c == _T_107[7:0] ? 4'h0 : _GEN_2032; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2034 = 8'h5d == _T_107[7:0] ? 4'h3 : _GEN_2033; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2035 = 8'h5e == _T_107[7:0] ? 4'hd : _GEN_2034; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2036 = 8'h5f == _T_107[7:0] ? 4'h3 : _GEN_2035; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2037 = 8'h60 == _T_107[7:0] ? 4'h0 : _GEN_2036; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2038 = 8'h61 == _T_107[7:0] ? 4'h6 : _GEN_2037; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2039 = 8'h62 == _T_107[7:0] ? 4'h0 : _GEN_2038; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2040 = 8'h63 == _T_107[7:0] ? 4'h2 : _GEN_2039; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2041 = 8'h64 == _T_107[7:0] ? 4'h0 : _GEN_2040; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2042 = 8'h65 == _T_107[7:0] ? 4'h0 : _GEN_2041; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2043 = 8'h66 == _T_107[7:0] ? 4'h0 : _GEN_2042; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2044 = 8'h67 == _T_107[7:0] ? 4'h0 : _GEN_2043; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2045 = 8'h68 == _T_107[7:0] ? 4'h0 : _GEN_2044; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2046 = 8'h69 == _T_107[7:0] ? 4'h0 : _GEN_2045; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2047 = 8'h6a == _T_107[7:0] ? 4'h0 : _GEN_2046; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2048 = 8'h6b == _T_107[7:0] ? 4'h0 : _GEN_2047; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2049 = 8'h6c == _T_107[7:0] ? 4'h0 : _GEN_2048; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2050 = 8'h6d == _T_107[7:0] ? 4'h0 : _GEN_2049; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2051 = 8'h6e == _T_107[7:0] ? 4'h2 : _GEN_2050; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2052 = 8'h6f == _T_107[7:0] ? 4'h0 : _GEN_2051; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2053 = 8'h70 == _T_107[7:0] ? 4'h0 : _GEN_2052; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2054 = 8'h71 == _T_107[7:0] ? 4'h0 : _GEN_2053; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2055 = 8'h72 == _T_107[7:0] ? 4'h6 : _GEN_2054; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2056 = 8'h73 == _T_107[7:0] ? 4'he : _GEN_2055; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2057 = 8'h74 == _T_107[7:0] ? 4'h6 : _GEN_2056; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2058 = 8'h75 == _T_107[7:0] ? 4'h0 : _GEN_2057; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2059 = 8'h76 == _T_107[7:0] ? 4'h6 : _GEN_2058; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2060 = 8'h77 == _T_107[7:0] ? 4'h3 : _GEN_2059; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2061 = 8'h78 == _T_107[7:0] ? 4'h4 : _GEN_2060; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2062 = 8'h79 == _T_107[7:0] ? 4'h1 : _GEN_2061; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2063 = 8'h7a == _T_107[7:0] ? 4'h0 : _GEN_2062; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2064 = 8'h7b == _T_107[7:0] ? 4'h0 : _GEN_2063; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2065 = 8'h7c == _T_107[7:0] ? 4'h0 : _GEN_2064; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2066 = 8'h7d == _T_107[7:0] ? 4'h0 : _GEN_2065; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2067 = 8'h7e == _T_107[7:0] ? 4'h0 : _GEN_2066; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2068 = 8'h7f == _T_107[7:0] ? 4'h0 : _GEN_2067; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2069 = 8'h80 == _T_107[7:0] ? 4'h0 : _GEN_2068; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2070 = 8'h81 == _T_107[7:0] ? 4'h0 : _GEN_2069; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2071 = 8'h82 == _T_107[7:0] ? 4'h2 : _GEN_2070; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2072 = 8'h83 == _T_107[7:0] ? 4'h3 : _GEN_2071; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2073 = 8'h84 == _T_107[7:0] ? 4'h6 : _GEN_2072; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2074 = 8'h85 == _T_107[7:0] ? 4'h6 : _GEN_2073; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2075 = 8'h86 == _T_107[7:0] ? 4'he : _GEN_2074; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2076 = 8'h87 == _T_107[7:0] ? 4'ha : _GEN_2075; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2077 = 8'h88 == _T_107[7:0] ? 4'h6 : _GEN_2076; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2078 = 8'h89 == _T_107[7:0] ? 4'ha : _GEN_2077; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2079 = 8'h8a == _T_107[7:0] ? 4'he : _GEN_2078; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2080 = 8'h8b == _T_107[7:0] ? 4'h3 : _GEN_2079; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2081 = 8'h8c == _T_107[7:0] ? 4'h3 : _GEN_2080; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2082 = 8'h8d == _T_107[7:0] ? 4'h0 : _GEN_2081; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2083 = 8'h8e == _T_107[7:0] ? 4'h2 : _GEN_2082; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2084 = 8'h8f == _T_107[7:0] ? 4'h0 : _GEN_2083; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2085 = 8'h90 == _T_107[7:0] ? 4'h0 : _GEN_2084; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2086 = 8'h91 == _T_107[7:0] ? 4'h0 : _GEN_2085; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2087 = 8'h92 == _T_107[7:0] ? 4'h0 : _GEN_2086; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2088 = 8'h93 == _T_107[7:0] ? 4'h0 : _GEN_2087; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2089 = 8'h94 == _T_107[7:0] ? 4'h0 : _GEN_2088; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2090 = 8'h95 == _T_107[7:0] ? 4'h0 : _GEN_2089; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2091 = 8'h96 == _T_107[7:0] ? 4'h0 : _GEN_2090; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2092 = 8'h97 == _T_107[7:0] ? 4'h2 : _GEN_2091; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2093 = 8'h98 == _T_107[7:0] ? 4'h2 : _GEN_2092; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2094 = 8'h99 == _T_107[7:0] ? 4'h1 : _GEN_2093; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2095 = 8'h9a == _T_107[7:0] ? 4'h3 : _GEN_2094; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2096 = 8'h9b == _T_107[7:0] ? 4'he : _GEN_2095; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2097 = 8'h9c == _T_107[7:0] ? 4'he : _GEN_2096; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2098 = 8'h9d == _T_107[7:0] ? 4'h0 : _GEN_2097; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2099 = 8'h9e == _T_107[7:0] ? 4'he : _GEN_2098; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2100 = 8'h9f == _T_107[7:0] ? 4'he : _GEN_2099; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2101 = 8'ha0 == _T_107[7:0] ? 4'h3 : _GEN_2100; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2102 = 8'ha1 == _T_107[7:0] ? 4'h1 : _GEN_2101; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2103 = 8'ha2 == _T_107[7:0] ? 4'h2 : _GEN_2102; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2104 = 8'ha3 == _T_107[7:0] ? 4'h2 : _GEN_2103; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2105 = 8'ha4 == _T_107[7:0] ? 4'h0 : _GEN_2104; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2106 = 8'ha5 == _T_107[7:0] ? 4'h0 : _GEN_2105; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2107 = 8'ha6 == _T_107[7:0] ? 4'h0 : _GEN_2106; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2108 = 8'ha7 == _T_107[7:0] ? 4'h0 : _GEN_2107; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2109 = 8'ha8 == _T_107[7:0] ? 4'h0 : _GEN_2108; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2110 = 8'ha9 == _T_107[7:0] ? 4'h0 : _GEN_2109; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2111 = 8'haa == _T_107[7:0] ? 4'h0 : _GEN_2110; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2112 = 8'hab == _T_107[7:0] ? 4'h0 : _GEN_2111; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2113 = 8'hac == _T_107[7:0] ? 4'h2 : _GEN_2112; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2114 = 8'had == _T_107[7:0] ? 4'h3 : _GEN_2113; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2115 = 8'hae == _T_107[7:0] ? 4'h4 : _GEN_2114; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2116 = 8'haf == _T_107[7:0] ? 4'h3 : _GEN_2115; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2117 = 8'hb0 == _T_107[7:0] ? 4'h4 : _GEN_2116; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2118 = 8'hb1 == _T_107[7:0] ? 4'h3 : _GEN_2117; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2119 = 8'hb2 == _T_107[7:0] ? 4'h0 : _GEN_2118; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2120 = 8'hb3 == _T_107[7:0] ? 4'h3 : _GEN_2119; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2121 = 8'hb4 == _T_107[7:0] ? 4'h4 : _GEN_2120; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2122 = 8'hb5 == _T_107[7:0] ? 4'h3 : _GEN_2121; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2123 = 8'hb6 == _T_107[7:0] ? 4'h4 : _GEN_2122; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2124 = 8'hb7 == _T_107[7:0] ? 4'h3 : _GEN_2123; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2125 = 8'hb8 == _T_107[7:0] ? 4'h2 : _GEN_2124; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2126 = 8'hb9 == _T_107[7:0] ? 4'h0 : _GEN_2125; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2127 = 8'hba == _T_107[7:0] ? 4'h0 : _GEN_2126; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2128 = 8'hbb == _T_107[7:0] ? 4'h0 : _GEN_2127; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2129 = 8'hbc == _T_107[7:0] ? 4'h0 : _GEN_2128; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2130 = 8'hbd == _T_107[7:0] ? 4'h0 : _GEN_2129; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2131 = 8'hbe == _T_107[7:0] ? 4'h0 : _GEN_2130; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2132 = 8'hbf == _T_107[7:0] ? 4'h0 : _GEN_2131; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2133 = 8'hc0 == _T_107[7:0] ? 4'h0 : _GEN_2132; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2134 = 8'hc1 == _T_107[7:0] ? 4'h0 : _GEN_2133; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2135 = 8'hc2 == _T_107[7:0] ? 4'h8 : _GEN_2134; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2136 = 8'hc3 == _T_107[7:0] ? 4'hc : _GEN_2135; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2137 = 8'hc4 == _T_107[7:0] ? 4'h0 : _GEN_2136; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2138 = 8'hc5 == _T_107[7:0] ? 4'h2 : _GEN_2137; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2139 = 8'hc6 == _T_107[7:0] ? 4'h3 : _GEN_2138; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2140 = 8'hc7 == _T_107[7:0] ? 4'h2 : _GEN_2139; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2141 = 8'hc8 == _T_107[7:0] ? 4'h3 : _GEN_2140; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2142 = 8'hc9 == _T_107[7:0] ? 4'h2 : _GEN_2141; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2143 = 8'hca == _T_107[7:0] ? 4'h0 : _GEN_2142; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2144 = 8'hcb == _T_107[7:0] ? 4'hc : _GEN_2143; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2145 = 8'hcc == _T_107[7:0] ? 4'h8 : _GEN_2144; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2146 = 8'hcd == _T_107[7:0] ? 4'h0 : _GEN_2145; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2147 = 8'hce == _T_107[7:0] ? 4'h0 : _GEN_2146; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2148 = 8'hcf == _T_107[7:0] ? 4'h0 : _GEN_2147; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2149 = 8'hd0 == _T_107[7:0] ? 4'h0 : _GEN_2148; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2150 = 8'hd1 == _T_107[7:0] ? 4'h0 : _GEN_2149; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2151 = 8'hd2 == _T_107[7:0] ? 4'h0 : _GEN_2150; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2152 = 8'hd3 == _T_107[7:0] ? 4'h0 : _GEN_2151; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2153 = 8'hd4 == _T_107[7:0] ? 4'h0 : _GEN_2152; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2154 = 8'hd5 == _T_107[7:0] ? 4'h0 : _GEN_2153; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2155 = 8'hd6 == _T_107[7:0] ? 4'h0 : _GEN_2154; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2156 = 8'hd7 == _T_107[7:0] ? 4'h3 : _GEN_2155; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2157 = 8'hd8 == _T_107[7:0] ? 4'h6 : _GEN_2156; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2158 = 8'hd9 == _T_107[7:0] ? 4'h0 : _GEN_2157; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2159 = 8'hda == _T_107[7:0] ? 4'hb : _GEN_2158; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2160 = 8'hdb == _T_107[7:0] ? 4'h1 : _GEN_2159; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2161 = 8'hdc == _T_107[7:0] ? 4'h4 : _GEN_2160; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2162 = 8'hdd == _T_107[7:0] ? 4'h1 : _GEN_2161; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2163 = 8'hde == _T_107[7:0] ? 4'hb : _GEN_2162; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2164 = 8'hdf == _T_107[7:0] ? 4'h0 : _GEN_2163; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2165 = 8'he0 == _T_107[7:0] ? 4'h6 : _GEN_2164; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2166 = 8'he1 == _T_107[7:0] ? 4'h3 : _GEN_2165; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2167 = 8'he2 == _T_107[7:0] ? 4'h0 : _GEN_2166; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2168 = 8'he3 == _T_107[7:0] ? 4'h0 : _GEN_2167; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2169 = 8'he4 == _T_107[7:0] ? 4'h0 : _GEN_2168; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2170 = 8'he5 == _T_107[7:0] ? 4'h0 : _GEN_2169; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2171 = 8'he6 == _T_107[7:0] ? 4'h0 : _GEN_2170; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2172 = 8'he7 == _T_107[7:0] ? 4'h0 : _GEN_2171; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2173 = 8'he8 == _T_107[7:0] ? 4'h0 : _GEN_2172; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2174 = 8'he9 == _T_107[7:0] ? 4'h0 : _GEN_2173; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2175 = 8'hea == _T_107[7:0] ? 4'h0 : _GEN_2174; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2176 = 8'heb == _T_107[7:0] ? 4'h0 : _GEN_2175; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2177 = 8'hec == _T_107[7:0] ? 4'h0 : _GEN_2176; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2178 = 8'hed == _T_107[7:0] ? 4'h0 : _GEN_2177; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2179 = 8'hee == _T_107[7:0] ? 4'h0 : _GEN_2178; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2180 = 8'hef == _T_107[7:0] ? 4'h0 : _GEN_2179; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2181 = 8'hf0 == _T_107[7:0] ? 4'h0 : _GEN_2180; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2182 = 8'hf1 == _T_107[7:0] ? 4'h0 : _GEN_2181; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2183 = 8'hf2 == _T_107[7:0] ? 4'h0 : _GEN_2182; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2184 = 8'hf3 == _T_107[7:0] ? 4'h0 : _GEN_2183; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2185 = 8'hf4 == _T_107[7:0] ? 4'h0 : _GEN_2184; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2186 = 8'hf5 == _T_107[7:0] ? 4'h0 : _GEN_2185; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2187 = 8'hf6 == _T_107[7:0] ? 4'h0 : _GEN_2186; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2188 = 8'hf7 == _T_107[7:0] ? 4'h0 : _GEN_2187; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2189 = 8'hf8 == _T_107[7:0] ? 4'h0 : _GEN_2188; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2190 = 8'hf9 == _T_107[7:0] ? 4'h0 : _GEN_2189; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2191 = 8'hfa == _T_107[7:0] ? 4'h0 : _GEN_2190; // @[Filter.scala 204:102]
  wire [3:0] _GEN_2192 = 8'hfb == _T_107[7:0] ? 4'h0 : _GEN_2191; // @[Filter.scala 204:102]
  wire [6:0] _GEN_11227 = {{3'd0}, _GEN_2192}; // @[Filter.scala 204:102]
  wire [10:0] _T_114 = _GEN_11227 * 7'h46; // @[Filter.scala 204:102]
  wire [10:0] _GEN_11228 = {{2'd0}, _T_109}; // @[Filter.scala 204:69]
  wire [10:0] _T_116 = _GEN_11228 + _T_114; // @[Filter.scala 204:69]
  wire [3:0] _GEN_2201 = 8'h8 == _T_107[7:0] ? 4'h3 : 4'h0; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2202 = 8'h9 == _T_107[7:0] ? 4'h6 : _GEN_2201; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2203 = 8'ha == _T_107[7:0] ? 4'h6 : _GEN_2202; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2204 = 8'hb == _T_107[7:0] ? 4'h6 : _GEN_2203; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2205 = 8'hc == _T_107[7:0] ? 4'h3 : _GEN_2204; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2206 = 8'hd == _T_107[7:0] ? 4'h0 : _GEN_2205; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2207 = 8'he == _T_107[7:0] ? 4'h0 : _GEN_2206; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2208 = 8'hf == _T_107[7:0] ? 4'h0 : _GEN_2207; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2209 = 8'h10 == _T_107[7:0] ? 4'h0 : _GEN_2208; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2210 = 8'h11 == _T_107[7:0] ? 4'h0 : _GEN_2209; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2211 = 8'h12 == _T_107[7:0] ? 4'h0 : _GEN_2210; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2212 = 8'h13 == _T_107[7:0] ? 4'h0 : _GEN_2211; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2213 = 8'h14 == _T_107[7:0] ? 4'h0 : _GEN_2212; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2214 = 8'h15 == _T_107[7:0] ? 4'h0 : _GEN_2213; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2215 = 8'h16 == _T_107[7:0] ? 4'h0 : _GEN_2214; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2216 = 8'h17 == _T_107[7:0] ? 4'h0 : _GEN_2215; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2217 = 8'h18 == _T_107[7:0] ? 4'h0 : _GEN_2216; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2218 = 8'h19 == _T_107[7:0] ? 4'h0 : _GEN_2217; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2219 = 8'h1a == _T_107[7:0] ? 4'h0 : _GEN_2218; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2220 = 8'h1b == _T_107[7:0] ? 4'h0 : _GEN_2219; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2221 = 8'h1c == _T_107[7:0] ? 4'h6 : _GEN_2220; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2222 = 8'h1d == _T_107[7:0] ? 4'h3 : _GEN_2221; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2223 = 8'h1e == _T_107[7:0] ? 4'h0 : _GEN_2222; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2224 = 8'h1f == _T_107[7:0] ? 4'h0 : _GEN_2223; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2225 = 8'h20 == _T_107[7:0] ? 4'h0 : _GEN_2224; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2226 = 8'h21 == _T_107[7:0] ? 4'h3 : _GEN_2225; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2227 = 8'h22 == _T_107[7:0] ? 4'h6 : _GEN_2226; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2228 = 8'h23 == _T_107[7:0] ? 4'h0 : _GEN_2227; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2229 = 8'h24 == _T_107[7:0] ? 4'h0 : _GEN_2228; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2230 = 8'h25 == _T_107[7:0] ? 4'h0 : _GEN_2229; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2231 = 8'h26 == _T_107[7:0] ? 4'h0 : _GEN_2230; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2232 = 8'h27 == _T_107[7:0] ? 4'h0 : _GEN_2231; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2233 = 8'h28 == _T_107[7:0] ? 4'h0 : _GEN_2232; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2234 = 8'h29 == _T_107[7:0] ? 4'h0 : _GEN_2233; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2235 = 8'h2a == _T_107[7:0] ? 4'h0 : _GEN_2234; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2236 = 8'h2b == _T_107[7:0] ? 4'h0 : _GEN_2235; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2237 = 8'h2c == _T_107[7:0] ? 4'h0 : _GEN_2236; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2238 = 8'h2d == _T_107[7:0] ? 4'h0 : _GEN_2237; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2239 = 8'h2e == _T_107[7:0] ? 4'h0 : _GEN_2238; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2240 = 8'h2f == _T_107[7:0] ? 4'h0 : _GEN_2239; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2241 = 8'h30 == _T_107[7:0] ? 4'h6 : _GEN_2240; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2242 = 8'h31 == _T_107[7:0] ? 4'h3 : _GEN_2241; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2243 = 8'h32 == _T_107[7:0] ? 4'h0 : _GEN_2242; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2244 = 8'h33 == _T_107[7:0] ? 4'h1 : _GEN_2243; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2245 = 8'h34 == _T_107[7:0] ? 4'h1 : _GEN_2244; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2246 = 8'h35 == _T_107[7:0] ? 4'h0 : _GEN_2245; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2247 = 8'h36 == _T_107[7:0] ? 4'h0 : _GEN_2246; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2248 = 8'h37 == _T_107[7:0] ? 4'h0 : _GEN_2247; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2249 = 8'h38 == _T_107[7:0] ? 4'h6 : _GEN_2248; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2250 = 8'h39 == _T_107[7:0] ? 4'h0 : _GEN_2249; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2251 = 8'h3a == _T_107[7:0] ? 4'h0 : _GEN_2250; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2252 = 8'h3b == _T_107[7:0] ? 4'h0 : _GEN_2251; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2253 = 8'h3c == _T_107[7:0] ? 4'h0 : _GEN_2252; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2254 = 8'h3d == _T_107[7:0] ? 4'h0 : _GEN_2253; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2255 = 8'h3e == _T_107[7:0] ? 4'h0 : _GEN_2254; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2256 = 8'h3f == _T_107[7:0] ? 4'h0 : _GEN_2255; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2257 = 8'h40 == _T_107[7:0] ? 4'h0 : _GEN_2256; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2258 = 8'h41 == _T_107[7:0] ? 4'h0 : _GEN_2257; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2259 = 8'h42 == _T_107[7:0] ? 4'h0 : _GEN_2258; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2260 = 8'h43 == _T_107[7:0] ? 4'h0 : _GEN_2259; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2261 = 8'h44 == _T_107[7:0] ? 4'h3 : _GEN_2260; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2262 = 8'h45 == _T_107[7:0] ? 4'h6 : _GEN_2261; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2263 = 8'h46 == _T_107[7:0] ? 4'h9 : _GEN_2262; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2264 = 8'h47 == _T_107[7:0] ? 4'h0 : _GEN_2263; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2265 = 8'h48 == _T_107[7:0] ? 4'h0 : _GEN_2264; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2266 = 8'h49 == _T_107[7:0] ? 4'h0 : _GEN_2265; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2267 = 8'h4a == _T_107[7:0] ? 4'h1 : _GEN_2266; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2268 = 8'h4b == _T_107[7:0] ? 4'h0 : _GEN_2267; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2269 = 8'h4c == _T_107[7:0] ? 4'h0 : _GEN_2268; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2270 = 8'h4d == _T_107[7:0] ? 4'h0 : _GEN_2269; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2271 = 8'h4e == _T_107[7:0] ? 4'h6 : _GEN_2270; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2272 = 8'h4f == _T_107[7:0] ? 4'h0 : _GEN_2271; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2273 = 8'h50 == _T_107[7:0] ? 4'h0 : _GEN_2272; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2274 = 8'h51 == _T_107[7:0] ? 4'h0 : _GEN_2273; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2275 = 8'h52 == _T_107[7:0] ? 4'h0 : _GEN_2274; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2276 = 8'h53 == _T_107[7:0] ? 4'h0 : _GEN_2275; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2277 = 8'h54 == _T_107[7:0] ? 4'h0 : _GEN_2276; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2278 = 8'h55 == _T_107[7:0] ? 4'h0 : _GEN_2277; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2279 = 8'h56 == _T_107[7:0] ? 4'h0 : _GEN_2278; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2280 = 8'h57 == _T_107[7:0] ? 4'h0 : _GEN_2279; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2281 = 8'h58 == _T_107[7:0] ? 4'h0 : _GEN_2280; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2282 = 8'h59 == _T_107[7:0] ? 4'h6 : _GEN_2281; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2283 = 8'h5a == _T_107[7:0] ? 4'h3 : _GEN_2282; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2284 = 8'h5b == _T_107[7:0] ? 4'h0 : _GEN_2283; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2285 = 8'h5c == _T_107[7:0] ? 4'h0 : _GEN_2284; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2286 = 8'h5d == _T_107[7:0] ? 4'h0 : _GEN_2285; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2287 = 8'h5e == _T_107[7:0] ? 4'h7 : _GEN_2286; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2288 = 8'h5f == _T_107[7:0] ? 4'h0 : _GEN_2287; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2289 = 8'h60 == _T_107[7:0] ? 4'h0 : _GEN_2288; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2290 = 8'h61 == _T_107[7:0] ? 4'h1 : _GEN_2289; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2291 = 8'h62 == _T_107[7:0] ? 4'h0 : _GEN_2290; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2292 = 8'h63 == _T_107[7:0] ? 4'h6 : _GEN_2291; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2293 = 8'h64 == _T_107[7:0] ? 4'h0 : _GEN_2292; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2294 = 8'h65 == _T_107[7:0] ? 4'h0 : _GEN_2293; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2295 = 8'h66 == _T_107[7:0] ? 4'h0 : _GEN_2294; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2296 = 8'h67 == _T_107[7:0] ? 4'h0 : _GEN_2295; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2297 = 8'h68 == _T_107[7:0] ? 4'h0 : _GEN_2296; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2298 = 8'h69 == _T_107[7:0] ? 4'h0 : _GEN_2297; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2299 = 8'h6a == _T_107[7:0] ? 4'h0 : _GEN_2298; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2300 = 8'h6b == _T_107[7:0] ? 4'h0 : _GEN_2299; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2301 = 8'h6c == _T_107[7:0] ? 4'h0 : _GEN_2300; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2302 = 8'h6d == _T_107[7:0] ? 4'h0 : _GEN_2301; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2303 = 8'h6e == _T_107[7:0] ? 4'h6 : _GEN_2302; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2304 = 8'h6f == _T_107[7:0] ? 4'h0 : _GEN_2303; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2305 = 8'h70 == _T_107[7:0] ? 4'h0 : _GEN_2304; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2306 = 8'h71 == _T_107[7:0] ? 4'h0 : _GEN_2305; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2307 = 8'h72 == _T_107[7:0] ? 4'h3 : _GEN_2306; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2308 = 8'h73 == _T_107[7:0] ? 4'hc : _GEN_2307; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2309 = 8'h74 == _T_107[7:0] ? 4'h3 : _GEN_2308; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2310 = 8'h75 == _T_107[7:0] ? 4'h0 : _GEN_2309; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2311 = 8'h76 == _T_107[7:0] ? 4'h1 : _GEN_2310; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2312 = 8'h77 == _T_107[7:0] ? 4'h0 : _GEN_2311; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2313 = 8'h78 == _T_107[7:0] ? 4'h3 : _GEN_2312; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2314 = 8'h79 == _T_107[7:0] ? 4'h3 : _GEN_2313; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2315 = 8'h7a == _T_107[7:0] ? 4'h0 : _GEN_2314; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2316 = 8'h7b == _T_107[7:0] ? 4'h0 : _GEN_2315; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2317 = 8'h7c == _T_107[7:0] ? 4'h0 : _GEN_2316; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2318 = 8'h7d == _T_107[7:0] ? 4'h0 : _GEN_2317; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2319 = 8'h7e == _T_107[7:0] ? 4'h0 : _GEN_2318; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2320 = 8'h7f == _T_107[7:0] ? 4'h0 : _GEN_2319; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2321 = 8'h80 == _T_107[7:0] ? 4'h0 : _GEN_2320; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2322 = 8'h81 == _T_107[7:0] ? 4'h0 : _GEN_2321; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2323 = 8'h82 == _T_107[7:0] ? 4'h6 : _GEN_2322; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2324 = 8'h83 == _T_107[7:0] ? 4'h0 : _GEN_2323; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2325 = 8'h84 == _T_107[7:0] ? 4'h1 : _GEN_2324; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2326 = 8'h85 == _T_107[7:0] ? 4'h1 : _GEN_2325; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2327 = 8'h86 == _T_107[7:0] ? 4'ha : _GEN_2326; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2328 = 8'h87 == _T_107[7:0] ? 4'h4 : _GEN_2327; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2329 = 8'h88 == _T_107[7:0] ? 4'h1 : _GEN_2328; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2330 = 8'h89 == _T_107[7:0] ? 4'h4 : _GEN_2329; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2331 = 8'h8a == _T_107[7:0] ? 4'ha : _GEN_2330; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2332 = 8'h8b == _T_107[7:0] ? 4'h0 : _GEN_2331; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2333 = 8'h8c == _T_107[7:0] ? 4'h0 : _GEN_2332; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2334 = 8'h8d == _T_107[7:0] ? 4'h0 : _GEN_2333; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2335 = 8'h8e == _T_107[7:0] ? 4'h6 : _GEN_2334; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2336 = 8'h8f == _T_107[7:0] ? 4'h0 : _GEN_2335; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2337 = 8'h90 == _T_107[7:0] ? 4'h0 : _GEN_2336; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2338 = 8'h91 == _T_107[7:0] ? 4'h0 : _GEN_2337; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2339 = 8'h92 == _T_107[7:0] ? 4'h0 : _GEN_2338; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2340 = 8'h93 == _T_107[7:0] ? 4'h0 : _GEN_2339; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2341 = 8'h94 == _T_107[7:0] ? 4'h0 : _GEN_2340; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2342 = 8'h95 == _T_107[7:0] ? 4'h0 : _GEN_2341; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2343 = 8'h96 == _T_107[7:0] ? 4'h0 : _GEN_2342; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2344 = 8'h97 == _T_107[7:0] ? 4'h6 : _GEN_2343; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2345 = 8'h98 == _T_107[7:0] ? 4'h6 : _GEN_2344; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2346 = 8'h99 == _T_107[7:0] ? 4'h3 : _GEN_2345; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2347 = 8'h9a == _T_107[7:0] ? 4'h0 : _GEN_2346; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2348 = 8'h9b == _T_107[7:0] ? 4'ha : _GEN_2347; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2349 = 8'h9c == _T_107[7:0] ? 4'ha : _GEN_2348; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2350 = 8'h9d == _T_107[7:0] ? 4'h0 : _GEN_2349; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2351 = 8'h9e == _T_107[7:0] ? 4'ha : _GEN_2350; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2352 = 8'h9f == _T_107[7:0] ? 4'ha : _GEN_2351; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2353 = 8'ha0 == _T_107[7:0] ? 4'h0 : _GEN_2352; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2354 = 8'ha1 == _T_107[7:0] ? 4'h3 : _GEN_2353; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2355 = 8'ha2 == _T_107[7:0] ? 4'h6 : _GEN_2354; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2356 = 8'ha3 == _T_107[7:0] ? 4'h6 : _GEN_2355; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2357 = 8'ha4 == _T_107[7:0] ? 4'h0 : _GEN_2356; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2358 = 8'ha5 == _T_107[7:0] ? 4'h0 : _GEN_2357; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2359 = 8'ha6 == _T_107[7:0] ? 4'h0 : _GEN_2358; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2360 = 8'ha7 == _T_107[7:0] ? 4'h0 : _GEN_2359; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2361 = 8'ha8 == _T_107[7:0] ? 4'h0 : _GEN_2360; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2362 = 8'ha9 == _T_107[7:0] ? 4'h0 : _GEN_2361; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2363 = 8'haa == _T_107[7:0] ? 4'h0 : _GEN_2362; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2364 = 8'hab == _T_107[7:0] ? 4'h0 : _GEN_2363; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2365 = 8'hac == _T_107[7:0] ? 4'h6 : _GEN_2364; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2366 = 8'had == _T_107[7:0] ? 4'h0 : _GEN_2365; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2367 = 8'hae == _T_107[7:0] ? 4'h3 : _GEN_2366; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2368 = 8'haf == _T_107[7:0] ? 4'h9 : _GEN_2367; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2369 = 8'hb0 == _T_107[7:0] ? 4'h3 : _GEN_2368; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2370 = 8'hb1 == _T_107[7:0] ? 4'h0 : _GEN_2369; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2371 = 8'hb2 == _T_107[7:0] ? 4'h0 : _GEN_2370; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2372 = 8'hb3 == _T_107[7:0] ? 4'h0 : _GEN_2371; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2373 = 8'hb4 == _T_107[7:0] ? 4'h3 : _GEN_2372; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2374 = 8'hb5 == _T_107[7:0] ? 4'h9 : _GEN_2373; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2375 = 8'hb6 == _T_107[7:0] ? 4'h3 : _GEN_2374; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2376 = 8'hb7 == _T_107[7:0] ? 4'h0 : _GEN_2375; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2377 = 8'hb8 == _T_107[7:0] ? 4'h6 : _GEN_2376; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2378 = 8'hb9 == _T_107[7:0] ? 4'h0 : _GEN_2377; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2379 = 8'hba == _T_107[7:0] ? 4'h0 : _GEN_2378; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2380 = 8'hbb == _T_107[7:0] ? 4'h0 : _GEN_2379; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2381 = 8'hbc == _T_107[7:0] ? 4'h0 : _GEN_2380; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2382 = 8'hbd == _T_107[7:0] ? 4'h0 : _GEN_2381; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2383 = 8'hbe == _T_107[7:0] ? 4'h0 : _GEN_2382; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2384 = 8'hbf == _T_107[7:0] ? 4'h0 : _GEN_2383; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2385 = 8'hc0 == _T_107[7:0] ? 4'h0 : _GEN_2384; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2386 = 8'hc1 == _T_107[7:0] ? 4'h0 : _GEN_2385; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2387 = 8'hc2 == _T_107[7:0] ? 4'h7 : _GEN_2386; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2388 = 8'hc3 == _T_107[7:0] ? 4'h2 : _GEN_2387; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2389 = 8'hc4 == _T_107[7:0] ? 4'h0 : _GEN_2388; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2390 = 8'hc5 == _T_107[7:0] ? 4'h6 : _GEN_2389; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2391 = 8'hc6 == _T_107[7:0] ? 4'h9 : _GEN_2390; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2392 = 8'hc7 == _T_107[7:0] ? 4'h6 : _GEN_2391; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2393 = 8'hc8 == _T_107[7:0] ? 4'h9 : _GEN_2392; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2394 = 8'hc9 == _T_107[7:0] ? 4'h6 : _GEN_2393; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2395 = 8'hca == _T_107[7:0] ? 4'h0 : _GEN_2394; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2396 = 8'hcb == _T_107[7:0] ? 4'h2 : _GEN_2395; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2397 = 8'hcc == _T_107[7:0] ? 4'h7 : _GEN_2396; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2398 = 8'hcd == _T_107[7:0] ? 4'h0 : _GEN_2397; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2399 = 8'hce == _T_107[7:0] ? 4'h0 : _GEN_2398; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2400 = 8'hcf == _T_107[7:0] ? 4'h0 : _GEN_2399; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2401 = 8'hd0 == _T_107[7:0] ? 4'h0 : _GEN_2400; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2402 = 8'hd1 == _T_107[7:0] ? 4'h0 : _GEN_2401; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2403 = 8'hd2 == _T_107[7:0] ? 4'h0 : _GEN_2402; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2404 = 8'hd3 == _T_107[7:0] ? 4'h0 : _GEN_2403; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2405 = 8'hd4 == _T_107[7:0] ? 4'h0 : _GEN_2404; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2406 = 8'hd5 == _T_107[7:0] ? 4'h0 : _GEN_2405; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2407 = 8'hd6 == _T_107[7:0] ? 4'h0 : _GEN_2406; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2408 = 8'hd7 == _T_107[7:0] ? 4'h3 : _GEN_2407; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2409 = 8'hd8 == _T_107[7:0] ? 4'h3 : _GEN_2408; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2410 = 8'hd9 == _T_107[7:0] ? 4'h0 : _GEN_2409; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2411 = 8'hda == _T_107[7:0] ? 4'h9 : _GEN_2410; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2412 = 8'hdb == _T_107[7:0] ? 4'h3 : _GEN_2411; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2413 = 8'hdc == _T_107[7:0] ? 4'hc : _GEN_2412; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2414 = 8'hdd == _T_107[7:0] ? 4'h3 : _GEN_2413; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2415 = 8'hde == _T_107[7:0] ? 4'h9 : _GEN_2414; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2416 = 8'hdf == _T_107[7:0] ? 4'h0 : _GEN_2415; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2417 = 8'he0 == _T_107[7:0] ? 4'h3 : _GEN_2416; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2418 = 8'he1 == _T_107[7:0] ? 4'h3 : _GEN_2417; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2419 = 8'he2 == _T_107[7:0] ? 4'h0 : _GEN_2418; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2420 = 8'he3 == _T_107[7:0] ? 4'h0 : _GEN_2419; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2421 = 8'he4 == _T_107[7:0] ? 4'h0 : _GEN_2420; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2422 = 8'he5 == _T_107[7:0] ? 4'h0 : _GEN_2421; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2423 = 8'he6 == _T_107[7:0] ? 4'h0 : _GEN_2422; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2424 = 8'he7 == _T_107[7:0] ? 4'h0 : _GEN_2423; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2425 = 8'he8 == _T_107[7:0] ? 4'h0 : _GEN_2424; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2426 = 8'he9 == _T_107[7:0] ? 4'h0 : _GEN_2425; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2427 = 8'hea == _T_107[7:0] ? 4'h0 : _GEN_2426; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2428 = 8'heb == _T_107[7:0] ? 4'h0 : _GEN_2427; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2429 = 8'hec == _T_107[7:0] ? 4'h0 : _GEN_2428; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2430 = 8'hed == _T_107[7:0] ? 4'h0 : _GEN_2429; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2431 = 8'hee == _T_107[7:0] ? 4'h0 : _GEN_2430; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2432 = 8'hef == _T_107[7:0] ? 4'h0 : _GEN_2431; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2433 = 8'hf0 == _T_107[7:0] ? 4'h0 : _GEN_2432; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2434 = 8'hf1 == _T_107[7:0] ? 4'h0 : _GEN_2433; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2435 = 8'hf2 == _T_107[7:0] ? 4'h0 : _GEN_2434; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2436 = 8'hf3 == _T_107[7:0] ? 4'h0 : _GEN_2435; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2437 = 8'hf4 == _T_107[7:0] ? 4'h0 : _GEN_2436; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2438 = 8'hf5 == _T_107[7:0] ? 4'h0 : _GEN_2437; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2439 = 8'hf6 == _T_107[7:0] ? 4'h0 : _GEN_2438; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2440 = 8'hf7 == _T_107[7:0] ? 4'h0 : _GEN_2439; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2441 = 8'hf8 == _T_107[7:0] ? 4'h0 : _GEN_2440; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2442 = 8'hf9 == _T_107[7:0] ? 4'h0 : _GEN_2441; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2443 = 8'hfa == _T_107[7:0] ? 4'h0 : _GEN_2442; // @[Filter.scala 204:142]
  wire [3:0] _GEN_2444 = 8'hfb == _T_107[7:0] ? 4'h0 : _GEN_2443; // @[Filter.scala 204:142]
  wire [7:0] _T_121 = _GEN_2444 * 4'ha; // @[Filter.scala 204:142]
  wire [10:0] _GEN_11230 = {{3'd0}, _T_121}; // @[Filter.scala 204:109]
  wire [10:0] _T_123 = _T_116 + _GEN_11230; // @[Filter.scala 204:109]
  wire [10:0] _T_124 = _T_123 / 11'h64; // @[Filter.scala 204:150]
  wire  _T_126 = _T_97 >= 5'h15; // @[Filter.scala 207:31]
  wire  _T_130 = _T_104 >= 32'hc; // @[Filter.scala 207:63]
  wire  _T_131 = _T_126 | _T_130; // @[Filter.scala 207:58]
  wire [10:0] _GEN_2697 = io_SPI_distort ? _T_124 : {{7'd0}, _GEN_1940}; // @[Filter.scala 209:35]
  wire [10:0] _GEN_2698 = _T_131 ? 11'h0 : _GEN_2697; // @[Filter.scala 207:80]
  wire [10:0] _GEN_2951 = io_SPI_distort ? _T_124 : {{7'd0}, _GEN_2192}; // @[Filter.scala 209:35]
  wire [10:0] _GEN_2952 = _T_131 ? 11'h0 : _GEN_2951; // @[Filter.scala 207:80]
  wire [10:0] _GEN_3205 = io_SPI_distort ? _T_124 : {{7'd0}, _GEN_2444}; // @[Filter.scala 209:35]
  wire [10:0] _GEN_3206 = _T_131 ? 11'h0 : _GEN_3205; // @[Filter.scala 207:80]
  wire [31:0] _T_159 = pixelIndex + 32'h2; // @[Filter.scala 202:31]
  wire [31:0] _GEN_2 = _T_159 % 32'h15; // @[Filter.scala 202:38]
  wire [4:0] _T_160 = _GEN_2[4:0]; // @[Filter.scala 202:38]
  wire [4:0] _T_162 = _T_160 + _GEN_11210; // @[Filter.scala 202:53]
  wire [4:0] _T_164 = _T_162 - 5'h1; // @[Filter.scala 202:69]
  wire [31:0] _T_167 = _T_159 / 32'h15; // @[Filter.scala 203:38]
  wire [31:0] _T_169 = _T_167 + _GEN_11211; // @[Filter.scala 203:53]
  wire [31:0] _T_171 = _T_169 - 32'h1; // @[Filter.scala 203:69]
  wire [36:0] _T_172 = _T_171 * 32'h15; // @[Filter.scala 204:42]
  wire [36:0] _GEN_11236 = {{32'd0}, _T_164}; // @[Filter.scala 204:57]
  wire [36:0] _T_174 = _T_172 + _GEN_11236; // @[Filter.scala 204:57]
  wire [3:0] _GEN_3215 = 8'h8 == _T_174[7:0] ? 4'h1 : 4'h0; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3216 = 8'h9 == _T_174[7:0] ? 4'h2 : _GEN_3215; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3217 = 8'ha == _T_174[7:0] ? 4'h2 : _GEN_3216; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3218 = 8'hb == _T_174[7:0] ? 4'h2 : _GEN_3217; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3219 = 8'hc == _T_174[7:0] ? 4'h1 : _GEN_3218; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3220 = 8'hd == _T_174[7:0] ? 4'h0 : _GEN_3219; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3221 = 8'he == _T_174[7:0] ? 4'h0 : _GEN_3220; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3222 = 8'hf == _T_174[7:0] ? 4'h0 : _GEN_3221; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3223 = 8'h10 == _T_174[7:0] ? 4'h0 : _GEN_3222; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3224 = 8'h11 == _T_174[7:0] ? 4'h0 : _GEN_3223; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3225 = 8'h12 == _T_174[7:0] ? 4'h0 : _GEN_3224; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3226 = 8'h13 == _T_174[7:0] ? 4'h0 : _GEN_3225; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3227 = 8'h14 == _T_174[7:0] ? 4'h0 : _GEN_3226; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3228 = 8'h15 == _T_174[7:0] ? 4'h0 : _GEN_3227; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3229 = 8'h16 == _T_174[7:0] ? 4'h0 : _GEN_3228; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3230 = 8'h17 == _T_174[7:0] ? 4'h0 : _GEN_3229; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3231 = 8'h18 == _T_174[7:0] ? 4'h0 : _GEN_3230; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3232 = 8'h19 == _T_174[7:0] ? 4'h0 : _GEN_3231; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3233 = 8'h1a == _T_174[7:0] ? 4'h0 : _GEN_3232; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3234 = 8'h1b == _T_174[7:0] ? 4'h0 : _GEN_3233; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3235 = 8'h1c == _T_174[7:0] ? 4'h2 : _GEN_3234; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3236 = 8'h1d == _T_174[7:0] ? 4'h1 : _GEN_3235; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3237 = 8'h1e == _T_174[7:0] ? 4'h0 : _GEN_3236; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3238 = 8'h1f == _T_174[7:0] ? 4'h0 : _GEN_3237; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3239 = 8'h20 == _T_174[7:0] ? 4'h0 : _GEN_3238; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3240 = 8'h21 == _T_174[7:0] ? 4'h1 : _GEN_3239; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3241 = 8'h22 == _T_174[7:0] ? 4'h2 : _GEN_3240; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3242 = 8'h23 == _T_174[7:0] ? 4'h0 : _GEN_3241; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3243 = 8'h24 == _T_174[7:0] ? 4'h0 : _GEN_3242; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3244 = 8'h25 == _T_174[7:0] ? 4'h0 : _GEN_3243; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3245 = 8'h26 == _T_174[7:0] ? 4'h0 : _GEN_3244; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3246 = 8'h27 == _T_174[7:0] ? 4'h0 : _GEN_3245; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3247 = 8'h28 == _T_174[7:0] ? 4'h0 : _GEN_3246; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3248 = 8'h29 == _T_174[7:0] ? 4'h0 : _GEN_3247; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3249 = 8'h2a == _T_174[7:0] ? 4'h0 : _GEN_3248; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3250 = 8'h2b == _T_174[7:0] ? 4'h0 : _GEN_3249; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3251 = 8'h2c == _T_174[7:0] ? 4'h0 : _GEN_3250; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3252 = 8'h2d == _T_174[7:0] ? 4'h0 : _GEN_3251; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3253 = 8'h2e == _T_174[7:0] ? 4'h0 : _GEN_3252; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3254 = 8'h2f == _T_174[7:0] ? 4'h0 : _GEN_3253; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3255 = 8'h30 == _T_174[7:0] ? 4'h2 : _GEN_3254; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3256 = 8'h31 == _T_174[7:0] ? 4'h2 : _GEN_3255; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3257 = 8'h32 == _T_174[7:0] ? 4'h0 : _GEN_3256; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3258 = 8'h33 == _T_174[7:0] ? 4'h0 : _GEN_3257; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3259 = 8'h34 == _T_174[7:0] ? 4'h0 : _GEN_3258; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3260 = 8'h35 == _T_174[7:0] ? 4'h0 : _GEN_3259; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3261 = 8'h36 == _T_174[7:0] ? 4'h0 : _GEN_3260; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3262 = 8'h37 == _T_174[7:0] ? 4'h0 : _GEN_3261; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3263 = 8'h38 == _T_174[7:0] ? 4'h2 : _GEN_3262; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3264 = 8'h39 == _T_174[7:0] ? 4'h0 : _GEN_3263; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3265 = 8'h3a == _T_174[7:0] ? 4'h0 : _GEN_3264; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3266 = 8'h3b == _T_174[7:0] ? 4'h0 : _GEN_3265; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3267 = 8'h3c == _T_174[7:0] ? 4'h0 : _GEN_3266; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3268 = 8'h3d == _T_174[7:0] ? 4'h0 : _GEN_3267; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3269 = 8'h3e == _T_174[7:0] ? 4'h0 : _GEN_3268; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3270 = 8'h3f == _T_174[7:0] ? 4'h0 : _GEN_3269; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3271 = 8'h40 == _T_174[7:0] ? 4'h0 : _GEN_3270; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3272 = 8'h41 == _T_174[7:0] ? 4'h0 : _GEN_3271; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3273 = 8'h42 == _T_174[7:0] ? 4'h0 : _GEN_3272; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3274 = 8'h43 == _T_174[7:0] ? 4'h0 : _GEN_3273; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3275 = 8'h44 == _T_174[7:0] ? 4'h1 : _GEN_3274; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3276 = 8'h45 == _T_174[7:0] ? 4'h3 : _GEN_3275; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3277 = 8'h46 == _T_174[7:0] ? 4'h7 : _GEN_3276; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3278 = 8'h47 == _T_174[7:0] ? 4'h0 : _GEN_3277; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3279 = 8'h48 == _T_174[7:0] ? 4'h0 : _GEN_3278; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3280 = 8'h49 == _T_174[7:0] ? 4'h0 : _GEN_3279; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3281 = 8'h4a == _T_174[7:0] ? 4'h0 : _GEN_3280; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3282 = 8'h4b == _T_174[7:0] ? 4'h0 : _GEN_3281; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3283 = 8'h4c == _T_174[7:0] ? 4'h0 : _GEN_3282; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3284 = 8'h4d == _T_174[7:0] ? 4'h0 : _GEN_3283; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3285 = 8'h4e == _T_174[7:0] ? 4'h2 : _GEN_3284; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3286 = 8'h4f == _T_174[7:0] ? 4'h0 : _GEN_3285; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3287 = 8'h50 == _T_174[7:0] ? 4'h0 : _GEN_3286; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3288 = 8'h51 == _T_174[7:0] ? 4'h0 : _GEN_3287; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3289 = 8'h52 == _T_174[7:0] ? 4'h0 : _GEN_3288; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3290 = 8'h53 == _T_174[7:0] ? 4'h0 : _GEN_3289; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3291 = 8'h54 == _T_174[7:0] ? 4'h0 : _GEN_3290; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3292 = 8'h55 == _T_174[7:0] ? 4'h0 : _GEN_3291; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3293 = 8'h56 == _T_174[7:0] ? 4'h0 : _GEN_3292; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3294 = 8'h57 == _T_174[7:0] ? 4'h0 : _GEN_3293; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3295 = 8'h58 == _T_174[7:0] ? 4'h0 : _GEN_3294; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3296 = 8'h59 == _T_174[7:0] ? 4'h2 : _GEN_3295; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3297 = 8'h5a == _T_174[7:0] ? 4'h2 : _GEN_3296; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3298 = 8'h5b == _T_174[7:0] ? 4'h0 : _GEN_3297; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3299 = 8'h5c == _T_174[7:0] ? 4'h0 : _GEN_3298; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3300 = 8'h5d == _T_174[7:0] ? 4'h0 : _GEN_3299; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3301 = 8'h5e == _T_174[7:0] ? 4'h4 : _GEN_3300; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3302 = 8'h5f == _T_174[7:0] ? 4'h0 : _GEN_3301; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3303 = 8'h60 == _T_174[7:0] ? 4'h0 : _GEN_3302; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3304 = 8'h61 == _T_174[7:0] ? 4'h0 : _GEN_3303; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3305 = 8'h62 == _T_174[7:0] ? 4'h0 : _GEN_3304; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3306 = 8'h63 == _T_174[7:0] ? 4'h2 : _GEN_3305; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3307 = 8'h64 == _T_174[7:0] ? 4'h0 : _GEN_3306; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3308 = 8'h65 == _T_174[7:0] ? 4'h0 : _GEN_3307; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3309 = 8'h66 == _T_174[7:0] ? 4'h0 : _GEN_3308; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3310 = 8'h67 == _T_174[7:0] ? 4'h0 : _GEN_3309; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3311 = 8'h68 == _T_174[7:0] ? 4'h0 : _GEN_3310; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3312 = 8'h69 == _T_174[7:0] ? 4'h0 : _GEN_3311; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3313 = 8'h6a == _T_174[7:0] ? 4'h0 : _GEN_3312; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3314 = 8'h6b == _T_174[7:0] ? 4'h0 : _GEN_3313; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3315 = 8'h6c == _T_174[7:0] ? 4'h0 : _GEN_3314; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3316 = 8'h6d == _T_174[7:0] ? 4'h0 : _GEN_3315; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3317 = 8'h6e == _T_174[7:0] ? 4'h2 : _GEN_3316; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3318 = 8'h6f == _T_174[7:0] ? 4'h0 : _GEN_3317; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3319 = 8'h70 == _T_174[7:0] ? 4'h0 : _GEN_3318; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3320 = 8'h71 == _T_174[7:0] ? 4'h0 : _GEN_3319; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3321 = 8'h72 == _T_174[7:0] ? 4'h2 : _GEN_3320; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3322 = 8'h73 == _T_174[7:0] ? 4'h9 : _GEN_3321; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3323 = 8'h74 == _T_174[7:0] ? 4'h2 : _GEN_3322; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3324 = 8'h75 == _T_174[7:0] ? 4'h0 : _GEN_3323; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3325 = 8'h76 == _T_174[7:0] ? 4'h0 : _GEN_3324; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3326 = 8'h77 == _T_174[7:0] ? 4'h0 : _GEN_3325; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3327 = 8'h78 == _T_174[7:0] ? 4'h1 : _GEN_3326; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3328 = 8'h79 == _T_174[7:0] ? 4'h1 : _GEN_3327; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3329 = 8'h7a == _T_174[7:0] ? 4'h0 : _GEN_3328; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3330 = 8'h7b == _T_174[7:0] ? 4'h0 : _GEN_3329; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3331 = 8'h7c == _T_174[7:0] ? 4'h0 : _GEN_3330; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3332 = 8'h7d == _T_174[7:0] ? 4'h0 : _GEN_3331; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3333 = 8'h7e == _T_174[7:0] ? 4'h0 : _GEN_3332; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3334 = 8'h7f == _T_174[7:0] ? 4'h0 : _GEN_3333; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3335 = 8'h80 == _T_174[7:0] ? 4'h0 : _GEN_3334; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3336 = 8'h81 == _T_174[7:0] ? 4'h0 : _GEN_3335; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3337 = 8'h82 == _T_174[7:0] ? 4'h2 : _GEN_3336; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3338 = 8'h83 == _T_174[7:0] ? 4'h0 : _GEN_3337; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3339 = 8'h84 == _T_174[7:0] ? 4'h0 : _GEN_3338; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3340 = 8'h85 == _T_174[7:0] ? 4'h0 : _GEN_3339; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3341 = 8'h86 == _T_174[7:0] ? 4'h7 : _GEN_3340; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3342 = 8'h87 == _T_174[7:0] ? 4'h2 : _GEN_3341; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3343 = 8'h88 == _T_174[7:0] ? 4'h0 : _GEN_3342; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3344 = 8'h89 == _T_174[7:0] ? 4'h2 : _GEN_3343; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3345 = 8'h8a == _T_174[7:0] ? 4'h7 : _GEN_3344; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3346 = 8'h8b == _T_174[7:0] ? 4'h0 : _GEN_3345; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3347 = 8'h8c == _T_174[7:0] ? 4'h0 : _GEN_3346; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3348 = 8'h8d == _T_174[7:0] ? 4'h0 : _GEN_3347; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3349 = 8'h8e == _T_174[7:0] ? 4'h2 : _GEN_3348; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3350 = 8'h8f == _T_174[7:0] ? 4'h0 : _GEN_3349; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3351 = 8'h90 == _T_174[7:0] ? 4'h0 : _GEN_3350; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3352 = 8'h91 == _T_174[7:0] ? 4'h0 : _GEN_3351; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3353 = 8'h92 == _T_174[7:0] ? 4'h0 : _GEN_3352; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3354 = 8'h93 == _T_174[7:0] ? 4'h0 : _GEN_3353; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3355 = 8'h94 == _T_174[7:0] ? 4'h0 : _GEN_3354; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3356 = 8'h95 == _T_174[7:0] ? 4'h0 : _GEN_3355; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3357 = 8'h96 == _T_174[7:0] ? 4'h0 : _GEN_3356; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3358 = 8'h97 == _T_174[7:0] ? 4'h2 : _GEN_3357; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3359 = 8'h98 == _T_174[7:0] ? 4'h2 : _GEN_3358; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3360 = 8'h99 == _T_174[7:0] ? 4'h1 : _GEN_3359; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3361 = 8'h9a == _T_174[7:0] ? 4'h0 : _GEN_3360; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3362 = 8'h9b == _T_174[7:0] ? 4'h7 : _GEN_3361; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3363 = 8'h9c == _T_174[7:0] ? 4'h7 : _GEN_3362; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3364 = 8'h9d == _T_174[7:0] ? 4'h0 : _GEN_3363; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3365 = 8'h9e == _T_174[7:0] ? 4'h7 : _GEN_3364; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3366 = 8'h9f == _T_174[7:0] ? 4'h7 : _GEN_3365; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3367 = 8'ha0 == _T_174[7:0] ? 4'h0 : _GEN_3366; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3368 = 8'ha1 == _T_174[7:0] ? 4'h1 : _GEN_3367; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3369 = 8'ha2 == _T_174[7:0] ? 4'h2 : _GEN_3368; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3370 = 8'ha3 == _T_174[7:0] ? 4'h2 : _GEN_3369; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3371 = 8'ha4 == _T_174[7:0] ? 4'h0 : _GEN_3370; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3372 = 8'ha5 == _T_174[7:0] ? 4'h0 : _GEN_3371; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3373 = 8'ha6 == _T_174[7:0] ? 4'h0 : _GEN_3372; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3374 = 8'ha7 == _T_174[7:0] ? 4'h0 : _GEN_3373; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3375 = 8'ha8 == _T_174[7:0] ? 4'h0 : _GEN_3374; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3376 = 8'ha9 == _T_174[7:0] ? 4'h0 : _GEN_3375; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3377 = 8'haa == _T_174[7:0] ? 4'h0 : _GEN_3376; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3378 = 8'hab == _T_174[7:0] ? 4'h0 : _GEN_3377; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3379 = 8'hac == _T_174[7:0] ? 4'h2 : _GEN_3378; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3380 = 8'had == _T_174[7:0] ? 4'h0 : _GEN_3379; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3381 = 8'hae == _T_174[7:0] ? 4'h1 : _GEN_3380; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3382 = 8'haf == _T_174[7:0] ? 4'h3 : _GEN_3381; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3383 = 8'hb0 == _T_174[7:0] ? 4'h1 : _GEN_3382; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3384 = 8'hb1 == _T_174[7:0] ? 4'h0 : _GEN_3383; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3385 = 8'hb2 == _T_174[7:0] ? 4'h0 : _GEN_3384; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3386 = 8'hb3 == _T_174[7:0] ? 4'h0 : _GEN_3385; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3387 = 8'hb4 == _T_174[7:0] ? 4'h1 : _GEN_3386; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3388 = 8'hb5 == _T_174[7:0] ? 4'h3 : _GEN_3387; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3389 = 8'hb6 == _T_174[7:0] ? 4'h1 : _GEN_3388; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3390 = 8'hb7 == _T_174[7:0] ? 4'h0 : _GEN_3389; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3391 = 8'hb8 == _T_174[7:0] ? 4'h2 : _GEN_3390; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3392 = 8'hb9 == _T_174[7:0] ? 4'h0 : _GEN_3391; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3393 = 8'hba == _T_174[7:0] ? 4'h0 : _GEN_3392; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3394 = 8'hbb == _T_174[7:0] ? 4'h0 : _GEN_3393; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3395 = 8'hbc == _T_174[7:0] ? 4'h0 : _GEN_3394; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3396 = 8'hbd == _T_174[7:0] ? 4'h0 : _GEN_3395; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3397 = 8'hbe == _T_174[7:0] ? 4'h0 : _GEN_3396; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3398 = 8'hbf == _T_174[7:0] ? 4'h0 : _GEN_3397; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3399 = 8'hc0 == _T_174[7:0] ? 4'h0 : _GEN_3398; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3400 = 8'hc1 == _T_174[7:0] ? 4'h0 : _GEN_3399; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3401 = 8'hc2 == _T_174[7:0] ? 4'h3 : _GEN_3400; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3402 = 8'hc3 == _T_174[7:0] ? 4'h0 : _GEN_3401; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3403 = 8'hc4 == _T_174[7:0] ? 4'h0 : _GEN_3402; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3404 = 8'hc5 == _T_174[7:0] ? 4'h2 : _GEN_3403; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3405 = 8'hc6 == _T_174[7:0] ? 4'h3 : _GEN_3404; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3406 = 8'hc7 == _T_174[7:0] ? 4'h2 : _GEN_3405; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3407 = 8'hc8 == _T_174[7:0] ? 4'h3 : _GEN_3406; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3408 = 8'hc9 == _T_174[7:0] ? 4'h2 : _GEN_3407; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3409 = 8'hca == _T_174[7:0] ? 4'h0 : _GEN_3408; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3410 = 8'hcb == _T_174[7:0] ? 4'h0 : _GEN_3409; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3411 = 8'hcc == _T_174[7:0] ? 4'h3 : _GEN_3410; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3412 = 8'hcd == _T_174[7:0] ? 4'h0 : _GEN_3411; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3413 = 8'hce == _T_174[7:0] ? 4'h0 : _GEN_3412; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3414 = 8'hcf == _T_174[7:0] ? 4'h0 : _GEN_3413; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3415 = 8'hd0 == _T_174[7:0] ? 4'h0 : _GEN_3414; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3416 = 8'hd1 == _T_174[7:0] ? 4'h0 : _GEN_3415; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3417 = 8'hd2 == _T_174[7:0] ? 4'h0 : _GEN_3416; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3418 = 8'hd3 == _T_174[7:0] ? 4'h0 : _GEN_3417; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3419 = 8'hd4 == _T_174[7:0] ? 4'h0 : _GEN_3418; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3420 = 8'hd5 == _T_174[7:0] ? 4'h0 : _GEN_3419; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3421 = 8'hd6 == _T_174[7:0] ? 4'h0 : _GEN_3420; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3422 = 8'hd7 == _T_174[7:0] ? 4'h2 : _GEN_3421; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3423 = 8'hd8 == _T_174[7:0] ? 4'h2 : _GEN_3422; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3424 = 8'hd9 == _T_174[7:0] ? 4'h0 : _GEN_3423; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3425 = 8'hda == _T_174[7:0] ? 4'h7 : _GEN_3424; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3426 = 8'hdb == _T_174[7:0] ? 4'h1 : _GEN_3425; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3427 = 8'hdc == _T_174[7:0] ? 4'h4 : _GEN_3426; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3428 = 8'hdd == _T_174[7:0] ? 4'h1 : _GEN_3427; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3429 = 8'hde == _T_174[7:0] ? 4'h7 : _GEN_3428; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3430 = 8'hdf == _T_174[7:0] ? 4'h0 : _GEN_3429; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3431 = 8'he0 == _T_174[7:0] ? 4'h2 : _GEN_3430; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3432 = 8'he1 == _T_174[7:0] ? 4'h2 : _GEN_3431; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3433 = 8'he2 == _T_174[7:0] ? 4'h0 : _GEN_3432; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3434 = 8'he3 == _T_174[7:0] ? 4'h0 : _GEN_3433; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3435 = 8'he4 == _T_174[7:0] ? 4'h0 : _GEN_3434; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3436 = 8'he5 == _T_174[7:0] ? 4'h0 : _GEN_3435; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3437 = 8'he6 == _T_174[7:0] ? 4'h0 : _GEN_3436; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3438 = 8'he7 == _T_174[7:0] ? 4'h0 : _GEN_3437; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3439 = 8'he8 == _T_174[7:0] ? 4'h0 : _GEN_3438; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3440 = 8'he9 == _T_174[7:0] ? 4'h0 : _GEN_3439; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3441 = 8'hea == _T_174[7:0] ? 4'h0 : _GEN_3440; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3442 = 8'heb == _T_174[7:0] ? 4'h0 : _GEN_3441; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3443 = 8'hec == _T_174[7:0] ? 4'h0 : _GEN_3442; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3444 = 8'hed == _T_174[7:0] ? 4'h0 : _GEN_3443; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3445 = 8'hee == _T_174[7:0] ? 4'h0 : _GEN_3444; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3446 = 8'hef == _T_174[7:0] ? 4'h0 : _GEN_3445; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3447 = 8'hf0 == _T_174[7:0] ? 4'h0 : _GEN_3446; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3448 = 8'hf1 == _T_174[7:0] ? 4'h0 : _GEN_3447; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3449 = 8'hf2 == _T_174[7:0] ? 4'h0 : _GEN_3448; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3450 = 8'hf3 == _T_174[7:0] ? 4'h0 : _GEN_3449; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3451 = 8'hf4 == _T_174[7:0] ? 4'h0 : _GEN_3450; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3452 = 8'hf5 == _T_174[7:0] ? 4'h0 : _GEN_3451; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3453 = 8'hf6 == _T_174[7:0] ? 4'h0 : _GEN_3452; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3454 = 8'hf7 == _T_174[7:0] ? 4'h0 : _GEN_3453; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3455 = 8'hf8 == _T_174[7:0] ? 4'h0 : _GEN_3454; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3456 = 8'hf9 == _T_174[7:0] ? 4'h0 : _GEN_3455; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3457 = 8'hfa == _T_174[7:0] ? 4'h0 : _GEN_3456; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3458 = 8'hfb == _T_174[7:0] ? 4'h0 : _GEN_3457; // @[Filter.scala 204:62]
  wire [4:0] _GEN_11237 = {{1'd0}, _GEN_3458}; // @[Filter.scala 204:62]
  wire [8:0] _T_176 = _GEN_11237 * 5'h14; // @[Filter.scala 204:62]
  wire [3:0] _GEN_3508 = 8'h31 == _T_174[7:0] ? 4'h3 : _GEN_3255; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3509 = 8'h32 == _T_174[7:0] ? 4'h3 : _GEN_3508; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3510 = 8'h33 == _T_174[7:0] ? 4'h6 : _GEN_3509; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3511 = 8'h34 == _T_174[7:0] ? 4'h6 : _GEN_3510; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3512 = 8'h35 == _T_174[7:0] ? 4'h0 : _GEN_3511; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3513 = 8'h36 == _T_174[7:0] ? 4'h0 : _GEN_3512; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3514 = 8'h37 == _T_174[7:0] ? 4'h0 : _GEN_3513; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3515 = 8'h38 == _T_174[7:0] ? 4'h2 : _GEN_3514; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3516 = 8'h39 == _T_174[7:0] ? 4'h0 : _GEN_3515; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3517 = 8'h3a == _T_174[7:0] ? 4'h0 : _GEN_3516; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3518 = 8'h3b == _T_174[7:0] ? 4'h0 : _GEN_3517; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3519 = 8'h3c == _T_174[7:0] ? 4'h0 : _GEN_3518; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3520 = 8'h3d == _T_174[7:0] ? 4'h0 : _GEN_3519; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3521 = 8'h3e == _T_174[7:0] ? 4'h0 : _GEN_3520; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3522 = 8'h3f == _T_174[7:0] ? 4'h0 : _GEN_3521; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3523 = 8'h40 == _T_174[7:0] ? 4'h0 : _GEN_3522; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3524 = 8'h41 == _T_174[7:0] ? 4'h0 : _GEN_3523; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3525 = 8'h42 == _T_174[7:0] ? 4'h0 : _GEN_3524; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3526 = 8'h43 == _T_174[7:0] ? 4'h0 : _GEN_3525; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3527 = 8'h44 == _T_174[7:0] ? 4'h1 : _GEN_3526; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3528 = 8'h45 == _T_174[7:0] ? 4'h4 : _GEN_3527; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3529 = 8'h46 == _T_174[7:0] ? 4'hb : _GEN_3528; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3530 = 8'h47 == _T_174[7:0] ? 4'h0 : _GEN_3529; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3531 = 8'h48 == _T_174[7:0] ? 4'h0 : _GEN_3530; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3532 = 8'h49 == _T_174[7:0] ? 4'h0 : _GEN_3531; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3533 = 8'h4a == _T_174[7:0] ? 4'h6 : _GEN_3532; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3534 = 8'h4b == _T_174[7:0] ? 4'h0 : _GEN_3533; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3535 = 8'h4c == _T_174[7:0] ? 4'h3 : _GEN_3534; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3536 = 8'h4d == _T_174[7:0] ? 4'h3 : _GEN_3535; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3537 = 8'h4e == _T_174[7:0] ? 4'h2 : _GEN_3536; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3538 = 8'h4f == _T_174[7:0] ? 4'h0 : _GEN_3537; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3539 = 8'h50 == _T_174[7:0] ? 4'h0 : _GEN_3538; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3540 = 8'h51 == _T_174[7:0] ? 4'h0 : _GEN_3539; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3541 = 8'h52 == _T_174[7:0] ? 4'h0 : _GEN_3540; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3542 = 8'h53 == _T_174[7:0] ? 4'h0 : _GEN_3541; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3543 = 8'h54 == _T_174[7:0] ? 4'h0 : _GEN_3542; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3544 = 8'h55 == _T_174[7:0] ? 4'h0 : _GEN_3543; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3545 = 8'h56 == _T_174[7:0] ? 4'h0 : _GEN_3544; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3546 = 8'h57 == _T_174[7:0] ? 4'h0 : _GEN_3545; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3547 = 8'h58 == _T_174[7:0] ? 4'h0 : _GEN_3546; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3548 = 8'h59 == _T_174[7:0] ? 4'h2 : _GEN_3547; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3549 = 8'h5a == _T_174[7:0] ? 4'h3 : _GEN_3548; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3550 = 8'h5b == _T_174[7:0] ? 4'h0 : _GEN_3549; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3551 = 8'h5c == _T_174[7:0] ? 4'h0 : _GEN_3550; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3552 = 8'h5d == _T_174[7:0] ? 4'h3 : _GEN_3551; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3553 = 8'h5e == _T_174[7:0] ? 4'hd : _GEN_3552; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3554 = 8'h5f == _T_174[7:0] ? 4'h3 : _GEN_3553; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3555 = 8'h60 == _T_174[7:0] ? 4'h0 : _GEN_3554; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3556 = 8'h61 == _T_174[7:0] ? 4'h6 : _GEN_3555; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3557 = 8'h62 == _T_174[7:0] ? 4'h0 : _GEN_3556; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3558 = 8'h63 == _T_174[7:0] ? 4'h2 : _GEN_3557; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3559 = 8'h64 == _T_174[7:0] ? 4'h0 : _GEN_3558; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3560 = 8'h65 == _T_174[7:0] ? 4'h0 : _GEN_3559; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3561 = 8'h66 == _T_174[7:0] ? 4'h0 : _GEN_3560; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3562 = 8'h67 == _T_174[7:0] ? 4'h0 : _GEN_3561; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3563 = 8'h68 == _T_174[7:0] ? 4'h0 : _GEN_3562; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3564 = 8'h69 == _T_174[7:0] ? 4'h0 : _GEN_3563; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3565 = 8'h6a == _T_174[7:0] ? 4'h0 : _GEN_3564; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3566 = 8'h6b == _T_174[7:0] ? 4'h0 : _GEN_3565; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3567 = 8'h6c == _T_174[7:0] ? 4'h0 : _GEN_3566; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3568 = 8'h6d == _T_174[7:0] ? 4'h0 : _GEN_3567; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3569 = 8'h6e == _T_174[7:0] ? 4'h2 : _GEN_3568; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3570 = 8'h6f == _T_174[7:0] ? 4'h0 : _GEN_3569; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3571 = 8'h70 == _T_174[7:0] ? 4'h0 : _GEN_3570; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3572 = 8'h71 == _T_174[7:0] ? 4'h0 : _GEN_3571; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3573 = 8'h72 == _T_174[7:0] ? 4'h6 : _GEN_3572; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3574 = 8'h73 == _T_174[7:0] ? 4'he : _GEN_3573; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3575 = 8'h74 == _T_174[7:0] ? 4'h6 : _GEN_3574; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3576 = 8'h75 == _T_174[7:0] ? 4'h0 : _GEN_3575; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3577 = 8'h76 == _T_174[7:0] ? 4'h6 : _GEN_3576; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3578 = 8'h77 == _T_174[7:0] ? 4'h3 : _GEN_3577; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3579 = 8'h78 == _T_174[7:0] ? 4'h4 : _GEN_3578; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3580 = 8'h79 == _T_174[7:0] ? 4'h1 : _GEN_3579; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3581 = 8'h7a == _T_174[7:0] ? 4'h0 : _GEN_3580; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3582 = 8'h7b == _T_174[7:0] ? 4'h0 : _GEN_3581; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3583 = 8'h7c == _T_174[7:0] ? 4'h0 : _GEN_3582; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3584 = 8'h7d == _T_174[7:0] ? 4'h0 : _GEN_3583; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3585 = 8'h7e == _T_174[7:0] ? 4'h0 : _GEN_3584; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3586 = 8'h7f == _T_174[7:0] ? 4'h0 : _GEN_3585; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3587 = 8'h80 == _T_174[7:0] ? 4'h0 : _GEN_3586; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3588 = 8'h81 == _T_174[7:0] ? 4'h0 : _GEN_3587; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3589 = 8'h82 == _T_174[7:0] ? 4'h2 : _GEN_3588; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3590 = 8'h83 == _T_174[7:0] ? 4'h3 : _GEN_3589; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3591 = 8'h84 == _T_174[7:0] ? 4'h6 : _GEN_3590; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3592 = 8'h85 == _T_174[7:0] ? 4'h6 : _GEN_3591; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3593 = 8'h86 == _T_174[7:0] ? 4'he : _GEN_3592; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3594 = 8'h87 == _T_174[7:0] ? 4'ha : _GEN_3593; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3595 = 8'h88 == _T_174[7:0] ? 4'h6 : _GEN_3594; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3596 = 8'h89 == _T_174[7:0] ? 4'ha : _GEN_3595; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3597 = 8'h8a == _T_174[7:0] ? 4'he : _GEN_3596; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3598 = 8'h8b == _T_174[7:0] ? 4'h3 : _GEN_3597; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3599 = 8'h8c == _T_174[7:0] ? 4'h3 : _GEN_3598; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3600 = 8'h8d == _T_174[7:0] ? 4'h0 : _GEN_3599; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3601 = 8'h8e == _T_174[7:0] ? 4'h2 : _GEN_3600; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3602 = 8'h8f == _T_174[7:0] ? 4'h0 : _GEN_3601; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3603 = 8'h90 == _T_174[7:0] ? 4'h0 : _GEN_3602; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3604 = 8'h91 == _T_174[7:0] ? 4'h0 : _GEN_3603; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3605 = 8'h92 == _T_174[7:0] ? 4'h0 : _GEN_3604; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3606 = 8'h93 == _T_174[7:0] ? 4'h0 : _GEN_3605; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3607 = 8'h94 == _T_174[7:0] ? 4'h0 : _GEN_3606; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3608 = 8'h95 == _T_174[7:0] ? 4'h0 : _GEN_3607; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3609 = 8'h96 == _T_174[7:0] ? 4'h0 : _GEN_3608; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3610 = 8'h97 == _T_174[7:0] ? 4'h2 : _GEN_3609; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3611 = 8'h98 == _T_174[7:0] ? 4'h2 : _GEN_3610; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3612 = 8'h99 == _T_174[7:0] ? 4'h1 : _GEN_3611; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3613 = 8'h9a == _T_174[7:0] ? 4'h3 : _GEN_3612; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3614 = 8'h9b == _T_174[7:0] ? 4'he : _GEN_3613; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3615 = 8'h9c == _T_174[7:0] ? 4'he : _GEN_3614; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3616 = 8'h9d == _T_174[7:0] ? 4'h0 : _GEN_3615; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3617 = 8'h9e == _T_174[7:0] ? 4'he : _GEN_3616; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3618 = 8'h9f == _T_174[7:0] ? 4'he : _GEN_3617; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3619 = 8'ha0 == _T_174[7:0] ? 4'h3 : _GEN_3618; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3620 = 8'ha1 == _T_174[7:0] ? 4'h1 : _GEN_3619; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3621 = 8'ha2 == _T_174[7:0] ? 4'h2 : _GEN_3620; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3622 = 8'ha3 == _T_174[7:0] ? 4'h2 : _GEN_3621; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3623 = 8'ha4 == _T_174[7:0] ? 4'h0 : _GEN_3622; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3624 = 8'ha5 == _T_174[7:0] ? 4'h0 : _GEN_3623; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3625 = 8'ha6 == _T_174[7:0] ? 4'h0 : _GEN_3624; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3626 = 8'ha7 == _T_174[7:0] ? 4'h0 : _GEN_3625; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3627 = 8'ha8 == _T_174[7:0] ? 4'h0 : _GEN_3626; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3628 = 8'ha9 == _T_174[7:0] ? 4'h0 : _GEN_3627; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3629 = 8'haa == _T_174[7:0] ? 4'h0 : _GEN_3628; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3630 = 8'hab == _T_174[7:0] ? 4'h0 : _GEN_3629; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3631 = 8'hac == _T_174[7:0] ? 4'h2 : _GEN_3630; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3632 = 8'had == _T_174[7:0] ? 4'h3 : _GEN_3631; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3633 = 8'hae == _T_174[7:0] ? 4'h4 : _GEN_3632; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3634 = 8'haf == _T_174[7:0] ? 4'h3 : _GEN_3633; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3635 = 8'hb0 == _T_174[7:0] ? 4'h4 : _GEN_3634; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3636 = 8'hb1 == _T_174[7:0] ? 4'h3 : _GEN_3635; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3637 = 8'hb2 == _T_174[7:0] ? 4'h0 : _GEN_3636; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3638 = 8'hb3 == _T_174[7:0] ? 4'h3 : _GEN_3637; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3639 = 8'hb4 == _T_174[7:0] ? 4'h4 : _GEN_3638; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3640 = 8'hb5 == _T_174[7:0] ? 4'h3 : _GEN_3639; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3641 = 8'hb6 == _T_174[7:0] ? 4'h4 : _GEN_3640; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3642 = 8'hb7 == _T_174[7:0] ? 4'h3 : _GEN_3641; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3643 = 8'hb8 == _T_174[7:0] ? 4'h2 : _GEN_3642; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3644 = 8'hb9 == _T_174[7:0] ? 4'h0 : _GEN_3643; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3645 = 8'hba == _T_174[7:0] ? 4'h0 : _GEN_3644; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3646 = 8'hbb == _T_174[7:0] ? 4'h0 : _GEN_3645; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3647 = 8'hbc == _T_174[7:0] ? 4'h0 : _GEN_3646; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3648 = 8'hbd == _T_174[7:0] ? 4'h0 : _GEN_3647; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3649 = 8'hbe == _T_174[7:0] ? 4'h0 : _GEN_3648; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3650 = 8'hbf == _T_174[7:0] ? 4'h0 : _GEN_3649; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3651 = 8'hc0 == _T_174[7:0] ? 4'h0 : _GEN_3650; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3652 = 8'hc1 == _T_174[7:0] ? 4'h0 : _GEN_3651; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3653 = 8'hc2 == _T_174[7:0] ? 4'h8 : _GEN_3652; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3654 = 8'hc3 == _T_174[7:0] ? 4'hc : _GEN_3653; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3655 = 8'hc4 == _T_174[7:0] ? 4'h0 : _GEN_3654; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3656 = 8'hc5 == _T_174[7:0] ? 4'h2 : _GEN_3655; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3657 = 8'hc6 == _T_174[7:0] ? 4'h3 : _GEN_3656; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3658 = 8'hc7 == _T_174[7:0] ? 4'h2 : _GEN_3657; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3659 = 8'hc8 == _T_174[7:0] ? 4'h3 : _GEN_3658; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3660 = 8'hc9 == _T_174[7:0] ? 4'h2 : _GEN_3659; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3661 = 8'hca == _T_174[7:0] ? 4'h0 : _GEN_3660; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3662 = 8'hcb == _T_174[7:0] ? 4'hc : _GEN_3661; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3663 = 8'hcc == _T_174[7:0] ? 4'h8 : _GEN_3662; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3664 = 8'hcd == _T_174[7:0] ? 4'h0 : _GEN_3663; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3665 = 8'hce == _T_174[7:0] ? 4'h0 : _GEN_3664; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3666 = 8'hcf == _T_174[7:0] ? 4'h0 : _GEN_3665; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3667 = 8'hd0 == _T_174[7:0] ? 4'h0 : _GEN_3666; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3668 = 8'hd1 == _T_174[7:0] ? 4'h0 : _GEN_3667; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3669 = 8'hd2 == _T_174[7:0] ? 4'h0 : _GEN_3668; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3670 = 8'hd3 == _T_174[7:0] ? 4'h0 : _GEN_3669; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3671 = 8'hd4 == _T_174[7:0] ? 4'h0 : _GEN_3670; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3672 = 8'hd5 == _T_174[7:0] ? 4'h0 : _GEN_3671; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3673 = 8'hd6 == _T_174[7:0] ? 4'h0 : _GEN_3672; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3674 = 8'hd7 == _T_174[7:0] ? 4'h3 : _GEN_3673; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3675 = 8'hd8 == _T_174[7:0] ? 4'h6 : _GEN_3674; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3676 = 8'hd9 == _T_174[7:0] ? 4'h0 : _GEN_3675; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3677 = 8'hda == _T_174[7:0] ? 4'hb : _GEN_3676; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3678 = 8'hdb == _T_174[7:0] ? 4'h1 : _GEN_3677; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3679 = 8'hdc == _T_174[7:0] ? 4'h4 : _GEN_3678; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3680 = 8'hdd == _T_174[7:0] ? 4'h1 : _GEN_3679; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3681 = 8'hde == _T_174[7:0] ? 4'hb : _GEN_3680; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3682 = 8'hdf == _T_174[7:0] ? 4'h0 : _GEN_3681; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3683 = 8'he0 == _T_174[7:0] ? 4'h6 : _GEN_3682; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3684 = 8'he1 == _T_174[7:0] ? 4'h3 : _GEN_3683; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3685 = 8'he2 == _T_174[7:0] ? 4'h0 : _GEN_3684; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3686 = 8'he3 == _T_174[7:0] ? 4'h0 : _GEN_3685; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3687 = 8'he4 == _T_174[7:0] ? 4'h0 : _GEN_3686; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3688 = 8'he5 == _T_174[7:0] ? 4'h0 : _GEN_3687; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3689 = 8'he6 == _T_174[7:0] ? 4'h0 : _GEN_3688; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3690 = 8'he7 == _T_174[7:0] ? 4'h0 : _GEN_3689; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3691 = 8'he8 == _T_174[7:0] ? 4'h0 : _GEN_3690; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3692 = 8'he9 == _T_174[7:0] ? 4'h0 : _GEN_3691; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3693 = 8'hea == _T_174[7:0] ? 4'h0 : _GEN_3692; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3694 = 8'heb == _T_174[7:0] ? 4'h0 : _GEN_3693; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3695 = 8'hec == _T_174[7:0] ? 4'h0 : _GEN_3694; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3696 = 8'hed == _T_174[7:0] ? 4'h0 : _GEN_3695; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3697 = 8'hee == _T_174[7:0] ? 4'h0 : _GEN_3696; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3698 = 8'hef == _T_174[7:0] ? 4'h0 : _GEN_3697; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3699 = 8'hf0 == _T_174[7:0] ? 4'h0 : _GEN_3698; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3700 = 8'hf1 == _T_174[7:0] ? 4'h0 : _GEN_3699; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3701 = 8'hf2 == _T_174[7:0] ? 4'h0 : _GEN_3700; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3702 = 8'hf3 == _T_174[7:0] ? 4'h0 : _GEN_3701; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3703 = 8'hf4 == _T_174[7:0] ? 4'h0 : _GEN_3702; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3704 = 8'hf5 == _T_174[7:0] ? 4'h0 : _GEN_3703; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3705 = 8'hf6 == _T_174[7:0] ? 4'h0 : _GEN_3704; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3706 = 8'hf7 == _T_174[7:0] ? 4'h0 : _GEN_3705; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3707 = 8'hf8 == _T_174[7:0] ? 4'h0 : _GEN_3706; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3708 = 8'hf9 == _T_174[7:0] ? 4'h0 : _GEN_3707; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3709 = 8'hfa == _T_174[7:0] ? 4'h0 : _GEN_3708; // @[Filter.scala 204:102]
  wire [3:0] _GEN_3710 = 8'hfb == _T_174[7:0] ? 4'h0 : _GEN_3709; // @[Filter.scala 204:102]
  wire [6:0] _GEN_11239 = {{3'd0}, _GEN_3710}; // @[Filter.scala 204:102]
  wire [10:0] _T_181 = _GEN_11239 * 7'h46; // @[Filter.scala 204:102]
  wire [10:0] _GEN_11240 = {{2'd0}, _T_176}; // @[Filter.scala 204:69]
  wire [10:0] _T_183 = _GEN_11240 + _T_181; // @[Filter.scala 204:69]
  wire [3:0] _GEN_3719 = 8'h8 == _T_174[7:0] ? 4'h3 : 4'h0; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3720 = 8'h9 == _T_174[7:0] ? 4'h6 : _GEN_3719; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3721 = 8'ha == _T_174[7:0] ? 4'h6 : _GEN_3720; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3722 = 8'hb == _T_174[7:0] ? 4'h6 : _GEN_3721; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3723 = 8'hc == _T_174[7:0] ? 4'h3 : _GEN_3722; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3724 = 8'hd == _T_174[7:0] ? 4'h0 : _GEN_3723; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3725 = 8'he == _T_174[7:0] ? 4'h0 : _GEN_3724; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3726 = 8'hf == _T_174[7:0] ? 4'h0 : _GEN_3725; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3727 = 8'h10 == _T_174[7:0] ? 4'h0 : _GEN_3726; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3728 = 8'h11 == _T_174[7:0] ? 4'h0 : _GEN_3727; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3729 = 8'h12 == _T_174[7:0] ? 4'h0 : _GEN_3728; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3730 = 8'h13 == _T_174[7:0] ? 4'h0 : _GEN_3729; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3731 = 8'h14 == _T_174[7:0] ? 4'h0 : _GEN_3730; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3732 = 8'h15 == _T_174[7:0] ? 4'h0 : _GEN_3731; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3733 = 8'h16 == _T_174[7:0] ? 4'h0 : _GEN_3732; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3734 = 8'h17 == _T_174[7:0] ? 4'h0 : _GEN_3733; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3735 = 8'h18 == _T_174[7:0] ? 4'h0 : _GEN_3734; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3736 = 8'h19 == _T_174[7:0] ? 4'h0 : _GEN_3735; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3737 = 8'h1a == _T_174[7:0] ? 4'h0 : _GEN_3736; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3738 = 8'h1b == _T_174[7:0] ? 4'h0 : _GEN_3737; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3739 = 8'h1c == _T_174[7:0] ? 4'h6 : _GEN_3738; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3740 = 8'h1d == _T_174[7:0] ? 4'h3 : _GEN_3739; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3741 = 8'h1e == _T_174[7:0] ? 4'h0 : _GEN_3740; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3742 = 8'h1f == _T_174[7:0] ? 4'h0 : _GEN_3741; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3743 = 8'h20 == _T_174[7:0] ? 4'h0 : _GEN_3742; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3744 = 8'h21 == _T_174[7:0] ? 4'h3 : _GEN_3743; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3745 = 8'h22 == _T_174[7:0] ? 4'h6 : _GEN_3744; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3746 = 8'h23 == _T_174[7:0] ? 4'h0 : _GEN_3745; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3747 = 8'h24 == _T_174[7:0] ? 4'h0 : _GEN_3746; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3748 = 8'h25 == _T_174[7:0] ? 4'h0 : _GEN_3747; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3749 = 8'h26 == _T_174[7:0] ? 4'h0 : _GEN_3748; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3750 = 8'h27 == _T_174[7:0] ? 4'h0 : _GEN_3749; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3751 = 8'h28 == _T_174[7:0] ? 4'h0 : _GEN_3750; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3752 = 8'h29 == _T_174[7:0] ? 4'h0 : _GEN_3751; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3753 = 8'h2a == _T_174[7:0] ? 4'h0 : _GEN_3752; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3754 = 8'h2b == _T_174[7:0] ? 4'h0 : _GEN_3753; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3755 = 8'h2c == _T_174[7:0] ? 4'h0 : _GEN_3754; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3756 = 8'h2d == _T_174[7:0] ? 4'h0 : _GEN_3755; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3757 = 8'h2e == _T_174[7:0] ? 4'h0 : _GEN_3756; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3758 = 8'h2f == _T_174[7:0] ? 4'h0 : _GEN_3757; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3759 = 8'h30 == _T_174[7:0] ? 4'h6 : _GEN_3758; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3760 = 8'h31 == _T_174[7:0] ? 4'h3 : _GEN_3759; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3761 = 8'h32 == _T_174[7:0] ? 4'h0 : _GEN_3760; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3762 = 8'h33 == _T_174[7:0] ? 4'h1 : _GEN_3761; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3763 = 8'h34 == _T_174[7:0] ? 4'h1 : _GEN_3762; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3764 = 8'h35 == _T_174[7:0] ? 4'h0 : _GEN_3763; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3765 = 8'h36 == _T_174[7:0] ? 4'h0 : _GEN_3764; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3766 = 8'h37 == _T_174[7:0] ? 4'h0 : _GEN_3765; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3767 = 8'h38 == _T_174[7:0] ? 4'h6 : _GEN_3766; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3768 = 8'h39 == _T_174[7:0] ? 4'h0 : _GEN_3767; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3769 = 8'h3a == _T_174[7:0] ? 4'h0 : _GEN_3768; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3770 = 8'h3b == _T_174[7:0] ? 4'h0 : _GEN_3769; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3771 = 8'h3c == _T_174[7:0] ? 4'h0 : _GEN_3770; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3772 = 8'h3d == _T_174[7:0] ? 4'h0 : _GEN_3771; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3773 = 8'h3e == _T_174[7:0] ? 4'h0 : _GEN_3772; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3774 = 8'h3f == _T_174[7:0] ? 4'h0 : _GEN_3773; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3775 = 8'h40 == _T_174[7:0] ? 4'h0 : _GEN_3774; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3776 = 8'h41 == _T_174[7:0] ? 4'h0 : _GEN_3775; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3777 = 8'h42 == _T_174[7:0] ? 4'h0 : _GEN_3776; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3778 = 8'h43 == _T_174[7:0] ? 4'h0 : _GEN_3777; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3779 = 8'h44 == _T_174[7:0] ? 4'h3 : _GEN_3778; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3780 = 8'h45 == _T_174[7:0] ? 4'h6 : _GEN_3779; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3781 = 8'h46 == _T_174[7:0] ? 4'h9 : _GEN_3780; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3782 = 8'h47 == _T_174[7:0] ? 4'h0 : _GEN_3781; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3783 = 8'h48 == _T_174[7:0] ? 4'h0 : _GEN_3782; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3784 = 8'h49 == _T_174[7:0] ? 4'h0 : _GEN_3783; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3785 = 8'h4a == _T_174[7:0] ? 4'h1 : _GEN_3784; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3786 = 8'h4b == _T_174[7:0] ? 4'h0 : _GEN_3785; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3787 = 8'h4c == _T_174[7:0] ? 4'h0 : _GEN_3786; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3788 = 8'h4d == _T_174[7:0] ? 4'h0 : _GEN_3787; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3789 = 8'h4e == _T_174[7:0] ? 4'h6 : _GEN_3788; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3790 = 8'h4f == _T_174[7:0] ? 4'h0 : _GEN_3789; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3791 = 8'h50 == _T_174[7:0] ? 4'h0 : _GEN_3790; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3792 = 8'h51 == _T_174[7:0] ? 4'h0 : _GEN_3791; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3793 = 8'h52 == _T_174[7:0] ? 4'h0 : _GEN_3792; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3794 = 8'h53 == _T_174[7:0] ? 4'h0 : _GEN_3793; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3795 = 8'h54 == _T_174[7:0] ? 4'h0 : _GEN_3794; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3796 = 8'h55 == _T_174[7:0] ? 4'h0 : _GEN_3795; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3797 = 8'h56 == _T_174[7:0] ? 4'h0 : _GEN_3796; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3798 = 8'h57 == _T_174[7:0] ? 4'h0 : _GEN_3797; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3799 = 8'h58 == _T_174[7:0] ? 4'h0 : _GEN_3798; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3800 = 8'h59 == _T_174[7:0] ? 4'h6 : _GEN_3799; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3801 = 8'h5a == _T_174[7:0] ? 4'h3 : _GEN_3800; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3802 = 8'h5b == _T_174[7:0] ? 4'h0 : _GEN_3801; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3803 = 8'h5c == _T_174[7:0] ? 4'h0 : _GEN_3802; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3804 = 8'h5d == _T_174[7:0] ? 4'h0 : _GEN_3803; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3805 = 8'h5e == _T_174[7:0] ? 4'h7 : _GEN_3804; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3806 = 8'h5f == _T_174[7:0] ? 4'h0 : _GEN_3805; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3807 = 8'h60 == _T_174[7:0] ? 4'h0 : _GEN_3806; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3808 = 8'h61 == _T_174[7:0] ? 4'h1 : _GEN_3807; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3809 = 8'h62 == _T_174[7:0] ? 4'h0 : _GEN_3808; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3810 = 8'h63 == _T_174[7:0] ? 4'h6 : _GEN_3809; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3811 = 8'h64 == _T_174[7:0] ? 4'h0 : _GEN_3810; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3812 = 8'h65 == _T_174[7:0] ? 4'h0 : _GEN_3811; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3813 = 8'h66 == _T_174[7:0] ? 4'h0 : _GEN_3812; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3814 = 8'h67 == _T_174[7:0] ? 4'h0 : _GEN_3813; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3815 = 8'h68 == _T_174[7:0] ? 4'h0 : _GEN_3814; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3816 = 8'h69 == _T_174[7:0] ? 4'h0 : _GEN_3815; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3817 = 8'h6a == _T_174[7:0] ? 4'h0 : _GEN_3816; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3818 = 8'h6b == _T_174[7:0] ? 4'h0 : _GEN_3817; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3819 = 8'h6c == _T_174[7:0] ? 4'h0 : _GEN_3818; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3820 = 8'h6d == _T_174[7:0] ? 4'h0 : _GEN_3819; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3821 = 8'h6e == _T_174[7:0] ? 4'h6 : _GEN_3820; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3822 = 8'h6f == _T_174[7:0] ? 4'h0 : _GEN_3821; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3823 = 8'h70 == _T_174[7:0] ? 4'h0 : _GEN_3822; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3824 = 8'h71 == _T_174[7:0] ? 4'h0 : _GEN_3823; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3825 = 8'h72 == _T_174[7:0] ? 4'h3 : _GEN_3824; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3826 = 8'h73 == _T_174[7:0] ? 4'hc : _GEN_3825; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3827 = 8'h74 == _T_174[7:0] ? 4'h3 : _GEN_3826; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3828 = 8'h75 == _T_174[7:0] ? 4'h0 : _GEN_3827; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3829 = 8'h76 == _T_174[7:0] ? 4'h1 : _GEN_3828; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3830 = 8'h77 == _T_174[7:0] ? 4'h0 : _GEN_3829; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3831 = 8'h78 == _T_174[7:0] ? 4'h3 : _GEN_3830; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3832 = 8'h79 == _T_174[7:0] ? 4'h3 : _GEN_3831; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3833 = 8'h7a == _T_174[7:0] ? 4'h0 : _GEN_3832; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3834 = 8'h7b == _T_174[7:0] ? 4'h0 : _GEN_3833; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3835 = 8'h7c == _T_174[7:0] ? 4'h0 : _GEN_3834; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3836 = 8'h7d == _T_174[7:0] ? 4'h0 : _GEN_3835; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3837 = 8'h7e == _T_174[7:0] ? 4'h0 : _GEN_3836; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3838 = 8'h7f == _T_174[7:0] ? 4'h0 : _GEN_3837; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3839 = 8'h80 == _T_174[7:0] ? 4'h0 : _GEN_3838; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3840 = 8'h81 == _T_174[7:0] ? 4'h0 : _GEN_3839; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3841 = 8'h82 == _T_174[7:0] ? 4'h6 : _GEN_3840; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3842 = 8'h83 == _T_174[7:0] ? 4'h0 : _GEN_3841; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3843 = 8'h84 == _T_174[7:0] ? 4'h1 : _GEN_3842; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3844 = 8'h85 == _T_174[7:0] ? 4'h1 : _GEN_3843; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3845 = 8'h86 == _T_174[7:0] ? 4'ha : _GEN_3844; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3846 = 8'h87 == _T_174[7:0] ? 4'h4 : _GEN_3845; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3847 = 8'h88 == _T_174[7:0] ? 4'h1 : _GEN_3846; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3848 = 8'h89 == _T_174[7:0] ? 4'h4 : _GEN_3847; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3849 = 8'h8a == _T_174[7:0] ? 4'ha : _GEN_3848; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3850 = 8'h8b == _T_174[7:0] ? 4'h0 : _GEN_3849; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3851 = 8'h8c == _T_174[7:0] ? 4'h0 : _GEN_3850; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3852 = 8'h8d == _T_174[7:0] ? 4'h0 : _GEN_3851; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3853 = 8'h8e == _T_174[7:0] ? 4'h6 : _GEN_3852; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3854 = 8'h8f == _T_174[7:0] ? 4'h0 : _GEN_3853; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3855 = 8'h90 == _T_174[7:0] ? 4'h0 : _GEN_3854; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3856 = 8'h91 == _T_174[7:0] ? 4'h0 : _GEN_3855; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3857 = 8'h92 == _T_174[7:0] ? 4'h0 : _GEN_3856; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3858 = 8'h93 == _T_174[7:0] ? 4'h0 : _GEN_3857; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3859 = 8'h94 == _T_174[7:0] ? 4'h0 : _GEN_3858; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3860 = 8'h95 == _T_174[7:0] ? 4'h0 : _GEN_3859; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3861 = 8'h96 == _T_174[7:0] ? 4'h0 : _GEN_3860; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3862 = 8'h97 == _T_174[7:0] ? 4'h6 : _GEN_3861; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3863 = 8'h98 == _T_174[7:0] ? 4'h6 : _GEN_3862; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3864 = 8'h99 == _T_174[7:0] ? 4'h3 : _GEN_3863; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3865 = 8'h9a == _T_174[7:0] ? 4'h0 : _GEN_3864; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3866 = 8'h9b == _T_174[7:0] ? 4'ha : _GEN_3865; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3867 = 8'h9c == _T_174[7:0] ? 4'ha : _GEN_3866; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3868 = 8'h9d == _T_174[7:0] ? 4'h0 : _GEN_3867; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3869 = 8'h9e == _T_174[7:0] ? 4'ha : _GEN_3868; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3870 = 8'h9f == _T_174[7:0] ? 4'ha : _GEN_3869; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3871 = 8'ha0 == _T_174[7:0] ? 4'h0 : _GEN_3870; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3872 = 8'ha1 == _T_174[7:0] ? 4'h3 : _GEN_3871; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3873 = 8'ha2 == _T_174[7:0] ? 4'h6 : _GEN_3872; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3874 = 8'ha3 == _T_174[7:0] ? 4'h6 : _GEN_3873; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3875 = 8'ha4 == _T_174[7:0] ? 4'h0 : _GEN_3874; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3876 = 8'ha5 == _T_174[7:0] ? 4'h0 : _GEN_3875; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3877 = 8'ha6 == _T_174[7:0] ? 4'h0 : _GEN_3876; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3878 = 8'ha7 == _T_174[7:0] ? 4'h0 : _GEN_3877; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3879 = 8'ha8 == _T_174[7:0] ? 4'h0 : _GEN_3878; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3880 = 8'ha9 == _T_174[7:0] ? 4'h0 : _GEN_3879; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3881 = 8'haa == _T_174[7:0] ? 4'h0 : _GEN_3880; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3882 = 8'hab == _T_174[7:0] ? 4'h0 : _GEN_3881; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3883 = 8'hac == _T_174[7:0] ? 4'h6 : _GEN_3882; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3884 = 8'had == _T_174[7:0] ? 4'h0 : _GEN_3883; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3885 = 8'hae == _T_174[7:0] ? 4'h3 : _GEN_3884; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3886 = 8'haf == _T_174[7:0] ? 4'h9 : _GEN_3885; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3887 = 8'hb0 == _T_174[7:0] ? 4'h3 : _GEN_3886; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3888 = 8'hb1 == _T_174[7:0] ? 4'h0 : _GEN_3887; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3889 = 8'hb2 == _T_174[7:0] ? 4'h0 : _GEN_3888; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3890 = 8'hb3 == _T_174[7:0] ? 4'h0 : _GEN_3889; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3891 = 8'hb4 == _T_174[7:0] ? 4'h3 : _GEN_3890; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3892 = 8'hb5 == _T_174[7:0] ? 4'h9 : _GEN_3891; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3893 = 8'hb6 == _T_174[7:0] ? 4'h3 : _GEN_3892; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3894 = 8'hb7 == _T_174[7:0] ? 4'h0 : _GEN_3893; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3895 = 8'hb8 == _T_174[7:0] ? 4'h6 : _GEN_3894; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3896 = 8'hb9 == _T_174[7:0] ? 4'h0 : _GEN_3895; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3897 = 8'hba == _T_174[7:0] ? 4'h0 : _GEN_3896; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3898 = 8'hbb == _T_174[7:0] ? 4'h0 : _GEN_3897; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3899 = 8'hbc == _T_174[7:0] ? 4'h0 : _GEN_3898; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3900 = 8'hbd == _T_174[7:0] ? 4'h0 : _GEN_3899; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3901 = 8'hbe == _T_174[7:0] ? 4'h0 : _GEN_3900; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3902 = 8'hbf == _T_174[7:0] ? 4'h0 : _GEN_3901; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3903 = 8'hc0 == _T_174[7:0] ? 4'h0 : _GEN_3902; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3904 = 8'hc1 == _T_174[7:0] ? 4'h0 : _GEN_3903; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3905 = 8'hc2 == _T_174[7:0] ? 4'h7 : _GEN_3904; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3906 = 8'hc3 == _T_174[7:0] ? 4'h2 : _GEN_3905; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3907 = 8'hc4 == _T_174[7:0] ? 4'h0 : _GEN_3906; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3908 = 8'hc5 == _T_174[7:0] ? 4'h6 : _GEN_3907; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3909 = 8'hc6 == _T_174[7:0] ? 4'h9 : _GEN_3908; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3910 = 8'hc7 == _T_174[7:0] ? 4'h6 : _GEN_3909; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3911 = 8'hc8 == _T_174[7:0] ? 4'h9 : _GEN_3910; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3912 = 8'hc9 == _T_174[7:0] ? 4'h6 : _GEN_3911; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3913 = 8'hca == _T_174[7:0] ? 4'h0 : _GEN_3912; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3914 = 8'hcb == _T_174[7:0] ? 4'h2 : _GEN_3913; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3915 = 8'hcc == _T_174[7:0] ? 4'h7 : _GEN_3914; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3916 = 8'hcd == _T_174[7:0] ? 4'h0 : _GEN_3915; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3917 = 8'hce == _T_174[7:0] ? 4'h0 : _GEN_3916; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3918 = 8'hcf == _T_174[7:0] ? 4'h0 : _GEN_3917; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3919 = 8'hd0 == _T_174[7:0] ? 4'h0 : _GEN_3918; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3920 = 8'hd1 == _T_174[7:0] ? 4'h0 : _GEN_3919; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3921 = 8'hd2 == _T_174[7:0] ? 4'h0 : _GEN_3920; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3922 = 8'hd3 == _T_174[7:0] ? 4'h0 : _GEN_3921; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3923 = 8'hd4 == _T_174[7:0] ? 4'h0 : _GEN_3922; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3924 = 8'hd5 == _T_174[7:0] ? 4'h0 : _GEN_3923; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3925 = 8'hd6 == _T_174[7:0] ? 4'h0 : _GEN_3924; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3926 = 8'hd7 == _T_174[7:0] ? 4'h3 : _GEN_3925; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3927 = 8'hd8 == _T_174[7:0] ? 4'h3 : _GEN_3926; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3928 = 8'hd9 == _T_174[7:0] ? 4'h0 : _GEN_3927; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3929 = 8'hda == _T_174[7:0] ? 4'h9 : _GEN_3928; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3930 = 8'hdb == _T_174[7:0] ? 4'h3 : _GEN_3929; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3931 = 8'hdc == _T_174[7:0] ? 4'hc : _GEN_3930; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3932 = 8'hdd == _T_174[7:0] ? 4'h3 : _GEN_3931; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3933 = 8'hde == _T_174[7:0] ? 4'h9 : _GEN_3932; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3934 = 8'hdf == _T_174[7:0] ? 4'h0 : _GEN_3933; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3935 = 8'he0 == _T_174[7:0] ? 4'h3 : _GEN_3934; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3936 = 8'he1 == _T_174[7:0] ? 4'h3 : _GEN_3935; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3937 = 8'he2 == _T_174[7:0] ? 4'h0 : _GEN_3936; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3938 = 8'he3 == _T_174[7:0] ? 4'h0 : _GEN_3937; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3939 = 8'he4 == _T_174[7:0] ? 4'h0 : _GEN_3938; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3940 = 8'he5 == _T_174[7:0] ? 4'h0 : _GEN_3939; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3941 = 8'he6 == _T_174[7:0] ? 4'h0 : _GEN_3940; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3942 = 8'he7 == _T_174[7:0] ? 4'h0 : _GEN_3941; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3943 = 8'he8 == _T_174[7:0] ? 4'h0 : _GEN_3942; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3944 = 8'he9 == _T_174[7:0] ? 4'h0 : _GEN_3943; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3945 = 8'hea == _T_174[7:0] ? 4'h0 : _GEN_3944; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3946 = 8'heb == _T_174[7:0] ? 4'h0 : _GEN_3945; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3947 = 8'hec == _T_174[7:0] ? 4'h0 : _GEN_3946; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3948 = 8'hed == _T_174[7:0] ? 4'h0 : _GEN_3947; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3949 = 8'hee == _T_174[7:0] ? 4'h0 : _GEN_3948; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3950 = 8'hef == _T_174[7:0] ? 4'h0 : _GEN_3949; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3951 = 8'hf0 == _T_174[7:0] ? 4'h0 : _GEN_3950; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3952 = 8'hf1 == _T_174[7:0] ? 4'h0 : _GEN_3951; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3953 = 8'hf2 == _T_174[7:0] ? 4'h0 : _GEN_3952; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3954 = 8'hf3 == _T_174[7:0] ? 4'h0 : _GEN_3953; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3955 = 8'hf4 == _T_174[7:0] ? 4'h0 : _GEN_3954; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3956 = 8'hf5 == _T_174[7:0] ? 4'h0 : _GEN_3955; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3957 = 8'hf6 == _T_174[7:0] ? 4'h0 : _GEN_3956; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3958 = 8'hf7 == _T_174[7:0] ? 4'h0 : _GEN_3957; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3959 = 8'hf8 == _T_174[7:0] ? 4'h0 : _GEN_3958; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3960 = 8'hf9 == _T_174[7:0] ? 4'h0 : _GEN_3959; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3961 = 8'hfa == _T_174[7:0] ? 4'h0 : _GEN_3960; // @[Filter.scala 204:142]
  wire [3:0] _GEN_3962 = 8'hfb == _T_174[7:0] ? 4'h0 : _GEN_3961; // @[Filter.scala 204:142]
  wire [7:0] _T_188 = _GEN_3962 * 4'ha; // @[Filter.scala 204:142]
  wire [10:0] _GEN_11242 = {{3'd0}, _T_188}; // @[Filter.scala 204:109]
  wire [10:0] _T_190 = _T_183 + _GEN_11242; // @[Filter.scala 204:109]
  wire [10:0] _T_191 = _T_190 / 11'h64; // @[Filter.scala 204:150]
  wire  _T_193 = _T_164 >= 5'h15; // @[Filter.scala 207:31]
  wire  _T_197 = _T_171 >= 32'hc; // @[Filter.scala 207:63]
  wire  _T_198 = _T_193 | _T_197; // @[Filter.scala 207:58]
  wire [10:0] _GEN_4215 = io_SPI_distort ? _T_191 : {{7'd0}, _GEN_3458}; // @[Filter.scala 209:35]
  wire [10:0] _GEN_4216 = _T_198 ? 11'h0 : _GEN_4215; // @[Filter.scala 207:80]
  wire [10:0] _GEN_4469 = io_SPI_distort ? _T_191 : {{7'd0}, _GEN_3710}; // @[Filter.scala 209:35]
  wire [10:0] _GEN_4470 = _T_198 ? 11'h0 : _GEN_4469; // @[Filter.scala 207:80]
  wire [10:0] _GEN_4723 = io_SPI_distort ? _T_191 : {{7'd0}, _GEN_3962}; // @[Filter.scala 209:35]
  wire [10:0] _GEN_4724 = _T_198 ? 11'h0 : _GEN_4723; // @[Filter.scala 207:80]
  wire [31:0] _T_226 = pixelIndex + 32'h3; // @[Filter.scala 202:31]
  wire [31:0] _GEN_3 = _T_226 % 32'h15; // @[Filter.scala 202:38]
  wire [4:0] _T_227 = _GEN_3[4:0]; // @[Filter.scala 202:38]
  wire [4:0] _T_229 = _T_227 + _GEN_11210; // @[Filter.scala 202:53]
  wire [4:0] _T_231 = _T_229 - 5'h1; // @[Filter.scala 202:69]
  wire [31:0] _T_234 = _T_226 / 32'h15; // @[Filter.scala 203:38]
  wire [31:0] _T_236 = _T_234 + _GEN_11211; // @[Filter.scala 203:53]
  wire [31:0] _T_238 = _T_236 - 32'h1; // @[Filter.scala 203:69]
  wire [36:0] _T_239 = _T_238 * 32'h15; // @[Filter.scala 204:42]
  wire [36:0] _GEN_11248 = {{32'd0}, _T_231}; // @[Filter.scala 204:57]
  wire [36:0] _T_241 = _T_239 + _GEN_11248; // @[Filter.scala 204:57]
  wire [3:0] _GEN_4733 = 8'h8 == _T_241[7:0] ? 4'h1 : 4'h0; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4734 = 8'h9 == _T_241[7:0] ? 4'h2 : _GEN_4733; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4735 = 8'ha == _T_241[7:0] ? 4'h2 : _GEN_4734; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4736 = 8'hb == _T_241[7:0] ? 4'h2 : _GEN_4735; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4737 = 8'hc == _T_241[7:0] ? 4'h1 : _GEN_4736; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4738 = 8'hd == _T_241[7:0] ? 4'h0 : _GEN_4737; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4739 = 8'he == _T_241[7:0] ? 4'h0 : _GEN_4738; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4740 = 8'hf == _T_241[7:0] ? 4'h0 : _GEN_4739; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4741 = 8'h10 == _T_241[7:0] ? 4'h0 : _GEN_4740; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4742 = 8'h11 == _T_241[7:0] ? 4'h0 : _GEN_4741; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4743 = 8'h12 == _T_241[7:0] ? 4'h0 : _GEN_4742; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4744 = 8'h13 == _T_241[7:0] ? 4'h0 : _GEN_4743; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4745 = 8'h14 == _T_241[7:0] ? 4'h0 : _GEN_4744; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4746 = 8'h15 == _T_241[7:0] ? 4'h0 : _GEN_4745; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4747 = 8'h16 == _T_241[7:0] ? 4'h0 : _GEN_4746; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4748 = 8'h17 == _T_241[7:0] ? 4'h0 : _GEN_4747; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4749 = 8'h18 == _T_241[7:0] ? 4'h0 : _GEN_4748; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4750 = 8'h19 == _T_241[7:0] ? 4'h0 : _GEN_4749; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4751 = 8'h1a == _T_241[7:0] ? 4'h0 : _GEN_4750; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4752 = 8'h1b == _T_241[7:0] ? 4'h0 : _GEN_4751; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4753 = 8'h1c == _T_241[7:0] ? 4'h2 : _GEN_4752; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4754 = 8'h1d == _T_241[7:0] ? 4'h1 : _GEN_4753; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4755 = 8'h1e == _T_241[7:0] ? 4'h0 : _GEN_4754; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4756 = 8'h1f == _T_241[7:0] ? 4'h0 : _GEN_4755; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4757 = 8'h20 == _T_241[7:0] ? 4'h0 : _GEN_4756; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4758 = 8'h21 == _T_241[7:0] ? 4'h1 : _GEN_4757; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4759 = 8'h22 == _T_241[7:0] ? 4'h2 : _GEN_4758; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4760 = 8'h23 == _T_241[7:0] ? 4'h0 : _GEN_4759; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4761 = 8'h24 == _T_241[7:0] ? 4'h0 : _GEN_4760; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4762 = 8'h25 == _T_241[7:0] ? 4'h0 : _GEN_4761; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4763 = 8'h26 == _T_241[7:0] ? 4'h0 : _GEN_4762; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4764 = 8'h27 == _T_241[7:0] ? 4'h0 : _GEN_4763; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4765 = 8'h28 == _T_241[7:0] ? 4'h0 : _GEN_4764; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4766 = 8'h29 == _T_241[7:0] ? 4'h0 : _GEN_4765; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4767 = 8'h2a == _T_241[7:0] ? 4'h0 : _GEN_4766; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4768 = 8'h2b == _T_241[7:0] ? 4'h0 : _GEN_4767; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4769 = 8'h2c == _T_241[7:0] ? 4'h0 : _GEN_4768; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4770 = 8'h2d == _T_241[7:0] ? 4'h0 : _GEN_4769; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4771 = 8'h2e == _T_241[7:0] ? 4'h0 : _GEN_4770; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4772 = 8'h2f == _T_241[7:0] ? 4'h0 : _GEN_4771; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4773 = 8'h30 == _T_241[7:0] ? 4'h2 : _GEN_4772; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4774 = 8'h31 == _T_241[7:0] ? 4'h2 : _GEN_4773; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4775 = 8'h32 == _T_241[7:0] ? 4'h0 : _GEN_4774; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4776 = 8'h33 == _T_241[7:0] ? 4'h0 : _GEN_4775; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4777 = 8'h34 == _T_241[7:0] ? 4'h0 : _GEN_4776; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4778 = 8'h35 == _T_241[7:0] ? 4'h0 : _GEN_4777; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4779 = 8'h36 == _T_241[7:0] ? 4'h0 : _GEN_4778; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4780 = 8'h37 == _T_241[7:0] ? 4'h0 : _GEN_4779; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4781 = 8'h38 == _T_241[7:0] ? 4'h2 : _GEN_4780; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4782 = 8'h39 == _T_241[7:0] ? 4'h0 : _GEN_4781; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4783 = 8'h3a == _T_241[7:0] ? 4'h0 : _GEN_4782; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4784 = 8'h3b == _T_241[7:0] ? 4'h0 : _GEN_4783; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4785 = 8'h3c == _T_241[7:0] ? 4'h0 : _GEN_4784; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4786 = 8'h3d == _T_241[7:0] ? 4'h0 : _GEN_4785; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4787 = 8'h3e == _T_241[7:0] ? 4'h0 : _GEN_4786; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4788 = 8'h3f == _T_241[7:0] ? 4'h0 : _GEN_4787; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4789 = 8'h40 == _T_241[7:0] ? 4'h0 : _GEN_4788; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4790 = 8'h41 == _T_241[7:0] ? 4'h0 : _GEN_4789; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4791 = 8'h42 == _T_241[7:0] ? 4'h0 : _GEN_4790; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4792 = 8'h43 == _T_241[7:0] ? 4'h0 : _GEN_4791; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4793 = 8'h44 == _T_241[7:0] ? 4'h1 : _GEN_4792; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4794 = 8'h45 == _T_241[7:0] ? 4'h3 : _GEN_4793; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4795 = 8'h46 == _T_241[7:0] ? 4'h7 : _GEN_4794; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4796 = 8'h47 == _T_241[7:0] ? 4'h0 : _GEN_4795; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4797 = 8'h48 == _T_241[7:0] ? 4'h0 : _GEN_4796; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4798 = 8'h49 == _T_241[7:0] ? 4'h0 : _GEN_4797; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4799 = 8'h4a == _T_241[7:0] ? 4'h0 : _GEN_4798; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4800 = 8'h4b == _T_241[7:0] ? 4'h0 : _GEN_4799; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4801 = 8'h4c == _T_241[7:0] ? 4'h0 : _GEN_4800; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4802 = 8'h4d == _T_241[7:0] ? 4'h0 : _GEN_4801; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4803 = 8'h4e == _T_241[7:0] ? 4'h2 : _GEN_4802; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4804 = 8'h4f == _T_241[7:0] ? 4'h0 : _GEN_4803; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4805 = 8'h50 == _T_241[7:0] ? 4'h0 : _GEN_4804; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4806 = 8'h51 == _T_241[7:0] ? 4'h0 : _GEN_4805; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4807 = 8'h52 == _T_241[7:0] ? 4'h0 : _GEN_4806; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4808 = 8'h53 == _T_241[7:0] ? 4'h0 : _GEN_4807; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4809 = 8'h54 == _T_241[7:0] ? 4'h0 : _GEN_4808; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4810 = 8'h55 == _T_241[7:0] ? 4'h0 : _GEN_4809; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4811 = 8'h56 == _T_241[7:0] ? 4'h0 : _GEN_4810; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4812 = 8'h57 == _T_241[7:0] ? 4'h0 : _GEN_4811; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4813 = 8'h58 == _T_241[7:0] ? 4'h0 : _GEN_4812; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4814 = 8'h59 == _T_241[7:0] ? 4'h2 : _GEN_4813; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4815 = 8'h5a == _T_241[7:0] ? 4'h2 : _GEN_4814; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4816 = 8'h5b == _T_241[7:0] ? 4'h0 : _GEN_4815; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4817 = 8'h5c == _T_241[7:0] ? 4'h0 : _GEN_4816; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4818 = 8'h5d == _T_241[7:0] ? 4'h0 : _GEN_4817; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4819 = 8'h5e == _T_241[7:0] ? 4'h4 : _GEN_4818; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4820 = 8'h5f == _T_241[7:0] ? 4'h0 : _GEN_4819; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4821 = 8'h60 == _T_241[7:0] ? 4'h0 : _GEN_4820; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4822 = 8'h61 == _T_241[7:0] ? 4'h0 : _GEN_4821; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4823 = 8'h62 == _T_241[7:0] ? 4'h0 : _GEN_4822; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4824 = 8'h63 == _T_241[7:0] ? 4'h2 : _GEN_4823; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4825 = 8'h64 == _T_241[7:0] ? 4'h0 : _GEN_4824; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4826 = 8'h65 == _T_241[7:0] ? 4'h0 : _GEN_4825; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4827 = 8'h66 == _T_241[7:0] ? 4'h0 : _GEN_4826; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4828 = 8'h67 == _T_241[7:0] ? 4'h0 : _GEN_4827; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4829 = 8'h68 == _T_241[7:0] ? 4'h0 : _GEN_4828; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4830 = 8'h69 == _T_241[7:0] ? 4'h0 : _GEN_4829; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4831 = 8'h6a == _T_241[7:0] ? 4'h0 : _GEN_4830; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4832 = 8'h6b == _T_241[7:0] ? 4'h0 : _GEN_4831; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4833 = 8'h6c == _T_241[7:0] ? 4'h0 : _GEN_4832; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4834 = 8'h6d == _T_241[7:0] ? 4'h0 : _GEN_4833; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4835 = 8'h6e == _T_241[7:0] ? 4'h2 : _GEN_4834; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4836 = 8'h6f == _T_241[7:0] ? 4'h0 : _GEN_4835; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4837 = 8'h70 == _T_241[7:0] ? 4'h0 : _GEN_4836; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4838 = 8'h71 == _T_241[7:0] ? 4'h0 : _GEN_4837; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4839 = 8'h72 == _T_241[7:0] ? 4'h2 : _GEN_4838; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4840 = 8'h73 == _T_241[7:0] ? 4'h9 : _GEN_4839; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4841 = 8'h74 == _T_241[7:0] ? 4'h2 : _GEN_4840; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4842 = 8'h75 == _T_241[7:0] ? 4'h0 : _GEN_4841; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4843 = 8'h76 == _T_241[7:0] ? 4'h0 : _GEN_4842; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4844 = 8'h77 == _T_241[7:0] ? 4'h0 : _GEN_4843; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4845 = 8'h78 == _T_241[7:0] ? 4'h1 : _GEN_4844; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4846 = 8'h79 == _T_241[7:0] ? 4'h1 : _GEN_4845; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4847 = 8'h7a == _T_241[7:0] ? 4'h0 : _GEN_4846; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4848 = 8'h7b == _T_241[7:0] ? 4'h0 : _GEN_4847; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4849 = 8'h7c == _T_241[7:0] ? 4'h0 : _GEN_4848; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4850 = 8'h7d == _T_241[7:0] ? 4'h0 : _GEN_4849; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4851 = 8'h7e == _T_241[7:0] ? 4'h0 : _GEN_4850; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4852 = 8'h7f == _T_241[7:0] ? 4'h0 : _GEN_4851; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4853 = 8'h80 == _T_241[7:0] ? 4'h0 : _GEN_4852; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4854 = 8'h81 == _T_241[7:0] ? 4'h0 : _GEN_4853; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4855 = 8'h82 == _T_241[7:0] ? 4'h2 : _GEN_4854; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4856 = 8'h83 == _T_241[7:0] ? 4'h0 : _GEN_4855; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4857 = 8'h84 == _T_241[7:0] ? 4'h0 : _GEN_4856; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4858 = 8'h85 == _T_241[7:0] ? 4'h0 : _GEN_4857; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4859 = 8'h86 == _T_241[7:0] ? 4'h7 : _GEN_4858; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4860 = 8'h87 == _T_241[7:0] ? 4'h2 : _GEN_4859; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4861 = 8'h88 == _T_241[7:0] ? 4'h0 : _GEN_4860; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4862 = 8'h89 == _T_241[7:0] ? 4'h2 : _GEN_4861; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4863 = 8'h8a == _T_241[7:0] ? 4'h7 : _GEN_4862; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4864 = 8'h8b == _T_241[7:0] ? 4'h0 : _GEN_4863; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4865 = 8'h8c == _T_241[7:0] ? 4'h0 : _GEN_4864; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4866 = 8'h8d == _T_241[7:0] ? 4'h0 : _GEN_4865; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4867 = 8'h8e == _T_241[7:0] ? 4'h2 : _GEN_4866; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4868 = 8'h8f == _T_241[7:0] ? 4'h0 : _GEN_4867; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4869 = 8'h90 == _T_241[7:0] ? 4'h0 : _GEN_4868; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4870 = 8'h91 == _T_241[7:0] ? 4'h0 : _GEN_4869; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4871 = 8'h92 == _T_241[7:0] ? 4'h0 : _GEN_4870; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4872 = 8'h93 == _T_241[7:0] ? 4'h0 : _GEN_4871; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4873 = 8'h94 == _T_241[7:0] ? 4'h0 : _GEN_4872; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4874 = 8'h95 == _T_241[7:0] ? 4'h0 : _GEN_4873; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4875 = 8'h96 == _T_241[7:0] ? 4'h0 : _GEN_4874; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4876 = 8'h97 == _T_241[7:0] ? 4'h2 : _GEN_4875; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4877 = 8'h98 == _T_241[7:0] ? 4'h2 : _GEN_4876; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4878 = 8'h99 == _T_241[7:0] ? 4'h1 : _GEN_4877; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4879 = 8'h9a == _T_241[7:0] ? 4'h0 : _GEN_4878; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4880 = 8'h9b == _T_241[7:0] ? 4'h7 : _GEN_4879; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4881 = 8'h9c == _T_241[7:0] ? 4'h7 : _GEN_4880; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4882 = 8'h9d == _T_241[7:0] ? 4'h0 : _GEN_4881; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4883 = 8'h9e == _T_241[7:0] ? 4'h7 : _GEN_4882; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4884 = 8'h9f == _T_241[7:0] ? 4'h7 : _GEN_4883; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4885 = 8'ha0 == _T_241[7:0] ? 4'h0 : _GEN_4884; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4886 = 8'ha1 == _T_241[7:0] ? 4'h1 : _GEN_4885; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4887 = 8'ha2 == _T_241[7:0] ? 4'h2 : _GEN_4886; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4888 = 8'ha3 == _T_241[7:0] ? 4'h2 : _GEN_4887; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4889 = 8'ha4 == _T_241[7:0] ? 4'h0 : _GEN_4888; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4890 = 8'ha5 == _T_241[7:0] ? 4'h0 : _GEN_4889; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4891 = 8'ha6 == _T_241[7:0] ? 4'h0 : _GEN_4890; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4892 = 8'ha7 == _T_241[7:0] ? 4'h0 : _GEN_4891; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4893 = 8'ha8 == _T_241[7:0] ? 4'h0 : _GEN_4892; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4894 = 8'ha9 == _T_241[7:0] ? 4'h0 : _GEN_4893; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4895 = 8'haa == _T_241[7:0] ? 4'h0 : _GEN_4894; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4896 = 8'hab == _T_241[7:0] ? 4'h0 : _GEN_4895; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4897 = 8'hac == _T_241[7:0] ? 4'h2 : _GEN_4896; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4898 = 8'had == _T_241[7:0] ? 4'h0 : _GEN_4897; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4899 = 8'hae == _T_241[7:0] ? 4'h1 : _GEN_4898; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4900 = 8'haf == _T_241[7:0] ? 4'h3 : _GEN_4899; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4901 = 8'hb0 == _T_241[7:0] ? 4'h1 : _GEN_4900; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4902 = 8'hb1 == _T_241[7:0] ? 4'h0 : _GEN_4901; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4903 = 8'hb2 == _T_241[7:0] ? 4'h0 : _GEN_4902; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4904 = 8'hb3 == _T_241[7:0] ? 4'h0 : _GEN_4903; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4905 = 8'hb4 == _T_241[7:0] ? 4'h1 : _GEN_4904; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4906 = 8'hb5 == _T_241[7:0] ? 4'h3 : _GEN_4905; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4907 = 8'hb6 == _T_241[7:0] ? 4'h1 : _GEN_4906; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4908 = 8'hb7 == _T_241[7:0] ? 4'h0 : _GEN_4907; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4909 = 8'hb8 == _T_241[7:0] ? 4'h2 : _GEN_4908; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4910 = 8'hb9 == _T_241[7:0] ? 4'h0 : _GEN_4909; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4911 = 8'hba == _T_241[7:0] ? 4'h0 : _GEN_4910; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4912 = 8'hbb == _T_241[7:0] ? 4'h0 : _GEN_4911; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4913 = 8'hbc == _T_241[7:0] ? 4'h0 : _GEN_4912; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4914 = 8'hbd == _T_241[7:0] ? 4'h0 : _GEN_4913; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4915 = 8'hbe == _T_241[7:0] ? 4'h0 : _GEN_4914; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4916 = 8'hbf == _T_241[7:0] ? 4'h0 : _GEN_4915; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4917 = 8'hc0 == _T_241[7:0] ? 4'h0 : _GEN_4916; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4918 = 8'hc1 == _T_241[7:0] ? 4'h0 : _GEN_4917; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4919 = 8'hc2 == _T_241[7:0] ? 4'h3 : _GEN_4918; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4920 = 8'hc3 == _T_241[7:0] ? 4'h0 : _GEN_4919; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4921 = 8'hc4 == _T_241[7:0] ? 4'h0 : _GEN_4920; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4922 = 8'hc5 == _T_241[7:0] ? 4'h2 : _GEN_4921; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4923 = 8'hc6 == _T_241[7:0] ? 4'h3 : _GEN_4922; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4924 = 8'hc7 == _T_241[7:0] ? 4'h2 : _GEN_4923; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4925 = 8'hc8 == _T_241[7:0] ? 4'h3 : _GEN_4924; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4926 = 8'hc9 == _T_241[7:0] ? 4'h2 : _GEN_4925; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4927 = 8'hca == _T_241[7:0] ? 4'h0 : _GEN_4926; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4928 = 8'hcb == _T_241[7:0] ? 4'h0 : _GEN_4927; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4929 = 8'hcc == _T_241[7:0] ? 4'h3 : _GEN_4928; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4930 = 8'hcd == _T_241[7:0] ? 4'h0 : _GEN_4929; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4931 = 8'hce == _T_241[7:0] ? 4'h0 : _GEN_4930; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4932 = 8'hcf == _T_241[7:0] ? 4'h0 : _GEN_4931; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4933 = 8'hd0 == _T_241[7:0] ? 4'h0 : _GEN_4932; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4934 = 8'hd1 == _T_241[7:0] ? 4'h0 : _GEN_4933; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4935 = 8'hd2 == _T_241[7:0] ? 4'h0 : _GEN_4934; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4936 = 8'hd3 == _T_241[7:0] ? 4'h0 : _GEN_4935; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4937 = 8'hd4 == _T_241[7:0] ? 4'h0 : _GEN_4936; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4938 = 8'hd5 == _T_241[7:0] ? 4'h0 : _GEN_4937; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4939 = 8'hd6 == _T_241[7:0] ? 4'h0 : _GEN_4938; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4940 = 8'hd7 == _T_241[7:0] ? 4'h2 : _GEN_4939; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4941 = 8'hd8 == _T_241[7:0] ? 4'h2 : _GEN_4940; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4942 = 8'hd9 == _T_241[7:0] ? 4'h0 : _GEN_4941; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4943 = 8'hda == _T_241[7:0] ? 4'h7 : _GEN_4942; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4944 = 8'hdb == _T_241[7:0] ? 4'h1 : _GEN_4943; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4945 = 8'hdc == _T_241[7:0] ? 4'h4 : _GEN_4944; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4946 = 8'hdd == _T_241[7:0] ? 4'h1 : _GEN_4945; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4947 = 8'hde == _T_241[7:0] ? 4'h7 : _GEN_4946; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4948 = 8'hdf == _T_241[7:0] ? 4'h0 : _GEN_4947; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4949 = 8'he0 == _T_241[7:0] ? 4'h2 : _GEN_4948; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4950 = 8'he1 == _T_241[7:0] ? 4'h2 : _GEN_4949; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4951 = 8'he2 == _T_241[7:0] ? 4'h0 : _GEN_4950; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4952 = 8'he3 == _T_241[7:0] ? 4'h0 : _GEN_4951; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4953 = 8'he4 == _T_241[7:0] ? 4'h0 : _GEN_4952; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4954 = 8'he5 == _T_241[7:0] ? 4'h0 : _GEN_4953; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4955 = 8'he6 == _T_241[7:0] ? 4'h0 : _GEN_4954; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4956 = 8'he7 == _T_241[7:0] ? 4'h0 : _GEN_4955; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4957 = 8'he8 == _T_241[7:0] ? 4'h0 : _GEN_4956; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4958 = 8'he9 == _T_241[7:0] ? 4'h0 : _GEN_4957; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4959 = 8'hea == _T_241[7:0] ? 4'h0 : _GEN_4958; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4960 = 8'heb == _T_241[7:0] ? 4'h0 : _GEN_4959; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4961 = 8'hec == _T_241[7:0] ? 4'h0 : _GEN_4960; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4962 = 8'hed == _T_241[7:0] ? 4'h0 : _GEN_4961; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4963 = 8'hee == _T_241[7:0] ? 4'h0 : _GEN_4962; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4964 = 8'hef == _T_241[7:0] ? 4'h0 : _GEN_4963; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4965 = 8'hf0 == _T_241[7:0] ? 4'h0 : _GEN_4964; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4966 = 8'hf1 == _T_241[7:0] ? 4'h0 : _GEN_4965; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4967 = 8'hf2 == _T_241[7:0] ? 4'h0 : _GEN_4966; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4968 = 8'hf3 == _T_241[7:0] ? 4'h0 : _GEN_4967; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4969 = 8'hf4 == _T_241[7:0] ? 4'h0 : _GEN_4968; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4970 = 8'hf5 == _T_241[7:0] ? 4'h0 : _GEN_4969; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4971 = 8'hf6 == _T_241[7:0] ? 4'h0 : _GEN_4970; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4972 = 8'hf7 == _T_241[7:0] ? 4'h0 : _GEN_4971; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4973 = 8'hf8 == _T_241[7:0] ? 4'h0 : _GEN_4972; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4974 = 8'hf9 == _T_241[7:0] ? 4'h0 : _GEN_4973; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4975 = 8'hfa == _T_241[7:0] ? 4'h0 : _GEN_4974; // @[Filter.scala 204:62]
  wire [3:0] _GEN_4976 = 8'hfb == _T_241[7:0] ? 4'h0 : _GEN_4975; // @[Filter.scala 204:62]
  wire [4:0] _GEN_11249 = {{1'd0}, _GEN_4976}; // @[Filter.scala 204:62]
  wire [8:0] _T_243 = _GEN_11249 * 5'h14; // @[Filter.scala 204:62]
  wire [3:0] _GEN_5026 = 8'h31 == _T_241[7:0] ? 4'h3 : _GEN_4773; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5027 = 8'h32 == _T_241[7:0] ? 4'h3 : _GEN_5026; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5028 = 8'h33 == _T_241[7:0] ? 4'h6 : _GEN_5027; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5029 = 8'h34 == _T_241[7:0] ? 4'h6 : _GEN_5028; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5030 = 8'h35 == _T_241[7:0] ? 4'h0 : _GEN_5029; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5031 = 8'h36 == _T_241[7:0] ? 4'h0 : _GEN_5030; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5032 = 8'h37 == _T_241[7:0] ? 4'h0 : _GEN_5031; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5033 = 8'h38 == _T_241[7:0] ? 4'h2 : _GEN_5032; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5034 = 8'h39 == _T_241[7:0] ? 4'h0 : _GEN_5033; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5035 = 8'h3a == _T_241[7:0] ? 4'h0 : _GEN_5034; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5036 = 8'h3b == _T_241[7:0] ? 4'h0 : _GEN_5035; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5037 = 8'h3c == _T_241[7:0] ? 4'h0 : _GEN_5036; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5038 = 8'h3d == _T_241[7:0] ? 4'h0 : _GEN_5037; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5039 = 8'h3e == _T_241[7:0] ? 4'h0 : _GEN_5038; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5040 = 8'h3f == _T_241[7:0] ? 4'h0 : _GEN_5039; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5041 = 8'h40 == _T_241[7:0] ? 4'h0 : _GEN_5040; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5042 = 8'h41 == _T_241[7:0] ? 4'h0 : _GEN_5041; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5043 = 8'h42 == _T_241[7:0] ? 4'h0 : _GEN_5042; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5044 = 8'h43 == _T_241[7:0] ? 4'h0 : _GEN_5043; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5045 = 8'h44 == _T_241[7:0] ? 4'h1 : _GEN_5044; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5046 = 8'h45 == _T_241[7:0] ? 4'h4 : _GEN_5045; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5047 = 8'h46 == _T_241[7:0] ? 4'hb : _GEN_5046; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5048 = 8'h47 == _T_241[7:0] ? 4'h0 : _GEN_5047; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5049 = 8'h48 == _T_241[7:0] ? 4'h0 : _GEN_5048; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5050 = 8'h49 == _T_241[7:0] ? 4'h0 : _GEN_5049; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5051 = 8'h4a == _T_241[7:0] ? 4'h6 : _GEN_5050; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5052 = 8'h4b == _T_241[7:0] ? 4'h0 : _GEN_5051; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5053 = 8'h4c == _T_241[7:0] ? 4'h3 : _GEN_5052; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5054 = 8'h4d == _T_241[7:0] ? 4'h3 : _GEN_5053; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5055 = 8'h4e == _T_241[7:0] ? 4'h2 : _GEN_5054; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5056 = 8'h4f == _T_241[7:0] ? 4'h0 : _GEN_5055; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5057 = 8'h50 == _T_241[7:0] ? 4'h0 : _GEN_5056; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5058 = 8'h51 == _T_241[7:0] ? 4'h0 : _GEN_5057; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5059 = 8'h52 == _T_241[7:0] ? 4'h0 : _GEN_5058; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5060 = 8'h53 == _T_241[7:0] ? 4'h0 : _GEN_5059; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5061 = 8'h54 == _T_241[7:0] ? 4'h0 : _GEN_5060; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5062 = 8'h55 == _T_241[7:0] ? 4'h0 : _GEN_5061; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5063 = 8'h56 == _T_241[7:0] ? 4'h0 : _GEN_5062; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5064 = 8'h57 == _T_241[7:0] ? 4'h0 : _GEN_5063; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5065 = 8'h58 == _T_241[7:0] ? 4'h0 : _GEN_5064; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5066 = 8'h59 == _T_241[7:0] ? 4'h2 : _GEN_5065; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5067 = 8'h5a == _T_241[7:0] ? 4'h3 : _GEN_5066; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5068 = 8'h5b == _T_241[7:0] ? 4'h0 : _GEN_5067; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5069 = 8'h5c == _T_241[7:0] ? 4'h0 : _GEN_5068; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5070 = 8'h5d == _T_241[7:0] ? 4'h3 : _GEN_5069; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5071 = 8'h5e == _T_241[7:0] ? 4'hd : _GEN_5070; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5072 = 8'h5f == _T_241[7:0] ? 4'h3 : _GEN_5071; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5073 = 8'h60 == _T_241[7:0] ? 4'h0 : _GEN_5072; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5074 = 8'h61 == _T_241[7:0] ? 4'h6 : _GEN_5073; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5075 = 8'h62 == _T_241[7:0] ? 4'h0 : _GEN_5074; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5076 = 8'h63 == _T_241[7:0] ? 4'h2 : _GEN_5075; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5077 = 8'h64 == _T_241[7:0] ? 4'h0 : _GEN_5076; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5078 = 8'h65 == _T_241[7:0] ? 4'h0 : _GEN_5077; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5079 = 8'h66 == _T_241[7:0] ? 4'h0 : _GEN_5078; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5080 = 8'h67 == _T_241[7:0] ? 4'h0 : _GEN_5079; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5081 = 8'h68 == _T_241[7:0] ? 4'h0 : _GEN_5080; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5082 = 8'h69 == _T_241[7:0] ? 4'h0 : _GEN_5081; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5083 = 8'h6a == _T_241[7:0] ? 4'h0 : _GEN_5082; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5084 = 8'h6b == _T_241[7:0] ? 4'h0 : _GEN_5083; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5085 = 8'h6c == _T_241[7:0] ? 4'h0 : _GEN_5084; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5086 = 8'h6d == _T_241[7:0] ? 4'h0 : _GEN_5085; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5087 = 8'h6e == _T_241[7:0] ? 4'h2 : _GEN_5086; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5088 = 8'h6f == _T_241[7:0] ? 4'h0 : _GEN_5087; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5089 = 8'h70 == _T_241[7:0] ? 4'h0 : _GEN_5088; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5090 = 8'h71 == _T_241[7:0] ? 4'h0 : _GEN_5089; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5091 = 8'h72 == _T_241[7:0] ? 4'h6 : _GEN_5090; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5092 = 8'h73 == _T_241[7:0] ? 4'he : _GEN_5091; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5093 = 8'h74 == _T_241[7:0] ? 4'h6 : _GEN_5092; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5094 = 8'h75 == _T_241[7:0] ? 4'h0 : _GEN_5093; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5095 = 8'h76 == _T_241[7:0] ? 4'h6 : _GEN_5094; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5096 = 8'h77 == _T_241[7:0] ? 4'h3 : _GEN_5095; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5097 = 8'h78 == _T_241[7:0] ? 4'h4 : _GEN_5096; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5098 = 8'h79 == _T_241[7:0] ? 4'h1 : _GEN_5097; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5099 = 8'h7a == _T_241[7:0] ? 4'h0 : _GEN_5098; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5100 = 8'h7b == _T_241[7:0] ? 4'h0 : _GEN_5099; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5101 = 8'h7c == _T_241[7:0] ? 4'h0 : _GEN_5100; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5102 = 8'h7d == _T_241[7:0] ? 4'h0 : _GEN_5101; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5103 = 8'h7e == _T_241[7:0] ? 4'h0 : _GEN_5102; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5104 = 8'h7f == _T_241[7:0] ? 4'h0 : _GEN_5103; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5105 = 8'h80 == _T_241[7:0] ? 4'h0 : _GEN_5104; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5106 = 8'h81 == _T_241[7:0] ? 4'h0 : _GEN_5105; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5107 = 8'h82 == _T_241[7:0] ? 4'h2 : _GEN_5106; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5108 = 8'h83 == _T_241[7:0] ? 4'h3 : _GEN_5107; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5109 = 8'h84 == _T_241[7:0] ? 4'h6 : _GEN_5108; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5110 = 8'h85 == _T_241[7:0] ? 4'h6 : _GEN_5109; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5111 = 8'h86 == _T_241[7:0] ? 4'he : _GEN_5110; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5112 = 8'h87 == _T_241[7:0] ? 4'ha : _GEN_5111; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5113 = 8'h88 == _T_241[7:0] ? 4'h6 : _GEN_5112; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5114 = 8'h89 == _T_241[7:0] ? 4'ha : _GEN_5113; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5115 = 8'h8a == _T_241[7:0] ? 4'he : _GEN_5114; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5116 = 8'h8b == _T_241[7:0] ? 4'h3 : _GEN_5115; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5117 = 8'h8c == _T_241[7:0] ? 4'h3 : _GEN_5116; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5118 = 8'h8d == _T_241[7:0] ? 4'h0 : _GEN_5117; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5119 = 8'h8e == _T_241[7:0] ? 4'h2 : _GEN_5118; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5120 = 8'h8f == _T_241[7:0] ? 4'h0 : _GEN_5119; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5121 = 8'h90 == _T_241[7:0] ? 4'h0 : _GEN_5120; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5122 = 8'h91 == _T_241[7:0] ? 4'h0 : _GEN_5121; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5123 = 8'h92 == _T_241[7:0] ? 4'h0 : _GEN_5122; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5124 = 8'h93 == _T_241[7:0] ? 4'h0 : _GEN_5123; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5125 = 8'h94 == _T_241[7:0] ? 4'h0 : _GEN_5124; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5126 = 8'h95 == _T_241[7:0] ? 4'h0 : _GEN_5125; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5127 = 8'h96 == _T_241[7:0] ? 4'h0 : _GEN_5126; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5128 = 8'h97 == _T_241[7:0] ? 4'h2 : _GEN_5127; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5129 = 8'h98 == _T_241[7:0] ? 4'h2 : _GEN_5128; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5130 = 8'h99 == _T_241[7:0] ? 4'h1 : _GEN_5129; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5131 = 8'h9a == _T_241[7:0] ? 4'h3 : _GEN_5130; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5132 = 8'h9b == _T_241[7:0] ? 4'he : _GEN_5131; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5133 = 8'h9c == _T_241[7:0] ? 4'he : _GEN_5132; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5134 = 8'h9d == _T_241[7:0] ? 4'h0 : _GEN_5133; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5135 = 8'h9e == _T_241[7:0] ? 4'he : _GEN_5134; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5136 = 8'h9f == _T_241[7:0] ? 4'he : _GEN_5135; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5137 = 8'ha0 == _T_241[7:0] ? 4'h3 : _GEN_5136; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5138 = 8'ha1 == _T_241[7:0] ? 4'h1 : _GEN_5137; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5139 = 8'ha2 == _T_241[7:0] ? 4'h2 : _GEN_5138; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5140 = 8'ha3 == _T_241[7:0] ? 4'h2 : _GEN_5139; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5141 = 8'ha4 == _T_241[7:0] ? 4'h0 : _GEN_5140; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5142 = 8'ha5 == _T_241[7:0] ? 4'h0 : _GEN_5141; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5143 = 8'ha6 == _T_241[7:0] ? 4'h0 : _GEN_5142; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5144 = 8'ha7 == _T_241[7:0] ? 4'h0 : _GEN_5143; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5145 = 8'ha8 == _T_241[7:0] ? 4'h0 : _GEN_5144; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5146 = 8'ha9 == _T_241[7:0] ? 4'h0 : _GEN_5145; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5147 = 8'haa == _T_241[7:0] ? 4'h0 : _GEN_5146; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5148 = 8'hab == _T_241[7:0] ? 4'h0 : _GEN_5147; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5149 = 8'hac == _T_241[7:0] ? 4'h2 : _GEN_5148; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5150 = 8'had == _T_241[7:0] ? 4'h3 : _GEN_5149; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5151 = 8'hae == _T_241[7:0] ? 4'h4 : _GEN_5150; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5152 = 8'haf == _T_241[7:0] ? 4'h3 : _GEN_5151; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5153 = 8'hb0 == _T_241[7:0] ? 4'h4 : _GEN_5152; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5154 = 8'hb1 == _T_241[7:0] ? 4'h3 : _GEN_5153; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5155 = 8'hb2 == _T_241[7:0] ? 4'h0 : _GEN_5154; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5156 = 8'hb3 == _T_241[7:0] ? 4'h3 : _GEN_5155; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5157 = 8'hb4 == _T_241[7:0] ? 4'h4 : _GEN_5156; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5158 = 8'hb5 == _T_241[7:0] ? 4'h3 : _GEN_5157; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5159 = 8'hb6 == _T_241[7:0] ? 4'h4 : _GEN_5158; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5160 = 8'hb7 == _T_241[7:0] ? 4'h3 : _GEN_5159; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5161 = 8'hb8 == _T_241[7:0] ? 4'h2 : _GEN_5160; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5162 = 8'hb9 == _T_241[7:0] ? 4'h0 : _GEN_5161; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5163 = 8'hba == _T_241[7:0] ? 4'h0 : _GEN_5162; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5164 = 8'hbb == _T_241[7:0] ? 4'h0 : _GEN_5163; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5165 = 8'hbc == _T_241[7:0] ? 4'h0 : _GEN_5164; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5166 = 8'hbd == _T_241[7:0] ? 4'h0 : _GEN_5165; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5167 = 8'hbe == _T_241[7:0] ? 4'h0 : _GEN_5166; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5168 = 8'hbf == _T_241[7:0] ? 4'h0 : _GEN_5167; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5169 = 8'hc0 == _T_241[7:0] ? 4'h0 : _GEN_5168; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5170 = 8'hc1 == _T_241[7:0] ? 4'h0 : _GEN_5169; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5171 = 8'hc2 == _T_241[7:0] ? 4'h8 : _GEN_5170; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5172 = 8'hc3 == _T_241[7:0] ? 4'hc : _GEN_5171; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5173 = 8'hc4 == _T_241[7:0] ? 4'h0 : _GEN_5172; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5174 = 8'hc5 == _T_241[7:0] ? 4'h2 : _GEN_5173; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5175 = 8'hc6 == _T_241[7:0] ? 4'h3 : _GEN_5174; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5176 = 8'hc7 == _T_241[7:0] ? 4'h2 : _GEN_5175; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5177 = 8'hc8 == _T_241[7:0] ? 4'h3 : _GEN_5176; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5178 = 8'hc9 == _T_241[7:0] ? 4'h2 : _GEN_5177; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5179 = 8'hca == _T_241[7:0] ? 4'h0 : _GEN_5178; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5180 = 8'hcb == _T_241[7:0] ? 4'hc : _GEN_5179; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5181 = 8'hcc == _T_241[7:0] ? 4'h8 : _GEN_5180; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5182 = 8'hcd == _T_241[7:0] ? 4'h0 : _GEN_5181; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5183 = 8'hce == _T_241[7:0] ? 4'h0 : _GEN_5182; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5184 = 8'hcf == _T_241[7:0] ? 4'h0 : _GEN_5183; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5185 = 8'hd0 == _T_241[7:0] ? 4'h0 : _GEN_5184; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5186 = 8'hd1 == _T_241[7:0] ? 4'h0 : _GEN_5185; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5187 = 8'hd2 == _T_241[7:0] ? 4'h0 : _GEN_5186; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5188 = 8'hd3 == _T_241[7:0] ? 4'h0 : _GEN_5187; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5189 = 8'hd4 == _T_241[7:0] ? 4'h0 : _GEN_5188; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5190 = 8'hd5 == _T_241[7:0] ? 4'h0 : _GEN_5189; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5191 = 8'hd6 == _T_241[7:0] ? 4'h0 : _GEN_5190; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5192 = 8'hd7 == _T_241[7:0] ? 4'h3 : _GEN_5191; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5193 = 8'hd8 == _T_241[7:0] ? 4'h6 : _GEN_5192; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5194 = 8'hd9 == _T_241[7:0] ? 4'h0 : _GEN_5193; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5195 = 8'hda == _T_241[7:0] ? 4'hb : _GEN_5194; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5196 = 8'hdb == _T_241[7:0] ? 4'h1 : _GEN_5195; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5197 = 8'hdc == _T_241[7:0] ? 4'h4 : _GEN_5196; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5198 = 8'hdd == _T_241[7:0] ? 4'h1 : _GEN_5197; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5199 = 8'hde == _T_241[7:0] ? 4'hb : _GEN_5198; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5200 = 8'hdf == _T_241[7:0] ? 4'h0 : _GEN_5199; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5201 = 8'he0 == _T_241[7:0] ? 4'h6 : _GEN_5200; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5202 = 8'he1 == _T_241[7:0] ? 4'h3 : _GEN_5201; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5203 = 8'he2 == _T_241[7:0] ? 4'h0 : _GEN_5202; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5204 = 8'he3 == _T_241[7:0] ? 4'h0 : _GEN_5203; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5205 = 8'he4 == _T_241[7:0] ? 4'h0 : _GEN_5204; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5206 = 8'he5 == _T_241[7:0] ? 4'h0 : _GEN_5205; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5207 = 8'he6 == _T_241[7:0] ? 4'h0 : _GEN_5206; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5208 = 8'he7 == _T_241[7:0] ? 4'h0 : _GEN_5207; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5209 = 8'he8 == _T_241[7:0] ? 4'h0 : _GEN_5208; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5210 = 8'he9 == _T_241[7:0] ? 4'h0 : _GEN_5209; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5211 = 8'hea == _T_241[7:0] ? 4'h0 : _GEN_5210; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5212 = 8'heb == _T_241[7:0] ? 4'h0 : _GEN_5211; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5213 = 8'hec == _T_241[7:0] ? 4'h0 : _GEN_5212; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5214 = 8'hed == _T_241[7:0] ? 4'h0 : _GEN_5213; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5215 = 8'hee == _T_241[7:0] ? 4'h0 : _GEN_5214; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5216 = 8'hef == _T_241[7:0] ? 4'h0 : _GEN_5215; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5217 = 8'hf0 == _T_241[7:0] ? 4'h0 : _GEN_5216; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5218 = 8'hf1 == _T_241[7:0] ? 4'h0 : _GEN_5217; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5219 = 8'hf2 == _T_241[7:0] ? 4'h0 : _GEN_5218; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5220 = 8'hf3 == _T_241[7:0] ? 4'h0 : _GEN_5219; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5221 = 8'hf4 == _T_241[7:0] ? 4'h0 : _GEN_5220; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5222 = 8'hf5 == _T_241[7:0] ? 4'h0 : _GEN_5221; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5223 = 8'hf6 == _T_241[7:0] ? 4'h0 : _GEN_5222; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5224 = 8'hf7 == _T_241[7:0] ? 4'h0 : _GEN_5223; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5225 = 8'hf8 == _T_241[7:0] ? 4'h0 : _GEN_5224; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5226 = 8'hf9 == _T_241[7:0] ? 4'h0 : _GEN_5225; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5227 = 8'hfa == _T_241[7:0] ? 4'h0 : _GEN_5226; // @[Filter.scala 204:102]
  wire [3:0] _GEN_5228 = 8'hfb == _T_241[7:0] ? 4'h0 : _GEN_5227; // @[Filter.scala 204:102]
  wire [6:0] _GEN_11251 = {{3'd0}, _GEN_5228}; // @[Filter.scala 204:102]
  wire [10:0] _T_248 = _GEN_11251 * 7'h46; // @[Filter.scala 204:102]
  wire [10:0] _GEN_11252 = {{2'd0}, _T_243}; // @[Filter.scala 204:69]
  wire [10:0] _T_250 = _GEN_11252 + _T_248; // @[Filter.scala 204:69]
  wire [3:0] _GEN_5237 = 8'h8 == _T_241[7:0] ? 4'h3 : 4'h0; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5238 = 8'h9 == _T_241[7:0] ? 4'h6 : _GEN_5237; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5239 = 8'ha == _T_241[7:0] ? 4'h6 : _GEN_5238; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5240 = 8'hb == _T_241[7:0] ? 4'h6 : _GEN_5239; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5241 = 8'hc == _T_241[7:0] ? 4'h3 : _GEN_5240; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5242 = 8'hd == _T_241[7:0] ? 4'h0 : _GEN_5241; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5243 = 8'he == _T_241[7:0] ? 4'h0 : _GEN_5242; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5244 = 8'hf == _T_241[7:0] ? 4'h0 : _GEN_5243; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5245 = 8'h10 == _T_241[7:0] ? 4'h0 : _GEN_5244; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5246 = 8'h11 == _T_241[7:0] ? 4'h0 : _GEN_5245; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5247 = 8'h12 == _T_241[7:0] ? 4'h0 : _GEN_5246; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5248 = 8'h13 == _T_241[7:0] ? 4'h0 : _GEN_5247; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5249 = 8'h14 == _T_241[7:0] ? 4'h0 : _GEN_5248; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5250 = 8'h15 == _T_241[7:0] ? 4'h0 : _GEN_5249; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5251 = 8'h16 == _T_241[7:0] ? 4'h0 : _GEN_5250; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5252 = 8'h17 == _T_241[7:0] ? 4'h0 : _GEN_5251; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5253 = 8'h18 == _T_241[7:0] ? 4'h0 : _GEN_5252; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5254 = 8'h19 == _T_241[7:0] ? 4'h0 : _GEN_5253; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5255 = 8'h1a == _T_241[7:0] ? 4'h0 : _GEN_5254; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5256 = 8'h1b == _T_241[7:0] ? 4'h0 : _GEN_5255; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5257 = 8'h1c == _T_241[7:0] ? 4'h6 : _GEN_5256; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5258 = 8'h1d == _T_241[7:0] ? 4'h3 : _GEN_5257; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5259 = 8'h1e == _T_241[7:0] ? 4'h0 : _GEN_5258; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5260 = 8'h1f == _T_241[7:0] ? 4'h0 : _GEN_5259; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5261 = 8'h20 == _T_241[7:0] ? 4'h0 : _GEN_5260; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5262 = 8'h21 == _T_241[7:0] ? 4'h3 : _GEN_5261; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5263 = 8'h22 == _T_241[7:0] ? 4'h6 : _GEN_5262; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5264 = 8'h23 == _T_241[7:0] ? 4'h0 : _GEN_5263; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5265 = 8'h24 == _T_241[7:0] ? 4'h0 : _GEN_5264; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5266 = 8'h25 == _T_241[7:0] ? 4'h0 : _GEN_5265; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5267 = 8'h26 == _T_241[7:0] ? 4'h0 : _GEN_5266; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5268 = 8'h27 == _T_241[7:0] ? 4'h0 : _GEN_5267; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5269 = 8'h28 == _T_241[7:0] ? 4'h0 : _GEN_5268; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5270 = 8'h29 == _T_241[7:0] ? 4'h0 : _GEN_5269; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5271 = 8'h2a == _T_241[7:0] ? 4'h0 : _GEN_5270; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5272 = 8'h2b == _T_241[7:0] ? 4'h0 : _GEN_5271; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5273 = 8'h2c == _T_241[7:0] ? 4'h0 : _GEN_5272; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5274 = 8'h2d == _T_241[7:0] ? 4'h0 : _GEN_5273; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5275 = 8'h2e == _T_241[7:0] ? 4'h0 : _GEN_5274; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5276 = 8'h2f == _T_241[7:0] ? 4'h0 : _GEN_5275; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5277 = 8'h30 == _T_241[7:0] ? 4'h6 : _GEN_5276; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5278 = 8'h31 == _T_241[7:0] ? 4'h3 : _GEN_5277; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5279 = 8'h32 == _T_241[7:0] ? 4'h0 : _GEN_5278; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5280 = 8'h33 == _T_241[7:0] ? 4'h1 : _GEN_5279; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5281 = 8'h34 == _T_241[7:0] ? 4'h1 : _GEN_5280; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5282 = 8'h35 == _T_241[7:0] ? 4'h0 : _GEN_5281; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5283 = 8'h36 == _T_241[7:0] ? 4'h0 : _GEN_5282; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5284 = 8'h37 == _T_241[7:0] ? 4'h0 : _GEN_5283; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5285 = 8'h38 == _T_241[7:0] ? 4'h6 : _GEN_5284; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5286 = 8'h39 == _T_241[7:0] ? 4'h0 : _GEN_5285; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5287 = 8'h3a == _T_241[7:0] ? 4'h0 : _GEN_5286; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5288 = 8'h3b == _T_241[7:0] ? 4'h0 : _GEN_5287; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5289 = 8'h3c == _T_241[7:0] ? 4'h0 : _GEN_5288; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5290 = 8'h3d == _T_241[7:0] ? 4'h0 : _GEN_5289; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5291 = 8'h3e == _T_241[7:0] ? 4'h0 : _GEN_5290; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5292 = 8'h3f == _T_241[7:0] ? 4'h0 : _GEN_5291; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5293 = 8'h40 == _T_241[7:0] ? 4'h0 : _GEN_5292; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5294 = 8'h41 == _T_241[7:0] ? 4'h0 : _GEN_5293; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5295 = 8'h42 == _T_241[7:0] ? 4'h0 : _GEN_5294; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5296 = 8'h43 == _T_241[7:0] ? 4'h0 : _GEN_5295; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5297 = 8'h44 == _T_241[7:0] ? 4'h3 : _GEN_5296; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5298 = 8'h45 == _T_241[7:0] ? 4'h6 : _GEN_5297; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5299 = 8'h46 == _T_241[7:0] ? 4'h9 : _GEN_5298; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5300 = 8'h47 == _T_241[7:0] ? 4'h0 : _GEN_5299; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5301 = 8'h48 == _T_241[7:0] ? 4'h0 : _GEN_5300; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5302 = 8'h49 == _T_241[7:0] ? 4'h0 : _GEN_5301; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5303 = 8'h4a == _T_241[7:0] ? 4'h1 : _GEN_5302; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5304 = 8'h4b == _T_241[7:0] ? 4'h0 : _GEN_5303; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5305 = 8'h4c == _T_241[7:0] ? 4'h0 : _GEN_5304; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5306 = 8'h4d == _T_241[7:0] ? 4'h0 : _GEN_5305; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5307 = 8'h4e == _T_241[7:0] ? 4'h6 : _GEN_5306; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5308 = 8'h4f == _T_241[7:0] ? 4'h0 : _GEN_5307; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5309 = 8'h50 == _T_241[7:0] ? 4'h0 : _GEN_5308; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5310 = 8'h51 == _T_241[7:0] ? 4'h0 : _GEN_5309; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5311 = 8'h52 == _T_241[7:0] ? 4'h0 : _GEN_5310; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5312 = 8'h53 == _T_241[7:0] ? 4'h0 : _GEN_5311; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5313 = 8'h54 == _T_241[7:0] ? 4'h0 : _GEN_5312; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5314 = 8'h55 == _T_241[7:0] ? 4'h0 : _GEN_5313; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5315 = 8'h56 == _T_241[7:0] ? 4'h0 : _GEN_5314; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5316 = 8'h57 == _T_241[7:0] ? 4'h0 : _GEN_5315; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5317 = 8'h58 == _T_241[7:0] ? 4'h0 : _GEN_5316; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5318 = 8'h59 == _T_241[7:0] ? 4'h6 : _GEN_5317; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5319 = 8'h5a == _T_241[7:0] ? 4'h3 : _GEN_5318; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5320 = 8'h5b == _T_241[7:0] ? 4'h0 : _GEN_5319; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5321 = 8'h5c == _T_241[7:0] ? 4'h0 : _GEN_5320; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5322 = 8'h5d == _T_241[7:0] ? 4'h0 : _GEN_5321; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5323 = 8'h5e == _T_241[7:0] ? 4'h7 : _GEN_5322; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5324 = 8'h5f == _T_241[7:0] ? 4'h0 : _GEN_5323; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5325 = 8'h60 == _T_241[7:0] ? 4'h0 : _GEN_5324; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5326 = 8'h61 == _T_241[7:0] ? 4'h1 : _GEN_5325; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5327 = 8'h62 == _T_241[7:0] ? 4'h0 : _GEN_5326; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5328 = 8'h63 == _T_241[7:0] ? 4'h6 : _GEN_5327; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5329 = 8'h64 == _T_241[7:0] ? 4'h0 : _GEN_5328; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5330 = 8'h65 == _T_241[7:0] ? 4'h0 : _GEN_5329; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5331 = 8'h66 == _T_241[7:0] ? 4'h0 : _GEN_5330; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5332 = 8'h67 == _T_241[7:0] ? 4'h0 : _GEN_5331; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5333 = 8'h68 == _T_241[7:0] ? 4'h0 : _GEN_5332; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5334 = 8'h69 == _T_241[7:0] ? 4'h0 : _GEN_5333; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5335 = 8'h6a == _T_241[7:0] ? 4'h0 : _GEN_5334; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5336 = 8'h6b == _T_241[7:0] ? 4'h0 : _GEN_5335; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5337 = 8'h6c == _T_241[7:0] ? 4'h0 : _GEN_5336; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5338 = 8'h6d == _T_241[7:0] ? 4'h0 : _GEN_5337; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5339 = 8'h6e == _T_241[7:0] ? 4'h6 : _GEN_5338; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5340 = 8'h6f == _T_241[7:0] ? 4'h0 : _GEN_5339; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5341 = 8'h70 == _T_241[7:0] ? 4'h0 : _GEN_5340; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5342 = 8'h71 == _T_241[7:0] ? 4'h0 : _GEN_5341; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5343 = 8'h72 == _T_241[7:0] ? 4'h3 : _GEN_5342; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5344 = 8'h73 == _T_241[7:0] ? 4'hc : _GEN_5343; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5345 = 8'h74 == _T_241[7:0] ? 4'h3 : _GEN_5344; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5346 = 8'h75 == _T_241[7:0] ? 4'h0 : _GEN_5345; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5347 = 8'h76 == _T_241[7:0] ? 4'h1 : _GEN_5346; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5348 = 8'h77 == _T_241[7:0] ? 4'h0 : _GEN_5347; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5349 = 8'h78 == _T_241[7:0] ? 4'h3 : _GEN_5348; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5350 = 8'h79 == _T_241[7:0] ? 4'h3 : _GEN_5349; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5351 = 8'h7a == _T_241[7:0] ? 4'h0 : _GEN_5350; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5352 = 8'h7b == _T_241[7:0] ? 4'h0 : _GEN_5351; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5353 = 8'h7c == _T_241[7:0] ? 4'h0 : _GEN_5352; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5354 = 8'h7d == _T_241[7:0] ? 4'h0 : _GEN_5353; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5355 = 8'h7e == _T_241[7:0] ? 4'h0 : _GEN_5354; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5356 = 8'h7f == _T_241[7:0] ? 4'h0 : _GEN_5355; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5357 = 8'h80 == _T_241[7:0] ? 4'h0 : _GEN_5356; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5358 = 8'h81 == _T_241[7:0] ? 4'h0 : _GEN_5357; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5359 = 8'h82 == _T_241[7:0] ? 4'h6 : _GEN_5358; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5360 = 8'h83 == _T_241[7:0] ? 4'h0 : _GEN_5359; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5361 = 8'h84 == _T_241[7:0] ? 4'h1 : _GEN_5360; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5362 = 8'h85 == _T_241[7:0] ? 4'h1 : _GEN_5361; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5363 = 8'h86 == _T_241[7:0] ? 4'ha : _GEN_5362; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5364 = 8'h87 == _T_241[7:0] ? 4'h4 : _GEN_5363; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5365 = 8'h88 == _T_241[7:0] ? 4'h1 : _GEN_5364; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5366 = 8'h89 == _T_241[7:0] ? 4'h4 : _GEN_5365; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5367 = 8'h8a == _T_241[7:0] ? 4'ha : _GEN_5366; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5368 = 8'h8b == _T_241[7:0] ? 4'h0 : _GEN_5367; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5369 = 8'h8c == _T_241[7:0] ? 4'h0 : _GEN_5368; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5370 = 8'h8d == _T_241[7:0] ? 4'h0 : _GEN_5369; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5371 = 8'h8e == _T_241[7:0] ? 4'h6 : _GEN_5370; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5372 = 8'h8f == _T_241[7:0] ? 4'h0 : _GEN_5371; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5373 = 8'h90 == _T_241[7:0] ? 4'h0 : _GEN_5372; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5374 = 8'h91 == _T_241[7:0] ? 4'h0 : _GEN_5373; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5375 = 8'h92 == _T_241[7:0] ? 4'h0 : _GEN_5374; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5376 = 8'h93 == _T_241[7:0] ? 4'h0 : _GEN_5375; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5377 = 8'h94 == _T_241[7:0] ? 4'h0 : _GEN_5376; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5378 = 8'h95 == _T_241[7:0] ? 4'h0 : _GEN_5377; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5379 = 8'h96 == _T_241[7:0] ? 4'h0 : _GEN_5378; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5380 = 8'h97 == _T_241[7:0] ? 4'h6 : _GEN_5379; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5381 = 8'h98 == _T_241[7:0] ? 4'h6 : _GEN_5380; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5382 = 8'h99 == _T_241[7:0] ? 4'h3 : _GEN_5381; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5383 = 8'h9a == _T_241[7:0] ? 4'h0 : _GEN_5382; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5384 = 8'h9b == _T_241[7:0] ? 4'ha : _GEN_5383; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5385 = 8'h9c == _T_241[7:0] ? 4'ha : _GEN_5384; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5386 = 8'h9d == _T_241[7:0] ? 4'h0 : _GEN_5385; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5387 = 8'h9e == _T_241[7:0] ? 4'ha : _GEN_5386; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5388 = 8'h9f == _T_241[7:0] ? 4'ha : _GEN_5387; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5389 = 8'ha0 == _T_241[7:0] ? 4'h0 : _GEN_5388; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5390 = 8'ha1 == _T_241[7:0] ? 4'h3 : _GEN_5389; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5391 = 8'ha2 == _T_241[7:0] ? 4'h6 : _GEN_5390; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5392 = 8'ha3 == _T_241[7:0] ? 4'h6 : _GEN_5391; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5393 = 8'ha4 == _T_241[7:0] ? 4'h0 : _GEN_5392; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5394 = 8'ha5 == _T_241[7:0] ? 4'h0 : _GEN_5393; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5395 = 8'ha6 == _T_241[7:0] ? 4'h0 : _GEN_5394; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5396 = 8'ha7 == _T_241[7:0] ? 4'h0 : _GEN_5395; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5397 = 8'ha8 == _T_241[7:0] ? 4'h0 : _GEN_5396; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5398 = 8'ha9 == _T_241[7:0] ? 4'h0 : _GEN_5397; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5399 = 8'haa == _T_241[7:0] ? 4'h0 : _GEN_5398; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5400 = 8'hab == _T_241[7:0] ? 4'h0 : _GEN_5399; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5401 = 8'hac == _T_241[7:0] ? 4'h6 : _GEN_5400; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5402 = 8'had == _T_241[7:0] ? 4'h0 : _GEN_5401; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5403 = 8'hae == _T_241[7:0] ? 4'h3 : _GEN_5402; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5404 = 8'haf == _T_241[7:0] ? 4'h9 : _GEN_5403; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5405 = 8'hb0 == _T_241[7:0] ? 4'h3 : _GEN_5404; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5406 = 8'hb1 == _T_241[7:0] ? 4'h0 : _GEN_5405; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5407 = 8'hb2 == _T_241[7:0] ? 4'h0 : _GEN_5406; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5408 = 8'hb3 == _T_241[7:0] ? 4'h0 : _GEN_5407; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5409 = 8'hb4 == _T_241[7:0] ? 4'h3 : _GEN_5408; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5410 = 8'hb5 == _T_241[7:0] ? 4'h9 : _GEN_5409; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5411 = 8'hb6 == _T_241[7:0] ? 4'h3 : _GEN_5410; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5412 = 8'hb7 == _T_241[7:0] ? 4'h0 : _GEN_5411; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5413 = 8'hb8 == _T_241[7:0] ? 4'h6 : _GEN_5412; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5414 = 8'hb9 == _T_241[7:0] ? 4'h0 : _GEN_5413; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5415 = 8'hba == _T_241[7:0] ? 4'h0 : _GEN_5414; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5416 = 8'hbb == _T_241[7:0] ? 4'h0 : _GEN_5415; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5417 = 8'hbc == _T_241[7:0] ? 4'h0 : _GEN_5416; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5418 = 8'hbd == _T_241[7:0] ? 4'h0 : _GEN_5417; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5419 = 8'hbe == _T_241[7:0] ? 4'h0 : _GEN_5418; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5420 = 8'hbf == _T_241[7:0] ? 4'h0 : _GEN_5419; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5421 = 8'hc0 == _T_241[7:0] ? 4'h0 : _GEN_5420; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5422 = 8'hc1 == _T_241[7:0] ? 4'h0 : _GEN_5421; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5423 = 8'hc2 == _T_241[7:0] ? 4'h7 : _GEN_5422; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5424 = 8'hc3 == _T_241[7:0] ? 4'h2 : _GEN_5423; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5425 = 8'hc4 == _T_241[7:0] ? 4'h0 : _GEN_5424; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5426 = 8'hc5 == _T_241[7:0] ? 4'h6 : _GEN_5425; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5427 = 8'hc6 == _T_241[7:0] ? 4'h9 : _GEN_5426; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5428 = 8'hc7 == _T_241[7:0] ? 4'h6 : _GEN_5427; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5429 = 8'hc8 == _T_241[7:0] ? 4'h9 : _GEN_5428; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5430 = 8'hc9 == _T_241[7:0] ? 4'h6 : _GEN_5429; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5431 = 8'hca == _T_241[7:0] ? 4'h0 : _GEN_5430; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5432 = 8'hcb == _T_241[7:0] ? 4'h2 : _GEN_5431; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5433 = 8'hcc == _T_241[7:0] ? 4'h7 : _GEN_5432; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5434 = 8'hcd == _T_241[7:0] ? 4'h0 : _GEN_5433; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5435 = 8'hce == _T_241[7:0] ? 4'h0 : _GEN_5434; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5436 = 8'hcf == _T_241[7:0] ? 4'h0 : _GEN_5435; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5437 = 8'hd0 == _T_241[7:0] ? 4'h0 : _GEN_5436; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5438 = 8'hd1 == _T_241[7:0] ? 4'h0 : _GEN_5437; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5439 = 8'hd2 == _T_241[7:0] ? 4'h0 : _GEN_5438; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5440 = 8'hd3 == _T_241[7:0] ? 4'h0 : _GEN_5439; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5441 = 8'hd4 == _T_241[7:0] ? 4'h0 : _GEN_5440; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5442 = 8'hd5 == _T_241[7:0] ? 4'h0 : _GEN_5441; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5443 = 8'hd6 == _T_241[7:0] ? 4'h0 : _GEN_5442; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5444 = 8'hd7 == _T_241[7:0] ? 4'h3 : _GEN_5443; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5445 = 8'hd8 == _T_241[7:0] ? 4'h3 : _GEN_5444; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5446 = 8'hd9 == _T_241[7:0] ? 4'h0 : _GEN_5445; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5447 = 8'hda == _T_241[7:0] ? 4'h9 : _GEN_5446; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5448 = 8'hdb == _T_241[7:0] ? 4'h3 : _GEN_5447; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5449 = 8'hdc == _T_241[7:0] ? 4'hc : _GEN_5448; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5450 = 8'hdd == _T_241[7:0] ? 4'h3 : _GEN_5449; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5451 = 8'hde == _T_241[7:0] ? 4'h9 : _GEN_5450; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5452 = 8'hdf == _T_241[7:0] ? 4'h0 : _GEN_5451; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5453 = 8'he0 == _T_241[7:0] ? 4'h3 : _GEN_5452; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5454 = 8'he1 == _T_241[7:0] ? 4'h3 : _GEN_5453; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5455 = 8'he2 == _T_241[7:0] ? 4'h0 : _GEN_5454; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5456 = 8'he3 == _T_241[7:0] ? 4'h0 : _GEN_5455; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5457 = 8'he4 == _T_241[7:0] ? 4'h0 : _GEN_5456; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5458 = 8'he5 == _T_241[7:0] ? 4'h0 : _GEN_5457; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5459 = 8'he6 == _T_241[7:0] ? 4'h0 : _GEN_5458; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5460 = 8'he7 == _T_241[7:0] ? 4'h0 : _GEN_5459; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5461 = 8'he8 == _T_241[7:0] ? 4'h0 : _GEN_5460; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5462 = 8'he9 == _T_241[7:0] ? 4'h0 : _GEN_5461; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5463 = 8'hea == _T_241[7:0] ? 4'h0 : _GEN_5462; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5464 = 8'heb == _T_241[7:0] ? 4'h0 : _GEN_5463; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5465 = 8'hec == _T_241[7:0] ? 4'h0 : _GEN_5464; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5466 = 8'hed == _T_241[7:0] ? 4'h0 : _GEN_5465; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5467 = 8'hee == _T_241[7:0] ? 4'h0 : _GEN_5466; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5468 = 8'hef == _T_241[7:0] ? 4'h0 : _GEN_5467; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5469 = 8'hf0 == _T_241[7:0] ? 4'h0 : _GEN_5468; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5470 = 8'hf1 == _T_241[7:0] ? 4'h0 : _GEN_5469; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5471 = 8'hf2 == _T_241[7:0] ? 4'h0 : _GEN_5470; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5472 = 8'hf3 == _T_241[7:0] ? 4'h0 : _GEN_5471; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5473 = 8'hf4 == _T_241[7:0] ? 4'h0 : _GEN_5472; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5474 = 8'hf5 == _T_241[7:0] ? 4'h0 : _GEN_5473; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5475 = 8'hf6 == _T_241[7:0] ? 4'h0 : _GEN_5474; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5476 = 8'hf7 == _T_241[7:0] ? 4'h0 : _GEN_5475; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5477 = 8'hf8 == _T_241[7:0] ? 4'h0 : _GEN_5476; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5478 = 8'hf9 == _T_241[7:0] ? 4'h0 : _GEN_5477; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5479 = 8'hfa == _T_241[7:0] ? 4'h0 : _GEN_5478; // @[Filter.scala 204:142]
  wire [3:0] _GEN_5480 = 8'hfb == _T_241[7:0] ? 4'h0 : _GEN_5479; // @[Filter.scala 204:142]
  wire [7:0] _T_255 = _GEN_5480 * 4'ha; // @[Filter.scala 204:142]
  wire [10:0] _GEN_11254 = {{3'd0}, _T_255}; // @[Filter.scala 204:109]
  wire [10:0] _T_257 = _T_250 + _GEN_11254; // @[Filter.scala 204:109]
  wire [10:0] _T_258 = _T_257 / 11'h64; // @[Filter.scala 204:150]
  wire  _T_260 = _T_231 >= 5'h15; // @[Filter.scala 207:31]
  wire  _T_264 = _T_238 >= 32'hc; // @[Filter.scala 207:63]
  wire  _T_265 = _T_260 | _T_264; // @[Filter.scala 207:58]
  wire [10:0] _GEN_5733 = io_SPI_distort ? _T_258 : {{7'd0}, _GEN_4976}; // @[Filter.scala 209:35]
  wire [10:0] _GEN_5734 = _T_265 ? 11'h0 : _GEN_5733; // @[Filter.scala 207:80]
  wire [10:0] _GEN_5987 = io_SPI_distort ? _T_258 : {{7'd0}, _GEN_5228}; // @[Filter.scala 209:35]
  wire [10:0] _GEN_5988 = _T_265 ? 11'h0 : _GEN_5987; // @[Filter.scala 207:80]
  wire [10:0] _GEN_6241 = io_SPI_distort ? _T_258 : {{7'd0}, _GEN_5480}; // @[Filter.scala 209:35]
  wire [10:0] _GEN_6242 = _T_265 ? 11'h0 : _GEN_6241; // @[Filter.scala 207:80]
  wire [31:0] _T_293 = pixelIndex + 32'h4; // @[Filter.scala 202:31]
  wire [31:0] _GEN_4 = _T_293 % 32'h15; // @[Filter.scala 202:38]
  wire [4:0] _T_294 = _GEN_4[4:0]; // @[Filter.scala 202:38]
  wire [4:0] _T_296 = _T_294 + _GEN_11210; // @[Filter.scala 202:53]
  wire [4:0] _T_298 = _T_296 - 5'h1; // @[Filter.scala 202:69]
  wire [31:0] _T_301 = _T_293 / 32'h15; // @[Filter.scala 203:38]
  wire [31:0] _T_303 = _T_301 + _GEN_11211; // @[Filter.scala 203:53]
  wire [31:0] _T_305 = _T_303 - 32'h1; // @[Filter.scala 203:69]
  wire [36:0] _T_306 = _T_305 * 32'h15; // @[Filter.scala 204:42]
  wire [36:0] _GEN_11260 = {{32'd0}, _T_298}; // @[Filter.scala 204:57]
  wire [36:0] _T_308 = _T_306 + _GEN_11260; // @[Filter.scala 204:57]
  wire [3:0] _GEN_6251 = 8'h8 == _T_308[7:0] ? 4'h1 : 4'h0; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6252 = 8'h9 == _T_308[7:0] ? 4'h2 : _GEN_6251; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6253 = 8'ha == _T_308[7:0] ? 4'h2 : _GEN_6252; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6254 = 8'hb == _T_308[7:0] ? 4'h2 : _GEN_6253; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6255 = 8'hc == _T_308[7:0] ? 4'h1 : _GEN_6254; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6256 = 8'hd == _T_308[7:0] ? 4'h0 : _GEN_6255; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6257 = 8'he == _T_308[7:0] ? 4'h0 : _GEN_6256; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6258 = 8'hf == _T_308[7:0] ? 4'h0 : _GEN_6257; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6259 = 8'h10 == _T_308[7:0] ? 4'h0 : _GEN_6258; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6260 = 8'h11 == _T_308[7:0] ? 4'h0 : _GEN_6259; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6261 = 8'h12 == _T_308[7:0] ? 4'h0 : _GEN_6260; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6262 = 8'h13 == _T_308[7:0] ? 4'h0 : _GEN_6261; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6263 = 8'h14 == _T_308[7:0] ? 4'h0 : _GEN_6262; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6264 = 8'h15 == _T_308[7:0] ? 4'h0 : _GEN_6263; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6265 = 8'h16 == _T_308[7:0] ? 4'h0 : _GEN_6264; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6266 = 8'h17 == _T_308[7:0] ? 4'h0 : _GEN_6265; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6267 = 8'h18 == _T_308[7:0] ? 4'h0 : _GEN_6266; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6268 = 8'h19 == _T_308[7:0] ? 4'h0 : _GEN_6267; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6269 = 8'h1a == _T_308[7:0] ? 4'h0 : _GEN_6268; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6270 = 8'h1b == _T_308[7:0] ? 4'h0 : _GEN_6269; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6271 = 8'h1c == _T_308[7:0] ? 4'h2 : _GEN_6270; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6272 = 8'h1d == _T_308[7:0] ? 4'h1 : _GEN_6271; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6273 = 8'h1e == _T_308[7:0] ? 4'h0 : _GEN_6272; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6274 = 8'h1f == _T_308[7:0] ? 4'h0 : _GEN_6273; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6275 = 8'h20 == _T_308[7:0] ? 4'h0 : _GEN_6274; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6276 = 8'h21 == _T_308[7:0] ? 4'h1 : _GEN_6275; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6277 = 8'h22 == _T_308[7:0] ? 4'h2 : _GEN_6276; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6278 = 8'h23 == _T_308[7:0] ? 4'h0 : _GEN_6277; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6279 = 8'h24 == _T_308[7:0] ? 4'h0 : _GEN_6278; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6280 = 8'h25 == _T_308[7:0] ? 4'h0 : _GEN_6279; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6281 = 8'h26 == _T_308[7:0] ? 4'h0 : _GEN_6280; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6282 = 8'h27 == _T_308[7:0] ? 4'h0 : _GEN_6281; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6283 = 8'h28 == _T_308[7:0] ? 4'h0 : _GEN_6282; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6284 = 8'h29 == _T_308[7:0] ? 4'h0 : _GEN_6283; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6285 = 8'h2a == _T_308[7:0] ? 4'h0 : _GEN_6284; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6286 = 8'h2b == _T_308[7:0] ? 4'h0 : _GEN_6285; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6287 = 8'h2c == _T_308[7:0] ? 4'h0 : _GEN_6286; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6288 = 8'h2d == _T_308[7:0] ? 4'h0 : _GEN_6287; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6289 = 8'h2e == _T_308[7:0] ? 4'h0 : _GEN_6288; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6290 = 8'h2f == _T_308[7:0] ? 4'h0 : _GEN_6289; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6291 = 8'h30 == _T_308[7:0] ? 4'h2 : _GEN_6290; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6292 = 8'h31 == _T_308[7:0] ? 4'h2 : _GEN_6291; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6293 = 8'h32 == _T_308[7:0] ? 4'h0 : _GEN_6292; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6294 = 8'h33 == _T_308[7:0] ? 4'h0 : _GEN_6293; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6295 = 8'h34 == _T_308[7:0] ? 4'h0 : _GEN_6294; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6296 = 8'h35 == _T_308[7:0] ? 4'h0 : _GEN_6295; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6297 = 8'h36 == _T_308[7:0] ? 4'h0 : _GEN_6296; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6298 = 8'h37 == _T_308[7:0] ? 4'h0 : _GEN_6297; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6299 = 8'h38 == _T_308[7:0] ? 4'h2 : _GEN_6298; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6300 = 8'h39 == _T_308[7:0] ? 4'h0 : _GEN_6299; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6301 = 8'h3a == _T_308[7:0] ? 4'h0 : _GEN_6300; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6302 = 8'h3b == _T_308[7:0] ? 4'h0 : _GEN_6301; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6303 = 8'h3c == _T_308[7:0] ? 4'h0 : _GEN_6302; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6304 = 8'h3d == _T_308[7:0] ? 4'h0 : _GEN_6303; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6305 = 8'h3e == _T_308[7:0] ? 4'h0 : _GEN_6304; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6306 = 8'h3f == _T_308[7:0] ? 4'h0 : _GEN_6305; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6307 = 8'h40 == _T_308[7:0] ? 4'h0 : _GEN_6306; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6308 = 8'h41 == _T_308[7:0] ? 4'h0 : _GEN_6307; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6309 = 8'h42 == _T_308[7:0] ? 4'h0 : _GEN_6308; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6310 = 8'h43 == _T_308[7:0] ? 4'h0 : _GEN_6309; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6311 = 8'h44 == _T_308[7:0] ? 4'h1 : _GEN_6310; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6312 = 8'h45 == _T_308[7:0] ? 4'h3 : _GEN_6311; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6313 = 8'h46 == _T_308[7:0] ? 4'h7 : _GEN_6312; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6314 = 8'h47 == _T_308[7:0] ? 4'h0 : _GEN_6313; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6315 = 8'h48 == _T_308[7:0] ? 4'h0 : _GEN_6314; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6316 = 8'h49 == _T_308[7:0] ? 4'h0 : _GEN_6315; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6317 = 8'h4a == _T_308[7:0] ? 4'h0 : _GEN_6316; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6318 = 8'h4b == _T_308[7:0] ? 4'h0 : _GEN_6317; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6319 = 8'h4c == _T_308[7:0] ? 4'h0 : _GEN_6318; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6320 = 8'h4d == _T_308[7:0] ? 4'h0 : _GEN_6319; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6321 = 8'h4e == _T_308[7:0] ? 4'h2 : _GEN_6320; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6322 = 8'h4f == _T_308[7:0] ? 4'h0 : _GEN_6321; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6323 = 8'h50 == _T_308[7:0] ? 4'h0 : _GEN_6322; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6324 = 8'h51 == _T_308[7:0] ? 4'h0 : _GEN_6323; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6325 = 8'h52 == _T_308[7:0] ? 4'h0 : _GEN_6324; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6326 = 8'h53 == _T_308[7:0] ? 4'h0 : _GEN_6325; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6327 = 8'h54 == _T_308[7:0] ? 4'h0 : _GEN_6326; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6328 = 8'h55 == _T_308[7:0] ? 4'h0 : _GEN_6327; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6329 = 8'h56 == _T_308[7:0] ? 4'h0 : _GEN_6328; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6330 = 8'h57 == _T_308[7:0] ? 4'h0 : _GEN_6329; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6331 = 8'h58 == _T_308[7:0] ? 4'h0 : _GEN_6330; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6332 = 8'h59 == _T_308[7:0] ? 4'h2 : _GEN_6331; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6333 = 8'h5a == _T_308[7:0] ? 4'h2 : _GEN_6332; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6334 = 8'h5b == _T_308[7:0] ? 4'h0 : _GEN_6333; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6335 = 8'h5c == _T_308[7:0] ? 4'h0 : _GEN_6334; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6336 = 8'h5d == _T_308[7:0] ? 4'h0 : _GEN_6335; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6337 = 8'h5e == _T_308[7:0] ? 4'h4 : _GEN_6336; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6338 = 8'h5f == _T_308[7:0] ? 4'h0 : _GEN_6337; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6339 = 8'h60 == _T_308[7:0] ? 4'h0 : _GEN_6338; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6340 = 8'h61 == _T_308[7:0] ? 4'h0 : _GEN_6339; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6341 = 8'h62 == _T_308[7:0] ? 4'h0 : _GEN_6340; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6342 = 8'h63 == _T_308[7:0] ? 4'h2 : _GEN_6341; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6343 = 8'h64 == _T_308[7:0] ? 4'h0 : _GEN_6342; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6344 = 8'h65 == _T_308[7:0] ? 4'h0 : _GEN_6343; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6345 = 8'h66 == _T_308[7:0] ? 4'h0 : _GEN_6344; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6346 = 8'h67 == _T_308[7:0] ? 4'h0 : _GEN_6345; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6347 = 8'h68 == _T_308[7:0] ? 4'h0 : _GEN_6346; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6348 = 8'h69 == _T_308[7:0] ? 4'h0 : _GEN_6347; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6349 = 8'h6a == _T_308[7:0] ? 4'h0 : _GEN_6348; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6350 = 8'h6b == _T_308[7:0] ? 4'h0 : _GEN_6349; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6351 = 8'h6c == _T_308[7:0] ? 4'h0 : _GEN_6350; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6352 = 8'h6d == _T_308[7:0] ? 4'h0 : _GEN_6351; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6353 = 8'h6e == _T_308[7:0] ? 4'h2 : _GEN_6352; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6354 = 8'h6f == _T_308[7:0] ? 4'h0 : _GEN_6353; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6355 = 8'h70 == _T_308[7:0] ? 4'h0 : _GEN_6354; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6356 = 8'h71 == _T_308[7:0] ? 4'h0 : _GEN_6355; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6357 = 8'h72 == _T_308[7:0] ? 4'h2 : _GEN_6356; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6358 = 8'h73 == _T_308[7:0] ? 4'h9 : _GEN_6357; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6359 = 8'h74 == _T_308[7:0] ? 4'h2 : _GEN_6358; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6360 = 8'h75 == _T_308[7:0] ? 4'h0 : _GEN_6359; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6361 = 8'h76 == _T_308[7:0] ? 4'h0 : _GEN_6360; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6362 = 8'h77 == _T_308[7:0] ? 4'h0 : _GEN_6361; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6363 = 8'h78 == _T_308[7:0] ? 4'h1 : _GEN_6362; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6364 = 8'h79 == _T_308[7:0] ? 4'h1 : _GEN_6363; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6365 = 8'h7a == _T_308[7:0] ? 4'h0 : _GEN_6364; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6366 = 8'h7b == _T_308[7:0] ? 4'h0 : _GEN_6365; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6367 = 8'h7c == _T_308[7:0] ? 4'h0 : _GEN_6366; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6368 = 8'h7d == _T_308[7:0] ? 4'h0 : _GEN_6367; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6369 = 8'h7e == _T_308[7:0] ? 4'h0 : _GEN_6368; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6370 = 8'h7f == _T_308[7:0] ? 4'h0 : _GEN_6369; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6371 = 8'h80 == _T_308[7:0] ? 4'h0 : _GEN_6370; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6372 = 8'h81 == _T_308[7:0] ? 4'h0 : _GEN_6371; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6373 = 8'h82 == _T_308[7:0] ? 4'h2 : _GEN_6372; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6374 = 8'h83 == _T_308[7:0] ? 4'h0 : _GEN_6373; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6375 = 8'h84 == _T_308[7:0] ? 4'h0 : _GEN_6374; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6376 = 8'h85 == _T_308[7:0] ? 4'h0 : _GEN_6375; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6377 = 8'h86 == _T_308[7:0] ? 4'h7 : _GEN_6376; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6378 = 8'h87 == _T_308[7:0] ? 4'h2 : _GEN_6377; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6379 = 8'h88 == _T_308[7:0] ? 4'h0 : _GEN_6378; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6380 = 8'h89 == _T_308[7:0] ? 4'h2 : _GEN_6379; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6381 = 8'h8a == _T_308[7:0] ? 4'h7 : _GEN_6380; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6382 = 8'h8b == _T_308[7:0] ? 4'h0 : _GEN_6381; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6383 = 8'h8c == _T_308[7:0] ? 4'h0 : _GEN_6382; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6384 = 8'h8d == _T_308[7:0] ? 4'h0 : _GEN_6383; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6385 = 8'h8e == _T_308[7:0] ? 4'h2 : _GEN_6384; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6386 = 8'h8f == _T_308[7:0] ? 4'h0 : _GEN_6385; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6387 = 8'h90 == _T_308[7:0] ? 4'h0 : _GEN_6386; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6388 = 8'h91 == _T_308[7:0] ? 4'h0 : _GEN_6387; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6389 = 8'h92 == _T_308[7:0] ? 4'h0 : _GEN_6388; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6390 = 8'h93 == _T_308[7:0] ? 4'h0 : _GEN_6389; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6391 = 8'h94 == _T_308[7:0] ? 4'h0 : _GEN_6390; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6392 = 8'h95 == _T_308[7:0] ? 4'h0 : _GEN_6391; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6393 = 8'h96 == _T_308[7:0] ? 4'h0 : _GEN_6392; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6394 = 8'h97 == _T_308[7:0] ? 4'h2 : _GEN_6393; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6395 = 8'h98 == _T_308[7:0] ? 4'h2 : _GEN_6394; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6396 = 8'h99 == _T_308[7:0] ? 4'h1 : _GEN_6395; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6397 = 8'h9a == _T_308[7:0] ? 4'h0 : _GEN_6396; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6398 = 8'h9b == _T_308[7:0] ? 4'h7 : _GEN_6397; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6399 = 8'h9c == _T_308[7:0] ? 4'h7 : _GEN_6398; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6400 = 8'h9d == _T_308[7:0] ? 4'h0 : _GEN_6399; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6401 = 8'h9e == _T_308[7:0] ? 4'h7 : _GEN_6400; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6402 = 8'h9f == _T_308[7:0] ? 4'h7 : _GEN_6401; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6403 = 8'ha0 == _T_308[7:0] ? 4'h0 : _GEN_6402; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6404 = 8'ha1 == _T_308[7:0] ? 4'h1 : _GEN_6403; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6405 = 8'ha2 == _T_308[7:0] ? 4'h2 : _GEN_6404; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6406 = 8'ha3 == _T_308[7:0] ? 4'h2 : _GEN_6405; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6407 = 8'ha4 == _T_308[7:0] ? 4'h0 : _GEN_6406; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6408 = 8'ha5 == _T_308[7:0] ? 4'h0 : _GEN_6407; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6409 = 8'ha6 == _T_308[7:0] ? 4'h0 : _GEN_6408; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6410 = 8'ha7 == _T_308[7:0] ? 4'h0 : _GEN_6409; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6411 = 8'ha8 == _T_308[7:0] ? 4'h0 : _GEN_6410; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6412 = 8'ha9 == _T_308[7:0] ? 4'h0 : _GEN_6411; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6413 = 8'haa == _T_308[7:0] ? 4'h0 : _GEN_6412; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6414 = 8'hab == _T_308[7:0] ? 4'h0 : _GEN_6413; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6415 = 8'hac == _T_308[7:0] ? 4'h2 : _GEN_6414; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6416 = 8'had == _T_308[7:0] ? 4'h0 : _GEN_6415; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6417 = 8'hae == _T_308[7:0] ? 4'h1 : _GEN_6416; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6418 = 8'haf == _T_308[7:0] ? 4'h3 : _GEN_6417; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6419 = 8'hb0 == _T_308[7:0] ? 4'h1 : _GEN_6418; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6420 = 8'hb1 == _T_308[7:0] ? 4'h0 : _GEN_6419; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6421 = 8'hb2 == _T_308[7:0] ? 4'h0 : _GEN_6420; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6422 = 8'hb3 == _T_308[7:0] ? 4'h0 : _GEN_6421; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6423 = 8'hb4 == _T_308[7:0] ? 4'h1 : _GEN_6422; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6424 = 8'hb5 == _T_308[7:0] ? 4'h3 : _GEN_6423; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6425 = 8'hb6 == _T_308[7:0] ? 4'h1 : _GEN_6424; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6426 = 8'hb7 == _T_308[7:0] ? 4'h0 : _GEN_6425; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6427 = 8'hb8 == _T_308[7:0] ? 4'h2 : _GEN_6426; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6428 = 8'hb9 == _T_308[7:0] ? 4'h0 : _GEN_6427; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6429 = 8'hba == _T_308[7:0] ? 4'h0 : _GEN_6428; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6430 = 8'hbb == _T_308[7:0] ? 4'h0 : _GEN_6429; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6431 = 8'hbc == _T_308[7:0] ? 4'h0 : _GEN_6430; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6432 = 8'hbd == _T_308[7:0] ? 4'h0 : _GEN_6431; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6433 = 8'hbe == _T_308[7:0] ? 4'h0 : _GEN_6432; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6434 = 8'hbf == _T_308[7:0] ? 4'h0 : _GEN_6433; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6435 = 8'hc0 == _T_308[7:0] ? 4'h0 : _GEN_6434; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6436 = 8'hc1 == _T_308[7:0] ? 4'h0 : _GEN_6435; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6437 = 8'hc2 == _T_308[7:0] ? 4'h3 : _GEN_6436; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6438 = 8'hc3 == _T_308[7:0] ? 4'h0 : _GEN_6437; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6439 = 8'hc4 == _T_308[7:0] ? 4'h0 : _GEN_6438; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6440 = 8'hc5 == _T_308[7:0] ? 4'h2 : _GEN_6439; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6441 = 8'hc6 == _T_308[7:0] ? 4'h3 : _GEN_6440; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6442 = 8'hc7 == _T_308[7:0] ? 4'h2 : _GEN_6441; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6443 = 8'hc8 == _T_308[7:0] ? 4'h3 : _GEN_6442; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6444 = 8'hc9 == _T_308[7:0] ? 4'h2 : _GEN_6443; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6445 = 8'hca == _T_308[7:0] ? 4'h0 : _GEN_6444; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6446 = 8'hcb == _T_308[7:0] ? 4'h0 : _GEN_6445; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6447 = 8'hcc == _T_308[7:0] ? 4'h3 : _GEN_6446; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6448 = 8'hcd == _T_308[7:0] ? 4'h0 : _GEN_6447; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6449 = 8'hce == _T_308[7:0] ? 4'h0 : _GEN_6448; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6450 = 8'hcf == _T_308[7:0] ? 4'h0 : _GEN_6449; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6451 = 8'hd0 == _T_308[7:0] ? 4'h0 : _GEN_6450; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6452 = 8'hd1 == _T_308[7:0] ? 4'h0 : _GEN_6451; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6453 = 8'hd2 == _T_308[7:0] ? 4'h0 : _GEN_6452; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6454 = 8'hd3 == _T_308[7:0] ? 4'h0 : _GEN_6453; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6455 = 8'hd4 == _T_308[7:0] ? 4'h0 : _GEN_6454; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6456 = 8'hd5 == _T_308[7:0] ? 4'h0 : _GEN_6455; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6457 = 8'hd6 == _T_308[7:0] ? 4'h0 : _GEN_6456; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6458 = 8'hd7 == _T_308[7:0] ? 4'h2 : _GEN_6457; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6459 = 8'hd8 == _T_308[7:0] ? 4'h2 : _GEN_6458; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6460 = 8'hd9 == _T_308[7:0] ? 4'h0 : _GEN_6459; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6461 = 8'hda == _T_308[7:0] ? 4'h7 : _GEN_6460; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6462 = 8'hdb == _T_308[7:0] ? 4'h1 : _GEN_6461; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6463 = 8'hdc == _T_308[7:0] ? 4'h4 : _GEN_6462; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6464 = 8'hdd == _T_308[7:0] ? 4'h1 : _GEN_6463; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6465 = 8'hde == _T_308[7:0] ? 4'h7 : _GEN_6464; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6466 = 8'hdf == _T_308[7:0] ? 4'h0 : _GEN_6465; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6467 = 8'he0 == _T_308[7:0] ? 4'h2 : _GEN_6466; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6468 = 8'he1 == _T_308[7:0] ? 4'h2 : _GEN_6467; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6469 = 8'he2 == _T_308[7:0] ? 4'h0 : _GEN_6468; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6470 = 8'he3 == _T_308[7:0] ? 4'h0 : _GEN_6469; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6471 = 8'he4 == _T_308[7:0] ? 4'h0 : _GEN_6470; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6472 = 8'he5 == _T_308[7:0] ? 4'h0 : _GEN_6471; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6473 = 8'he6 == _T_308[7:0] ? 4'h0 : _GEN_6472; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6474 = 8'he7 == _T_308[7:0] ? 4'h0 : _GEN_6473; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6475 = 8'he8 == _T_308[7:0] ? 4'h0 : _GEN_6474; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6476 = 8'he9 == _T_308[7:0] ? 4'h0 : _GEN_6475; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6477 = 8'hea == _T_308[7:0] ? 4'h0 : _GEN_6476; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6478 = 8'heb == _T_308[7:0] ? 4'h0 : _GEN_6477; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6479 = 8'hec == _T_308[7:0] ? 4'h0 : _GEN_6478; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6480 = 8'hed == _T_308[7:0] ? 4'h0 : _GEN_6479; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6481 = 8'hee == _T_308[7:0] ? 4'h0 : _GEN_6480; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6482 = 8'hef == _T_308[7:0] ? 4'h0 : _GEN_6481; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6483 = 8'hf0 == _T_308[7:0] ? 4'h0 : _GEN_6482; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6484 = 8'hf1 == _T_308[7:0] ? 4'h0 : _GEN_6483; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6485 = 8'hf2 == _T_308[7:0] ? 4'h0 : _GEN_6484; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6486 = 8'hf3 == _T_308[7:0] ? 4'h0 : _GEN_6485; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6487 = 8'hf4 == _T_308[7:0] ? 4'h0 : _GEN_6486; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6488 = 8'hf5 == _T_308[7:0] ? 4'h0 : _GEN_6487; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6489 = 8'hf6 == _T_308[7:0] ? 4'h0 : _GEN_6488; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6490 = 8'hf7 == _T_308[7:0] ? 4'h0 : _GEN_6489; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6491 = 8'hf8 == _T_308[7:0] ? 4'h0 : _GEN_6490; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6492 = 8'hf9 == _T_308[7:0] ? 4'h0 : _GEN_6491; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6493 = 8'hfa == _T_308[7:0] ? 4'h0 : _GEN_6492; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6494 = 8'hfb == _T_308[7:0] ? 4'h0 : _GEN_6493; // @[Filter.scala 204:62]
  wire [4:0] _GEN_11261 = {{1'd0}, _GEN_6494}; // @[Filter.scala 204:62]
  wire [8:0] _T_310 = _GEN_11261 * 5'h14; // @[Filter.scala 204:62]
  wire [3:0] _GEN_6544 = 8'h31 == _T_308[7:0] ? 4'h3 : _GEN_6291; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6545 = 8'h32 == _T_308[7:0] ? 4'h3 : _GEN_6544; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6546 = 8'h33 == _T_308[7:0] ? 4'h6 : _GEN_6545; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6547 = 8'h34 == _T_308[7:0] ? 4'h6 : _GEN_6546; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6548 = 8'h35 == _T_308[7:0] ? 4'h0 : _GEN_6547; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6549 = 8'h36 == _T_308[7:0] ? 4'h0 : _GEN_6548; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6550 = 8'h37 == _T_308[7:0] ? 4'h0 : _GEN_6549; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6551 = 8'h38 == _T_308[7:0] ? 4'h2 : _GEN_6550; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6552 = 8'h39 == _T_308[7:0] ? 4'h0 : _GEN_6551; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6553 = 8'h3a == _T_308[7:0] ? 4'h0 : _GEN_6552; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6554 = 8'h3b == _T_308[7:0] ? 4'h0 : _GEN_6553; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6555 = 8'h3c == _T_308[7:0] ? 4'h0 : _GEN_6554; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6556 = 8'h3d == _T_308[7:0] ? 4'h0 : _GEN_6555; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6557 = 8'h3e == _T_308[7:0] ? 4'h0 : _GEN_6556; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6558 = 8'h3f == _T_308[7:0] ? 4'h0 : _GEN_6557; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6559 = 8'h40 == _T_308[7:0] ? 4'h0 : _GEN_6558; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6560 = 8'h41 == _T_308[7:0] ? 4'h0 : _GEN_6559; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6561 = 8'h42 == _T_308[7:0] ? 4'h0 : _GEN_6560; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6562 = 8'h43 == _T_308[7:0] ? 4'h0 : _GEN_6561; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6563 = 8'h44 == _T_308[7:0] ? 4'h1 : _GEN_6562; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6564 = 8'h45 == _T_308[7:0] ? 4'h4 : _GEN_6563; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6565 = 8'h46 == _T_308[7:0] ? 4'hb : _GEN_6564; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6566 = 8'h47 == _T_308[7:0] ? 4'h0 : _GEN_6565; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6567 = 8'h48 == _T_308[7:0] ? 4'h0 : _GEN_6566; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6568 = 8'h49 == _T_308[7:0] ? 4'h0 : _GEN_6567; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6569 = 8'h4a == _T_308[7:0] ? 4'h6 : _GEN_6568; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6570 = 8'h4b == _T_308[7:0] ? 4'h0 : _GEN_6569; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6571 = 8'h4c == _T_308[7:0] ? 4'h3 : _GEN_6570; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6572 = 8'h4d == _T_308[7:0] ? 4'h3 : _GEN_6571; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6573 = 8'h4e == _T_308[7:0] ? 4'h2 : _GEN_6572; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6574 = 8'h4f == _T_308[7:0] ? 4'h0 : _GEN_6573; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6575 = 8'h50 == _T_308[7:0] ? 4'h0 : _GEN_6574; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6576 = 8'h51 == _T_308[7:0] ? 4'h0 : _GEN_6575; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6577 = 8'h52 == _T_308[7:0] ? 4'h0 : _GEN_6576; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6578 = 8'h53 == _T_308[7:0] ? 4'h0 : _GEN_6577; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6579 = 8'h54 == _T_308[7:0] ? 4'h0 : _GEN_6578; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6580 = 8'h55 == _T_308[7:0] ? 4'h0 : _GEN_6579; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6581 = 8'h56 == _T_308[7:0] ? 4'h0 : _GEN_6580; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6582 = 8'h57 == _T_308[7:0] ? 4'h0 : _GEN_6581; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6583 = 8'h58 == _T_308[7:0] ? 4'h0 : _GEN_6582; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6584 = 8'h59 == _T_308[7:0] ? 4'h2 : _GEN_6583; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6585 = 8'h5a == _T_308[7:0] ? 4'h3 : _GEN_6584; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6586 = 8'h5b == _T_308[7:0] ? 4'h0 : _GEN_6585; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6587 = 8'h5c == _T_308[7:0] ? 4'h0 : _GEN_6586; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6588 = 8'h5d == _T_308[7:0] ? 4'h3 : _GEN_6587; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6589 = 8'h5e == _T_308[7:0] ? 4'hd : _GEN_6588; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6590 = 8'h5f == _T_308[7:0] ? 4'h3 : _GEN_6589; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6591 = 8'h60 == _T_308[7:0] ? 4'h0 : _GEN_6590; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6592 = 8'h61 == _T_308[7:0] ? 4'h6 : _GEN_6591; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6593 = 8'h62 == _T_308[7:0] ? 4'h0 : _GEN_6592; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6594 = 8'h63 == _T_308[7:0] ? 4'h2 : _GEN_6593; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6595 = 8'h64 == _T_308[7:0] ? 4'h0 : _GEN_6594; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6596 = 8'h65 == _T_308[7:0] ? 4'h0 : _GEN_6595; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6597 = 8'h66 == _T_308[7:0] ? 4'h0 : _GEN_6596; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6598 = 8'h67 == _T_308[7:0] ? 4'h0 : _GEN_6597; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6599 = 8'h68 == _T_308[7:0] ? 4'h0 : _GEN_6598; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6600 = 8'h69 == _T_308[7:0] ? 4'h0 : _GEN_6599; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6601 = 8'h6a == _T_308[7:0] ? 4'h0 : _GEN_6600; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6602 = 8'h6b == _T_308[7:0] ? 4'h0 : _GEN_6601; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6603 = 8'h6c == _T_308[7:0] ? 4'h0 : _GEN_6602; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6604 = 8'h6d == _T_308[7:0] ? 4'h0 : _GEN_6603; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6605 = 8'h6e == _T_308[7:0] ? 4'h2 : _GEN_6604; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6606 = 8'h6f == _T_308[7:0] ? 4'h0 : _GEN_6605; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6607 = 8'h70 == _T_308[7:0] ? 4'h0 : _GEN_6606; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6608 = 8'h71 == _T_308[7:0] ? 4'h0 : _GEN_6607; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6609 = 8'h72 == _T_308[7:0] ? 4'h6 : _GEN_6608; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6610 = 8'h73 == _T_308[7:0] ? 4'he : _GEN_6609; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6611 = 8'h74 == _T_308[7:0] ? 4'h6 : _GEN_6610; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6612 = 8'h75 == _T_308[7:0] ? 4'h0 : _GEN_6611; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6613 = 8'h76 == _T_308[7:0] ? 4'h6 : _GEN_6612; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6614 = 8'h77 == _T_308[7:0] ? 4'h3 : _GEN_6613; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6615 = 8'h78 == _T_308[7:0] ? 4'h4 : _GEN_6614; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6616 = 8'h79 == _T_308[7:0] ? 4'h1 : _GEN_6615; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6617 = 8'h7a == _T_308[7:0] ? 4'h0 : _GEN_6616; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6618 = 8'h7b == _T_308[7:0] ? 4'h0 : _GEN_6617; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6619 = 8'h7c == _T_308[7:0] ? 4'h0 : _GEN_6618; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6620 = 8'h7d == _T_308[7:0] ? 4'h0 : _GEN_6619; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6621 = 8'h7e == _T_308[7:0] ? 4'h0 : _GEN_6620; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6622 = 8'h7f == _T_308[7:0] ? 4'h0 : _GEN_6621; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6623 = 8'h80 == _T_308[7:0] ? 4'h0 : _GEN_6622; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6624 = 8'h81 == _T_308[7:0] ? 4'h0 : _GEN_6623; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6625 = 8'h82 == _T_308[7:0] ? 4'h2 : _GEN_6624; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6626 = 8'h83 == _T_308[7:0] ? 4'h3 : _GEN_6625; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6627 = 8'h84 == _T_308[7:0] ? 4'h6 : _GEN_6626; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6628 = 8'h85 == _T_308[7:0] ? 4'h6 : _GEN_6627; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6629 = 8'h86 == _T_308[7:0] ? 4'he : _GEN_6628; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6630 = 8'h87 == _T_308[7:0] ? 4'ha : _GEN_6629; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6631 = 8'h88 == _T_308[7:0] ? 4'h6 : _GEN_6630; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6632 = 8'h89 == _T_308[7:0] ? 4'ha : _GEN_6631; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6633 = 8'h8a == _T_308[7:0] ? 4'he : _GEN_6632; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6634 = 8'h8b == _T_308[7:0] ? 4'h3 : _GEN_6633; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6635 = 8'h8c == _T_308[7:0] ? 4'h3 : _GEN_6634; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6636 = 8'h8d == _T_308[7:0] ? 4'h0 : _GEN_6635; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6637 = 8'h8e == _T_308[7:0] ? 4'h2 : _GEN_6636; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6638 = 8'h8f == _T_308[7:0] ? 4'h0 : _GEN_6637; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6639 = 8'h90 == _T_308[7:0] ? 4'h0 : _GEN_6638; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6640 = 8'h91 == _T_308[7:0] ? 4'h0 : _GEN_6639; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6641 = 8'h92 == _T_308[7:0] ? 4'h0 : _GEN_6640; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6642 = 8'h93 == _T_308[7:0] ? 4'h0 : _GEN_6641; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6643 = 8'h94 == _T_308[7:0] ? 4'h0 : _GEN_6642; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6644 = 8'h95 == _T_308[7:0] ? 4'h0 : _GEN_6643; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6645 = 8'h96 == _T_308[7:0] ? 4'h0 : _GEN_6644; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6646 = 8'h97 == _T_308[7:0] ? 4'h2 : _GEN_6645; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6647 = 8'h98 == _T_308[7:0] ? 4'h2 : _GEN_6646; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6648 = 8'h99 == _T_308[7:0] ? 4'h1 : _GEN_6647; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6649 = 8'h9a == _T_308[7:0] ? 4'h3 : _GEN_6648; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6650 = 8'h9b == _T_308[7:0] ? 4'he : _GEN_6649; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6651 = 8'h9c == _T_308[7:0] ? 4'he : _GEN_6650; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6652 = 8'h9d == _T_308[7:0] ? 4'h0 : _GEN_6651; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6653 = 8'h9e == _T_308[7:0] ? 4'he : _GEN_6652; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6654 = 8'h9f == _T_308[7:0] ? 4'he : _GEN_6653; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6655 = 8'ha0 == _T_308[7:0] ? 4'h3 : _GEN_6654; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6656 = 8'ha1 == _T_308[7:0] ? 4'h1 : _GEN_6655; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6657 = 8'ha2 == _T_308[7:0] ? 4'h2 : _GEN_6656; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6658 = 8'ha3 == _T_308[7:0] ? 4'h2 : _GEN_6657; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6659 = 8'ha4 == _T_308[7:0] ? 4'h0 : _GEN_6658; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6660 = 8'ha5 == _T_308[7:0] ? 4'h0 : _GEN_6659; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6661 = 8'ha6 == _T_308[7:0] ? 4'h0 : _GEN_6660; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6662 = 8'ha7 == _T_308[7:0] ? 4'h0 : _GEN_6661; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6663 = 8'ha8 == _T_308[7:0] ? 4'h0 : _GEN_6662; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6664 = 8'ha9 == _T_308[7:0] ? 4'h0 : _GEN_6663; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6665 = 8'haa == _T_308[7:0] ? 4'h0 : _GEN_6664; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6666 = 8'hab == _T_308[7:0] ? 4'h0 : _GEN_6665; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6667 = 8'hac == _T_308[7:0] ? 4'h2 : _GEN_6666; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6668 = 8'had == _T_308[7:0] ? 4'h3 : _GEN_6667; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6669 = 8'hae == _T_308[7:0] ? 4'h4 : _GEN_6668; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6670 = 8'haf == _T_308[7:0] ? 4'h3 : _GEN_6669; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6671 = 8'hb0 == _T_308[7:0] ? 4'h4 : _GEN_6670; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6672 = 8'hb1 == _T_308[7:0] ? 4'h3 : _GEN_6671; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6673 = 8'hb2 == _T_308[7:0] ? 4'h0 : _GEN_6672; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6674 = 8'hb3 == _T_308[7:0] ? 4'h3 : _GEN_6673; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6675 = 8'hb4 == _T_308[7:0] ? 4'h4 : _GEN_6674; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6676 = 8'hb5 == _T_308[7:0] ? 4'h3 : _GEN_6675; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6677 = 8'hb6 == _T_308[7:0] ? 4'h4 : _GEN_6676; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6678 = 8'hb7 == _T_308[7:0] ? 4'h3 : _GEN_6677; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6679 = 8'hb8 == _T_308[7:0] ? 4'h2 : _GEN_6678; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6680 = 8'hb9 == _T_308[7:0] ? 4'h0 : _GEN_6679; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6681 = 8'hba == _T_308[7:0] ? 4'h0 : _GEN_6680; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6682 = 8'hbb == _T_308[7:0] ? 4'h0 : _GEN_6681; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6683 = 8'hbc == _T_308[7:0] ? 4'h0 : _GEN_6682; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6684 = 8'hbd == _T_308[7:0] ? 4'h0 : _GEN_6683; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6685 = 8'hbe == _T_308[7:0] ? 4'h0 : _GEN_6684; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6686 = 8'hbf == _T_308[7:0] ? 4'h0 : _GEN_6685; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6687 = 8'hc0 == _T_308[7:0] ? 4'h0 : _GEN_6686; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6688 = 8'hc1 == _T_308[7:0] ? 4'h0 : _GEN_6687; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6689 = 8'hc2 == _T_308[7:0] ? 4'h8 : _GEN_6688; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6690 = 8'hc3 == _T_308[7:0] ? 4'hc : _GEN_6689; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6691 = 8'hc4 == _T_308[7:0] ? 4'h0 : _GEN_6690; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6692 = 8'hc5 == _T_308[7:0] ? 4'h2 : _GEN_6691; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6693 = 8'hc6 == _T_308[7:0] ? 4'h3 : _GEN_6692; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6694 = 8'hc7 == _T_308[7:0] ? 4'h2 : _GEN_6693; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6695 = 8'hc8 == _T_308[7:0] ? 4'h3 : _GEN_6694; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6696 = 8'hc9 == _T_308[7:0] ? 4'h2 : _GEN_6695; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6697 = 8'hca == _T_308[7:0] ? 4'h0 : _GEN_6696; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6698 = 8'hcb == _T_308[7:0] ? 4'hc : _GEN_6697; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6699 = 8'hcc == _T_308[7:0] ? 4'h8 : _GEN_6698; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6700 = 8'hcd == _T_308[7:0] ? 4'h0 : _GEN_6699; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6701 = 8'hce == _T_308[7:0] ? 4'h0 : _GEN_6700; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6702 = 8'hcf == _T_308[7:0] ? 4'h0 : _GEN_6701; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6703 = 8'hd0 == _T_308[7:0] ? 4'h0 : _GEN_6702; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6704 = 8'hd1 == _T_308[7:0] ? 4'h0 : _GEN_6703; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6705 = 8'hd2 == _T_308[7:0] ? 4'h0 : _GEN_6704; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6706 = 8'hd3 == _T_308[7:0] ? 4'h0 : _GEN_6705; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6707 = 8'hd4 == _T_308[7:0] ? 4'h0 : _GEN_6706; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6708 = 8'hd5 == _T_308[7:0] ? 4'h0 : _GEN_6707; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6709 = 8'hd6 == _T_308[7:0] ? 4'h0 : _GEN_6708; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6710 = 8'hd7 == _T_308[7:0] ? 4'h3 : _GEN_6709; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6711 = 8'hd8 == _T_308[7:0] ? 4'h6 : _GEN_6710; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6712 = 8'hd9 == _T_308[7:0] ? 4'h0 : _GEN_6711; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6713 = 8'hda == _T_308[7:0] ? 4'hb : _GEN_6712; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6714 = 8'hdb == _T_308[7:0] ? 4'h1 : _GEN_6713; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6715 = 8'hdc == _T_308[7:0] ? 4'h4 : _GEN_6714; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6716 = 8'hdd == _T_308[7:0] ? 4'h1 : _GEN_6715; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6717 = 8'hde == _T_308[7:0] ? 4'hb : _GEN_6716; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6718 = 8'hdf == _T_308[7:0] ? 4'h0 : _GEN_6717; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6719 = 8'he0 == _T_308[7:0] ? 4'h6 : _GEN_6718; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6720 = 8'he1 == _T_308[7:0] ? 4'h3 : _GEN_6719; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6721 = 8'he2 == _T_308[7:0] ? 4'h0 : _GEN_6720; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6722 = 8'he3 == _T_308[7:0] ? 4'h0 : _GEN_6721; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6723 = 8'he4 == _T_308[7:0] ? 4'h0 : _GEN_6722; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6724 = 8'he5 == _T_308[7:0] ? 4'h0 : _GEN_6723; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6725 = 8'he6 == _T_308[7:0] ? 4'h0 : _GEN_6724; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6726 = 8'he7 == _T_308[7:0] ? 4'h0 : _GEN_6725; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6727 = 8'he8 == _T_308[7:0] ? 4'h0 : _GEN_6726; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6728 = 8'he9 == _T_308[7:0] ? 4'h0 : _GEN_6727; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6729 = 8'hea == _T_308[7:0] ? 4'h0 : _GEN_6728; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6730 = 8'heb == _T_308[7:0] ? 4'h0 : _GEN_6729; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6731 = 8'hec == _T_308[7:0] ? 4'h0 : _GEN_6730; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6732 = 8'hed == _T_308[7:0] ? 4'h0 : _GEN_6731; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6733 = 8'hee == _T_308[7:0] ? 4'h0 : _GEN_6732; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6734 = 8'hef == _T_308[7:0] ? 4'h0 : _GEN_6733; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6735 = 8'hf0 == _T_308[7:0] ? 4'h0 : _GEN_6734; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6736 = 8'hf1 == _T_308[7:0] ? 4'h0 : _GEN_6735; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6737 = 8'hf2 == _T_308[7:0] ? 4'h0 : _GEN_6736; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6738 = 8'hf3 == _T_308[7:0] ? 4'h0 : _GEN_6737; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6739 = 8'hf4 == _T_308[7:0] ? 4'h0 : _GEN_6738; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6740 = 8'hf5 == _T_308[7:0] ? 4'h0 : _GEN_6739; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6741 = 8'hf6 == _T_308[7:0] ? 4'h0 : _GEN_6740; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6742 = 8'hf7 == _T_308[7:0] ? 4'h0 : _GEN_6741; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6743 = 8'hf8 == _T_308[7:0] ? 4'h0 : _GEN_6742; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6744 = 8'hf9 == _T_308[7:0] ? 4'h0 : _GEN_6743; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6745 = 8'hfa == _T_308[7:0] ? 4'h0 : _GEN_6744; // @[Filter.scala 204:102]
  wire [3:0] _GEN_6746 = 8'hfb == _T_308[7:0] ? 4'h0 : _GEN_6745; // @[Filter.scala 204:102]
  wire [6:0] _GEN_11263 = {{3'd0}, _GEN_6746}; // @[Filter.scala 204:102]
  wire [10:0] _T_315 = _GEN_11263 * 7'h46; // @[Filter.scala 204:102]
  wire [10:0] _GEN_11264 = {{2'd0}, _T_310}; // @[Filter.scala 204:69]
  wire [10:0] _T_317 = _GEN_11264 + _T_315; // @[Filter.scala 204:69]
  wire [3:0] _GEN_6755 = 8'h8 == _T_308[7:0] ? 4'h3 : 4'h0; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6756 = 8'h9 == _T_308[7:0] ? 4'h6 : _GEN_6755; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6757 = 8'ha == _T_308[7:0] ? 4'h6 : _GEN_6756; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6758 = 8'hb == _T_308[7:0] ? 4'h6 : _GEN_6757; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6759 = 8'hc == _T_308[7:0] ? 4'h3 : _GEN_6758; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6760 = 8'hd == _T_308[7:0] ? 4'h0 : _GEN_6759; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6761 = 8'he == _T_308[7:0] ? 4'h0 : _GEN_6760; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6762 = 8'hf == _T_308[7:0] ? 4'h0 : _GEN_6761; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6763 = 8'h10 == _T_308[7:0] ? 4'h0 : _GEN_6762; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6764 = 8'h11 == _T_308[7:0] ? 4'h0 : _GEN_6763; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6765 = 8'h12 == _T_308[7:0] ? 4'h0 : _GEN_6764; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6766 = 8'h13 == _T_308[7:0] ? 4'h0 : _GEN_6765; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6767 = 8'h14 == _T_308[7:0] ? 4'h0 : _GEN_6766; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6768 = 8'h15 == _T_308[7:0] ? 4'h0 : _GEN_6767; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6769 = 8'h16 == _T_308[7:0] ? 4'h0 : _GEN_6768; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6770 = 8'h17 == _T_308[7:0] ? 4'h0 : _GEN_6769; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6771 = 8'h18 == _T_308[7:0] ? 4'h0 : _GEN_6770; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6772 = 8'h19 == _T_308[7:0] ? 4'h0 : _GEN_6771; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6773 = 8'h1a == _T_308[7:0] ? 4'h0 : _GEN_6772; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6774 = 8'h1b == _T_308[7:0] ? 4'h0 : _GEN_6773; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6775 = 8'h1c == _T_308[7:0] ? 4'h6 : _GEN_6774; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6776 = 8'h1d == _T_308[7:0] ? 4'h3 : _GEN_6775; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6777 = 8'h1e == _T_308[7:0] ? 4'h0 : _GEN_6776; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6778 = 8'h1f == _T_308[7:0] ? 4'h0 : _GEN_6777; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6779 = 8'h20 == _T_308[7:0] ? 4'h0 : _GEN_6778; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6780 = 8'h21 == _T_308[7:0] ? 4'h3 : _GEN_6779; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6781 = 8'h22 == _T_308[7:0] ? 4'h6 : _GEN_6780; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6782 = 8'h23 == _T_308[7:0] ? 4'h0 : _GEN_6781; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6783 = 8'h24 == _T_308[7:0] ? 4'h0 : _GEN_6782; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6784 = 8'h25 == _T_308[7:0] ? 4'h0 : _GEN_6783; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6785 = 8'h26 == _T_308[7:0] ? 4'h0 : _GEN_6784; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6786 = 8'h27 == _T_308[7:0] ? 4'h0 : _GEN_6785; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6787 = 8'h28 == _T_308[7:0] ? 4'h0 : _GEN_6786; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6788 = 8'h29 == _T_308[7:0] ? 4'h0 : _GEN_6787; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6789 = 8'h2a == _T_308[7:0] ? 4'h0 : _GEN_6788; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6790 = 8'h2b == _T_308[7:0] ? 4'h0 : _GEN_6789; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6791 = 8'h2c == _T_308[7:0] ? 4'h0 : _GEN_6790; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6792 = 8'h2d == _T_308[7:0] ? 4'h0 : _GEN_6791; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6793 = 8'h2e == _T_308[7:0] ? 4'h0 : _GEN_6792; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6794 = 8'h2f == _T_308[7:0] ? 4'h0 : _GEN_6793; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6795 = 8'h30 == _T_308[7:0] ? 4'h6 : _GEN_6794; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6796 = 8'h31 == _T_308[7:0] ? 4'h3 : _GEN_6795; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6797 = 8'h32 == _T_308[7:0] ? 4'h0 : _GEN_6796; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6798 = 8'h33 == _T_308[7:0] ? 4'h1 : _GEN_6797; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6799 = 8'h34 == _T_308[7:0] ? 4'h1 : _GEN_6798; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6800 = 8'h35 == _T_308[7:0] ? 4'h0 : _GEN_6799; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6801 = 8'h36 == _T_308[7:0] ? 4'h0 : _GEN_6800; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6802 = 8'h37 == _T_308[7:0] ? 4'h0 : _GEN_6801; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6803 = 8'h38 == _T_308[7:0] ? 4'h6 : _GEN_6802; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6804 = 8'h39 == _T_308[7:0] ? 4'h0 : _GEN_6803; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6805 = 8'h3a == _T_308[7:0] ? 4'h0 : _GEN_6804; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6806 = 8'h3b == _T_308[7:0] ? 4'h0 : _GEN_6805; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6807 = 8'h3c == _T_308[7:0] ? 4'h0 : _GEN_6806; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6808 = 8'h3d == _T_308[7:0] ? 4'h0 : _GEN_6807; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6809 = 8'h3e == _T_308[7:0] ? 4'h0 : _GEN_6808; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6810 = 8'h3f == _T_308[7:0] ? 4'h0 : _GEN_6809; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6811 = 8'h40 == _T_308[7:0] ? 4'h0 : _GEN_6810; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6812 = 8'h41 == _T_308[7:0] ? 4'h0 : _GEN_6811; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6813 = 8'h42 == _T_308[7:0] ? 4'h0 : _GEN_6812; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6814 = 8'h43 == _T_308[7:0] ? 4'h0 : _GEN_6813; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6815 = 8'h44 == _T_308[7:0] ? 4'h3 : _GEN_6814; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6816 = 8'h45 == _T_308[7:0] ? 4'h6 : _GEN_6815; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6817 = 8'h46 == _T_308[7:0] ? 4'h9 : _GEN_6816; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6818 = 8'h47 == _T_308[7:0] ? 4'h0 : _GEN_6817; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6819 = 8'h48 == _T_308[7:0] ? 4'h0 : _GEN_6818; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6820 = 8'h49 == _T_308[7:0] ? 4'h0 : _GEN_6819; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6821 = 8'h4a == _T_308[7:0] ? 4'h1 : _GEN_6820; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6822 = 8'h4b == _T_308[7:0] ? 4'h0 : _GEN_6821; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6823 = 8'h4c == _T_308[7:0] ? 4'h0 : _GEN_6822; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6824 = 8'h4d == _T_308[7:0] ? 4'h0 : _GEN_6823; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6825 = 8'h4e == _T_308[7:0] ? 4'h6 : _GEN_6824; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6826 = 8'h4f == _T_308[7:0] ? 4'h0 : _GEN_6825; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6827 = 8'h50 == _T_308[7:0] ? 4'h0 : _GEN_6826; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6828 = 8'h51 == _T_308[7:0] ? 4'h0 : _GEN_6827; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6829 = 8'h52 == _T_308[7:0] ? 4'h0 : _GEN_6828; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6830 = 8'h53 == _T_308[7:0] ? 4'h0 : _GEN_6829; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6831 = 8'h54 == _T_308[7:0] ? 4'h0 : _GEN_6830; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6832 = 8'h55 == _T_308[7:0] ? 4'h0 : _GEN_6831; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6833 = 8'h56 == _T_308[7:0] ? 4'h0 : _GEN_6832; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6834 = 8'h57 == _T_308[7:0] ? 4'h0 : _GEN_6833; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6835 = 8'h58 == _T_308[7:0] ? 4'h0 : _GEN_6834; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6836 = 8'h59 == _T_308[7:0] ? 4'h6 : _GEN_6835; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6837 = 8'h5a == _T_308[7:0] ? 4'h3 : _GEN_6836; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6838 = 8'h5b == _T_308[7:0] ? 4'h0 : _GEN_6837; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6839 = 8'h5c == _T_308[7:0] ? 4'h0 : _GEN_6838; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6840 = 8'h5d == _T_308[7:0] ? 4'h0 : _GEN_6839; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6841 = 8'h5e == _T_308[7:0] ? 4'h7 : _GEN_6840; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6842 = 8'h5f == _T_308[7:0] ? 4'h0 : _GEN_6841; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6843 = 8'h60 == _T_308[7:0] ? 4'h0 : _GEN_6842; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6844 = 8'h61 == _T_308[7:0] ? 4'h1 : _GEN_6843; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6845 = 8'h62 == _T_308[7:0] ? 4'h0 : _GEN_6844; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6846 = 8'h63 == _T_308[7:0] ? 4'h6 : _GEN_6845; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6847 = 8'h64 == _T_308[7:0] ? 4'h0 : _GEN_6846; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6848 = 8'h65 == _T_308[7:0] ? 4'h0 : _GEN_6847; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6849 = 8'h66 == _T_308[7:0] ? 4'h0 : _GEN_6848; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6850 = 8'h67 == _T_308[7:0] ? 4'h0 : _GEN_6849; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6851 = 8'h68 == _T_308[7:0] ? 4'h0 : _GEN_6850; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6852 = 8'h69 == _T_308[7:0] ? 4'h0 : _GEN_6851; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6853 = 8'h6a == _T_308[7:0] ? 4'h0 : _GEN_6852; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6854 = 8'h6b == _T_308[7:0] ? 4'h0 : _GEN_6853; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6855 = 8'h6c == _T_308[7:0] ? 4'h0 : _GEN_6854; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6856 = 8'h6d == _T_308[7:0] ? 4'h0 : _GEN_6855; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6857 = 8'h6e == _T_308[7:0] ? 4'h6 : _GEN_6856; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6858 = 8'h6f == _T_308[7:0] ? 4'h0 : _GEN_6857; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6859 = 8'h70 == _T_308[7:0] ? 4'h0 : _GEN_6858; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6860 = 8'h71 == _T_308[7:0] ? 4'h0 : _GEN_6859; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6861 = 8'h72 == _T_308[7:0] ? 4'h3 : _GEN_6860; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6862 = 8'h73 == _T_308[7:0] ? 4'hc : _GEN_6861; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6863 = 8'h74 == _T_308[7:0] ? 4'h3 : _GEN_6862; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6864 = 8'h75 == _T_308[7:0] ? 4'h0 : _GEN_6863; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6865 = 8'h76 == _T_308[7:0] ? 4'h1 : _GEN_6864; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6866 = 8'h77 == _T_308[7:0] ? 4'h0 : _GEN_6865; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6867 = 8'h78 == _T_308[7:0] ? 4'h3 : _GEN_6866; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6868 = 8'h79 == _T_308[7:0] ? 4'h3 : _GEN_6867; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6869 = 8'h7a == _T_308[7:0] ? 4'h0 : _GEN_6868; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6870 = 8'h7b == _T_308[7:0] ? 4'h0 : _GEN_6869; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6871 = 8'h7c == _T_308[7:0] ? 4'h0 : _GEN_6870; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6872 = 8'h7d == _T_308[7:0] ? 4'h0 : _GEN_6871; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6873 = 8'h7e == _T_308[7:0] ? 4'h0 : _GEN_6872; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6874 = 8'h7f == _T_308[7:0] ? 4'h0 : _GEN_6873; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6875 = 8'h80 == _T_308[7:0] ? 4'h0 : _GEN_6874; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6876 = 8'h81 == _T_308[7:0] ? 4'h0 : _GEN_6875; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6877 = 8'h82 == _T_308[7:0] ? 4'h6 : _GEN_6876; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6878 = 8'h83 == _T_308[7:0] ? 4'h0 : _GEN_6877; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6879 = 8'h84 == _T_308[7:0] ? 4'h1 : _GEN_6878; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6880 = 8'h85 == _T_308[7:0] ? 4'h1 : _GEN_6879; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6881 = 8'h86 == _T_308[7:0] ? 4'ha : _GEN_6880; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6882 = 8'h87 == _T_308[7:0] ? 4'h4 : _GEN_6881; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6883 = 8'h88 == _T_308[7:0] ? 4'h1 : _GEN_6882; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6884 = 8'h89 == _T_308[7:0] ? 4'h4 : _GEN_6883; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6885 = 8'h8a == _T_308[7:0] ? 4'ha : _GEN_6884; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6886 = 8'h8b == _T_308[7:0] ? 4'h0 : _GEN_6885; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6887 = 8'h8c == _T_308[7:0] ? 4'h0 : _GEN_6886; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6888 = 8'h8d == _T_308[7:0] ? 4'h0 : _GEN_6887; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6889 = 8'h8e == _T_308[7:0] ? 4'h6 : _GEN_6888; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6890 = 8'h8f == _T_308[7:0] ? 4'h0 : _GEN_6889; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6891 = 8'h90 == _T_308[7:0] ? 4'h0 : _GEN_6890; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6892 = 8'h91 == _T_308[7:0] ? 4'h0 : _GEN_6891; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6893 = 8'h92 == _T_308[7:0] ? 4'h0 : _GEN_6892; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6894 = 8'h93 == _T_308[7:0] ? 4'h0 : _GEN_6893; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6895 = 8'h94 == _T_308[7:0] ? 4'h0 : _GEN_6894; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6896 = 8'h95 == _T_308[7:0] ? 4'h0 : _GEN_6895; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6897 = 8'h96 == _T_308[7:0] ? 4'h0 : _GEN_6896; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6898 = 8'h97 == _T_308[7:0] ? 4'h6 : _GEN_6897; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6899 = 8'h98 == _T_308[7:0] ? 4'h6 : _GEN_6898; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6900 = 8'h99 == _T_308[7:0] ? 4'h3 : _GEN_6899; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6901 = 8'h9a == _T_308[7:0] ? 4'h0 : _GEN_6900; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6902 = 8'h9b == _T_308[7:0] ? 4'ha : _GEN_6901; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6903 = 8'h9c == _T_308[7:0] ? 4'ha : _GEN_6902; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6904 = 8'h9d == _T_308[7:0] ? 4'h0 : _GEN_6903; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6905 = 8'h9e == _T_308[7:0] ? 4'ha : _GEN_6904; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6906 = 8'h9f == _T_308[7:0] ? 4'ha : _GEN_6905; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6907 = 8'ha0 == _T_308[7:0] ? 4'h0 : _GEN_6906; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6908 = 8'ha1 == _T_308[7:0] ? 4'h3 : _GEN_6907; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6909 = 8'ha2 == _T_308[7:0] ? 4'h6 : _GEN_6908; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6910 = 8'ha3 == _T_308[7:0] ? 4'h6 : _GEN_6909; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6911 = 8'ha4 == _T_308[7:0] ? 4'h0 : _GEN_6910; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6912 = 8'ha5 == _T_308[7:0] ? 4'h0 : _GEN_6911; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6913 = 8'ha6 == _T_308[7:0] ? 4'h0 : _GEN_6912; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6914 = 8'ha7 == _T_308[7:0] ? 4'h0 : _GEN_6913; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6915 = 8'ha8 == _T_308[7:0] ? 4'h0 : _GEN_6914; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6916 = 8'ha9 == _T_308[7:0] ? 4'h0 : _GEN_6915; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6917 = 8'haa == _T_308[7:0] ? 4'h0 : _GEN_6916; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6918 = 8'hab == _T_308[7:0] ? 4'h0 : _GEN_6917; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6919 = 8'hac == _T_308[7:0] ? 4'h6 : _GEN_6918; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6920 = 8'had == _T_308[7:0] ? 4'h0 : _GEN_6919; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6921 = 8'hae == _T_308[7:0] ? 4'h3 : _GEN_6920; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6922 = 8'haf == _T_308[7:0] ? 4'h9 : _GEN_6921; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6923 = 8'hb0 == _T_308[7:0] ? 4'h3 : _GEN_6922; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6924 = 8'hb1 == _T_308[7:0] ? 4'h0 : _GEN_6923; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6925 = 8'hb2 == _T_308[7:0] ? 4'h0 : _GEN_6924; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6926 = 8'hb3 == _T_308[7:0] ? 4'h0 : _GEN_6925; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6927 = 8'hb4 == _T_308[7:0] ? 4'h3 : _GEN_6926; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6928 = 8'hb5 == _T_308[7:0] ? 4'h9 : _GEN_6927; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6929 = 8'hb6 == _T_308[7:0] ? 4'h3 : _GEN_6928; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6930 = 8'hb7 == _T_308[7:0] ? 4'h0 : _GEN_6929; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6931 = 8'hb8 == _T_308[7:0] ? 4'h6 : _GEN_6930; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6932 = 8'hb9 == _T_308[7:0] ? 4'h0 : _GEN_6931; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6933 = 8'hba == _T_308[7:0] ? 4'h0 : _GEN_6932; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6934 = 8'hbb == _T_308[7:0] ? 4'h0 : _GEN_6933; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6935 = 8'hbc == _T_308[7:0] ? 4'h0 : _GEN_6934; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6936 = 8'hbd == _T_308[7:0] ? 4'h0 : _GEN_6935; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6937 = 8'hbe == _T_308[7:0] ? 4'h0 : _GEN_6936; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6938 = 8'hbf == _T_308[7:0] ? 4'h0 : _GEN_6937; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6939 = 8'hc0 == _T_308[7:0] ? 4'h0 : _GEN_6938; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6940 = 8'hc1 == _T_308[7:0] ? 4'h0 : _GEN_6939; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6941 = 8'hc2 == _T_308[7:0] ? 4'h7 : _GEN_6940; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6942 = 8'hc3 == _T_308[7:0] ? 4'h2 : _GEN_6941; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6943 = 8'hc4 == _T_308[7:0] ? 4'h0 : _GEN_6942; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6944 = 8'hc5 == _T_308[7:0] ? 4'h6 : _GEN_6943; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6945 = 8'hc6 == _T_308[7:0] ? 4'h9 : _GEN_6944; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6946 = 8'hc7 == _T_308[7:0] ? 4'h6 : _GEN_6945; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6947 = 8'hc8 == _T_308[7:0] ? 4'h9 : _GEN_6946; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6948 = 8'hc9 == _T_308[7:0] ? 4'h6 : _GEN_6947; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6949 = 8'hca == _T_308[7:0] ? 4'h0 : _GEN_6948; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6950 = 8'hcb == _T_308[7:0] ? 4'h2 : _GEN_6949; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6951 = 8'hcc == _T_308[7:0] ? 4'h7 : _GEN_6950; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6952 = 8'hcd == _T_308[7:0] ? 4'h0 : _GEN_6951; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6953 = 8'hce == _T_308[7:0] ? 4'h0 : _GEN_6952; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6954 = 8'hcf == _T_308[7:0] ? 4'h0 : _GEN_6953; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6955 = 8'hd0 == _T_308[7:0] ? 4'h0 : _GEN_6954; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6956 = 8'hd1 == _T_308[7:0] ? 4'h0 : _GEN_6955; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6957 = 8'hd2 == _T_308[7:0] ? 4'h0 : _GEN_6956; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6958 = 8'hd3 == _T_308[7:0] ? 4'h0 : _GEN_6957; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6959 = 8'hd4 == _T_308[7:0] ? 4'h0 : _GEN_6958; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6960 = 8'hd5 == _T_308[7:0] ? 4'h0 : _GEN_6959; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6961 = 8'hd6 == _T_308[7:0] ? 4'h0 : _GEN_6960; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6962 = 8'hd7 == _T_308[7:0] ? 4'h3 : _GEN_6961; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6963 = 8'hd8 == _T_308[7:0] ? 4'h3 : _GEN_6962; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6964 = 8'hd9 == _T_308[7:0] ? 4'h0 : _GEN_6963; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6965 = 8'hda == _T_308[7:0] ? 4'h9 : _GEN_6964; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6966 = 8'hdb == _T_308[7:0] ? 4'h3 : _GEN_6965; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6967 = 8'hdc == _T_308[7:0] ? 4'hc : _GEN_6966; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6968 = 8'hdd == _T_308[7:0] ? 4'h3 : _GEN_6967; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6969 = 8'hde == _T_308[7:0] ? 4'h9 : _GEN_6968; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6970 = 8'hdf == _T_308[7:0] ? 4'h0 : _GEN_6969; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6971 = 8'he0 == _T_308[7:0] ? 4'h3 : _GEN_6970; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6972 = 8'he1 == _T_308[7:0] ? 4'h3 : _GEN_6971; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6973 = 8'he2 == _T_308[7:0] ? 4'h0 : _GEN_6972; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6974 = 8'he3 == _T_308[7:0] ? 4'h0 : _GEN_6973; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6975 = 8'he4 == _T_308[7:0] ? 4'h0 : _GEN_6974; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6976 = 8'he5 == _T_308[7:0] ? 4'h0 : _GEN_6975; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6977 = 8'he6 == _T_308[7:0] ? 4'h0 : _GEN_6976; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6978 = 8'he7 == _T_308[7:0] ? 4'h0 : _GEN_6977; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6979 = 8'he8 == _T_308[7:0] ? 4'h0 : _GEN_6978; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6980 = 8'he9 == _T_308[7:0] ? 4'h0 : _GEN_6979; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6981 = 8'hea == _T_308[7:0] ? 4'h0 : _GEN_6980; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6982 = 8'heb == _T_308[7:0] ? 4'h0 : _GEN_6981; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6983 = 8'hec == _T_308[7:0] ? 4'h0 : _GEN_6982; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6984 = 8'hed == _T_308[7:0] ? 4'h0 : _GEN_6983; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6985 = 8'hee == _T_308[7:0] ? 4'h0 : _GEN_6984; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6986 = 8'hef == _T_308[7:0] ? 4'h0 : _GEN_6985; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6987 = 8'hf0 == _T_308[7:0] ? 4'h0 : _GEN_6986; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6988 = 8'hf1 == _T_308[7:0] ? 4'h0 : _GEN_6987; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6989 = 8'hf2 == _T_308[7:0] ? 4'h0 : _GEN_6988; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6990 = 8'hf3 == _T_308[7:0] ? 4'h0 : _GEN_6989; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6991 = 8'hf4 == _T_308[7:0] ? 4'h0 : _GEN_6990; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6992 = 8'hf5 == _T_308[7:0] ? 4'h0 : _GEN_6991; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6993 = 8'hf6 == _T_308[7:0] ? 4'h0 : _GEN_6992; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6994 = 8'hf7 == _T_308[7:0] ? 4'h0 : _GEN_6993; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6995 = 8'hf8 == _T_308[7:0] ? 4'h0 : _GEN_6994; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6996 = 8'hf9 == _T_308[7:0] ? 4'h0 : _GEN_6995; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6997 = 8'hfa == _T_308[7:0] ? 4'h0 : _GEN_6996; // @[Filter.scala 204:142]
  wire [3:0] _GEN_6998 = 8'hfb == _T_308[7:0] ? 4'h0 : _GEN_6997; // @[Filter.scala 204:142]
  wire [7:0] _T_322 = _GEN_6998 * 4'ha; // @[Filter.scala 204:142]
  wire [10:0] _GEN_11266 = {{3'd0}, _T_322}; // @[Filter.scala 204:109]
  wire [10:0] _T_324 = _T_317 + _GEN_11266; // @[Filter.scala 204:109]
  wire [10:0] _T_325 = _T_324 / 11'h64; // @[Filter.scala 204:150]
  wire  _T_327 = _T_298 >= 5'h15; // @[Filter.scala 207:31]
  wire  _T_331 = _T_305 >= 32'hc; // @[Filter.scala 207:63]
  wire  _T_332 = _T_327 | _T_331; // @[Filter.scala 207:58]
  wire [10:0] _GEN_7251 = io_SPI_distort ? _T_325 : {{7'd0}, _GEN_6494}; // @[Filter.scala 209:35]
  wire [10:0] _GEN_7252 = _T_332 ? 11'h0 : _GEN_7251; // @[Filter.scala 207:80]
  wire [10:0] _GEN_7505 = io_SPI_distort ? _T_325 : {{7'd0}, _GEN_6746}; // @[Filter.scala 209:35]
  wire [10:0] _GEN_7506 = _T_332 ? 11'h0 : _GEN_7505; // @[Filter.scala 207:80]
  wire [10:0] _GEN_7759 = io_SPI_distort ? _T_325 : {{7'd0}, _GEN_6998}; // @[Filter.scala 209:35]
  wire [10:0] _GEN_7760 = _T_332 ? 11'h0 : _GEN_7759; // @[Filter.scala 207:80]
  wire [31:0] _T_360 = pixelIndex + 32'h5; // @[Filter.scala 202:31]
  wire [31:0] _GEN_5 = _T_360 % 32'h15; // @[Filter.scala 202:38]
  wire [4:0] _T_361 = _GEN_5[4:0]; // @[Filter.scala 202:38]
  wire [4:0] _T_363 = _T_361 + _GEN_11210; // @[Filter.scala 202:53]
  wire [4:0] _T_365 = _T_363 - 5'h1; // @[Filter.scala 202:69]
  wire [31:0] _T_368 = _T_360 / 32'h15; // @[Filter.scala 203:38]
  wire [31:0] _T_370 = _T_368 + _GEN_11211; // @[Filter.scala 203:53]
  wire [31:0] _T_372 = _T_370 - 32'h1; // @[Filter.scala 203:69]
  wire [36:0] _T_373 = _T_372 * 32'h15; // @[Filter.scala 204:42]
  wire [36:0] _GEN_11272 = {{32'd0}, _T_365}; // @[Filter.scala 204:57]
  wire [36:0] _T_375 = _T_373 + _GEN_11272; // @[Filter.scala 204:57]
  wire [3:0] _GEN_7769 = 8'h8 == _T_375[7:0] ? 4'h1 : 4'h0; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7770 = 8'h9 == _T_375[7:0] ? 4'h2 : _GEN_7769; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7771 = 8'ha == _T_375[7:0] ? 4'h2 : _GEN_7770; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7772 = 8'hb == _T_375[7:0] ? 4'h2 : _GEN_7771; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7773 = 8'hc == _T_375[7:0] ? 4'h1 : _GEN_7772; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7774 = 8'hd == _T_375[7:0] ? 4'h0 : _GEN_7773; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7775 = 8'he == _T_375[7:0] ? 4'h0 : _GEN_7774; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7776 = 8'hf == _T_375[7:0] ? 4'h0 : _GEN_7775; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7777 = 8'h10 == _T_375[7:0] ? 4'h0 : _GEN_7776; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7778 = 8'h11 == _T_375[7:0] ? 4'h0 : _GEN_7777; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7779 = 8'h12 == _T_375[7:0] ? 4'h0 : _GEN_7778; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7780 = 8'h13 == _T_375[7:0] ? 4'h0 : _GEN_7779; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7781 = 8'h14 == _T_375[7:0] ? 4'h0 : _GEN_7780; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7782 = 8'h15 == _T_375[7:0] ? 4'h0 : _GEN_7781; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7783 = 8'h16 == _T_375[7:0] ? 4'h0 : _GEN_7782; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7784 = 8'h17 == _T_375[7:0] ? 4'h0 : _GEN_7783; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7785 = 8'h18 == _T_375[7:0] ? 4'h0 : _GEN_7784; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7786 = 8'h19 == _T_375[7:0] ? 4'h0 : _GEN_7785; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7787 = 8'h1a == _T_375[7:0] ? 4'h0 : _GEN_7786; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7788 = 8'h1b == _T_375[7:0] ? 4'h0 : _GEN_7787; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7789 = 8'h1c == _T_375[7:0] ? 4'h2 : _GEN_7788; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7790 = 8'h1d == _T_375[7:0] ? 4'h1 : _GEN_7789; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7791 = 8'h1e == _T_375[7:0] ? 4'h0 : _GEN_7790; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7792 = 8'h1f == _T_375[7:0] ? 4'h0 : _GEN_7791; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7793 = 8'h20 == _T_375[7:0] ? 4'h0 : _GEN_7792; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7794 = 8'h21 == _T_375[7:0] ? 4'h1 : _GEN_7793; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7795 = 8'h22 == _T_375[7:0] ? 4'h2 : _GEN_7794; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7796 = 8'h23 == _T_375[7:0] ? 4'h0 : _GEN_7795; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7797 = 8'h24 == _T_375[7:0] ? 4'h0 : _GEN_7796; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7798 = 8'h25 == _T_375[7:0] ? 4'h0 : _GEN_7797; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7799 = 8'h26 == _T_375[7:0] ? 4'h0 : _GEN_7798; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7800 = 8'h27 == _T_375[7:0] ? 4'h0 : _GEN_7799; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7801 = 8'h28 == _T_375[7:0] ? 4'h0 : _GEN_7800; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7802 = 8'h29 == _T_375[7:0] ? 4'h0 : _GEN_7801; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7803 = 8'h2a == _T_375[7:0] ? 4'h0 : _GEN_7802; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7804 = 8'h2b == _T_375[7:0] ? 4'h0 : _GEN_7803; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7805 = 8'h2c == _T_375[7:0] ? 4'h0 : _GEN_7804; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7806 = 8'h2d == _T_375[7:0] ? 4'h0 : _GEN_7805; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7807 = 8'h2e == _T_375[7:0] ? 4'h0 : _GEN_7806; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7808 = 8'h2f == _T_375[7:0] ? 4'h0 : _GEN_7807; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7809 = 8'h30 == _T_375[7:0] ? 4'h2 : _GEN_7808; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7810 = 8'h31 == _T_375[7:0] ? 4'h2 : _GEN_7809; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7811 = 8'h32 == _T_375[7:0] ? 4'h0 : _GEN_7810; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7812 = 8'h33 == _T_375[7:0] ? 4'h0 : _GEN_7811; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7813 = 8'h34 == _T_375[7:0] ? 4'h0 : _GEN_7812; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7814 = 8'h35 == _T_375[7:0] ? 4'h0 : _GEN_7813; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7815 = 8'h36 == _T_375[7:0] ? 4'h0 : _GEN_7814; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7816 = 8'h37 == _T_375[7:0] ? 4'h0 : _GEN_7815; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7817 = 8'h38 == _T_375[7:0] ? 4'h2 : _GEN_7816; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7818 = 8'h39 == _T_375[7:0] ? 4'h0 : _GEN_7817; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7819 = 8'h3a == _T_375[7:0] ? 4'h0 : _GEN_7818; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7820 = 8'h3b == _T_375[7:0] ? 4'h0 : _GEN_7819; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7821 = 8'h3c == _T_375[7:0] ? 4'h0 : _GEN_7820; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7822 = 8'h3d == _T_375[7:0] ? 4'h0 : _GEN_7821; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7823 = 8'h3e == _T_375[7:0] ? 4'h0 : _GEN_7822; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7824 = 8'h3f == _T_375[7:0] ? 4'h0 : _GEN_7823; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7825 = 8'h40 == _T_375[7:0] ? 4'h0 : _GEN_7824; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7826 = 8'h41 == _T_375[7:0] ? 4'h0 : _GEN_7825; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7827 = 8'h42 == _T_375[7:0] ? 4'h0 : _GEN_7826; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7828 = 8'h43 == _T_375[7:0] ? 4'h0 : _GEN_7827; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7829 = 8'h44 == _T_375[7:0] ? 4'h1 : _GEN_7828; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7830 = 8'h45 == _T_375[7:0] ? 4'h3 : _GEN_7829; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7831 = 8'h46 == _T_375[7:0] ? 4'h7 : _GEN_7830; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7832 = 8'h47 == _T_375[7:0] ? 4'h0 : _GEN_7831; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7833 = 8'h48 == _T_375[7:0] ? 4'h0 : _GEN_7832; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7834 = 8'h49 == _T_375[7:0] ? 4'h0 : _GEN_7833; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7835 = 8'h4a == _T_375[7:0] ? 4'h0 : _GEN_7834; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7836 = 8'h4b == _T_375[7:0] ? 4'h0 : _GEN_7835; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7837 = 8'h4c == _T_375[7:0] ? 4'h0 : _GEN_7836; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7838 = 8'h4d == _T_375[7:0] ? 4'h0 : _GEN_7837; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7839 = 8'h4e == _T_375[7:0] ? 4'h2 : _GEN_7838; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7840 = 8'h4f == _T_375[7:0] ? 4'h0 : _GEN_7839; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7841 = 8'h50 == _T_375[7:0] ? 4'h0 : _GEN_7840; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7842 = 8'h51 == _T_375[7:0] ? 4'h0 : _GEN_7841; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7843 = 8'h52 == _T_375[7:0] ? 4'h0 : _GEN_7842; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7844 = 8'h53 == _T_375[7:0] ? 4'h0 : _GEN_7843; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7845 = 8'h54 == _T_375[7:0] ? 4'h0 : _GEN_7844; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7846 = 8'h55 == _T_375[7:0] ? 4'h0 : _GEN_7845; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7847 = 8'h56 == _T_375[7:0] ? 4'h0 : _GEN_7846; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7848 = 8'h57 == _T_375[7:0] ? 4'h0 : _GEN_7847; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7849 = 8'h58 == _T_375[7:0] ? 4'h0 : _GEN_7848; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7850 = 8'h59 == _T_375[7:0] ? 4'h2 : _GEN_7849; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7851 = 8'h5a == _T_375[7:0] ? 4'h2 : _GEN_7850; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7852 = 8'h5b == _T_375[7:0] ? 4'h0 : _GEN_7851; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7853 = 8'h5c == _T_375[7:0] ? 4'h0 : _GEN_7852; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7854 = 8'h5d == _T_375[7:0] ? 4'h0 : _GEN_7853; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7855 = 8'h5e == _T_375[7:0] ? 4'h4 : _GEN_7854; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7856 = 8'h5f == _T_375[7:0] ? 4'h0 : _GEN_7855; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7857 = 8'h60 == _T_375[7:0] ? 4'h0 : _GEN_7856; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7858 = 8'h61 == _T_375[7:0] ? 4'h0 : _GEN_7857; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7859 = 8'h62 == _T_375[7:0] ? 4'h0 : _GEN_7858; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7860 = 8'h63 == _T_375[7:0] ? 4'h2 : _GEN_7859; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7861 = 8'h64 == _T_375[7:0] ? 4'h0 : _GEN_7860; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7862 = 8'h65 == _T_375[7:0] ? 4'h0 : _GEN_7861; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7863 = 8'h66 == _T_375[7:0] ? 4'h0 : _GEN_7862; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7864 = 8'h67 == _T_375[7:0] ? 4'h0 : _GEN_7863; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7865 = 8'h68 == _T_375[7:0] ? 4'h0 : _GEN_7864; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7866 = 8'h69 == _T_375[7:0] ? 4'h0 : _GEN_7865; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7867 = 8'h6a == _T_375[7:0] ? 4'h0 : _GEN_7866; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7868 = 8'h6b == _T_375[7:0] ? 4'h0 : _GEN_7867; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7869 = 8'h6c == _T_375[7:0] ? 4'h0 : _GEN_7868; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7870 = 8'h6d == _T_375[7:0] ? 4'h0 : _GEN_7869; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7871 = 8'h6e == _T_375[7:0] ? 4'h2 : _GEN_7870; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7872 = 8'h6f == _T_375[7:0] ? 4'h0 : _GEN_7871; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7873 = 8'h70 == _T_375[7:0] ? 4'h0 : _GEN_7872; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7874 = 8'h71 == _T_375[7:0] ? 4'h0 : _GEN_7873; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7875 = 8'h72 == _T_375[7:0] ? 4'h2 : _GEN_7874; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7876 = 8'h73 == _T_375[7:0] ? 4'h9 : _GEN_7875; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7877 = 8'h74 == _T_375[7:0] ? 4'h2 : _GEN_7876; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7878 = 8'h75 == _T_375[7:0] ? 4'h0 : _GEN_7877; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7879 = 8'h76 == _T_375[7:0] ? 4'h0 : _GEN_7878; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7880 = 8'h77 == _T_375[7:0] ? 4'h0 : _GEN_7879; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7881 = 8'h78 == _T_375[7:0] ? 4'h1 : _GEN_7880; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7882 = 8'h79 == _T_375[7:0] ? 4'h1 : _GEN_7881; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7883 = 8'h7a == _T_375[7:0] ? 4'h0 : _GEN_7882; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7884 = 8'h7b == _T_375[7:0] ? 4'h0 : _GEN_7883; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7885 = 8'h7c == _T_375[7:0] ? 4'h0 : _GEN_7884; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7886 = 8'h7d == _T_375[7:0] ? 4'h0 : _GEN_7885; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7887 = 8'h7e == _T_375[7:0] ? 4'h0 : _GEN_7886; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7888 = 8'h7f == _T_375[7:0] ? 4'h0 : _GEN_7887; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7889 = 8'h80 == _T_375[7:0] ? 4'h0 : _GEN_7888; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7890 = 8'h81 == _T_375[7:0] ? 4'h0 : _GEN_7889; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7891 = 8'h82 == _T_375[7:0] ? 4'h2 : _GEN_7890; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7892 = 8'h83 == _T_375[7:0] ? 4'h0 : _GEN_7891; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7893 = 8'h84 == _T_375[7:0] ? 4'h0 : _GEN_7892; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7894 = 8'h85 == _T_375[7:0] ? 4'h0 : _GEN_7893; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7895 = 8'h86 == _T_375[7:0] ? 4'h7 : _GEN_7894; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7896 = 8'h87 == _T_375[7:0] ? 4'h2 : _GEN_7895; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7897 = 8'h88 == _T_375[7:0] ? 4'h0 : _GEN_7896; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7898 = 8'h89 == _T_375[7:0] ? 4'h2 : _GEN_7897; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7899 = 8'h8a == _T_375[7:0] ? 4'h7 : _GEN_7898; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7900 = 8'h8b == _T_375[7:0] ? 4'h0 : _GEN_7899; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7901 = 8'h8c == _T_375[7:0] ? 4'h0 : _GEN_7900; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7902 = 8'h8d == _T_375[7:0] ? 4'h0 : _GEN_7901; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7903 = 8'h8e == _T_375[7:0] ? 4'h2 : _GEN_7902; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7904 = 8'h8f == _T_375[7:0] ? 4'h0 : _GEN_7903; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7905 = 8'h90 == _T_375[7:0] ? 4'h0 : _GEN_7904; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7906 = 8'h91 == _T_375[7:0] ? 4'h0 : _GEN_7905; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7907 = 8'h92 == _T_375[7:0] ? 4'h0 : _GEN_7906; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7908 = 8'h93 == _T_375[7:0] ? 4'h0 : _GEN_7907; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7909 = 8'h94 == _T_375[7:0] ? 4'h0 : _GEN_7908; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7910 = 8'h95 == _T_375[7:0] ? 4'h0 : _GEN_7909; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7911 = 8'h96 == _T_375[7:0] ? 4'h0 : _GEN_7910; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7912 = 8'h97 == _T_375[7:0] ? 4'h2 : _GEN_7911; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7913 = 8'h98 == _T_375[7:0] ? 4'h2 : _GEN_7912; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7914 = 8'h99 == _T_375[7:0] ? 4'h1 : _GEN_7913; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7915 = 8'h9a == _T_375[7:0] ? 4'h0 : _GEN_7914; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7916 = 8'h9b == _T_375[7:0] ? 4'h7 : _GEN_7915; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7917 = 8'h9c == _T_375[7:0] ? 4'h7 : _GEN_7916; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7918 = 8'h9d == _T_375[7:0] ? 4'h0 : _GEN_7917; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7919 = 8'h9e == _T_375[7:0] ? 4'h7 : _GEN_7918; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7920 = 8'h9f == _T_375[7:0] ? 4'h7 : _GEN_7919; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7921 = 8'ha0 == _T_375[7:0] ? 4'h0 : _GEN_7920; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7922 = 8'ha1 == _T_375[7:0] ? 4'h1 : _GEN_7921; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7923 = 8'ha2 == _T_375[7:0] ? 4'h2 : _GEN_7922; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7924 = 8'ha3 == _T_375[7:0] ? 4'h2 : _GEN_7923; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7925 = 8'ha4 == _T_375[7:0] ? 4'h0 : _GEN_7924; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7926 = 8'ha5 == _T_375[7:0] ? 4'h0 : _GEN_7925; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7927 = 8'ha6 == _T_375[7:0] ? 4'h0 : _GEN_7926; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7928 = 8'ha7 == _T_375[7:0] ? 4'h0 : _GEN_7927; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7929 = 8'ha8 == _T_375[7:0] ? 4'h0 : _GEN_7928; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7930 = 8'ha9 == _T_375[7:0] ? 4'h0 : _GEN_7929; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7931 = 8'haa == _T_375[7:0] ? 4'h0 : _GEN_7930; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7932 = 8'hab == _T_375[7:0] ? 4'h0 : _GEN_7931; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7933 = 8'hac == _T_375[7:0] ? 4'h2 : _GEN_7932; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7934 = 8'had == _T_375[7:0] ? 4'h0 : _GEN_7933; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7935 = 8'hae == _T_375[7:0] ? 4'h1 : _GEN_7934; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7936 = 8'haf == _T_375[7:0] ? 4'h3 : _GEN_7935; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7937 = 8'hb0 == _T_375[7:0] ? 4'h1 : _GEN_7936; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7938 = 8'hb1 == _T_375[7:0] ? 4'h0 : _GEN_7937; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7939 = 8'hb2 == _T_375[7:0] ? 4'h0 : _GEN_7938; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7940 = 8'hb3 == _T_375[7:0] ? 4'h0 : _GEN_7939; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7941 = 8'hb4 == _T_375[7:0] ? 4'h1 : _GEN_7940; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7942 = 8'hb5 == _T_375[7:0] ? 4'h3 : _GEN_7941; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7943 = 8'hb6 == _T_375[7:0] ? 4'h1 : _GEN_7942; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7944 = 8'hb7 == _T_375[7:0] ? 4'h0 : _GEN_7943; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7945 = 8'hb8 == _T_375[7:0] ? 4'h2 : _GEN_7944; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7946 = 8'hb9 == _T_375[7:0] ? 4'h0 : _GEN_7945; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7947 = 8'hba == _T_375[7:0] ? 4'h0 : _GEN_7946; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7948 = 8'hbb == _T_375[7:0] ? 4'h0 : _GEN_7947; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7949 = 8'hbc == _T_375[7:0] ? 4'h0 : _GEN_7948; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7950 = 8'hbd == _T_375[7:0] ? 4'h0 : _GEN_7949; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7951 = 8'hbe == _T_375[7:0] ? 4'h0 : _GEN_7950; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7952 = 8'hbf == _T_375[7:0] ? 4'h0 : _GEN_7951; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7953 = 8'hc0 == _T_375[7:0] ? 4'h0 : _GEN_7952; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7954 = 8'hc1 == _T_375[7:0] ? 4'h0 : _GEN_7953; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7955 = 8'hc2 == _T_375[7:0] ? 4'h3 : _GEN_7954; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7956 = 8'hc3 == _T_375[7:0] ? 4'h0 : _GEN_7955; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7957 = 8'hc4 == _T_375[7:0] ? 4'h0 : _GEN_7956; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7958 = 8'hc5 == _T_375[7:0] ? 4'h2 : _GEN_7957; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7959 = 8'hc6 == _T_375[7:0] ? 4'h3 : _GEN_7958; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7960 = 8'hc7 == _T_375[7:0] ? 4'h2 : _GEN_7959; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7961 = 8'hc8 == _T_375[7:0] ? 4'h3 : _GEN_7960; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7962 = 8'hc9 == _T_375[7:0] ? 4'h2 : _GEN_7961; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7963 = 8'hca == _T_375[7:0] ? 4'h0 : _GEN_7962; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7964 = 8'hcb == _T_375[7:0] ? 4'h0 : _GEN_7963; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7965 = 8'hcc == _T_375[7:0] ? 4'h3 : _GEN_7964; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7966 = 8'hcd == _T_375[7:0] ? 4'h0 : _GEN_7965; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7967 = 8'hce == _T_375[7:0] ? 4'h0 : _GEN_7966; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7968 = 8'hcf == _T_375[7:0] ? 4'h0 : _GEN_7967; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7969 = 8'hd0 == _T_375[7:0] ? 4'h0 : _GEN_7968; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7970 = 8'hd1 == _T_375[7:0] ? 4'h0 : _GEN_7969; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7971 = 8'hd2 == _T_375[7:0] ? 4'h0 : _GEN_7970; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7972 = 8'hd3 == _T_375[7:0] ? 4'h0 : _GEN_7971; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7973 = 8'hd4 == _T_375[7:0] ? 4'h0 : _GEN_7972; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7974 = 8'hd5 == _T_375[7:0] ? 4'h0 : _GEN_7973; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7975 = 8'hd6 == _T_375[7:0] ? 4'h0 : _GEN_7974; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7976 = 8'hd7 == _T_375[7:0] ? 4'h2 : _GEN_7975; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7977 = 8'hd8 == _T_375[7:0] ? 4'h2 : _GEN_7976; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7978 = 8'hd9 == _T_375[7:0] ? 4'h0 : _GEN_7977; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7979 = 8'hda == _T_375[7:0] ? 4'h7 : _GEN_7978; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7980 = 8'hdb == _T_375[7:0] ? 4'h1 : _GEN_7979; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7981 = 8'hdc == _T_375[7:0] ? 4'h4 : _GEN_7980; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7982 = 8'hdd == _T_375[7:0] ? 4'h1 : _GEN_7981; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7983 = 8'hde == _T_375[7:0] ? 4'h7 : _GEN_7982; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7984 = 8'hdf == _T_375[7:0] ? 4'h0 : _GEN_7983; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7985 = 8'he0 == _T_375[7:0] ? 4'h2 : _GEN_7984; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7986 = 8'he1 == _T_375[7:0] ? 4'h2 : _GEN_7985; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7987 = 8'he2 == _T_375[7:0] ? 4'h0 : _GEN_7986; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7988 = 8'he3 == _T_375[7:0] ? 4'h0 : _GEN_7987; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7989 = 8'he4 == _T_375[7:0] ? 4'h0 : _GEN_7988; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7990 = 8'he5 == _T_375[7:0] ? 4'h0 : _GEN_7989; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7991 = 8'he6 == _T_375[7:0] ? 4'h0 : _GEN_7990; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7992 = 8'he7 == _T_375[7:0] ? 4'h0 : _GEN_7991; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7993 = 8'he8 == _T_375[7:0] ? 4'h0 : _GEN_7992; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7994 = 8'he9 == _T_375[7:0] ? 4'h0 : _GEN_7993; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7995 = 8'hea == _T_375[7:0] ? 4'h0 : _GEN_7994; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7996 = 8'heb == _T_375[7:0] ? 4'h0 : _GEN_7995; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7997 = 8'hec == _T_375[7:0] ? 4'h0 : _GEN_7996; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7998 = 8'hed == _T_375[7:0] ? 4'h0 : _GEN_7997; // @[Filter.scala 204:62]
  wire [3:0] _GEN_7999 = 8'hee == _T_375[7:0] ? 4'h0 : _GEN_7998; // @[Filter.scala 204:62]
  wire [3:0] _GEN_8000 = 8'hef == _T_375[7:0] ? 4'h0 : _GEN_7999; // @[Filter.scala 204:62]
  wire [3:0] _GEN_8001 = 8'hf0 == _T_375[7:0] ? 4'h0 : _GEN_8000; // @[Filter.scala 204:62]
  wire [3:0] _GEN_8002 = 8'hf1 == _T_375[7:0] ? 4'h0 : _GEN_8001; // @[Filter.scala 204:62]
  wire [3:0] _GEN_8003 = 8'hf2 == _T_375[7:0] ? 4'h0 : _GEN_8002; // @[Filter.scala 204:62]
  wire [3:0] _GEN_8004 = 8'hf3 == _T_375[7:0] ? 4'h0 : _GEN_8003; // @[Filter.scala 204:62]
  wire [3:0] _GEN_8005 = 8'hf4 == _T_375[7:0] ? 4'h0 : _GEN_8004; // @[Filter.scala 204:62]
  wire [3:0] _GEN_8006 = 8'hf5 == _T_375[7:0] ? 4'h0 : _GEN_8005; // @[Filter.scala 204:62]
  wire [3:0] _GEN_8007 = 8'hf6 == _T_375[7:0] ? 4'h0 : _GEN_8006; // @[Filter.scala 204:62]
  wire [3:0] _GEN_8008 = 8'hf7 == _T_375[7:0] ? 4'h0 : _GEN_8007; // @[Filter.scala 204:62]
  wire [3:0] _GEN_8009 = 8'hf8 == _T_375[7:0] ? 4'h0 : _GEN_8008; // @[Filter.scala 204:62]
  wire [3:0] _GEN_8010 = 8'hf9 == _T_375[7:0] ? 4'h0 : _GEN_8009; // @[Filter.scala 204:62]
  wire [3:0] _GEN_8011 = 8'hfa == _T_375[7:0] ? 4'h0 : _GEN_8010; // @[Filter.scala 204:62]
  wire [3:0] _GEN_8012 = 8'hfb == _T_375[7:0] ? 4'h0 : _GEN_8011; // @[Filter.scala 204:62]
  wire [4:0] _GEN_11273 = {{1'd0}, _GEN_8012}; // @[Filter.scala 204:62]
  wire [8:0] _T_377 = _GEN_11273 * 5'h14; // @[Filter.scala 204:62]
  wire [3:0] _GEN_8062 = 8'h31 == _T_375[7:0] ? 4'h3 : _GEN_7809; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8063 = 8'h32 == _T_375[7:0] ? 4'h3 : _GEN_8062; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8064 = 8'h33 == _T_375[7:0] ? 4'h6 : _GEN_8063; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8065 = 8'h34 == _T_375[7:0] ? 4'h6 : _GEN_8064; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8066 = 8'h35 == _T_375[7:0] ? 4'h0 : _GEN_8065; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8067 = 8'h36 == _T_375[7:0] ? 4'h0 : _GEN_8066; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8068 = 8'h37 == _T_375[7:0] ? 4'h0 : _GEN_8067; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8069 = 8'h38 == _T_375[7:0] ? 4'h2 : _GEN_8068; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8070 = 8'h39 == _T_375[7:0] ? 4'h0 : _GEN_8069; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8071 = 8'h3a == _T_375[7:0] ? 4'h0 : _GEN_8070; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8072 = 8'h3b == _T_375[7:0] ? 4'h0 : _GEN_8071; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8073 = 8'h3c == _T_375[7:0] ? 4'h0 : _GEN_8072; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8074 = 8'h3d == _T_375[7:0] ? 4'h0 : _GEN_8073; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8075 = 8'h3e == _T_375[7:0] ? 4'h0 : _GEN_8074; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8076 = 8'h3f == _T_375[7:0] ? 4'h0 : _GEN_8075; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8077 = 8'h40 == _T_375[7:0] ? 4'h0 : _GEN_8076; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8078 = 8'h41 == _T_375[7:0] ? 4'h0 : _GEN_8077; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8079 = 8'h42 == _T_375[7:0] ? 4'h0 : _GEN_8078; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8080 = 8'h43 == _T_375[7:0] ? 4'h0 : _GEN_8079; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8081 = 8'h44 == _T_375[7:0] ? 4'h1 : _GEN_8080; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8082 = 8'h45 == _T_375[7:0] ? 4'h4 : _GEN_8081; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8083 = 8'h46 == _T_375[7:0] ? 4'hb : _GEN_8082; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8084 = 8'h47 == _T_375[7:0] ? 4'h0 : _GEN_8083; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8085 = 8'h48 == _T_375[7:0] ? 4'h0 : _GEN_8084; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8086 = 8'h49 == _T_375[7:0] ? 4'h0 : _GEN_8085; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8087 = 8'h4a == _T_375[7:0] ? 4'h6 : _GEN_8086; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8088 = 8'h4b == _T_375[7:0] ? 4'h0 : _GEN_8087; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8089 = 8'h4c == _T_375[7:0] ? 4'h3 : _GEN_8088; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8090 = 8'h4d == _T_375[7:0] ? 4'h3 : _GEN_8089; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8091 = 8'h4e == _T_375[7:0] ? 4'h2 : _GEN_8090; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8092 = 8'h4f == _T_375[7:0] ? 4'h0 : _GEN_8091; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8093 = 8'h50 == _T_375[7:0] ? 4'h0 : _GEN_8092; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8094 = 8'h51 == _T_375[7:0] ? 4'h0 : _GEN_8093; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8095 = 8'h52 == _T_375[7:0] ? 4'h0 : _GEN_8094; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8096 = 8'h53 == _T_375[7:0] ? 4'h0 : _GEN_8095; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8097 = 8'h54 == _T_375[7:0] ? 4'h0 : _GEN_8096; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8098 = 8'h55 == _T_375[7:0] ? 4'h0 : _GEN_8097; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8099 = 8'h56 == _T_375[7:0] ? 4'h0 : _GEN_8098; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8100 = 8'h57 == _T_375[7:0] ? 4'h0 : _GEN_8099; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8101 = 8'h58 == _T_375[7:0] ? 4'h0 : _GEN_8100; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8102 = 8'h59 == _T_375[7:0] ? 4'h2 : _GEN_8101; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8103 = 8'h5a == _T_375[7:0] ? 4'h3 : _GEN_8102; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8104 = 8'h5b == _T_375[7:0] ? 4'h0 : _GEN_8103; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8105 = 8'h5c == _T_375[7:0] ? 4'h0 : _GEN_8104; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8106 = 8'h5d == _T_375[7:0] ? 4'h3 : _GEN_8105; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8107 = 8'h5e == _T_375[7:0] ? 4'hd : _GEN_8106; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8108 = 8'h5f == _T_375[7:0] ? 4'h3 : _GEN_8107; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8109 = 8'h60 == _T_375[7:0] ? 4'h0 : _GEN_8108; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8110 = 8'h61 == _T_375[7:0] ? 4'h6 : _GEN_8109; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8111 = 8'h62 == _T_375[7:0] ? 4'h0 : _GEN_8110; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8112 = 8'h63 == _T_375[7:0] ? 4'h2 : _GEN_8111; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8113 = 8'h64 == _T_375[7:0] ? 4'h0 : _GEN_8112; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8114 = 8'h65 == _T_375[7:0] ? 4'h0 : _GEN_8113; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8115 = 8'h66 == _T_375[7:0] ? 4'h0 : _GEN_8114; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8116 = 8'h67 == _T_375[7:0] ? 4'h0 : _GEN_8115; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8117 = 8'h68 == _T_375[7:0] ? 4'h0 : _GEN_8116; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8118 = 8'h69 == _T_375[7:0] ? 4'h0 : _GEN_8117; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8119 = 8'h6a == _T_375[7:0] ? 4'h0 : _GEN_8118; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8120 = 8'h6b == _T_375[7:0] ? 4'h0 : _GEN_8119; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8121 = 8'h6c == _T_375[7:0] ? 4'h0 : _GEN_8120; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8122 = 8'h6d == _T_375[7:0] ? 4'h0 : _GEN_8121; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8123 = 8'h6e == _T_375[7:0] ? 4'h2 : _GEN_8122; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8124 = 8'h6f == _T_375[7:0] ? 4'h0 : _GEN_8123; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8125 = 8'h70 == _T_375[7:0] ? 4'h0 : _GEN_8124; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8126 = 8'h71 == _T_375[7:0] ? 4'h0 : _GEN_8125; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8127 = 8'h72 == _T_375[7:0] ? 4'h6 : _GEN_8126; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8128 = 8'h73 == _T_375[7:0] ? 4'he : _GEN_8127; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8129 = 8'h74 == _T_375[7:0] ? 4'h6 : _GEN_8128; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8130 = 8'h75 == _T_375[7:0] ? 4'h0 : _GEN_8129; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8131 = 8'h76 == _T_375[7:0] ? 4'h6 : _GEN_8130; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8132 = 8'h77 == _T_375[7:0] ? 4'h3 : _GEN_8131; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8133 = 8'h78 == _T_375[7:0] ? 4'h4 : _GEN_8132; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8134 = 8'h79 == _T_375[7:0] ? 4'h1 : _GEN_8133; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8135 = 8'h7a == _T_375[7:0] ? 4'h0 : _GEN_8134; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8136 = 8'h7b == _T_375[7:0] ? 4'h0 : _GEN_8135; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8137 = 8'h7c == _T_375[7:0] ? 4'h0 : _GEN_8136; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8138 = 8'h7d == _T_375[7:0] ? 4'h0 : _GEN_8137; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8139 = 8'h7e == _T_375[7:0] ? 4'h0 : _GEN_8138; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8140 = 8'h7f == _T_375[7:0] ? 4'h0 : _GEN_8139; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8141 = 8'h80 == _T_375[7:0] ? 4'h0 : _GEN_8140; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8142 = 8'h81 == _T_375[7:0] ? 4'h0 : _GEN_8141; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8143 = 8'h82 == _T_375[7:0] ? 4'h2 : _GEN_8142; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8144 = 8'h83 == _T_375[7:0] ? 4'h3 : _GEN_8143; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8145 = 8'h84 == _T_375[7:0] ? 4'h6 : _GEN_8144; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8146 = 8'h85 == _T_375[7:0] ? 4'h6 : _GEN_8145; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8147 = 8'h86 == _T_375[7:0] ? 4'he : _GEN_8146; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8148 = 8'h87 == _T_375[7:0] ? 4'ha : _GEN_8147; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8149 = 8'h88 == _T_375[7:0] ? 4'h6 : _GEN_8148; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8150 = 8'h89 == _T_375[7:0] ? 4'ha : _GEN_8149; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8151 = 8'h8a == _T_375[7:0] ? 4'he : _GEN_8150; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8152 = 8'h8b == _T_375[7:0] ? 4'h3 : _GEN_8151; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8153 = 8'h8c == _T_375[7:0] ? 4'h3 : _GEN_8152; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8154 = 8'h8d == _T_375[7:0] ? 4'h0 : _GEN_8153; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8155 = 8'h8e == _T_375[7:0] ? 4'h2 : _GEN_8154; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8156 = 8'h8f == _T_375[7:0] ? 4'h0 : _GEN_8155; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8157 = 8'h90 == _T_375[7:0] ? 4'h0 : _GEN_8156; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8158 = 8'h91 == _T_375[7:0] ? 4'h0 : _GEN_8157; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8159 = 8'h92 == _T_375[7:0] ? 4'h0 : _GEN_8158; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8160 = 8'h93 == _T_375[7:0] ? 4'h0 : _GEN_8159; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8161 = 8'h94 == _T_375[7:0] ? 4'h0 : _GEN_8160; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8162 = 8'h95 == _T_375[7:0] ? 4'h0 : _GEN_8161; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8163 = 8'h96 == _T_375[7:0] ? 4'h0 : _GEN_8162; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8164 = 8'h97 == _T_375[7:0] ? 4'h2 : _GEN_8163; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8165 = 8'h98 == _T_375[7:0] ? 4'h2 : _GEN_8164; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8166 = 8'h99 == _T_375[7:0] ? 4'h1 : _GEN_8165; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8167 = 8'h9a == _T_375[7:0] ? 4'h3 : _GEN_8166; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8168 = 8'h9b == _T_375[7:0] ? 4'he : _GEN_8167; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8169 = 8'h9c == _T_375[7:0] ? 4'he : _GEN_8168; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8170 = 8'h9d == _T_375[7:0] ? 4'h0 : _GEN_8169; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8171 = 8'h9e == _T_375[7:0] ? 4'he : _GEN_8170; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8172 = 8'h9f == _T_375[7:0] ? 4'he : _GEN_8171; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8173 = 8'ha0 == _T_375[7:0] ? 4'h3 : _GEN_8172; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8174 = 8'ha1 == _T_375[7:0] ? 4'h1 : _GEN_8173; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8175 = 8'ha2 == _T_375[7:0] ? 4'h2 : _GEN_8174; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8176 = 8'ha3 == _T_375[7:0] ? 4'h2 : _GEN_8175; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8177 = 8'ha4 == _T_375[7:0] ? 4'h0 : _GEN_8176; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8178 = 8'ha5 == _T_375[7:0] ? 4'h0 : _GEN_8177; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8179 = 8'ha6 == _T_375[7:0] ? 4'h0 : _GEN_8178; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8180 = 8'ha7 == _T_375[7:0] ? 4'h0 : _GEN_8179; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8181 = 8'ha8 == _T_375[7:0] ? 4'h0 : _GEN_8180; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8182 = 8'ha9 == _T_375[7:0] ? 4'h0 : _GEN_8181; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8183 = 8'haa == _T_375[7:0] ? 4'h0 : _GEN_8182; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8184 = 8'hab == _T_375[7:0] ? 4'h0 : _GEN_8183; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8185 = 8'hac == _T_375[7:0] ? 4'h2 : _GEN_8184; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8186 = 8'had == _T_375[7:0] ? 4'h3 : _GEN_8185; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8187 = 8'hae == _T_375[7:0] ? 4'h4 : _GEN_8186; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8188 = 8'haf == _T_375[7:0] ? 4'h3 : _GEN_8187; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8189 = 8'hb0 == _T_375[7:0] ? 4'h4 : _GEN_8188; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8190 = 8'hb1 == _T_375[7:0] ? 4'h3 : _GEN_8189; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8191 = 8'hb2 == _T_375[7:0] ? 4'h0 : _GEN_8190; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8192 = 8'hb3 == _T_375[7:0] ? 4'h3 : _GEN_8191; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8193 = 8'hb4 == _T_375[7:0] ? 4'h4 : _GEN_8192; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8194 = 8'hb5 == _T_375[7:0] ? 4'h3 : _GEN_8193; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8195 = 8'hb6 == _T_375[7:0] ? 4'h4 : _GEN_8194; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8196 = 8'hb7 == _T_375[7:0] ? 4'h3 : _GEN_8195; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8197 = 8'hb8 == _T_375[7:0] ? 4'h2 : _GEN_8196; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8198 = 8'hb9 == _T_375[7:0] ? 4'h0 : _GEN_8197; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8199 = 8'hba == _T_375[7:0] ? 4'h0 : _GEN_8198; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8200 = 8'hbb == _T_375[7:0] ? 4'h0 : _GEN_8199; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8201 = 8'hbc == _T_375[7:0] ? 4'h0 : _GEN_8200; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8202 = 8'hbd == _T_375[7:0] ? 4'h0 : _GEN_8201; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8203 = 8'hbe == _T_375[7:0] ? 4'h0 : _GEN_8202; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8204 = 8'hbf == _T_375[7:0] ? 4'h0 : _GEN_8203; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8205 = 8'hc0 == _T_375[7:0] ? 4'h0 : _GEN_8204; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8206 = 8'hc1 == _T_375[7:0] ? 4'h0 : _GEN_8205; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8207 = 8'hc2 == _T_375[7:0] ? 4'h8 : _GEN_8206; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8208 = 8'hc3 == _T_375[7:0] ? 4'hc : _GEN_8207; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8209 = 8'hc4 == _T_375[7:0] ? 4'h0 : _GEN_8208; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8210 = 8'hc5 == _T_375[7:0] ? 4'h2 : _GEN_8209; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8211 = 8'hc6 == _T_375[7:0] ? 4'h3 : _GEN_8210; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8212 = 8'hc7 == _T_375[7:0] ? 4'h2 : _GEN_8211; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8213 = 8'hc8 == _T_375[7:0] ? 4'h3 : _GEN_8212; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8214 = 8'hc9 == _T_375[7:0] ? 4'h2 : _GEN_8213; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8215 = 8'hca == _T_375[7:0] ? 4'h0 : _GEN_8214; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8216 = 8'hcb == _T_375[7:0] ? 4'hc : _GEN_8215; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8217 = 8'hcc == _T_375[7:0] ? 4'h8 : _GEN_8216; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8218 = 8'hcd == _T_375[7:0] ? 4'h0 : _GEN_8217; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8219 = 8'hce == _T_375[7:0] ? 4'h0 : _GEN_8218; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8220 = 8'hcf == _T_375[7:0] ? 4'h0 : _GEN_8219; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8221 = 8'hd0 == _T_375[7:0] ? 4'h0 : _GEN_8220; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8222 = 8'hd1 == _T_375[7:0] ? 4'h0 : _GEN_8221; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8223 = 8'hd2 == _T_375[7:0] ? 4'h0 : _GEN_8222; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8224 = 8'hd3 == _T_375[7:0] ? 4'h0 : _GEN_8223; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8225 = 8'hd4 == _T_375[7:0] ? 4'h0 : _GEN_8224; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8226 = 8'hd5 == _T_375[7:0] ? 4'h0 : _GEN_8225; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8227 = 8'hd6 == _T_375[7:0] ? 4'h0 : _GEN_8226; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8228 = 8'hd7 == _T_375[7:0] ? 4'h3 : _GEN_8227; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8229 = 8'hd8 == _T_375[7:0] ? 4'h6 : _GEN_8228; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8230 = 8'hd9 == _T_375[7:0] ? 4'h0 : _GEN_8229; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8231 = 8'hda == _T_375[7:0] ? 4'hb : _GEN_8230; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8232 = 8'hdb == _T_375[7:0] ? 4'h1 : _GEN_8231; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8233 = 8'hdc == _T_375[7:0] ? 4'h4 : _GEN_8232; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8234 = 8'hdd == _T_375[7:0] ? 4'h1 : _GEN_8233; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8235 = 8'hde == _T_375[7:0] ? 4'hb : _GEN_8234; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8236 = 8'hdf == _T_375[7:0] ? 4'h0 : _GEN_8235; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8237 = 8'he0 == _T_375[7:0] ? 4'h6 : _GEN_8236; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8238 = 8'he1 == _T_375[7:0] ? 4'h3 : _GEN_8237; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8239 = 8'he2 == _T_375[7:0] ? 4'h0 : _GEN_8238; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8240 = 8'he3 == _T_375[7:0] ? 4'h0 : _GEN_8239; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8241 = 8'he4 == _T_375[7:0] ? 4'h0 : _GEN_8240; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8242 = 8'he5 == _T_375[7:0] ? 4'h0 : _GEN_8241; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8243 = 8'he6 == _T_375[7:0] ? 4'h0 : _GEN_8242; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8244 = 8'he7 == _T_375[7:0] ? 4'h0 : _GEN_8243; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8245 = 8'he8 == _T_375[7:0] ? 4'h0 : _GEN_8244; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8246 = 8'he9 == _T_375[7:0] ? 4'h0 : _GEN_8245; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8247 = 8'hea == _T_375[7:0] ? 4'h0 : _GEN_8246; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8248 = 8'heb == _T_375[7:0] ? 4'h0 : _GEN_8247; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8249 = 8'hec == _T_375[7:0] ? 4'h0 : _GEN_8248; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8250 = 8'hed == _T_375[7:0] ? 4'h0 : _GEN_8249; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8251 = 8'hee == _T_375[7:0] ? 4'h0 : _GEN_8250; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8252 = 8'hef == _T_375[7:0] ? 4'h0 : _GEN_8251; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8253 = 8'hf0 == _T_375[7:0] ? 4'h0 : _GEN_8252; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8254 = 8'hf1 == _T_375[7:0] ? 4'h0 : _GEN_8253; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8255 = 8'hf2 == _T_375[7:0] ? 4'h0 : _GEN_8254; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8256 = 8'hf3 == _T_375[7:0] ? 4'h0 : _GEN_8255; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8257 = 8'hf4 == _T_375[7:0] ? 4'h0 : _GEN_8256; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8258 = 8'hf5 == _T_375[7:0] ? 4'h0 : _GEN_8257; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8259 = 8'hf6 == _T_375[7:0] ? 4'h0 : _GEN_8258; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8260 = 8'hf7 == _T_375[7:0] ? 4'h0 : _GEN_8259; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8261 = 8'hf8 == _T_375[7:0] ? 4'h0 : _GEN_8260; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8262 = 8'hf9 == _T_375[7:0] ? 4'h0 : _GEN_8261; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8263 = 8'hfa == _T_375[7:0] ? 4'h0 : _GEN_8262; // @[Filter.scala 204:102]
  wire [3:0] _GEN_8264 = 8'hfb == _T_375[7:0] ? 4'h0 : _GEN_8263; // @[Filter.scala 204:102]
  wire [6:0] _GEN_11275 = {{3'd0}, _GEN_8264}; // @[Filter.scala 204:102]
  wire [10:0] _T_382 = _GEN_11275 * 7'h46; // @[Filter.scala 204:102]
  wire [10:0] _GEN_11276 = {{2'd0}, _T_377}; // @[Filter.scala 204:69]
  wire [10:0] _T_384 = _GEN_11276 + _T_382; // @[Filter.scala 204:69]
  wire [3:0] _GEN_8273 = 8'h8 == _T_375[7:0] ? 4'h3 : 4'h0; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8274 = 8'h9 == _T_375[7:0] ? 4'h6 : _GEN_8273; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8275 = 8'ha == _T_375[7:0] ? 4'h6 : _GEN_8274; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8276 = 8'hb == _T_375[7:0] ? 4'h6 : _GEN_8275; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8277 = 8'hc == _T_375[7:0] ? 4'h3 : _GEN_8276; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8278 = 8'hd == _T_375[7:0] ? 4'h0 : _GEN_8277; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8279 = 8'he == _T_375[7:0] ? 4'h0 : _GEN_8278; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8280 = 8'hf == _T_375[7:0] ? 4'h0 : _GEN_8279; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8281 = 8'h10 == _T_375[7:0] ? 4'h0 : _GEN_8280; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8282 = 8'h11 == _T_375[7:0] ? 4'h0 : _GEN_8281; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8283 = 8'h12 == _T_375[7:0] ? 4'h0 : _GEN_8282; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8284 = 8'h13 == _T_375[7:0] ? 4'h0 : _GEN_8283; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8285 = 8'h14 == _T_375[7:0] ? 4'h0 : _GEN_8284; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8286 = 8'h15 == _T_375[7:0] ? 4'h0 : _GEN_8285; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8287 = 8'h16 == _T_375[7:0] ? 4'h0 : _GEN_8286; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8288 = 8'h17 == _T_375[7:0] ? 4'h0 : _GEN_8287; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8289 = 8'h18 == _T_375[7:0] ? 4'h0 : _GEN_8288; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8290 = 8'h19 == _T_375[7:0] ? 4'h0 : _GEN_8289; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8291 = 8'h1a == _T_375[7:0] ? 4'h0 : _GEN_8290; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8292 = 8'h1b == _T_375[7:0] ? 4'h0 : _GEN_8291; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8293 = 8'h1c == _T_375[7:0] ? 4'h6 : _GEN_8292; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8294 = 8'h1d == _T_375[7:0] ? 4'h3 : _GEN_8293; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8295 = 8'h1e == _T_375[7:0] ? 4'h0 : _GEN_8294; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8296 = 8'h1f == _T_375[7:0] ? 4'h0 : _GEN_8295; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8297 = 8'h20 == _T_375[7:0] ? 4'h0 : _GEN_8296; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8298 = 8'h21 == _T_375[7:0] ? 4'h3 : _GEN_8297; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8299 = 8'h22 == _T_375[7:0] ? 4'h6 : _GEN_8298; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8300 = 8'h23 == _T_375[7:0] ? 4'h0 : _GEN_8299; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8301 = 8'h24 == _T_375[7:0] ? 4'h0 : _GEN_8300; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8302 = 8'h25 == _T_375[7:0] ? 4'h0 : _GEN_8301; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8303 = 8'h26 == _T_375[7:0] ? 4'h0 : _GEN_8302; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8304 = 8'h27 == _T_375[7:0] ? 4'h0 : _GEN_8303; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8305 = 8'h28 == _T_375[7:0] ? 4'h0 : _GEN_8304; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8306 = 8'h29 == _T_375[7:0] ? 4'h0 : _GEN_8305; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8307 = 8'h2a == _T_375[7:0] ? 4'h0 : _GEN_8306; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8308 = 8'h2b == _T_375[7:0] ? 4'h0 : _GEN_8307; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8309 = 8'h2c == _T_375[7:0] ? 4'h0 : _GEN_8308; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8310 = 8'h2d == _T_375[7:0] ? 4'h0 : _GEN_8309; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8311 = 8'h2e == _T_375[7:0] ? 4'h0 : _GEN_8310; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8312 = 8'h2f == _T_375[7:0] ? 4'h0 : _GEN_8311; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8313 = 8'h30 == _T_375[7:0] ? 4'h6 : _GEN_8312; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8314 = 8'h31 == _T_375[7:0] ? 4'h3 : _GEN_8313; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8315 = 8'h32 == _T_375[7:0] ? 4'h0 : _GEN_8314; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8316 = 8'h33 == _T_375[7:0] ? 4'h1 : _GEN_8315; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8317 = 8'h34 == _T_375[7:0] ? 4'h1 : _GEN_8316; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8318 = 8'h35 == _T_375[7:0] ? 4'h0 : _GEN_8317; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8319 = 8'h36 == _T_375[7:0] ? 4'h0 : _GEN_8318; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8320 = 8'h37 == _T_375[7:0] ? 4'h0 : _GEN_8319; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8321 = 8'h38 == _T_375[7:0] ? 4'h6 : _GEN_8320; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8322 = 8'h39 == _T_375[7:0] ? 4'h0 : _GEN_8321; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8323 = 8'h3a == _T_375[7:0] ? 4'h0 : _GEN_8322; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8324 = 8'h3b == _T_375[7:0] ? 4'h0 : _GEN_8323; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8325 = 8'h3c == _T_375[7:0] ? 4'h0 : _GEN_8324; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8326 = 8'h3d == _T_375[7:0] ? 4'h0 : _GEN_8325; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8327 = 8'h3e == _T_375[7:0] ? 4'h0 : _GEN_8326; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8328 = 8'h3f == _T_375[7:0] ? 4'h0 : _GEN_8327; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8329 = 8'h40 == _T_375[7:0] ? 4'h0 : _GEN_8328; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8330 = 8'h41 == _T_375[7:0] ? 4'h0 : _GEN_8329; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8331 = 8'h42 == _T_375[7:0] ? 4'h0 : _GEN_8330; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8332 = 8'h43 == _T_375[7:0] ? 4'h0 : _GEN_8331; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8333 = 8'h44 == _T_375[7:0] ? 4'h3 : _GEN_8332; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8334 = 8'h45 == _T_375[7:0] ? 4'h6 : _GEN_8333; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8335 = 8'h46 == _T_375[7:0] ? 4'h9 : _GEN_8334; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8336 = 8'h47 == _T_375[7:0] ? 4'h0 : _GEN_8335; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8337 = 8'h48 == _T_375[7:0] ? 4'h0 : _GEN_8336; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8338 = 8'h49 == _T_375[7:0] ? 4'h0 : _GEN_8337; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8339 = 8'h4a == _T_375[7:0] ? 4'h1 : _GEN_8338; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8340 = 8'h4b == _T_375[7:0] ? 4'h0 : _GEN_8339; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8341 = 8'h4c == _T_375[7:0] ? 4'h0 : _GEN_8340; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8342 = 8'h4d == _T_375[7:0] ? 4'h0 : _GEN_8341; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8343 = 8'h4e == _T_375[7:0] ? 4'h6 : _GEN_8342; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8344 = 8'h4f == _T_375[7:0] ? 4'h0 : _GEN_8343; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8345 = 8'h50 == _T_375[7:0] ? 4'h0 : _GEN_8344; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8346 = 8'h51 == _T_375[7:0] ? 4'h0 : _GEN_8345; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8347 = 8'h52 == _T_375[7:0] ? 4'h0 : _GEN_8346; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8348 = 8'h53 == _T_375[7:0] ? 4'h0 : _GEN_8347; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8349 = 8'h54 == _T_375[7:0] ? 4'h0 : _GEN_8348; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8350 = 8'h55 == _T_375[7:0] ? 4'h0 : _GEN_8349; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8351 = 8'h56 == _T_375[7:0] ? 4'h0 : _GEN_8350; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8352 = 8'h57 == _T_375[7:0] ? 4'h0 : _GEN_8351; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8353 = 8'h58 == _T_375[7:0] ? 4'h0 : _GEN_8352; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8354 = 8'h59 == _T_375[7:0] ? 4'h6 : _GEN_8353; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8355 = 8'h5a == _T_375[7:0] ? 4'h3 : _GEN_8354; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8356 = 8'h5b == _T_375[7:0] ? 4'h0 : _GEN_8355; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8357 = 8'h5c == _T_375[7:0] ? 4'h0 : _GEN_8356; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8358 = 8'h5d == _T_375[7:0] ? 4'h0 : _GEN_8357; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8359 = 8'h5e == _T_375[7:0] ? 4'h7 : _GEN_8358; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8360 = 8'h5f == _T_375[7:0] ? 4'h0 : _GEN_8359; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8361 = 8'h60 == _T_375[7:0] ? 4'h0 : _GEN_8360; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8362 = 8'h61 == _T_375[7:0] ? 4'h1 : _GEN_8361; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8363 = 8'h62 == _T_375[7:0] ? 4'h0 : _GEN_8362; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8364 = 8'h63 == _T_375[7:0] ? 4'h6 : _GEN_8363; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8365 = 8'h64 == _T_375[7:0] ? 4'h0 : _GEN_8364; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8366 = 8'h65 == _T_375[7:0] ? 4'h0 : _GEN_8365; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8367 = 8'h66 == _T_375[7:0] ? 4'h0 : _GEN_8366; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8368 = 8'h67 == _T_375[7:0] ? 4'h0 : _GEN_8367; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8369 = 8'h68 == _T_375[7:0] ? 4'h0 : _GEN_8368; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8370 = 8'h69 == _T_375[7:0] ? 4'h0 : _GEN_8369; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8371 = 8'h6a == _T_375[7:0] ? 4'h0 : _GEN_8370; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8372 = 8'h6b == _T_375[7:0] ? 4'h0 : _GEN_8371; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8373 = 8'h6c == _T_375[7:0] ? 4'h0 : _GEN_8372; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8374 = 8'h6d == _T_375[7:0] ? 4'h0 : _GEN_8373; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8375 = 8'h6e == _T_375[7:0] ? 4'h6 : _GEN_8374; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8376 = 8'h6f == _T_375[7:0] ? 4'h0 : _GEN_8375; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8377 = 8'h70 == _T_375[7:0] ? 4'h0 : _GEN_8376; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8378 = 8'h71 == _T_375[7:0] ? 4'h0 : _GEN_8377; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8379 = 8'h72 == _T_375[7:0] ? 4'h3 : _GEN_8378; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8380 = 8'h73 == _T_375[7:0] ? 4'hc : _GEN_8379; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8381 = 8'h74 == _T_375[7:0] ? 4'h3 : _GEN_8380; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8382 = 8'h75 == _T_375[7:0] ? 4'h0 : _GEN_8381; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8383 = 8'h76 == _T_375[7:0] ? 4'h1 : _GEN_8382; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8384 = 8'h77 == _T_375[7:0] ? 4'h0 : _GEN_8383; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8385 = 8'h78 == _T_375[7:0] ? 4'h3 : _GEN_8384; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8386 = 8'h79 == _T_375[7:0] ? 4'h3 : _GEN_8385; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8387 = 8'h7a == _T_375[7:0] ? 4'h0 : _GEN_8386; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8388 = 8'h7b == _T_375[7:0] ? 4'h0 : _GEN_8387; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8389 = 8'h7c == _T_375[7:0] ? 4'h0 : _GEN_8388; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8390 = 8'h7d == _T_375[7:0] ? 4'h0 : _GEN_8389; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8391 = 8'h7e == _T_375[7:0] ? 4'h0 : _GEN_8390; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8392 = 8'h7f == _T_375[7:0] ? 4'h0 : _GEN_8391; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8393 = 8'h80 == _T_375[7:0] ? 4'h0 : _GEN_8392; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8394 = 8'h81 == _T_375[7:0] ? 4'h0 : _GEN_8393; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8395 = 8'h82 == _T_375[7:0] ? 4'h6 : _GEN_8394; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8396 = 8'h83 == _T_375[7:0] ? 4'h0 : _GEN_8395; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8397 = 8'h84 == _T_375[7:0] ? 4'h1 : _GEN_8396; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8398 = 8'h85 == _T_375[7:0] ? 4'h1 : _GEN_8397; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8399 = 8'h86 == _T_375[7:0] ? 4'ha : _GEN_8398; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8400 = 8'h87 == _T_375[7:0] ? 4'h4 : _GEN_8399; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8401 = 8'h88 == _T_375[7:0] ? 4'h1 : _GEN_8400; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8402 = 8'h89 == _T_375[7:0] ? 4'h4 : _GEN_8401; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8403 = 8'h8a == _T_375[7:0] ? 4'ha : _GEN_8402; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8404 = 8'h8b == _T_375[7:0] ? 4'h0 : _GEN_8403; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8405 = 8'h8c == _T_375[7:0] ? 4'h0 : _GEN_8404; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8406 = 8'h8d == _T_375[7:0] ? 4'h0 : _GEN_8405; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8407 = 8'h8e == _T_375[7:0] ? 4'h6 : _GEN_8406; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8408 = 8'h8f == _T_375[7:0] ? 4'h0 : _GEN_8407; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8409 = 8'h90 == _T_375[7:0] ? 4'h0 : _GEN_8408; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8410 = 8'h91 == _T_375[7:0] ? 4'h0 : _GEN_8409; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8411 = 8'h92 == _T_375[7:0] ? 4'h0 : _GEN_8410; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8412 = 8'h93 == _T_375[7:0] ? 4'h0 : _GEN_8411; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8413 = 8'h94 == _T_375[7:0] ? 4'h0 : _GEN_8412; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8414 = 8'h95 == _T_375[7:0] ? 4'h0 : _GEN_8413; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8415 = 8'h96 == _T_375[7:0] ? 4'h0 : _GEN_8414; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8416 = 8'h97 == _T_375[7:0] ? 4'h6 : _GEN_8415; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8417 = 8'h98 == _T_375[7:0] ? 4'h6 : _GEN_8416; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8418 = 8'h99 == _T_375[7:0] ? 4'h3 : _GEN_8417; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8419 = 8'h9a == _T_375[7:0] ? 4'h0 : _GEN_8418; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8420 = 8'h9b == _T_375[7:0] ? 4'ha : _GEN_8419; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8421 = 8'h9c == _T_375[7:0] ? 4'ha : _GEN_8420; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8422 = 8'h9d == _T_375[7:0] ? 4'h0 : _GEN_8421; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8423 = 8'h9e == _T_375[7:0] ? 4'ha : _GEN_8422; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8424 = 8'h9f == _T_375[7:0] ? 4'ha : _GEN_8423; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8425 = 8'ha0 == _T_375[7:0] ? 4'h0 : _GEN_8424; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8426 = 8'ha1 == _T_375[7:0] ? 4'h3 : _GEN_8425; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8427 = 8'ha2 == _T_375[7:0] ? 4'h6 : _GEN_8426; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8428 = 8'ha3 == _T_375[7:0] ? 4'h6 : _GEN_8427; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8429 = 8'ha4 == _T_375[7:0] ? 4'h0 : _GEN_8428; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8430 = 8'ha5 == _T_375[7:0] ? 4'h0 : _GEN_8429; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8431 = 8'ha6 == _T_375[7:0] ? 4'h0 : _GEN_8430; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8432 = 8'ha7 == _T_375[7:0] ? 4'h0 : _GEN_8431; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8433 = 8'ha8 == _T_375[7:0] ? 4'h0 : _GEN_8432; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8434 = 8'ha9 == _T_375[7:0] ? 4'h0 : _GEN_8433; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8435 = 8'haa == _T_375[7:0] ? 4'h0 : _GEN_8434; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8436 = 8'hab == _T_375[7:0] ? 4'h0 : _GEN_8435; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8437 = 8'hac == _T_375[7:0] ? 4'h6 : _GEN_8436; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8438 = 8'had == _T_375[7:0] ? 4'h0 : _GEN_8437; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8439 = 8'hae == _T_375[7:0] ? 4'h3 : _GEN_8438; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8440 = 8'haf == _T_375[7:0] ? 4'h9 : _GEN_8439; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8441 = 8'hb0 == _T_375[7:0] ? 4'h3 : _GEN_8440; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8442 = 8'hb1 == _T_375[7:0] ? 4'h0 : _GEN_8441; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8443 = 8'hb2 == _T_375[7:0] ? 4'h0 : _GEN_8442; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8444 = 8'hb3 == _T_375[7:0] ? 4'h0 : _GEN_8443; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8445 = 8'hb4 == _T_375[7:0] ? 4'h3 : _GEN_8444; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8446 = 8'hb5 == _T_375[7:0] ? 4'h9 : _GEN_8445; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8447 = 8'hb6 == _T_375[7:0] ? 4'h3 : _GEN_8446; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8448 = 8'hb7 == _T_375[7:0] ? 4'h0 : _GEN_8447; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8449 = 8'hb8 == _T_375[7:0] ? 4'h6 : _GEN_8448; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8450 = 8'hb9 == _T_375[7:0] ? 4'h0 : _GEN_8449; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8451 = 8'hba == _T_375[7:0] ? 4'h0 : _GEN_8450; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8452 = 8'hbb == _T_375[7:0] ? 4'h0 : _GEN_8451; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8453 = 8'hbc == _T_375[7:0] ? 4'h0 : _GEN_8452; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8454 = 8'hbd == _T_375[7:0] ? 4'h0 : _GEN_8453; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8455 = 8'hbe == _T_375[7:0] ? 4'h0 : _GEN_8454; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8456 = 8'hbf == _T_375[7:0] ? 4'h0 : _GEN_8455; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8457 = 8'hc0 == _T_375[7:0] ? 4'h0 : _GEN_8456; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8458 = 8'hc1 == _T_375[7:0] ? 4'h0 : _GEN_8457; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8459 = 8'hc2 == _T_375[7:0] ? 4'h7 : _GEN_8458; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8460 = 8'hc3 == _T_375[7:0] ? 4'h2 : _GEN_8459; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8461 = 8'hc4 == _T_375[7:0] ? 4'h0 : _GEN_8460; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8462 = 8'hc5 == _T_375[7:0] ? 4'h6 : _GEN_8461; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8463 = 8'hc6 == _T_375[7:0] ? 4'h9 : _GEN_8462; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8464 = 8'hc7 == _T_375[7:0] ? 4'h6 : _GEN_8463; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8465 = 8'hc8 == _T_375[7:0] ? 4'h9 : _GEN_8464; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8466 = 8'hc9 == _T_375[7:0] ? 4'h6 : _GEN_8465; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8467 = 8'hca == _T_375[7:0] ? 4'h0 : _GEN_8466; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8468 = 8'hcb == _T_375[7:0] ? 4'h2 : _GEN_8467; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8469 = 8'hcc == _T_375[7:0] ? 4'h7 : _GEN_8468; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8470 = 8'hcd == _T_375[7:0] ? 4'h0 : _GEN_8469; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8471 = 8'hce == _T_375[7:0] ? 4'h0 : _GEN_8470; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8472 = 8'hcf == _T_375[7:0] ? 4'h0 : _GEN_8471; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8473 = 8'hd0 == _T_375[7:0] ? 4'h0 : _GEN_8472; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8474 = 8'hd1 == _T_375[7:0] ? 4'h0 : _GEN_8473; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8475 = 8'hd2 == _T_375[7:0] ? 4'h0 : _GEN_8474; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8476 = 8'hd3 == _T_375[7:0] ? 4'h0 : _GEN_8475; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8477 = 8'hd4 == _T_375[7:0] ? 4'h0 : _GEN_8476; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8478 = 8'hd5 == _T_375[7:0] ? 4'h0 : _GEN_8477; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8479 = 8'hd6 == _T_375[7:0] ? 4'h0 : _GEN_8478; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8480 = 8'hd7 == _T_375[7:0] ? 4'h3 : _GEN_8479; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8481 = 8'hd8 == _T_375[7:0] ? 4'h3 : _GEN_8480; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8482 = 8'hd9 == _T_375[7:0] ? 4'h0 : _GEN_8481; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8483 = 8'hda == _T_375[7:0] ? 4'h9 : _GEN_8482; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8484 = 8'hdb == _T_375[7:0] ? 4'h3 : _GEN_8483; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8485 = 8'hdc == _T_375[7:0] ? 4'hc : _GEN_8484; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8486 = 8'hdd == _T_375[7:0] ? 4'h3 : _GEN_8485; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8487 = 8'hde == _T_375[7:0] ? 4'h9 : _GEN_8486; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8488 = 8'hdf == _T_375[7:0] ? 4'h0 : _GEN_8487; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8489 = 8'he0 == _T_375[7:0] ? 4'h3 : _GEN_8488; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8490 = 8'he1 == _T_375[7:0] ? 4'h3 : _GEN_8489; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8491 = 8'he2 == _T_375[7:0] ? 4'h0 : _GEN_8490; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8492 = 8'he3 == _T_375[7:0] ? 4'h0 : _GEN_8491; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8493 = 8'he4 == _T_375[7:0] ? 4'h0 : _GEN_8492; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8494 = 8'he5 == _T_375[7:0] ? 4'h0 : _GEN_8493; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8495 = 8'he6 == _T_375[7:0] ? 4'h0 : _GEN_8494; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8496 = 8'he7 == _T_375[7:0] ? 4'h0 : _GEN_8495; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8497 = 8'he8 == _T_375[7:0] ? 4'h0 : _GEN_8496; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8498 = 8'he9 == _T_375[7:0] ? 4'h0 : _GEN_8497; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8499 = 8'hea == _T_375[7:0] ? 4'h0 : _GEN_8498; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8500 = 8'heb == _T_375[7:0] ? 4'h0 : _GEN_8499; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8501 = 8'hec == _T_375[7:0] ? 4'h0 : _GEN_8500; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8502 = 8'hed == _T_375[7:0] ? 4'h0 : _GEN_8501; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8503 = 8'hee == _T_375[7:0] ? 4'h0 : _GEN_8502; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8504 = 8'hef == _T_375[7:0] ? 4'h0 : _GEN_8503; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8505 = 8'hf0 == _T_375[7:0] ? 4'h0 : _GEN_8504; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8506 = 8'hf1 == _T_375[7:0] ? 4'h0 : _GEN_8505; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8507 = 8'hf2 == _T_375[7:0] ? 4'h0 : _GEN_8506; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8508 = 8'hf3 == _T_375[7:0] ? 4'h0 : _GEN_8507; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8509 = 8'hf4 == _T_375[7:0] ? 4'h0 : _GEN_8508; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8510 = 8'hf5 == _T_375[7:0] ? 4'h0 : _GEN_8509; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8511 = 8'hf6 == _T_375[7:0] ? 4'h0 : _GEN_8510; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8512 = 8'hf7 == _T_375[7:0] ? 4'h0 : _GEN_8511; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8513 = 8'hf8 == _T_375[7:0] ? 4'h0 : _GEN_8512; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8514 = 8'hf9 == _T_375[7:0] ? 4'h0 : _GEN_8513; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8515 = 8'hfa == _T_375[7:0] ? 4'h0 : _GEN_8514; // @[Filter.scala 204:142]
  wire [3:0] _GEN_8516 = 8'hfb == _T_375[7:0] ? 4'h0 : _GEN_8515; // @[Filter.scala 204:142]
  wire [7:0] _T_389 = _GEN_8516 * 4'ha; // @[Filter.scala 204:142]
  wire [10:0] _GEN_11278 = {{3'd0}, _T_389}; // @[Filter.scala 204:109]
  wire [10:0] _T_391 = _T_384 + _GEN_11278; // @[Filter.scala 204:109]
  wire [10:0] _T_392 = _T_391 / 11'h64; // @[Filter.scala 204:150]
  wire  _T_394 = _T_365 >= 5'h15; // @[Filter.scala 207:31]
  wire  _T_398 = _T_372 >= 32'hc; // @[Filter.scala 207:63]
  wire  _T_399 = _T_394 | _T_398; // @[Filter.scala 207:58]
  wire [10:0] _GEN_8769 = io_SPI_distort ? _T_392 : {{7'd0}, _GEN_8012}; // @[Filter.scala 209:35]
  wire [10:0] _GEN_8770 = _T_399 ? 11'h0 : _GEN_8769; // @[Filter.scala 207:80]
  wire [10:0] _GEN_9023 = io_SPI_distort ? _T_392 : {{7'd0}, _GEN_8264}; // @[Filter.scala 209:35]
  wire [10:0] _GEN_9024 = _T_399 ? 11'h0 : _GEN_9023; // @[Filter.scala 207:80]
  wire [10:0] _GEN_9277 = io_SPI_distort ? _T_392 : {{7'd0}, _GEN_8516}; // @[Filter.scala 209:35]
  wire [10:0] _GEN_9278 = _T_399 ? 11'h0 : _GEN_9277; // @[Filter.scala 207:80]
  wire [31:0] _T_427 = pixelIndex + 32'h6; // @[Filter.scala 202:31]
  wire [31:0] _GEN_6 = _T_427 % 32'h15; // @[Filter.scala 202:38]
  wire [4:0] _T_428 = _GEN_6[4:0]; // @[Filter.scala 202:38]
  wire [4:0] _T_430 = _T_428 + _GEN_11210; // @[Filter.scala 202:53]
  wire [4:0] _T_432 = _T_430 - 5'h1; // @[Filter.scala 202:69]
  wire [31:0] _T_435 = _T_427 / 32'h15; // @[Filter.scala 203:38]
  wire [31:0] _T_437 = _T_435 + _GEN_11211; // @[Filter.scala 203:53]
  wire [31:0] _T_439 = _T_437 - 32'h1; // @[Filter.scala 203:69]
  wire [36:0] _T_440 = _T_439 * 32'h15; // @[Filter.scala 204:42]
  wire [36:0] _GEN_11284 = {{32'd0}, _T_432}; // @[Filter.scala 204:57]
  wire [36:0] _T_442 = _T_440 + _GEN_11284; // @[Filter.scala 204:57]
  wire [3:0] _GEN_9287 = 8'h8 == _T_442[7:0] ? 4'h1 : 4'h0; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9288 = 8'h9 == _T_442[7:0] ? 4'h2 : _GEN_9287; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9289 = 8'ha == _T_442[7:0] ? 4'h2 : _GEN_9288; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9290 = 8'hb == _T_442[7:0] ? 4'h2 : _GEN_9289; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9291 = 8'hc == _T_442[7:0] ? 4'h1 : _GEN_9290; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9292 = 8'hd == _T_442[7:0] ? 4'h0 : _GEN_9291; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9293 = 8'he == _T_442[7:0] ? 4'h0 : _GEN_9292; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9294 = 8'hf == _T_442[7:0] ? 4'h0 : _GEN_9293; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9295 = 8'h10 == _T_442[7:0] ? 4'h0 : _GEN_9294; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9296 = 8'h11 == _T_442[7:0] ? 4'h0 : _GEN_9295; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9297 = 8'h12 == _T_442[7:0] ? 4'h0 : _GEN_9296; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9298 = 8'h13 == _T_442[7:0] ? 4'h0 : _GEN_9297; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9299 = 8'h14 == _T_442[7:0] ? 4'h0 : _GEN_9298; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9300 = 8'h15 == _T_442[7:0] ? 4'h0 : _GEN_9299; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9301 = 8'h16 == _T_442[7:0] ? 4'h0 : _GEN_9300; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9302 = 8'h17 == _T_442[7:0] ? 4'h0 : _GEN_9301; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9303 = 8'h18 == _T_442[7:0] ? 4'h0 : _GEN_9302; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9304 = 8'h19 == _T_442[7:0] ? 4'h0 : _GEN_9303; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9305 = 8'h1a == _T_442[7:0] ? 4'h0 : _GEN_9304; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9306 = 8'h1b == _T_442[7:0] ? 4'h0 : _GEN_9305; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9307 = 8'h1c == _T_442[7:0] ? 4'h2 : _GEN_9306; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9308 = 8'h1d == _T_442[7:0] ? 4'h1 : _GEN_9307; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9309 = 8'h1e == _T_442[7:0] ? 4'h0 : _GEN_9308; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9310 = 8'h1f == _T_442[7:0] ? 4'h0 : _GEN_9309; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9311 = 8'h20 == _T_442[7:0] ? 4'h0 : _GEN_9310; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9312 = 8'h21 == _T_442[7:0] ? 4'h1 : _GEN_9311; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9313 = 8'h22 == _T_442[7:0] ? 4'h2 : _GEN_9312; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9314 = 8'h23 == _T_442[7:0] ? 4'h0 : _GEN_9313; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9315 = 8'h24 == _T_442[7:0] ? 4'h0 : _GEN_9314; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9316 = 8'h25 == _T_442[7:0] ? 4'h0 : _GEN_9315; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9317 = 8'h26 == _T_442[7:0] ? 4'h0 : _GEN_9316; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9318 = 8'h27 == _T_442[7:0] ? 4'h0 : _GEN_9317; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9319 = 8'h28 == _T_442[7:0] ? 4'h0 : _GEN_9318; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9320 = 8'h29 == _T_442[7:0] ? 4'h0 : _GEN_9319; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9321 = 8'h2a == _T_442[7:0] ? 4'h0 : _GEN_9320; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9322 = 8'h2b == _T_442[7:0] ? 4'h0 : _GEN_9321; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9323 = 8'h2c == _T_442[7:0] ? 4'h0 : _GEN_9322; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9324 = 8'h2d == _T_442[7:0] ? 4'h0 : _GEN_9323; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9325 = 8'h2e == _T_442[7:0] ? 4'h0 : _GEN_9324; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9326 = 8'h2f == _T_442[7:0] ? 4'h0 : _GEN_9325; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9327 = 8'h30 == _T_442[7:0] ? 4'h2 : _GEN_9326; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9328 = 8'h31 == _T_442[7:0] ? 4'h2 : _GEN_9327; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9329 = 8'h32 == _T_442[7:0] ? 4'h0 : _GEN_9328; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9330 = 8'h33 == _T_442[7:0] ? 4'h0 : _GEN_9329; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9331 = 8'h34 == _T_442[7:0] ? 4'h0 : _GEN_9330; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9332 = 8'h35 == _T_442[7:0] ? 4'h0 : _GEN_9331; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9333 = 8'h36 == _T_442[7:0] ? 4'h0 : _GEN_9332; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9334 = 8'h37 == _T_442[7:0] ? 4'h0 : _GEN_9333; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9335 = 8'h38 == _T_442[7:0] ? 4'h2 : _GEN_9334; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9336 = 8'h39 == _T_442[7:0] ? 4'h0 : _GEN_9335; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9337 = 8'h3a == _T_442[7:0] ? 4'h0 : _GEN_9336; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9338 = 8'h3b == _T_442[7:0] ? 4'h0 : _GEN_9337; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9339 = 8'h3c == _T_442[7:0] ? 4'h0 : _GEN_9338; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9340 = 8'h3d == _T_442[7:0] ? 4'h0 : _GEN_9339; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9341 = 8'h3e == _T_442[7:0] ? 4'h0 : _GEN_9340; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9342 = 8'h3f == _T_442[7:0] ? 4'h0 : _GEN_9341; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9343 = 8'h40 == _T_442[7:0] ? 4'h0 : _GEN_9342; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9344 = 8'h41 == _T_442[7:0] ? 4'h0 : _GEN_9343; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9345 = 8'h42 == _T_442[7:0] ? 4'h0 : _GEN_9344; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9346 = 8'h43 == _T_442[7:0] ? 4'h0 : _GEN_9345; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9347 = 8'h44 == _T_442[7:0] ? 4'h1 : _GEN_9346; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9348 = 8'h45 == _T_442[7:0] ? 4'h3 : _GEN_9347; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9349 = 8'h46 == _T_442[7:0] ? 4'h7 : _GEN_9348; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9350 = 8'h47 == _T_442[7:0] ? 4'h0 : _GEN_9349; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9351 = 8'h48 == _T_442[7:0] ? 4'h0 : _GEN_9350; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9352 = 8'h49 == _T_442[7:0] ? 4'h0 : _GEN_9351; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9353 = 8'h4a == _T_442[7:0] ? 4'h0 : _GEN_9352; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9354 = 8'h4b == _T_442[7:0] ? 4'h0 : _GEN_9353; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9355 = 8'h4c == _T_442[7:0] ? 4'h0 : _GEN_9354; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9356 = 8'h4d == _T_442[7:0] ? 4'h0 : _GEN_9355; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9357 = 8'h4e == _T_442[7:0] ? 4'h2 : _GEN_9356; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9358 = 8'h4f == _T_442[7:0] ? 4'h0 : _GEN_9357; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9359 = 8'h50 == _T_442[7:0] ? 4'h0 : _GEN_9358; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9360 = 8'h51 == _T_442[7:0] ? 4'h0 : _GEN_9359; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9361 = 8'h52 == _T_442[7:0] ? 4'h0 : _GEN_9360; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9362 = 8'h53 == _T_442[7:0] ? 4'h0 : _GEN_9361; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9363 = 8'h54 == _T_442[7:0] ? 4'h0 : _GEN_9362; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9364 = 8'h55 == _T_442[7:0] ? 4'h0 : _GEN_9363; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9365 = 8'h56 == _T_442[7:0] ? 4'h0 : _GEN_9364; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9366 = 8'h57 == _T_442[7:0] ? 4'h0 : _GEN_9365; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9367 = 8'h58 == _T_442[7:0] ? 4'h0 : _GEN_9366; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9368 = 8'h59 == _T_442[7:0] ? 4'h2 : _GEN_9367; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9369 = 8'h5a == _T_442[7:0] ? 4'h2 : _GEN_9368; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9370 = 8'h5b == _T_442[7:0] ? 4'h0 : _GEN_9369; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9371 = 8'h5c == _T_442[7:0] ? 4'h0 : _GEN_9370; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9372 = 8'h5d == _T_442[7:0] ? 4'h0 : _GEN_9371; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9373 = 8'h5e == _T_442[7:0] ? 4'h4 : _GEN_9372; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9374 = 8'h5f == _T_442[7:0] ? 4'h0 : _GEN_9373; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9375 = 8'h60 == _T_442[7:0] ? 4'h0 : _GEN_9374; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9376 = 8'h61 == _T_442[7:0] ? 4'h0 : _GEN_9375; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9377 = 8'h62 == _T_442[7:0] ? 4'h0 : _GEN_9376; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9378 = 8'h63 == _T_442[7:0] ? 4'h2 : _GEN_9377; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9379 = 8'h64 == _T_442[7:0] ? 4'h0 : _GEN_9378; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9380 = 8'h65 == _T_442[7:0] ? 4'h0 : _GEN_9379; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9381 = 8'h66 == _T_442[7:0] ? 4'h0 : _GEN_9380; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9382 = 8'h67 == _T_442[7:0] ? 4'h0 : _GEN_9381; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9383 = 8'h68 == _T_442[7:0] ? 4'h0 : _GEN_9382; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9384 = 8'h69 == _T_442[7:0] ? 4'h0 : _GEN_9383; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9385 = 8'h6a == _T_442[7:0] ? 4'h0 : _GEN_9384; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9386 = 8'h6b == _T_442[7:0] ? 4'h0 : _GEN_9385; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9387 = 8'h6c == _T_442[7:0] ? 4'h0 : _GEN_9386; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9388 = 8'h6d == _T_442[7:0] ? 4'h0 : _GEN_9387; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9389 = 8'h6e == _T_442[7:0] ? 4'h2 : _GEN_9388; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9390 = 8'h6f == _T_442[7:0] ? 4'h0 : _GEN_9389; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9391 = 8'h70 == _T_442[7:0] ? 4'h0 : _GEN_9390; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9392 = 8'h71 == _T_442[7:0] ? 4'h0 : _GEN_9391; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9393 = 8'h72 == _T_442[7:0] ? 4'h2 : _GEN_9392; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9394 = 8'h73 == _T_442[7:0] ? 4'h9 : _GEN_9393; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9395 = 8'h74 == _T_442[7:0] ? 4'h2 : _GEN_9394; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9396 = 8'h75 == _T_442[7:0] ? 4'h0 : _GEN_9395; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9397 = 8'h76 == _T_442[7:0] ? 4'h0 : _GEN_9396; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9398 = 8'h77 == _T_442[7:0] ? 4'h0 : _GEN_9397; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9399 = 8'h78 == _T_442[7:0] ? 4'h1 : _GEN_9398; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9400 = 8'h79 == _T_442[7:0] ? 4'h1 : _GEN_9399; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9401 = 8'h7a == _T_442[7:0] ? 4'h0 : _GEN_9400; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9402 = 8'h7b == _T_442[7:0] ? 4'h0 : _GEN_9401; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9403 = 8'h7c == _T_442[7:0] ? 4'h0 : _GEN_9402; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9404 = 8'h7d == _T_442[7:0] ? 4'h0 : _GEN_9403; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9405 = 8'h7e == _T_442[7:0] ? 4'h0 : _GEN_9404; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9406 = 8'h7f == _T_442[7:0] ? 4'h0 : _GEN_9405; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9407 = 8'h80 == _T_442[7:0] ? 4'h0 : _GEN_9406; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9408 = 8'h81 == _T_442[7:0] ? 4'h0 : _GEN_9407; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9409 = 8'h82 == _T_442[7:0] ? 4'h2 : _GEN_9408; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9410 = 8'h83 == _T_442[7:0] ? 4'h0 : _GEN_9409; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9411 = 8'h84 == _T_442[7:0] ? 4'h0 : _GEN_9410; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9412 = 8'h85 == _T_442[7:0] ? 4'h0 : _GEN_9411; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9413 = 8'h86 == _T_442[7:0] ? 4'h7 : _GEN_9412; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9414 = 8'h87 == _T_442[7:0] ? 4'h2 : _GEN_9413; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9415 = 8'h88 == _T_442[7:0] ? 4'h0 : _GEN_9414; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9416 = 8'h89 == _T_442[7:0] ? 4'h2 : _GEN_9415; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9417 = 8'h8a == _T_442[7:0] ? 4'h7 : _GEN_9416; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9418 = 8'h8b == _T_442[7:0] ? 4'h0 : _GEN_9417; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9419 = 8'h8c == _T_442[7:0] ? 4'h0 : _GEN_9418; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9420 = 8'h8d == _T_442[7:0] ? 4'h0 : _GEN_9419; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9421 = 8'h8e == _T_442[7:0] ? 4'h2 : _GEN_9420; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9422 = 8'h8f == _T_442[7:0] ? 4'h0 : _GEN_9421; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9423 = 8'h90 == _T_442[7:0] ? 4'h0 : _GEN_9422; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9424 = 8'h91 == _T_442[7:0] ? 4'h0 : _GEN_9423; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9425 = 8'h92 == _T_442[7:0] ? 4'h0 : _GEN_9424; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9426 = 8'h93 == _T_442[7:0] ? 4'h0 : _GEN_9425; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9427 = 8'h94 == _T_442[7:0] ? 4'h0 : _GEN_9426; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9428 = 8'h95 == _T_442[7:0] ? 4'h0 : _GEN_9427; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9429 = 8'h96 == _T_442[7:0] ? 4'h0 : _GEN_9428; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9430 = 8'h97 == _T_442[7:0] ? 4'h2 : _GEN_9429; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9431 = 8'h98 == _T_442[7:0] ? 4'h2 : _GEN_9430; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9432 = 8'h99 == _T_442[7:0] ? 4'h1 : _GEN_9431; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9433 = 8'h9a == _T_442[7:0] ? 4'h0 : _GEN_9432; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9434 = 8'h9b == _T_442[7:0] ? 4'h7 : _GEN_9433; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9435 = 8'h9c == _T_442[7:0] ? 4'h7 : _GEN_9434; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9436 = 8'h9d == _T_442[7:0] ? 4'h0 : _GEN_9435; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9437 = 8'h9e == _T_442[7:0] ? 4'h7 : _GEN_9436; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9438 = 8'h9f == _T_442[7:0] ? 4'h7 : _GEN_9437; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9439 = 8'ha0 == _T_442[7:0] ? 4'h0 : _GEN_9438; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9440 = 8'ha1 == _T_442[7:0] ? 4'h1 : _GEN_9439; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9441 = 8'ha2 == _T_442[7:0] ? 4'h2 : _GEN_9440; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9442 = 8'ha3 == _T_442[7:0] ? 4'h2 : _GEN_9441; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9443 = 8'ha4 == _T_442[7:0] ? 4'h0 : _GEN_9442; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9444 = 8'ha5 == _T_442[7:0] ? 4'h0 : _GEN_9443; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9445 = 8'ha6 == _T_442[7:0] ? 4'h0 : _GEN_9444; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9446 = 8'ha7 == _T_442[7:0] ? 4'h0 : _GEN_9445; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9447 = 8'ha8 == _T_442[7:0] ? 4'h0 : _GEN_9446; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9448 = 8'ha9 == _T_442[7:0] ? 4'h0 : _GEN_9447; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9449 = 8'haa == _T_442[7:0] ? 4'h0 : _GEN_9448; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9450 = 8'hab == _T_442[7:0] ? 4'h0 : _GEN_9449; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9451 = 8'hac == _T_442[7:0] ? 4'h2 : _GEN_9450; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9452 = 8'had == _T_442[7:0] ? 4'h0 : _GEN_9451; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9453 = 8'hae == _T_442[7:0] ? 4'h1 : _GEN_9452; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9454 = 8'haf == _T_442[7:0] ? 4'h3 : _GEN_9453; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9455 = 8'hb0 == _T_442[7:0] ? 4'h1 : _GEN_9454; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9456 = 8'hb1 == _T_442[7:0] ? 4'h0 : _GEN_9455; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9457 = 8'hb2 == _T_442[7:0] ? 4'h0 : _GEN_9456; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9458 = 8'hb3 == _T_442[7:0] ? 4'h0 : _GEN_9457; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9459 = 8'hb4 == _T_442[7:0] ? 4'h1 : _GEN_9458; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9460 = 8'hb5 == _T_442[7:0] ? 4'h3 : _GEN_9459; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9461 = 8'hb6 == _T_442[7:0] ? 4'h1 : _GEN_9460; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9462 = 8'hb7 == _T_442[7:0] ? 4'h0 : _GEN_9461; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9463 = 8'hb8 == _T_442[7:0] ? 4'h2 : _GEN_9462; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9464 = 8'hb9 == _T_442[7:0] ? 4'h0 : _GEN_9463; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9465 = 8'hba == _T_442[7:0] ? 4'h0 : _GEN_9464; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9466 = 8'hbb == _T_442[7:0] ? 4'h0 : _GEN_9465; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9467 = 8'hbc == _T_442[7:0] ? 4'h0 : _GEN_9466; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9468 = 8'hbd == _T_442[7:0] ? 4'h0 : _GEN_9467; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9469 = 8'hbe == _T_442[7:0] ? 4'h0 : _GEN_9468; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9470 = 8'hbf == _T_442[7:0] ? 4'h0 : _GEN_9469; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9471 = 8'hc0 == _T_442[7:0] ? 4'h0 : _GEN_9470; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9472 = 8'hc1 == _T_442[7:0] ? 4'h0 : _GEN_9471; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9473 = 8'hc2 == _T_442[7:0] ? 4'h3 : _GEN_9472; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9474 = 8'hc3 == _T_442[7:0] ? 4'h0 : _GEN_9473; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9475 = 8'hc4 == _T_442[7:0] ? 4'h0 : _GEN_9474; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9476 = 8'hc5 == _T_442[7:0] ? 4'h2 : _GEN_9475; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9477 = 8'hc6 == _T_442[7:0] ? 4'h3 : _GEN_9476; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9478 = 8'hc7 == _T_442[7:0] ? 4'h2 : _GEN_9477; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9479 = 8'hc8 == _T_442[7:0] ? 4'h3 : _GEN_9478; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9480 = 8'hc9 == _T_442[7:0] ? 4'h2 : _GEN_9479; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9481 = 8'hca == _T_442[7:0] ? 4'h0 : _GEN_9480; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9482 = 8'hcb == _T_442[7:0] ? 4'h0 : _GEN_9481; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9483 = 8'hcc == _T_442[7:0] ? 4'h3 : _GEN_9482; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9484 = 8'hcd == _T_442[7:0] ? 4'h0 : _GEN_9483; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9485 = 8'hce == _T_442[7:0] ? 4'h0 : _GEN_9484; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9486 = 8'hcf == _T_442[7:0] ? 4'h0 : _GEN_9485; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9487 = 8'hd0 == _T_442[7:0] ? 4'h0 : _GEN_9486; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9488 = 8'hd1 == _T_442[7:0] ? 4'h0 : _GEN_9487; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9489 = 8'hd2 == _T_442[7:0] ? 4'h0 : _GEN_9488; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9490 = 8'hd3 == _T_442[7:0] ? 4'h0 : _GEN_9489; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9491 = 8'hd4 == _T_442[7:0] ? 4'h0 : _GEN_9490; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9492 = 8'hd5 == _T_442[7:0] ? 4'h0 : _GEN_9491; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9493 = 8'hd6 == _T_442[7:0] ? 4'h0 : _GEN_9492; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9494 = 8'hd7 == _T_442[7:0] ? 4'h2 : _GEN_9493; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9495 = 8'hd8 == _T_442[7:0] ? 4'h2 : _GEN_9494; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9496 = 8'hd9 == _T_442[7:0] ? 4'h0 : _GEN_9495; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9497 = 8'hda == _T_442[7:0] ? 4'h7 : _GEN_9496; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9498 = 8'hdb == _T_442[7:0] ? 4'h1 : _GEN_9497; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9499 = 8'hdc == _T_442[7:0] ? 4'h4 : _GEN_9498; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9500 = 8'hdd == _T_442[7:0] ? 4'h1 : _GEN_9499; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9501 = 8'hde == _T_442[7:0] ? 4'h7 : _GEN_9500; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9502 = 8'hdf == _T_442[7:0] ? 4'h0 : _GEN_9501; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9503 = 8'he0 == _T_442[7:0] ? 4'h2 : _GEN_9502; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9504 = 8'he1 == _T_442[7:0] ? 4'h2 : _GEN_9503; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9505 = 8'he2 == _T_442[7:0] ? 4'h0 : _GEN_9504; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9506 = 8'he3 == _T_442[7:0] ? 4'h0 : _GEN_9505; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9507 = 8'he4 == _T_442[7:0] ? 4'h0 : _GEN_9506; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9508 = 8'he5 == _T_442[7:0] ? 4'h0 : _GEN_9507; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9509 = 8'he6 == _T_442[7:0] ? 4'h0 : _GEN_9508; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9510 = 8'he7 == _T_442[7:0] ? 4'h0 : _GEN_9509; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9511 = 8'he8 == _T_442[7:0] ? 4'h0 : _GEN_9510; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9512 = 8'he9 == _T_442[7:0] ? 4'h0 : _GEN_9511; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9513 = 8'hea == _T_442[7:0] ? 4'h0 : _GEN_9512; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9514 = 8'heb == _T_442[7:0] ? 4'h0 : _GEN_9513; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9515 = 8'hec == _T_442[7:0] ? 4'h0 : _GEN_9514; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9516 = 8'hed == _T_442[7:0] ? 4'h0 : _GEN_9515; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9517 = 8'hee == _T_442[7:0] ? 4'h0 : _GEN_9516; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9518 = 8'hef == _T_442[7:0] ? 4'h0 : _GEN_9517; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9519 = 8'hf0 == _T_442[7:0] ? 4'h0 : _GEN_9518; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9520 = 8'hf1 == _T_442[7:0] ? 4'h0 : _GEN_9519; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9521 = 8'hf2 == _T_442[7:0] ? 4'h0 : _GEN_9520; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9522 = 8'hf3 == _T_442[7:0] ? 4'h0 : _GEN_9521; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9523 = 8'hf4 == _T_442[7:0] ? 4'h0 : _GEN_9522; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9524 = 8'hf5 == _T_442[7:0] ? 4'h0 : _GEN_9523; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9525 = 8'hf6 == _T_442[7:0] ? 4'h0 : _GEN_9524; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9526 = 8'hf7 == _T_442[7:0] ? 4'h0 : _GEN_9525; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9527 = 8'hf8 == _T_442[7:0] ? 4'h0 : _GEN_9526; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9528 = 8'hf9 == _T_442[7:0] ? 4'h0 : _GEN_9527; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9529 = 8'hfa == _T_442[7:0] ? 4'h0 : _GEN_9528; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9530 = 8'hfb == _T_442[7:0] ? 4'h0 : _GEN_9529; // @[Filter.scala 204:62]
  wire [4:0] _GEN_11285 = {{1'd0}, _GEN_9530}; // @[Filter.scala 204:62]
  wire [8:0] _T_444 = _GEN_11285 * 5'h14; // @[Filter.scala 204:62]
  wire [3:0] _GEN_9580 = 8'h31 == _T_442[7:0] ? 4'h3 : _GEN_9327; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9581 = 8'h32 == _T_442[7:0] ? 4'h3 : _GEN_9580; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9582 = 8'h33 == _T_442[7:0] ? 4'h6 : _GEN_9581; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9583 = 8'h34 == _T_442[7:0] ? 4'h6 : _GEN_9582; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9584 = 8'h35 == _T_442[7:0] ? 4'h0 : _GEN_9583; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9585 = 8'h36 == _T_442[7:0] ? 4'h0 : _GEN_9584; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9586 = 8'h37 == _T_442[7:0] ? 4'h0 : _GEN_9585; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9587 = 8'h38 == _T_442[7:0] ? 4'h2 : _GEN_9586; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9588 = 8'h39 == _T_442[7:0] ? 4'h0 : _GEN_9587; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9589 = 8'h3a == _T_442[7:0] ? 4'h0 : _GEN_9588; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9590 = 8'h3b == _T_442[7:0] ? 4'h0 : _GEN_9589; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9591 = 8'h3c == _T_442[7:0] ? 4'h0 : _GEN_9590; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9592 = 8'h3d == _T_442[7:0] ? 4'h0 : _GEN_9591; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9593 = 8'h3e == _T_442[7:0] ? 4'h0 : _GEN_9592; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9594 = 8'h3f == _T_442[7:0] ? 4'h0 : _GEN_9593; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9595 = 8'h40 == _T_442[7:0] ? 4'h0 : _GEN_9594; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9596 = 8'h41 == _T_442[7:0] ? 4'h0 : _GEN_9595; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9597 = 8'h42 == _T_442[7:0] ? 4'h0 : _GEN_9596; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9598 = 8'h43 == _T_442[7:0] ? 4'h0 : _GEN_9597; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9599 = 8'h44 == _T_442[7:0] ? 4'h1 : _GEN_9598; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9600 = 8'h45 == _T_442[7:0] ? 4'h4 : _GEN_9599; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9601 = 8'h46 == _T_442[7:0] ? 4'hb : _GEN_9600; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9602 = 8'h47 == _T_442[7:0] ? 4'h0 : _GEN_9601; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9603 = 8'h48 == _T_442[7:0] ? 4'h0 : _GEN_9602; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9604 = 8'h49 == _T_442[7:0] ? 4'h0 : _GEN_9603; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9605 = 8'h4a == _T_442[7:0] ? 4'h6 : _GEN_9604; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9606 = 8'h4b == _T_442[7:0] ? 4'h0 : _GEN_9605; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9607 = 8'h4c == _T_442[7:0] ? 4'h3 : _GEN_9606; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9608 = 8'h4d == _T_442[7:0] ? 4'h3 : _GEN_9607; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9609 = 8'h4e == _T_442[7:0] ? 4'h2 : _GEN_9608; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9610 = 8'h4f == _T_442[7:0] ? 4'h0 : _GEN_9609; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9611 = 8'h50 == _T_442[7:0] ? 4'h0 : _GEN_9610; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9612 = 8'h51 == _T_442[7:0] ? 4'h0 : _GEN_9611; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9613 = 8'h52 == _T_442[7:0] ? 4'h0 : _GEN_9612; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9614 = 8'h53 == _T_442[7:0] ? 4'h0 : _GEN_9613; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9615 = 8'h54 == _T_442[7:0] ? 4'h0 : _GEN_9614; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9616 = 8'h55 == _T_442[7:0] ? 4'h0 : _GEN_9615; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9617 = 8'h56 == _T_442[7:0] ? 4'h0 : _GEN_9616; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9618 = 8'h57 == _T_442[7:0] ? 4'h0 : _GEN_9617; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9619 = 8'h58 == _T_442[7:0] ? 4'h0 : _GEN_9618; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9620 = 8'h59 == _T_442[7:0] ? 4'h2 : _GEN_9619; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9621 = 8'h5a == _T_442[7:0] ? 4'h3 : _GEN_9620; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9622 = 8'h5b == _T_442[7:0] ? 4'h0 : _GEN_9621; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9623 = 8'h5c == _T_442[7:0] ? 4'h0 : _GEN_9622; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9624 = 8'h5d == _T_442[7:0] ? 4'h3 : _GEN_9623; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9625 = 8'h5e == _T_442[7:0] ? 4'hd : _GEN_9624; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9626 = 8'h5f == _T_442[7:0] ? 4'h3 : _GEN_9625; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9627 = 8'h60 == _T_442[7:0] ? 4'h0 : _GEN_9626; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9628 = 8'h61 == _T_442[7:0] ? 4'h6 : _GEN_9627; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9629 = 8'h62 == _T_442[7:0] ? 4'h0 : _GEN_9628; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9630 = 8'h63 == _T_442[7:0] ? 4'h2 : _GEN_9629; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9631 = 8'h64 == _T_442[7:0] ? 4'h0 : _GEN_9630; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9632 = 8'h65 == _T_442[7:0] ? 4'h0 : _GEN_9631; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9633 = 8'h66 == _T_442[7:0] ? 4'h0 : _GEN_9632; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9634 = 8'h67 == _T_442[7:0] ? 4'h0 : _GEN_9633; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9635 = 8'h68 == _T_442[7:0] ? 4'h0 : _GEN_9634; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9636 = 8'h69 == _T_442[7:0] ? 4'h0 : _GEN_9635; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9637 = 8'h6a == _T_442[7:0] ? 4'h0 : _GEN_9636; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9638 = 8'h6b == _T_442[7:0] ? 4'h0 : _GEN_9637; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9639 = 8'h6c == _T_442[7:0] ? 4'h0 : _GEN_9638; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9640 = 8'h6d == _T_442[7:0] ? 4'h0 : _GEN_9639; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9641 = 8'h6e == _T_442[7:0] ? 4'h2 : _GEN_9640; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9642 = 8'h6f == _T_442[7:0] ? 4'h0 : _GEN_9641; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9643 = 8'h70 == _T_442[7:0] ? 4'h0 : _GEN_9642; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9644 = 8'h71 == _T_442[7:0] ? 4'h0 : _GEN_9643; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9645 = 8'h72 == _T_442[7:0] ? 4'h6 : _GEN_9644; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9646 = 8'h73 == _T_442[7:0] ? 4'he : _GEN_9645; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9647 = 8'h74 == _T_442[7:0] ? 4'h6 : _GEN_9646; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9648 = 8'h75 == _T_442[7:0] ? 4'h0 : _GEN_9647; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9649 = 8'h76 == _T_442[7:0] ? 4'h6 : _GEN_9648; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9650 = 8'h77 == _T_442[7:0] ? 4'h3 : _GEN_9649; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9651 = 8'h78 == _T_442[7:0] ? 4'h4 : _GEN_9650; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9652 = 8'h79 == _T_442[7:0] ? 4'h1 : _GEN_9651; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9653 = 8'h7a == _T_442[7:0] ? 4'h0 : _GEN_9652; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9654 = 8'h7b == _T_442[7:0] ? 4'h0 : _GEN_9653; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9655 = 8'h7c == _T_442[7:0] ? 4'h0 : _GEN_9654; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9656 = 8'h7d == _T_442[7:0] ? 4'h0 : _GEN_9655; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9657 = 8'h7e == _T_442[7:0] ? 4'h0 : _GEN_9656; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9658 = 8'h7f == _T_442[7:0] ? 4'h0 : _GEN_9657; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9659 = 8'h80 == _T_442[7:0] ? 4'h0 : _GEN_9658; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9660 = 8'h81 == _T_442[7:0] ? 4'h0 : _GEN_9659; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9661 = 8'h82 == _T_442[7:0] ? 4'h2 : _GEN_9660; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9662 = 8'h83 == _T_442[7:0] ? 4'h3 : _GEN_9661; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9663 = 8'h84 == _T_442[7:0] ? 4'h6 : _GEN_9662; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9664 = 8'h85 == _T_442[7:0] ? 4'h6 : _GEN_9663; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9665 = 8'h86 == _T_442[7:0] ? 4'he : _GEN_9664; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9666 = 8'h87 == _T_442[7:0] ? 4'ha : _GEN_9665; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9667 = 8'h88 == _T_442[7:0] ? 4'h6 : _GEN_9666; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9668 = 8'h89 == _T_442[7:0] ? 4'ha : _GEN_9667; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9669 = 8'h8a == _T_442[7:0] ? 4'he : _GEN_9668; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9670 = 8'h8b == _T_442[7:0] ? 4'h3 : _GEN_9669; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9671 = 8'h8c == _T_442[7:0] ? 4'h3 : _GEN_9670; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9672 = 8'h8d == _T_442[7:0] ? 4'h0 : _GEN_9671; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9673 = 8'h8e == _T_442[7:0] ? 4'h2 : _GEN_9672; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9674 = 8'h8f == _T_442[7:0] ? 4'h0 : _GEN_9673; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9675 = 8'h90 == _T_442[7:0] ? 4'h0 : _GEN_9674; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9676 = 8'h91 == _T_442[7:0] ? 4'h0 : _GEN_9675; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9677 = 8'h92 == _T_442[7:0] ? 4'h0 : _GEN_9676; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9678 = 8'h93 == _T_442[7:0] ? 4'h0 : _GEN_9677; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9679 = 8'h94 == _T_442[7:0] ? 4'h0 : _GEN_9678; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9680 = 8'h95 == _T_442[7:0] ? 4'h0 : _GEN_9679; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9681 = 8'h96 == _T_442[7:0] ? 4'h0 : _GEN_9680; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9682 = 8'h97 == _T_442[7:0] ? 4'h2 : _GEN_9681; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9683 = 8'h98 == _T_442[7:0] ? 4'h2 : _GEN_9682; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9684 = 8'h99 == _T_442[7:0] ? 4'h1 : _GEN_9683; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9685 = 8'h9a == _T_442[7:0] ? 4'h3 : _GEN_9684; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9686 = 8'h9b == _T_442[7:0] ? 4'he : _GEN_9685; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9687 = 8'h9c == _T_442[7:0] ? 4'he : _GEN_9686; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9688 = 8'h9d == _T_442[7:0] ? 4'h0 : _GEN_9687; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9689 = 8'h9e == _T_442[7:0] ? 4'he : _GEN_9688; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9690 = 8'h9f == _T_442[7:0] ? 4'he : _GEN_9689; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9691 = 8'ha0 == _T_442[7:0] ? 4'h3 : _GEN_9690; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9692 = 8'ha1 == _T_442[7:0] ? 4'h1 : _GEN_9691; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9693 = 8'ha2 == _T_442[7:0] ? 4'h2 : _GEN_9692; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9694 = 8'ha3 == _T_442[7:0] ? 4'h2 : _GEN_9693; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9695 = 8'ha4 == _T_442[7:0] ? 4'h0 : _GEN_9694; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9696 = 8'ha5 == _T_442[7:0] ? 4'h0 : _GEN_9695; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9697 = 8'ha6 == _T_442[7:0] ? 4'h0 : _GEN_9696; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9698 = 8'ha7 == _T_442[7:0] ? 4'h0 : _GEN_9697; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9699 = 8'ha8 == _T_442[7:0] ? 4'h0 : _GEN_9698; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9700 = 8'ha9 == _T_442[7:0] ? 4'h0 : _GEN_9699; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9701 = 8'haa == _T_442[7:0] ? 4'h0 : _GEN_9700; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9702 = 8'hab == _T_442[7:0] ? 4'h0 : _GEN_9701; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9703 = 8'hac == _T_442[7:0] ? 4'h2 : _GEN_9702; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9704 = 8'had == _T_442[7:0] ? 4'h3 : _GEN_9703; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9705 = 8'hae == _T_442[7:0] ? 4'h4 : _GEN_9704; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9706 = 8'haf == _T_442[7:0] ? 4'h3 : _GEN_9705; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9707 = 8'hb0 == _T_442[7:0] ? 4'h4 : _GEN_9706; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9708 = 8'hb1 == _T_442[7:0] ? 4'h3 : _GEN_9707; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9709 = 8'hb2 == _T_442[7:0] ? 4'h0 : _GEN_9708; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9710 = 8'hb3 == _T_442[7:0] ? 4'h3 : _GEN_9709; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9711 = 8'hb4 == _T_442[7:0] ? 4'h4 : _GEN_9710; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9712 = 8'hb5 == _T_442[7:0] ? 4'h3 : _GEN_9711; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9713 = 8'hb6 == _T_442[7:0] ? 4'h4 : _GEN_9712; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9714 = 8'hb7 == _T_442[7:0] ? 4'h3 : _GEN_9713; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9715 = 8'hb8 == _T_442[7:0] ? 4'h2 : _GEN_9714; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9716 = 8'hb9 == _T_442[7:0] ? 4'h0 : _GEN_9715; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9717 = 8'hba == _T_442[7:0] ? 4'h0 : _GEN_9716; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9718 = 8'hbb == _T_442[7:0] ? 4'h0 : _GEN_9717; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9719 = 8'hbc == _T_442[7:0] ? 4'h0 : _GEN_9718; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9720 = 8'hbd == _T_442[7:0] ? 4'h0 : _GEN_9719; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9721 = 8'hbe == _T_442[7:0] ? 4'h0 : _GEN_9720; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9722 = 8'hbf == _T_442[7:0] ? 4'h0 : _GEN_9721; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9723 = 8'hc0 == _T_442[7:0] ? 4'h0 : _GEN_9722; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9724 = 8'hc1 == _T_442[7:0] ? 4'h0 : _GEN_9723; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9725 = 8'hc2 == _T_442[7:0] ? 4'h8 : _GEN_9724; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9726 = 8'hc3 == _T_442[7:0] ? 4'hc : _GEN_9725; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9727 = 8'hc4 == _T_442[7:0] ? 4'h0 : _GEN_9726; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9728 = 8'hc5 == _T_442[7:0] ? 4'h2 : _GEN_9727; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9729 = 8'hc6 == _T_442[7:0] ? 4'h3 : _GEN_9728; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9730 = 8'hc7 == _T_442[7:0] ? 4'h2 : _GEN_9729; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9731 = 8'hc8 == _T_442[7:0] ? 4'h3 : _GEN_9730; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9732 = 8'hc9 == _T_442[7:0] ? 4'h2 : _GEN_9731; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9733 = 8'hca == _T_442[7:0] ? 4'h0 : _GEN_9732; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9734 = 8'hcb == _T_442[7:0] ? 4'hc : _GEN_9733; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9735 = 8'hcc == _T_442[7:0] ? 4'h8 : _GEN_9734; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9736 = 8'hcd == _T_442[7:0] ? 4'h0 : _GEN_9735; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9737 = 8'hce == _T_442[7:0] ? 4'h0 : _GEN_9736; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9738 = 8'hcf == _T_442[7:0] ? 4'h0 : _GEN_9737; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9739 = 8'hd0 == _T_442[7:0] ? 4'h0 : _GEN_9738; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9740 = 8'hd1 == _T_442[7:0] ? 4'h0 : _GEN_9739; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9741 = 8'hd2 == _T_442[7:0] ? 4'h0 : _GEN_9740; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9742 = 8'hd3 == _T_442[7:0] ? 4'h0 : _GEN_9741; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9743 = 8'hd4 == _T_442[7:0] ? 4'h0 : _GEN_9742; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9744 = 8'hd5 == _T_442[7:0] ? 4'h0 : _GEN_9743; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9745 = 8'hd6 == _T_442[7:0] ? 4'h0 : _GEN_9744; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9746 = 8'hd7 == _T_442[7:0] ? 4'h3 : _GEN_9745; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9747 = 8'hd8 == _T_442[7:0] ? 4'h6 : _GEN_9746; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9748 = 8'hd9 == _T_442[7:0] ? 4'h0 : _GEN_9747; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9749 = 8'hda == _T_442[7:0] ? 4'hb : _GEN_9748; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9750 = 8'hdb == _T_442[7:0] ? 4'h1 : _GEN_9749; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9751 = 8'hdc == _T_442[7:0] ? 4'h4 : _GEN_9750; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9752 = 8'hdd == _T_442[7:0] ? 4'h1 : _GEN_9751; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9753 = 8'hde == _T_442[7:0] ? 4'hb : _GEN_9752; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9754 = 8'hdf == _T_442[7:0] ? 4'h0 : _GEN_9753; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9755 = 8'he0 == _T_442[7:0] ? 4'h6 : _GEN_9754; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9756 = 8'he1 == _T_442[7:0] ? 4'h3 : _GEN_9755; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9757 = 8'he2 == _T_442[7:0] ? 4'h0 : _GEN_9756; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9758 = 8'he3 == _T_442[7:0] ? 4'h0 : _GEN_9757; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9759 = 8'he4 == _T_442[7:0] ? 4'h0 : _GEN_9758; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9760 = 8'he5 == _T_442[7:0] ? 4'h0 : _GEN_9759; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9761 = 8'he6 == _T_442[7:0] ? 4'h0 : _GEN_9760; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9762 = 8'he7 == _T_442[7:0] ? 4'h0 : _GEN_9761; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9763 = 8'he8 == _T_442[7:0] ? 4'h0 : _GEN_9762; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9764 = 8'he9 == _T_442[7:0] ? 4'h0 : _GEN_9763; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9765 = 8'hea == _T_442[7:0] ? 4'h0 : _GEN_9764; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9766 = 8'heb == _T_442[7:0] ? 4'h0 : _GEN_9765; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9767 = 8'hec == _T_442[7:0] ? 4'h0 : _GEN_9766; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9768 = 8'hed == _T_442[7:0] ? 4'h0 : _GEN_9767; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9769 = 8'hee == _T_442[7:0] ? 4'h0 : _GEN_9768; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9770 = 8'hef == _T_442[7:0] ? 4'h0 : _GEN_9769; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9771 = 8'hf0 == _T_442[7:0] ? 4'h0 : _GEN_9770; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9772 = 8'hf1 == _T_442[7:0] ? 4'h0 : _GEN_9771; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9773 = 8'hf2 == _T_442[7:0] ? 4'h0 : _GEN_9772; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9774 = 8'hf3 == _T_442[7:0] ? 4'h0 : _GEN_9773; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9775 = 8'hf4 == _T_442[7:0] ? 4'h0 : _GEN_9774; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9776 = 8'hf5 == _T_442[7:0] ? 4'h0 : _GEN_9775; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9777 = 8'hf6 == _T_442[7:0] ? 4'h0 : _GEN_9776; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9778 = 8'hf7 == _T_442[7:0] ? 4'h0 : _GEN_9777; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9779 = 8'hf8 == _T_442[7:0] ? 4'h0 : _GEN_9778; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9780 = 8'hf9 == _T_442[7:0] ? 4'h0 : _GEN_9779; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9781 = 8'hfa == _T_442[7:0] ? 4'h0 : _GEN_9780; // @[Filter.scala 204:102]
  wire [3:0] _GEN_9782 = 8'hfb == _T_442[7:0] ? 4'h0 : _GEN_9781; // @[Filter.scala 204:102]
  wire [6:0] _GEN_11287 = {{3'd0}, _GEN_9782}; // @[Filter.scala 204:102]
  wire [10:0] _T_449 = _GEN_11287 * 7'h46; // @[Filter.scala 204:102]
  wire [10:0] _GEN_11288 = {{2'd0}, _T_444}; // @[Filter.scala 204:69]
  wire [10:0] _T_451 = _GEN_11288 + _T_449; // @[Filter.scala 204:69]
  wire [3:0] _GEN_9791 = 8'h8 == _T_442[7:0] ? 4'h3 : 4'h0; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9792 = 8'h9 == _T_442[7:0] ? 4'h6 : _GEN_9791; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9793 = 8'ha == _T_442[7:0] ? 4'h6 : _GEN_9792; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9794 = 8'hb == _T_442[7:0] ? 4'h6 : _GEN_9793; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9795 = 8'hc == _T_442[7:0] ? 4'h3 : _GEN_9794; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9796 = 8'hd == _T_442[7:0] ? 4'h0 : _GEN_9795; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9797 = 8'he == _T_442[7:0] ? 4'h0 : _GEN_9796; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9798 = 8'hf == _T_442[7:0] ? 4'h0 : _GEN_9797; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9799 = 8'h10 == _T_442[7:0] ? 4'h0 : _GEN_9798; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9800 = 8'h11 == _T_442[7:0] ? 4'h0 : _GEN_9799; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9801 = 8'h12 == _T_442[7:0] ? 4'h0 : _GEN_9800; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9802 = 8'h13 == _T_442[7:0] ? 4'h0 : _GEN_9801; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9803 = 8'h14 == _T_442[7:0] ? 4'h0 : _GEN_9802; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9804 = 8'h15 == _T_442[7:0] ? 4'h0 : _GEN_9803; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9805 = 8'h16 == _T_442[7:0] ? 4'h0 : _GEN_9804; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9806 = 8'h17 == _T_442[7:0] ? 4'h0 : _GEN_9805; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9807 = 8'h18 == _T_442[7:0] ? 4'h0 : _GEN_9806; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9808 = 8'h19 == _T_442[7:0] ? 4'h0 : _GEN_9807; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9809 = 8'h1a == _T_442[7:0] ? 4'h0 : _GEN_9808; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9810 = 8'h1b == _T_442[7:0] ? 4'h0 : _GEN_9809; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9811 = 8'h1c == _T_442[7:0] ? 4'h6 : _GEN_9810; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9812 = 8'h1d == _T_442[7:0] ? 4'h3 : _GEN_9811; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9813 = 8'h1e == _T_442[7:0] ? 4'h0 : _GEN_9812; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9814 = 8'h1f == _T_442[7:0] ? 4'h0 : _GEN_9813; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9815 = 8'h20 == _T_442[7:0] ? 4'h0 : _GEN_9814; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9816 = 8'h21 == _T_442[7:0] ? 4'h3 : _GEN_9815; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9817 = 8'h22 == _T_442[7:0] ? 4'h6 : _GEN_9816; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9818 = 8'h23 == _T_442[7:0] ? 4'h0 : _GEN_9817; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9819 = 8'h24 == _T_442[7:0] ? 4'h0 : _GEN_9818; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9820 = 8'h25 == _T_442[7:0] ? 4'h0 : _GEN_9819; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9821 = 8'h26 == _T_442[7:0] ? 4'h0 : _GEN_9820; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9822 = 8'h27 == _T_442[7:0] ? 4'h0 : _GEN_9821; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9823 = 8'h28 == _T_442[7:0] ? 4'h0 : _GEN_9822; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9824 = 8'h29 == _T_442[7:0] ? 4'h0 : _GEN_9823; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9825 = 8'h2a == _T_442[7:0] ? 4'h0 : _GEN_9824; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9826 = 8'h2b == _T_442[7:0] ? 4'h0 : _GEN_9825; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9827 = 8'h2c == _T_442[7:0] ? 4'h0 : _GEN_9826; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9828 = 8'h2d == _T_442[7:0] ? 4'h0 : _GEN_9827; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9829 = 8'h2e == _T_442[7:0] ? 4'h0 : _GEN_9828; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9830 = 8'h2f == _T_442[7:0] ? 4'h0 : _GEN_9829; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9831 = 8'h30 == _T_442[7:0] ? 4'h6 : _GEN_9830; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9832 = 8'h31 == _T_442[7:0] ? 4'h3 : _GEN_9831; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9833 = 8'h32 == _T_442[7:0] ? 4'h0 : _GEN_9832; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9834 = 8'h33 == _T_442[7:0] ? 4'h1 : _GEN_9833; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9835 = 8'h34 == _T_442[7:0] ? 4'h1 : _GEN_9834; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9836 = 8'h35 == _T_442[7:0] ? 4'h0 : _GEN_9835; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9837 = 8'h36 == _T_442[7:0] ? 4'h0 : _GEN_9836; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9838 = 8'h37 == _T_442[7:0] ? 4'h0 : _GEN_9837; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9839 = 8'h38 == _T_442[7:0] ? 4'h6 : _GEN_9838; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9840 = 8'h39 == _T_442[7:0] ? 4'h0 : _GEN_9839; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9841 = 8'h3a == _T_442[7:0] ? 4'h0 : _GEN_9840; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9842 = 8'h3b == _T_442[7:0] ? 4'h0 : _GEN_9841; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9843 = 8'h3c == _T_442[7:0] ? 4'h0 : _GEN_9842; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9844 = 8'h3d == _T_442[7:0] ? 4'h0 : _GEN_9843; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9845 = 8'h3e == _T_442[7:0] ? 4'h0 : _GEN_9844; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9846 = 8'h3f == _T_442[7:0] ? 4'h0 : _GEN_9845; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9847 = 8'h40 == _T_442[7:0] ? 4'h0 : _GEN_9846; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9848 = 8'h41 == _T_442[7:0] ? 4'h0 : _GEN_9847; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9849 = 8'h42 == _T_442[7:0] ? 4'h0 : _GEN_9848; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9850 = 8'h43 == _T_442[7:0] ? 4'h0 : _GEN_9849; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9851 = 8'h44 == _T_442[7:0] ? 4'h3 : _GEN_9850; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9852 = 8'h45 == _T_442[7:0] ? 4'h6 : _GEN_9851; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9853 = 8'h46 == _T_442[7:0] ? 4'h9 : _GEN_9852; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9854 = 8'h47 == _T_442[7:0] ? 4'h0 : _GEN_9853; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9855 = 8'h48 == _T_442[7:0] ? 4'h0 : _GEN_9854; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9856 = 8'h49 == _T_442[7:0] ? 4'h0 : _GEN_9855; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9857 = 8'h4a == _T_442[7:0] ? 4'h1 : _GEN_9856; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9858 = 8'h4b == _T_442[7:0] ? 4'h0 : _GEN_9857; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9859 = 8'h4c == _T_442[7:0] ? 4'h0 : _GEN_9858; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9860 = 8'h4d == _T_442[7:0] ? 4'h0 : _GEN_9859; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9861 = 8'h4e == _T_442[7:0] ? 4'h6 : _GEN_9860; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9862 = 8'h4f == _T_442[7:0] ? 4'h0 : _GEN_9861; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9863 = 8'h50 == _T_442[7:0] ? 4'h0 : _GEN_9862; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9864 = 8'h51 == _T_442[7:0] ? 4'h0 : _GEN_9863; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9865 = 8'h52 == _T_442[7:0] ? 4'h0 : _GEN_9864; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9866 = 8'h53 == _T_442[7:0] ? 4'h0 : _GEN_9865; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9867 = 8'h54 == _T_442[7:0] ? 4'h0 : _GEN_9866; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9868 = 8'h55 == _T_442[7:0] ? 4'h0 : _GEN_9867; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9869 = 8'h56 == _T_442[7:0] ? 4'h0 : _GEN_9868; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9870 = 8'h57 == _T_442[7:0] ? 4'h0 : _GEN_9869; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9871 = 8'h58 == _T_442[7:0] ? 4'h0 : _GEN_9870; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9872 = 8'h59 == _T_442[7:0] ? 4'h6 : _GEN_9871; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9873 = 8'h5a == _T_442[7:0] ? 4'h3 : _GEN_9872; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9874 = 8'h5b == _T_442[7:0] ? 4'h0 : _GEN_9873; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9875 = 8'h5c == _T_442[7:0] ? 4'h0 : _GEN_9874; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9876 = 8'h5d == _T_442[7:0] ? 4'h0 : _GEN_9875; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9877 = 8'h5e == _T_442[7:0] ? 4'h7 : _GEN_9876; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9878 = 8'h5f == _T_442[7:0] ? 4'h0 : _GEN_9877; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9879 = 8'h60 == _T_442[7:0] ? 4'h0 : _GEN_9878; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9880 = 8'h61 == _T_442[7:0] ? 4'h1 : _GEN_9879; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9881 = 8'h62 == _T_442[7:0] ? 4'h0 : _GEN_9880; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9882 = 8'h63 == _T_442[7:0] ? 4'h6 : _GEN_9881; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9883 = 8'h64 == _T_442[7:0] ? 4'h0 : _GEN_9882; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9884 = 8'h65 == _T_442[7:0] ? 4'h0 : _GEN_9883; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9885 = 8'h66 == _T_442[7:0] ? 4'h0 : _GEN_9884; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9886 = 8'h67 == _T_442[7:0] ? 4'h0 : _GEN_9885; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9887 = 8'h68 == _T_442[7:0] ? 4'h0 : _GEN_9886; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9888 = 8'h69 == _T_442[7:0] ? 4'h0 : _GEN_9887; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9889 = 8'h6a == _T_442[7:0] ? 4'h0 : _GEN_9888; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9890 = 8'h6b == _T_442[7:0] ? 4'h0 : _GEN_9889; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9891 = 8'h6c == _T_442[7:0] ? 4'h0 : _GEN_9890; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9892 = 8'h6d == _T_442[7:0] ? 4'h0 : _GEN_9891; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9893 = 8'h6e == _T_442[7:0] ? 4'h6 : _GEN_9892; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9894 = 8'h6f == _T_442[7:0] ? 4'h0 : _GEN_9893; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9895 = 8'h70 == _T_442[7:0] ? 4'h0 : _GEN_9894; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9896 = 8'h71 == _T_442[7:0] ? 4'h0 : _GEN_9895; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9897 = 8'h72 == _T_442[7:0] ? 4'h3 : _GEN_9896; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9898 = 8'h73 == _T_442[7:0] ? 4'hc : _GEN_9897; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9899 = 8'h74 == _T_442[7:0] ? 4'h3 : _GEN_9898; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9900 = 8'h75 == _T_442[7:0] ? 4'h0 : _GEN_9899; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9901 = 8'h76 == _T_442[7:0] ? 4'h1 : _GEN_9900; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9902 = 8'h77 == _T_442[7:0] ? 4'h0 : _GEN_9901; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9903 = 8'h78 == _T_442[7:0] ? 4'h3 : _GEN_9902; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9904 = 8'h79 == _T_442[7:0] ? 4'h3 : _GEN_9903; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9905 = 8'h7a == _T_442[7:0] ? 4'h0 : _GEN_9904; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9906 = 8'h7b == _T_442[7:0] ? 4'h0 : _GEN_9905; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9907 = 8'h7c == _T_442[7:0] ? 4'h0 : _GEN_9906; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9908 = 8'h7d == _T_442[7:0] ? 4'h0 : _GEN_9907; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9909 = 8'h7e == _T_442[7:0] ? 4'h0 : _GEN_9908; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9910 = 8'h7f == _T_442[7:0] ? 4'h0 : _GEN_9909; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9911 = 8'h80 == _T_442[7:0] ? 4'h0 : _GEN_9910; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9912 = 8'h81 == _T_442[7:0] ? 4'h0 : _GEN_9911; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9913 = 8'h82 == _T_442[7:0] ? 4'h6 : _GEN_9912; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9914 = 8'h83 == _T_442[7:0] ? 4'h0 : _GEN_9913; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9915 = 8'h84 == _T_442[7:0] ? 4'h1 : _GEN_9914; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9916 = 8'h85 == _T_442[7:0] ? 4'h1 : _GEN_9915; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9917 = 8'h86 == _T_442[7:0] ? 4'ha : _GEN_9916; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9918 = 8'h87 == _T_442[7:0] ? 4'h4 : _GEN_9917; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9919 = 8'h88 == _T_442[7:0] ? 4'h1 : _GEN_9918; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9920 = 8'h89 == _T_442[7:0] ? 4'h4 : _GEN_9919; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9921 = 8'h8a == _T_442[7:0] ? 4'ha : _GEN_9920; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9922 = 8'h8b == _T_442[7:0] ? 4'h0 : _GEN_9921; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9923 = 8'h8c == _T_442[7:0] ? 4'h0 : _GEN_9922; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9924 = 8'h8d == _T_442[7:0] ? 4'h0 : _GEN_9923; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9925 = 8'h8e == _T_442[7:0] ? 4'h6 : _GEN_9924; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9926 = 8'h8f == _T_442[7:0] ? 4'h0 : _GEN_9925; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9927 = 8'h90 == _T_442[7:0] ? 4'h0 : _GEN_9926; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9928 = 8'h91 == _T_442[7:0] ? 4'h0 : _GEN_9927; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9929 = 8'h92 == _T_442[7:0] ? 4'h0 : _GEN_9928; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9930 = 8'h93 == _T_442[7:0] ? 4'h0 : _GEN_9929; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9931 = 8'h94 == _T_442[7:0] ? 4'h0 : _GEN_9930; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9932 = 8'h95 == _T_442[7:0] ? 4'h0 : _GEN_9931; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9933 = 8'h96 == _T_442[7:0] ? 4'h0 : _GEN_9932; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9934 = 8'h97 == _T_442[7:0] ? 4'h6 : _GEN_9933; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9935 = 8'h98 == _T_442[7:0] ? 4'h6 : _GEN_9934; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9936 = 8'h99 == _T_442[7:0] ? 4'h3 : _GEN_9935; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9937 = 8'h9a == _T_442[7:0] ? 4'h0 : _GEN_9936; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9938 = 8'h9b == _T_442[7:0] ? 4'ha : _GEN_9937; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9939 = 8'h9c == _T_442[7:0] ? 4'ha : _GEN_9938; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9940 = 8'h9d == _T_442[7:0] ? 4'h0 : _GEN_9939; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9941 = 8'h9e == _T_442[7:0] ? 4'ha : _GEN_9940; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9942 = 8'h9f == _T_442[7:0] ? 4'ha : _GEN_9941; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9943 = 8'ha0 == _T_442[7:0] ? 4'h0 : _GEN_9942; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9944 = 8'ha1 == _T_442[7:0] ? 4'h3 : _GEN_9943; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9945 = 8'ha2 == _T_442[7:0] ? 4'h6 : _GEN_9944; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9946 = 8'ha3 == _T_442[7:0] ? 4'h6 : _GEN_9945; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9947 = 8'ha4 == _T_442[7:0] ? 4'h0 : _GEN_9946; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9948 = 8'ha5 == _T_442[7:0] ? 4'h0 : _GEN_9947; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9949 = 8'ha6 == _T_442[7:0] ? 4'h0 : _GEN_9948; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9950 = 8'ha7 == _T_442[7:0] ? 4'h0 : _GEN_9949; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9951 = 8'ha8 == _T_442[7:0] ? 4'h0 : _GEN_9950; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9952 = 8'ha9 == _T_442[7:0] ? 4'h0 : _GEN_9951; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9953 = 8'haa == _T_442[7:0] ? 4'h0 : _GEN_9952; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9954 = 8'hab == _T_442[7:0] ? 4'h0 : _GEN_9953; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9955 = 8'hac == _T_442[7:0] ? 4'h6 : _GEN_9954; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9956 = 8'had == _T_442[7:0] ? 4'h0 : _GEN_9955; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9957 = 8'hae == _T_442[7:0] ? 4'h3 : _GEN_9956; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9958 = 8'haf == _T_442[7:0] ? 4'h9 : _GEN_9957; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9959 = 8'hb0 == _T_442[7:0] ? 4'h3 : _GEN_9958; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9960 = 8'hb1 == _T_442[7:0] ? 4'h0 : _GEN_9959; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9961 = 8'hb2 == _T_442[7:0] ? 4'h0 : _GEN_9960; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9962 = 8'hb3 == _T_442[7:0] ? 4'h0 : _GEN_9961; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9963 = 8'hb4 == _T_442[7:0] ? 4'h3 : _GEN_9962; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9964 = 8'hb5 == _T_442[7:0] ? 4'h9 : _GEN_9963; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9965 = 8'hb6 == _T_442[7:0] ? 4'h3 : _GEN_9964; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9966 = 8'hb7 == _T_442[7:0] ? 4'h0 : _GEN_9965; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9967 = 8'hb8 == _T_442[7:0] ? 4'h6 : _GEN_9966; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9968 = 8'hb9 == _T_442[7:0] ? 4'h0 : _GEN_9967; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9969 = 8'hba == _T_442[7:0] ? 4'h0 : _GEN_9968; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9970 = 8'hbb == _T_442[7:0] ? 4'h0 : _GEN_9969; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9971 = 8'hbc == _T_442[7:0] ? 4'h0 : _GEN_9970; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9972 = 8'hbd == _T_442[7:0] ? 4'h0 : _GEN_9971; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9973 = 8'hbe == _T_442[7:0] ? 4'h0 : _GEN_9972; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9974 = 8'hbf == _T_442[7:0] ? 4'h0 : _GEN_9973; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9975 = 8'hc0 == _T_442[7:0] ? 4'h0 : _GEN_9974; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9976 = 8'hc1 == _T_442[7:0] ? 4'h0 : _GEN_9975; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9977 = 8'hc2 == _T_442[7:0] ? 4'h7 : _GEN_9976; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9978 = 8'hc3 == _T_442[7:0] ? 4'h2 : _GEN_9977; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9979 = 8'hc4 == _T_442[7:0] ? 4'h0 : _GEN_9978; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9980 = 8'hc5 == _T_442[7:0] ? 4'h6 : _GEN_9979; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9981 = 8'hc6 == _T_442[7:0] ? 4'h9 : _GEN_9980; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9982 = 8'hc7 == _T_442[7:0] ? 4'h6 : _GEN_9981; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9983 = 8'hc8 == _T_442[7:0] ? 4'h9 : _GEN_9982; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9984 = 8'hc9 == _T_442[7:0] ? 4'h6 : _GEN_9983; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9985 = 8'hca == _T_442[7:0] ? 4'h0 : _GEN_9984; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9986 = 8'hcb == _T_442[7:0] ? 4'h2 : _GEN_9985; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9987 = 8'hcc == _T_442[7:0] ? 4'h7 : _GEN_9986; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9988 = 8'hcd == _T_442[7:0] ? 4'h0 : _GEN_9987; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9989 = 8'hce == _T_442[7:0] ? 4'h0 : _GEN_9988; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9990 = 8'hcf == _T_442[7:0] ? 4'h0 : _GEN_9989; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9991 = 8'hd0 == _T_442[7:0] ? 4'h0 : _GEN_9990; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9992 = 8'hd1 == _T_442[7:0] ? 4'h0 : _GEN_9991; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9993 = 8'hd2 == _T_442[7:0] ? 4'h0 : _GEN_9992; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9994 = 8'hd3 == _T_442[7:0] ? 4'h0 : _GEN_9993; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9995 = 8'hd4 == _T_442[7:0] ? 4'h0 : _GEN_9994; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9996 = 8'hd5 == _T_442[7:0] ? 4'h0 : _GEN_9995; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9997 = 8'hd6 == _T_442[7:0] ? 4'h0 : _GEN_9996; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9998 = 8'hd7 == _T_442[7:0] ? 4'h3 : _GEN_9997; // @[Filter.scala 204:142]
  wire [3:0] _GEN_9999 = 8'hd8 == _T_442[7:0] ? 4'h3 : _GEN_9998; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10000 = 8'hd9 == _T_442[7:0] ? 4'h0 : _GEN_9999; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10001 = 8'hda == _T_442[7:0] ? 4'h9 : _GEN_10000; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10002 = 8'hdb == _T_442[7:0] ? 4'h3 : _GEN_10001; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10003 = 8'hdc == _T_442[7:0] ? 4'hc : _GEN_10002; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10004 = 8'hdd == _T_442[7:0] ? 4'h3 : _GEN_10003; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10005 = 8'hde == _T_442[7:0] ? 4'h9 : _GEN_10004; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10006 = 8'hdf == _T_442[7:0] ? 4'h0 : _GEN_10005; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10007 = 8'he0 == _T_442[7:0] ? 4'h3 : _GEN_10006; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10008 = 8'he1 == _T_442[7:0] ? 4'h3 : _GEN_10007; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10009 = 8'he2 == _T_442[7:0] ? 4'h0 : _GEN_10008; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10010 = 8'he3 == _T_442[7:0] ? 4'h0 : _GEN_10009; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10011 = 8'he4 == _T_442[7:0] ? 4'h0 : _GEN_10010; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10012 = 8'he5 == _T_442[7:0] ? 4'h0 : _GEN_10011; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10013 = 8'he6 == _T_442[7:0] ? 4'h0 : _GEN_10012; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10014 = 8'he7 == _T_442[7:0] ? 4'h0 : _GEN_10013; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10015 = 8'he8 == _T_442[7:0] ? 4'h0 : _GEN_10014; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10016 = 8'he9 == _T_442[7:0] ? 4'h0 : _GEN_10015; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10017 = 8'hea == _T_442[7:0] ? 4'h0 : _GEN_10016; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10018 = 8'heb == _T_442[7:0] ? 4'h0 : _GEN_10017; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10019 = 8'hec == _T_442[7:0] ? 4'h0 : _GEN_10018; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10020 = 8'hed == _T_442[7:0] ? 4'h0 : _GEN_10019; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10021 = 8'hee == _T_442[7:0] ? 4'h0 : _GEN_10020; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10022 = 8'hef == _T_442[7:0] ? 4'h0 : _GEN_10021; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10023 = 8'hf0 == _T_442[7:0] ? 4'h0 : _GEN_10022; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10024 = 8'hf1 == _T_442[7:0] ? 4'h0 : _GEN_10023; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10025 = 8'hf2 == _T_442[7:0] ? 4'h0 : _GEN_10024; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10026 = 8'hf3 == _T_442[7:0] ? 4'h0 : _GEN_10025; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10027 = 8'hf4 == _T_442[7:0] ? 4'h0 : _GEN_10026; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10028 = 8'hf5 == _T_442[7:0] ? 4'h0 : _GEN_10027; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10029 = 8'hf6 == _T_442[7:0] ? 4'h0 : _GEN_10028; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10030 = 8'hf7 == _T_442[7:0] ? 4'h0 : _GEN_10029; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10031 = 8'hf8 == _T_442[7:0] ? 4'h0 : _GEN_10030; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10032 = 8'hf9 == _T_442[7:0] ? 4'h0 : _GEN_10031; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10033 = 8'hfa == _T_442[7:0] ? 4'h0 : _GEN_10032; // @[Filter.scala 204:142]
  wire [3:0] _GEN_10034 = 8'hfb == _T_442[7:0] ? 4'h0 : _GEN_10033; // @[Filter.scala 204:142]
  wire [7:0] _T_456 = _GEN_10034 * 4'ha; // @[Filter.scala 204:142]
  wire [10:0] _GEN_11290 = {{3'd0}, _T_456}; // @[Filter.scala 204:109]
  wire [10:0] _T_458 = _T_451 + _GEN_11290; // @[Filter.scala 204:109]
  wire [10:0] _T_459 = _T_458 / 11'h64; // @[Filter.scala 204:150]
  wire  _T_461 = _T_432 >= 5'h15; // @[Filter.scala 207:31]
  wire  _T_465 = _T_439 >= 32'hc; // @[Filter.scala 207:63]
  wire  _T_466 = _T_461 | _T_465; // @[Filter.scala 207:58]
  wire [10:0] _GEN_10287 = io_SPI_distort ? _T_459 : {{7'd0}, _GEN_9530}; // @[Filter.scala 209:35]
  wire [10:0] _GEN_10288 = _T_466 ? 11'h0 : _GEN_10287; // @[Filter.scala 207:80]
  wire [10:0] _GEN_10541 = io_SPI_distort ? _T_459 : {{7'd0}, _GEN_9782}; // @[Filter.scala 209:35]
  wire [10:0] _GEN_10542 = _T_466 ? 11'h0 : _GEN_10541; // @[Filter.scala 207:80]
  wire [10:0] _GEN_10795 = io_SPI_distort ? _T_459 : {{7'd0}, _GEN_10034}; // @[Filter.scala 209:35]
  wire [10:0] _GEN_10796 = _T_466 ? 11'h0 : _GEN_10795; // @[Filter.scala 207:80]
  reg [8:0] pixOut_0_0; // @[Filter.scala 218:32]
  reg [8:0] pixOut_0_1; // @[Filter.scala 218:32]
  reg [8:0] pixOut_0_2; // @[Filter.scala 218:32]
  reg [8:0] pixOut_0_3; // @[Filter.scala 218:32]
  reg [8:0] pixOut_0_4; // @[Filter.scala 218:32]
  reg [8:0] pixOut_0_5; // @[Filter.scala 218:32]
  reg [8:0] pixOut_0_6; // @[Filter.scala 218:32]
  reg [8:0] pixOut_1_0; // @[Filter.scala 218:87]
  reg [8:0] pixOut_1_1; // @[Filter.scala 218:87]
  reg [8:0] pixOut_1_2; // @[Filter.scala 218:87]
  reg [8:0] pixOut_1_3; // @[Filter.scala 218:87]
  reg [8:0] pixOut_1_4; // @[Filter.scala 218:87]
  reg [8:0] pixOut_1_5; // @[Filter.scala 218:87]
  reg [8:0] pixOut_1_6; // @[Filter.scala 218:87]
  reg [8:0] pixOut_2_0; // @[Filter.scala 218:142]
  reg [8:0] pixOut_2_1; // @[Filter.scala 218:142]
  reg [8:0] pixOut_2_2; // @[Filter.scala 218:142]
  reg [8:0] pixOut_2_3; // @[Filter.scala 218:142]
  reg [8:0] pixOut_2_4; // @[Filter.scala 218:142]
  reg [8:0] pixOut_2_5; // @[Filter.scala 218:142]
  reg [8:0] pixOut_2_6; // @[Filter.scala 218:142]
  reg  validOut; // @[Filter.scala 219:29]
  wire [7:0] _GEN_10798 = 3'h1 == io_SPI_filterIndex[2:0] ? $signed(8'sh9) : $signed(8'sh1); // @[Filter.scala 223:64]
  wire [7:0] _GEN_10799 = 3'h2 == io_SPI_filterIndex[2:0] ? $signed(8'sh10) : $signed(_GEN_10798); // @[Filter.scala 223:64]
  wire [7:0] _GEN_10800 = 3'h3 == io_SPI_filterIndex[2:0] ? $signed(8'sh1) : $signed(_GEN_10799); // @[Filter.scala 223:64]
  wire [7:0] _GEN_10801 = 3'h4 == io_SPI_filterIndex[2:0] ? $signed(8'sh1) : $signed(_GEN_10800); // @[Filter.scala 223:64]
  wire [7:0] _GEN_10802 = 3'h5 == io_SPI_filterIndex[2:0] ? $signed(8'sh1) : $signed(_GEN_10801); // @[Filter.scala 223:64]
  wire [8:0] _GEN_11294 = {{1{_GEN_10802[7]}},_GEN_10802}; // @[Filter.scala 223:64]
  wire [9:0] _T_497 = $signed(KernelConvolution_io_pixelVal_out_0) / $signed(_GEN_11294); // @[Filter.scala 223:64]
  wire  _T_498 = $signed(pixOut_0_0) < 9'sh0; // @[Filter.scala 225:30]
  wire  _T_499 = _T_498 & io_SPI_invert; // @[Filter.scala 225:36]
  wire  _T_501 = $signed(pixOut_0_0) > 9'shf; // @[Filter.scala 230:36]
  wire  _T_502 = _T_501 & io_SPI_invert; // @[Filter.scala 230:43]
  wire [8:0] _T_506 = 9'hf - pixOut_0_0; // @[Filter.scala 235:43]
  wire [8:0] _GEN_10803 = io_SPI_invert ? _T_506 : pixOut_0_0; // @[Filter.scala 234:36]
  wire [8:0] _GEN_10804 = _T_501 ? 9'hf : _GEN_10803; // @[Filter.scala 232:44]
  wire [8:0] _GEN_10805 = _T_502 ? 9'h0 : _GEN_10804; // @[Filter.scala 230:59]
  wire [8:0] _GEN_10806 = _T_498 ? 9'h0 : _GEN_10805; // @[Filter.scala 227:43]
  wire [8:0] _GEN_10807 = _T_499 ? 9'hf : _GEN_10806; // @[Filter.scala 225:52]
  wire [9:0] _T_508 = $signed(KernelConvolution_io_pixelVal_out_1) / $signed(_GEN_11294); // @[Filter.scala 223:64]
  wire  _T_509 = $signed(pixOut_0_1) < 9'sh0; // @[Filter.scala 225:30]
  wire  _T_510 = _T_509 & io_SPI_invert; // @[Filter.scala 225:36]
  wire  _T_512 = $signed(pixOut_0_1) > 9'shf; // @[Filter.scala 230:36]
  wire  _T_513 = _T_512 & io_SPI_invert; // @[Filter.scala 230:43]
  wire [8:0] _T_517 = 9'hf - pixOut_0_1; // @[Filter.scala 235:43]
  wire [8:0] _GEN_10808 = io_SPI_invert ? _T_517 : pixOut_0_1; // @[Filter.scala 234:36]
  wire [8:0] _GEN_10809 = _T_512 ? 9'hf : _GEN_10808; // @[Filter.scala 232:44]
  wire [8:0] _GEN_10810 = _T_513 ? 9'h0 : _GEN_10809; // @[Filter.scala 230:59]
  wire [8:0] _GEN_10811 = _T_509 ? 9'h0 : _GEN_10810; // @[Filter.scala 227:43]
  wire [8:0] _GEN_10812 = _T_510 ? 9'hf : _GEN_10811; // @[Filter.scala 225:52]
  wire [9:0] _T_519 = $signed(KernelConvolution_io_pixelVal_out_2) / $signed(_GEN_11294); // @[Filter.scala 223:64]
  wire  _T_520 = $signed(pixOut_0_2) < 9'sh0; // @[Filter.scala 225:30]
  wire  _T_521 = _T_520 & io_SPI_invert; // @[Filter.scala 225:36]
  wire  _T_523 = $signed(pixOut_0_2) > 9'shf; // @[Filter.scala 230:36]
  wire  _T_524 = _T_523 & io_SPI_invert; // @[Filter.scala 230:43]
  wire [8:0] _T_528 = 9'hf - pixOut_0_2; // @[Filter.scala 235:43]
  wire [8:0] _GEN_10813 = io_SPI_invert ? _T_528 : pixOut_0_2; // @[Filter.scala 234:36]
  wire [8:0] _GEN_10814 = _T_523 ? 9'hf : _GEN_10813; // @[Filter.scala 232:44]
  wire [8:0] _GEN_10815 = _T_524 ? 9'h0 : _GEN_10814; // @[Filter.scala 230:59]
  wire [8:0] _GEN_10816 = _T_520 ? 9'h0 : _GEN_10815; // @[Filter.scala 227:43]
  wire [8:0] _GEN_10817 = _T_521 ? 9'hf : _GEN_10816; // @[Filter.scala 225:52]
  wire [9:0] _T_530 = $signed(KernelConvolution_io_pixelVal_out_3) / $signed(_GEN_11294); // @[Filter.scala 223:64]
  wire  _T_531 = $signed(pixOut_0_3) < 9'sh0; // @[Filter.scala 225:30]
  wire  _T_532 = _T_531 & io_SPI_invert; // @[Filter.scala 225:36]
  wire  _T_534 = $signed(pixOut_0_3) > 9'shf; // @[Filter.scala 230:36]
  wire  _T_535 = _T_534 & io_SPI_invert; // @[Filter.scala 230:43]
  wire [8:0] _T_539 = 9'hf - pixOut_0_3; // @[Filter.scala 235:43]
  wire [8:0] _GEN_10818 = io_SPI_invert ? _T_539 : pixOut_0_3; // @[Filter.scala 234:36]
  wire [8:0] _GEN_10819 = _T_534 ? 9'hf : _GEN_10818; // @[Filter.scala 232:44]
  wire [8:0] _GEN_10820 = _T_535 ? 9'h0 : _GEN_10819; // @[Filter.scala 230:59]
  wire [8:0] _GEN_10821 = _T_531 ? 9'h0 : _GEN_10820; // @[Filter.scala 227:43]
  wire [8:0] _GEN_10822 = _T_532 ? 9'hf : _GEN_10821; // @[Filter.scala 225:52]
  wire [9:0] _T_541 = $signed(KernelConvolution_io_pixelVal_out_4) / $signed(_GEN_11294); // @[Filter.scala 223:64]
  wire  _T_542 = $signed(pixOut_0_4) < 9'sh0; // @[Filter.scala 225:30]
  wire  _T_543 = _T_542 & io_SPI_invert; // @[Filter.scala 225:36]
  wire  _T_545 = $signed(pixOut_0_4) > 9'shf; // @[Filter.scala 230:36]
  wire  _T_546 = _T_545 & io_SPI_invert; // @[Filter.scala 230:43]
  wire [8:0] _T_550 = 9'hf - pixOut_0_4; // @[Filter.scala 235:43]
  wire [8:0] _GEN_10823 = io_SPI_invert ? _T_550 : pixOut_0_4; // @[Filter.scala 234:36]
  wire [8:0] _GEN_10824 = _T_545 ? 9'hf : _GEN_10823; // @[Filter.scala 232:44]
  wire [8:0] _GEN_10825 = _T_546 ? 9'h0 : _GEN_10824; // @[Filter.scala 230:59]
  wire [8:0] _GEN_10826 = _T_542 ? 9'h0 : _GEN_10825; // @[Filter.scala 227:43]
  wire [8:0] _GEN_10827 = _T_543 ? 9'hf : _GEN_10826; // @[Filter.scala 225:52]
  wire [9:0] _T_552 = $signed(KernelConvolution_io_pixelVal_out_5) / $signed(_GEN_11294); // @[Filter.scala 223:64]
  wire  _T_553 = $signed(pixOut_0_5) < 9'sh0; // @[Filter.scala 225:30]
  wire  _T_554 = _T_553 & io_SPI_invert; // @[Filter.scala 225:36]
  wire  _T_556 = $signed(pixOut_0_5) > 9'shf; // @[Filter.scala 230:36]
  wire  _T_557 = _T_556 & io_SPI_invert; // @[Filter.scala 230:43]
  wire [8:0] _T_561 = 9'hf - pixOut_0_5; // @[Filter.scala 235:43]
  wire [8:0] _GEN_10828 = io_SPI_invert ? _T_561 : pixOut_0_5; // @[Filter.scala 234:36]
  wire [8:0] _GEN_10829 = _T_556 ? 9'hf : _GEN_10828; // @[Filter.scala 232:44]
  wire [8:0] _GEN_10830 = _T_557 ? 9'h0 : _GEN_10829; // @[Filter.scala 230:59]
  wire [8:0] _GEN_10831 = _T_553 ? 9'h0 : _GEN_10830; // @[Filter.scala 227:43]
  wire [8:0] _GEN_10832 = _T_554 ? 9'hf : _GEN_10831; // @[Filter.scala 225:52]
  wire [9:0] _T_563 = $signed(KernelConvolution_io_pixelVal_out_6) / $signed(_GEN_11294); // @[Filter.scala 223:64]
  wire  _T_564 = $signed(pixOut_0_6) < 9'sh0; // @[Filter.scala 225:30]
  wire  _T_565 = _T_564 & io_SPI_invert; // @[Filter.scala 225:36]
  wire  _T_567 = $signed(pixOut_0_6) > 9'shf; // @[Filter.scala 230:36]
  wire  _T_568 = _T_567 & io_SPI_invert; // @[Filter.scala 230:43]
  wire [8:0] _T_572 = 9'hf - pixOut_0_6; // @[Filter.scala 235:43]
  wire [8:0] _GEN_10833 = io_SPI_invert ? _T_572 : pixOut_0_6; // @[Filter.scala 234:36]
  wire [8:0] _GEN_10834 = _T_567 ? 9'hf : _GEN_10833; // @[Filter.scala 232:44]
  wire [8:0] _GEN_10835 = _T_568 ? 9'h0 : _GEN_10834; // @[Filter.scala 230:59]
  wire [8:0] _GEN_10836 = _T_564 ? 9'h0 : _GEN_10835; // @[Filter.scala 227:43]
  wire [8:0] _GEN_10837 = _T_565 ? 9'hf : _GEN_10836; // @[Filter.scala 225:52]
  wire [9:0] _T_574 = $signed(KernelConvolution_1_io_pixelVal_out_0) / $signed(_GEN_11294); // @[Filter.scala 223:64]
  wire  _T_575 = $signed(pixOut_1_0) < 9'sh0; // @[Filter.scala 225:30]
  wire  _T_576 = _T_575 & io_SPI_invert; // @[Filter.scala 225:36]
  wire  _T_578 = $signed(pixOut_1_0) > 9'shf; // @[Filter.scala 230:36]
  wire  _T_579 = _T_578 & io_SPI_invert; // @[Filter.scala 230:43]
  wire [8:0] _T_583 = 9'hf - pixOut_1_0; // @[Filter.scala 235:43]
  wire [8:0] _GEN_10838 = io_SPI_invert ? _T_583 : pixOut_1_0; // @[Filter.scala 234:36]
  wire [8:0] _GEN_10839 = _T_578 ? 9'hf : _GEN_10838; // @[Filter.scala 232:44]
  wire [8:0] _GEN_10840 = _T_579 ? 9'h0 : _GEN_10839; // @[Filter.scala 230:59]
  wire [8:0] _GEN_10841 = _T_575 ? 9'h0 : _GEN_10840; // @[Filter.scala 227:43]
  wire [8:0] _GEN_10842 = _T_576 ? 9'hf : _GEN_10841; // @[Filter.scala 225:52]
  wire [9:0] _T_585 = $signed(KernelConvolution_1_io_pixelVal_out_1) / $signed(_GEN_11294); // @[Filter.scala 223:64]
  wire  _T_586 = $signed(pixOut_1_1) < 9'sh0; // @[Filter.scala 225:30]
  wire  _T_587 = _T_586 & io_SPI_invert; // @[Filter.scala 225:36]
  wire  _T_589 = $signed(pixOut_1_1) > 9'shf; // @[Filter.scala 230:36]
  wire  _T_590 = _T_589 & io_SPI_invert; // @[Filter.scala 230:43]
  wire [8:0] _T_594 = 9'hf - pixOut_1_1; // @[Filter.scala 235:43]
  wire [8:0] _GEN_10843 = io_SPI_invert ? _T_594 : pixOut_1_1; // @[Filter.scala 234:36]
  wire [8:0] _GEN_10844 = _T_589 ? 9'hf : _GEN_10843; // @[Filter.scala 232:44]
  wire [8:0] _GEN_10845 = _T_590 ? 9'h0 : _GEN_10844; // @[Filter.scala 230:59]
  wire [8:0] _GEN_10846 = _T_586 ? 9'h0 : _GEN_10845; // @[Filter.scala 227:43]
  wire [8:0] _GEN_10847 = _T_587 ? 9'hf : _GEN_10846; // @[Filter.scala 225:52]
  wire [9:0] _T_596 = $signed(KernelConvolution_1_io_pixelVal_out_2) / $signed(_GEN_11294); // @[Filter.scala 223:64]
  wire  _T_597 = $signed(pixOut_1_2) < 9'sh0; // @[Filter.scala 225:30]
  wire  _T_598 = _T_597 & io_SPI_invert; // @[Filter.scala 225:36]
  wire  _T_600 = $signed(pixOut_1_2) > 9'shf; // @[Filter.scala 230:36]
  wire  _T_601 = _T_600 & io_SPI_invert; // @[Filter.scala 230:43]
  wire [8:0] _T_605 = 9'hf - pixOut_1_2; // @[Filter.scala 235:43]
  wire [8:0] _GEN_10848 = io_SPI_invert ? _T_605 : pixOut_1_2; // @[Filter.scala 234:36]
  wire [8:0] _GEN_10849 = _T_600 ? 9'hf : _GEN_10848; // @[Filter.scala 232:44]
  wire [8:0] _GEN_10850 = _T_601 ? 9'h0 : _GEN_10849; // @[Filter.scala 230:59]
  wire [8:0] _GEN_10851 = _T_597 ? 9'h0 : _GEN_10850; // @[Filter.scala 227:43]
  wire [8:0] _GEN_10852 = _T_598 ? 9'hf : _GEN_10851; // @[Filter.scala 225:52]
  wire [9:0] _T_607 = $signed(KernelConvolution_1_io_pixelVal_out_3) / $signed(_GEN_11294); // @[Filter.scala 223:64]
  wire  _T_608 = $signed(pixOut_1_3) < 9'sh0; // @[Filter.scala 225:30]
  wire  _T_609 = _T_608 & io_SPI_invert; // @[Filter.scala 225:36]
  wire  _T_611 = $signed(pixOut_1_3) > 9'shf; // @[Filter.scala 230:36]
  wire  _T_612 = _T_611 & io_SPI_invert; // @[Filter.scala 230:43]
  wire [8:0] _T_616 = 9'hf - pixOut_1_3; // @[Filter.scala 235:43]
  wire [8:0] _GEN_10853 = io_SPI_invert ? _T_616 : pixOut_1_3; // @[Filter.scala 234:36]
  wire [8:0] _GEN_10854 = _T_611 ? 9'hf : _GEN_10853; // @[Filter.scala 232:44]
  wire [8:0] _GEN_10855 = _T_612 ? 9'h0 : _GEN_10854; // @[Filter.scala 230:59]
  wire [8:0] _GEN_10856 = _T_608 ? 9'h0 : _GEN_10855; // @[Filter.scala 227:43]
  wire [8:0] _GEN_10857 = _T_609 ? 9'hf : _GEN_10856; // @[Filter.scala 225:52]
  wire [9:0] _T_618 = $signed(KernelConvolution_1_io_pixelVal_out_4) / $signed(_GEN_11294); // @[Filter.scala 223:64]
  wire  _T_619 = $signed(pixOut_1_4) < 9'sh0; // @[Filter.scala 225:30]
  wire  _T_620 = _T_619 & io_SPI_invert; // @[Filter.scala 225:36]
  wire  _T_622 = $signed(pixOut_1_4) > 9'shf; // @[Filter.scala 230:36]
  wire  _T_623 = _T_622 & io_SPI_invert; // @[Filter.scala 230:43]
  wire [8:0] _T_627 = 9'hf - pixOut_1_4; // @[Filter.scala 235:43]
  wire [8:0] _GEN_10858 = io_SPI_invert ? _T_627 : pixOut_1_4; // @[Filter.scala 234:36]
  wire [8:0] _GEN_10859 = _T_622 ? 9'hf : _GEN_10858; // @[Filter.scala 232:44]
  wire [8:0] _GEN_10860 = _T_623 ? 9'h0 : _GEN_10859; // @[Filter.scala 230:59]
  wire [8:0] _GEN_10861 = _T_619 ? 9'h0 : _GEN_10860; // @[Filter.scala 227:43]
  wire [8:0] _GEN_10862 = _T_620 ? 9'hf : _GEN_10861; // @[Filter.scala 225:52]
  wire [9:0] _T_629 = $signed(KernelConvolution_1_io_pixelVal_out_5) / $signed(_GEN_11294); // @[Filter.scala 223:64]
  wire  _T_630 = $signed(pixOut_1_5) < 9'sh0; // @[Filter.scala 225:30]
  wire  _T_631 = _T_630 & io_SPI_invert; // @[Filter.scala 225:36]
  wire  _T_633 = $signed(pixOut_1_5) > 9'shf; // @[Filter.scala 230:36]
  wire  _T_634 = _T_633 & io_SPI_invert; // @[Filter.scala 230:43]
  wire [8:0] _T_638 = 9'hf - pixOut_1_5; // @[Filter.scala 235:43]
  wire [8:0] _GEN_10863 = io_SPI_invert ? _T_638 : pixOut_1_5; // @[Filter.scala 234:36]
  wire [8:0] _GEN_10864 = _T_633 ? 9'hf : _GEN_10863; // @[Filter.scala 232:44]
  wire [8:0] _GEN_10865 = _T_634 ? 9'h0 : _GEN_10864; // @[Filter.scala 230:59]
  wire [8:0] _GEN_10866 = _T_630 ? 9'h0 : _GEN_10865; // @[Filter.scala 227:43]
  wire [8:0] _GEN_10867 = _T_631 ? 9'hf : _GEN_10866; // @[Filter.scala 225:52]
  wire [9:0] _T_640 = $signed(KernelConvolution_1_io_pixelVal_out_6) / $signed(_GEN_11294); // @[Filter.scala 223:64]
  wire  _T_641 = $signed(pixOut_1_6) < 9'sh0; // @[Filter.scala 225:30]
  wire  _T_642 = _T_641 & io_SPI_invert; // @[Filter.scala 225:36]
  wire  _T_644 = $signed(pixOut_1_6) > 9'shf; // @[Filter.scala 230:36]
  wire  _T_645 = _T_644 & io_SPI_invert; // @[Filter.scala 230:43]
  wire [8:0] _T_649 = 9'hf - pixOut_1_6; // @[Filter.scala 235:43]
  wire [8:0] _GEN_10868 = io_SPI_invert ? _T_649 : pixOut_1_6; // @[Filter.scala 234:36]
  wire [8:0] _GEN_10869 = _T_644 ? 9'hf : _GEN_10868; // @[Filter.scala 232:44]
  wire [8:0] _GEN_10870 = _T_645 ? 9'h0 : _GEN_10869; // @[Filter.scala 230:59]
  wire [8:0] _GEN_10871 = _T_641 ? 9'h0 : _GEN_10870; // @[Filter.scala 227:43]
  wire [8:0] _GEN_10872 = _T_642 ? 9'hf : _GEN_10871; // @[Filter.scala 225:52]
  wire [9:0] _T_651 = $signed(KernelConvolution_2_io_pixelVal_out_0) / $signed(_GEN_11294); // @[Filter.scala 223:64]
  wire  _T_652 = $signed(pixOut_2_0) < 9'sh0; // @[Filter.scala 225:30]
  wire  _T_653 = _T_652 & io_SPI_invert; // @[Filter.scala 225:36]
  wire  _T_655 = $signed(pixOut_2_0) > 9'shf; // @[Filter.scala 230:36]
  wire  _T_656 = _T_655 & io_SPI_invert; // @[Filter.scala 230:43]
  wire [8:0] _T_660 = 9'hf - pixOut_2_0; // @[Filter.scala 235:43]
  wire [8:0] _GEN_10873 = io_SPI_invert ? _T_660 : pixOut_2_0; // @[Filter.scala 234:36]
  wire [8:0] _GEN_10874 = _T_655 ? 9'hf : _GEN_10873; // @[Filter.scala 232:44]
  wire [8:0] _GEN_10875 = _T_656 ? 9'h0 : _GEN_10874; // @[Filter.scala 230:59]
  wire [8:0] _GEN_10876 = _T_652 ? 9'h0 : _GEN_10875; // @[Filter.scala 227:43]
  wire [8:0] _GEN_10877 = _T_653 ? 9'hf : _GEN_10876; // @[Filter.scala 225:52]
  wire [9:0] _T_662 = $signed(KernelConvolution_2_io_pixelVal_out_1) / $signed(_GEN_11294); // @[Filter.scala 223:64]
  wire  _T_663 = $signed(pixOut_2_1) < 9'sh0; // @[Filter.scala 225:30]
  wire  _T_664 = _T_663 & io_SPI_invert; // @[Filter.scala 225:36]
  wire  _T_666 = $signed(pixOut_2_1) > 9'shf; // @[Filter.scala 230:36]
  wire  _T_667 = _T_666 & io_SPI_invert; // @[Filter.scala 230:43]
  wire [8:0] _T_671 = 9'hf - pixOut_2_1; // @[Filter.scala 235:43]
  wire [8:0] _GEN_10878 = io_SPI_invert ? _T_671 : pixOut_2_1; // @[Filter.scala 234:36]
  wire [8:0] _GEN_10879 = _T_666 ? 9'hf : _GEN_10878; // @[Filter.scala 232:44]
  wire [8:0] _GEN_10880 = _T_667 ? 9'h0 : _GEN_10879; // @[Filter.scala 230:59]
  wire [8:0] _GEN_10881 = _T_663 ? 9'h0 : _GEN_10880; // @[Filter.scala 227:43]
  wire [8:0] _GEN_10882 = _T_664 ? 9'hf : _GEN_10881; // @[Filter.scala 225:52]
  wire [9:0] _T_673 = $signed(KernelConvolution_2_io_pixelVal_out_2) / $signed(_GEN_11294); // @[Filter.scala 223:64]
  wire  _T_674 = $signed(pixOut_2_2) < 9'sh0; // @[Filter.scala 225:30]
  wire  _T_675 = _T_674 & io_SPI_invert; // @[Filter.scala 225:36]
  wire  _T_677 = $signed(pixOut_2_2) > 9'shf; // @[Filter.scala 230:36]
  wire  _T_678 = _T_677 & io_SPI_invert; // @[Filter.scala 230:43]
  wire [8:0] _T_682 = 9'hf - pixOut_2_2; // @[Filter.scala 235:43]
  wire [8:0] _GEN_10883 = io_SPI_invert ? _T_682 : pixOut_2_2; // @[Filter.scala 234:36]
  wire [8:0] _GEN_10884 = _T_677 ? 9'hf : _GEN_10883; // @[Filter.scala 232:44]
  wire [8:0] _GEN_10885 = _T_678 ? 9'h0 : _GEN_10884; // @[Filter.scala 230:59]
  wire [8:0] _GEN_10886 = _T_674 ? 9'h0 : _GEN_10885; // @[Filter.scala 227:43]
  wire [8:0] _GEN_10887 = _T_675 ? 9'hf : _GEN_10886; // @[Filter.scala 225:52]
  wire [9:0] _T_684 = $signed(KernelConvolution_2_io_pixelVal_out_3) / $signed(_GEN_11294); // @[Filter.scala 223:64]
  wire  _T_685 = $signed(pixOut_2_3) < 9'sh0; // @[Filter.scala 225:30]
  wire  _T_686 = _T_685 & io_SPI_invert; // @[Filter.scala 225:36]
  wire  _T_688 = $signed(pixOut_2_3) > 9'shf; // @[Filter.scala 230:36]
  wire  _T_689 = _T_688 & io_SPI_invert; // @[Filter.scala 230:43]
  wire [8:0] _T_693 = 9'hf - pixOut_2_3; // @[Filter.scala 235:43]
  wire [8:0] _GEN_10888 = io_SPI_invert ? _T_693 : pixOut_2_3; // @[Filter.scala 234:36]
  wire [8:0] _GEN_10889 = _T_688 ? 9'hf : _GEN_10888; // @[Filter.scala 232:44]
  wire [8:0] _GEN_10890 = _T_689 ? 9'h0 : _GEN_10889; // @[Filter.scala 230:59]
  wire [8:0] _GEN_10891 = _T_685 ? 9'h0 : _GEN_10890; // @[Filter.scala 227:43]
  wire [8:0] _GEN_10892 = _T_686 ? 9'hf : _GEN_10891; // @[Filter.scala 225:52]
  wire [9:0] _T_695 = $signed(KernelConvolution_2_io_pixelVal_out_4) / $signed(_GEN_11294); // @[Filter.scala 223:64]
  wire  _T_696 = $signed(pixOut_2_4) < 9'sh0; // @[Filter.scala 225:30]
  wire  _T_697 = _T_696 & io_SPI_invert; // @[Filter.scala 225:36]
  wire  _T_699 = $signed(pixOut_2_4) > 9'shf; // @[Filter.scala 230:36]
  wire  _T_700 = _T_699 & io_SPI_invert; // @[Filter.scala 230:43]
  wire [8:0] _T_704 = 9'hf - pixOut_2_4; // @[Filter.scala 235:43]
  wire [8:0] _GEN_10893 = io_SPI_invert ? _T_704 : pixOut_2_4; // @[Filter.scala 234:36]
  wire [8:0] _GEN_10894 = _T_699 ? 9'hf : _GEN_10893; // @[Filter.scala 232:44]
  wire [8:0] _GEN_10895 = _T_700 ? 9'h0 : _GEN_10894; // @[Filter.scala 230:59]
  wire [8:0] _GEN_10896 = _T_696 ? 9'h0 : _GEN_10895; // @[Filter.scala 227:43]
  wire [8:0] _GEN_10897 = _T_697 ? 9'hf : _GEN_10896; // @[Filter.scala 225:52]
  wire [9:0] _T_706 = $signed(KernelConvolution_2_io_pixelVal_out_5) / $signed(_GEN_11294); // @[Filter.scala 223:64]
  wire  _T_707 = $signed(pixOut_2_5) < 9'sh0; // @[Filter.scala 225:30]
  wire  _T_708 = _T_707 & io_SPI_invert; // @[Filter.scala 225:36]
  wire  _T_710 = $signed(pixOut_2_5) > 9'shf; // @[Filter.scala 230:36]
  wire  _T_711 = _T_710 & io_SPI_invert; // @[Filter.scala 230:43]
  wire [8:0] _T_715 = 9'hf - pixOut_2_5; // @[Filter.scala 235:43]
  wire [8:0] _GEN_10898 = io_SPI_invert ? _T_715 : pixOut_2_5; // @[Filter.scala 234:36]
  wire [8:0] _GEN_10899 = _T_710 ? 9'hf : _GEN_10898; // @[Filter.scala 232:44]
  wire [8:0] _GEN_10900 = _T_711 ? 9'h0 : _GEN_10899; // @[Filter.scala 230:59]
  wire [8:0] _GEN_10901 = _T_707 ? 9'h0 : _GEN_10900; // @[Filter.scala 227:43]
  wire [8:0] _GEN_10902 = _T_708 ? 9'hf : _GEN_10901; // @[Filter.scala 225:52]
  wire [9:0] _T_717 = $signed(KernelConvolution_2_io_pixelVal_out_6) / $signed(_GEN_11294); // @[Filter.scala 223:64]
  wire  _T_718 = $signed(pixOut_2_6) < 9'sh0; // @[Filter.scala 225:30]
  wire  _T_719 = _T_718 & io_SPI_invert; // @[Filter.scala 225:36]
  wire  _T_721 = $signed(pixOut_2_6) > 9'shf; // @[Filter.scala 230:36]
  wire  _T_722 = _T_721 & io_SPI_invert; // @[Filter.scala 230:43]
  wire [8:0] _T_726 = 9'hf - pixOut_2_6; // @[Filter.scala 235:43]
  wire [8:0] _GEN_10903 = io_SPI_invert ? _T_726 : pixOut_2_6; // @[Filter.scala 234:36]
  wire [8:0] _GEN_10904 = _T_721 ? 9'hf : _GEN_10903; // @[Filter.scala 232:44]
  wire [8:0] _GEN_10905 = _T_722 ? 9'h0 : _GEN_10904; // @[Filter.scala 230:59]
  wire [8:0] _GEN_10906 = _T_718 ? 9'h0 : _GEN_10905; // @[Filter.scala 227:43]
  wire [8:0] _GEN_10907 = _T_719 ? 9'hf : _GEN_10906; // @[Filter.scala 225:52]
  wire [31:0] _T_729 = pixelIndex + 32'h7; // @[Filter.scala 247:34]
  wire [8:0] _T_730 = 5'h15 * 5'hc; // @[Filter.scala 248:42]
  wire [31:0] _GEN_11315 = {{23'd0}, _T_730}; // @[Filter.scala 248:25]
  wire  _T_731 = pixelIndex == _GEN_11315; // @[Filter.scala 248:25]
  KernelConvolution KernelConvolution ( // @[Filter.scala 186:36]
    .clock(KernelConvolution_clock),
    .reset(KernelConvolution_reset),
    .io_kernelVal_in(KernelConvolution_io_kernelVal_in),
    .io_pixelVal_in_0(KernelConvolution_io_pixelVal_in_0),
    .io_pixelVal_in_1(KernelConvolution_io_pixelVal_in_1),
    .io_pixelVal_in_2(KernelConvolution_io_pixelVal_in_2),
    .io_pixelVal_in_3(KernelConvolution_io_pixelVal_in_3),
    .io_pixelVal_in_4(KernelConvolution_io_pixelVal_in_4),
    .io_pixelVal_in_5(KernelConvolution_io_pixelVal_in_5),
    .io_pixelVal_in_6(KernelConvolution_io_pixelVal_in_6),
    .io_pixelVal_out_0(KernelConvolution_io_pixelVal_out_0),
    .io_pixelVal_out_1(KernelConvolution_io_pixelVal_out_1),
    .io_pixelVal_out_2(KernelConvolution_io_pixelVal_out_2),
    .io_pixelVal_out_3(KernelConvolution_io_pixelVal_out_3),
    .io_pixelVal_out_4(KernelConvolution_io_pixelVal_out_4),
    .io_pixelVal_out_5(KernelConvolution_io_pixelVal_out_5),
    .io_pixelVal_out_6(KernelConvolution_io_pixelVal_out_6),
    .io_valid_out(KernelConvolution_io_valid_out)
  );
  KernelConvolution KernelConvolution_1 ( // @[Filter.scala 187:36]
    .clock(KernelConvolution_1_clock),
    .reset(KernelConvolution_1_reset),
    .io_kernelVal_in(KernelConvolution_1_io_kernelVal_in),
    .io_pixelVal_in_0(KernelConvolution_1_io_pixelVal_in_0),
    .io_pixelVal_in_1(KernelConvolution_1_io_pixelVal_in_1),
    .io_pixelVal_in_2(KernelConvolution_1_io_pixelVal_in_2),
    .io_pixelVal_in_3(KernelConvolution_1_io_pixelVal_in_3),
    .io_pixelVal_in_4(KernelConvolution_1_io_pixelVal_in_4),
    .io_pixelVal_in_5(KernelConvolution_1_io_pixelVal_in_5),
    .io_pixelVal_in_6(KernelConvolution_1_io_pixelVal_in_6),
    .io_pixelVal_out_0(KernelConvolution_1_io_pixelVal_out_0),
    .io_pixelVal_out_1(KernelConvolution_1_io_pixelVal_out_1),
    .io_pixelVal_out_2(KernelConvolution_1_io_pixelVal_out_2),
    .io_pixelVal_out_3(KernelConvolution_1_io_pixelVal_out_3),
    .io_pixelVal_out_4(KernelConvolution_1_io_pixelVal_out_4),
    .io_pixelVal_out_5(KernelConvolution_1_io_pixelVal_out_5),
    .io_pixelVal_out_6(KernelConvolution_1_io_pixelVal_out_6),
    .io_valid_out(KernelConvolution_1_io_valid_out)
  );
  KernelConvolution KernelConvolution_2 ( // @[Filter.scala 188:36]
    .clock(KernelConvolution_2_clock),
    .reset(KernelConvolution_2_reset),
    .io_kernelVal_in(KernelConvolution_2_io_kernelVal_in),
    .io_pixelVal_in_0(KernelConvolution_2_io_pixelVal_in_0),
    .io_pixelVal_in_1(KernelConvolution_2_io_pixelVal_in_1),
    .io_pixelVal_in_2(KernelConvolution_2_io_pixelVal_in_2),
    .io_pixelVal_in_3(KernelConvolution_2_io_pixelVal_in_3),
    .io_pixelVal_in_4(KernelConvolution_2_io_pixelVal_in_4),
    .io_pixelVal_in_5(KernelConvolution_2_io_pixelVal_in_5),
    .io_pixelVal_in_6(KernelConvolution_2_io_pixelVal_in_6),
    .io_pixelVal_out_0(KernelConvolution_2_io_pixelVal_out_0),
    .io_pixelVal_out_1(KernelConvolution_2_io_pixelVal_out_1),
    .io_pixelVal_out_2(KernelConvolution_2_io_pixelVal_out_2),
    .io_pixelVal_out_3(KernelConvolution_2_io_pixelVal_out_3),
    .io_pixelVal_out_4(KernelConvolution_2_io_pixelVal_out_4),
    .io_pixelVal_out_5(KernelConvolution_2_io_pixelVal_out_5),
    .io_pixelVal_out_6(KernelConvolution_2_io_pixelVal_out_6),
    .io_valid_out(KernelConvolution_2_io_valid_out)
  );
  assign io_pixelVal_out_0_0 = _GEN_10807[3:0]; // @[Filter.scala 226:35 Filter.scala 228:37 Filter.scala 231:35 Filter.scala 233:35 Filter.scala 235:35 Filter.scala 237:35]
  assign io_pixelVal_out_0_1 = _GEN_10812[3:0]; // @[Filter.scala 226:35 Filter.scala 228:37 Filter.scala 231:35 Filter.scala 233:35 Filter.scala 235:35 Filter.scala 237:35]
  assign io_pixelVal_out_0_2 = _GEN_10817[3:0]; // @[Filter.scala 226:35 Filter.scala 228:37 Filter.scala 231:35 Filter.scala 233:35 Filter.scala 235:35 Filter.scala 237:35]
  assign io_pixelVal_out_0_3 = _GEN_10822[3:0]; // @[Filter.scala 226:35 Filter.scala 228:37 Filter.scala 231:35 Filter.scala 233:35 Filter.scala 235:35 Filter.scala 237:35]
  assign io_pixelVal_out_0_4 = _GEN_10827[3:0]; // @[Filter.scala 226:35 Filter.scala 228:37 Filter.scala 231:35 Filter.scala 233:35 Filter.scala 235:35 Filter.scala 237:35]
  assign io_pixelVal_out_0_5 = _GEN_10832[3:0]; // @[Filter.scala 226:35 Filter.scala 228:37 Filter.scala 231:35 Filter.scala 233:35 Filter.scala 235:35 Filter.scala 237:35]
  assign io_pixelVal_out_0_6 = _GEN_10837[3:0]; // @[Filter.scala 226:35 Filter.scala 228:37 Filter.scala 231:35 Filter.scala 233:35 Filter.scala 235:35 Filter.scala 237:35]
  assign io_pixelVal_out_1_0 = _GEN_10842[3:0]; // @[Filter.scala 226:35 Filter.scala 228:37 Filter.scala 231:35 Filter.scala 233:35 Filter.scala 235:35 Filter.scala 237:35]
  assign io_pixelVal_out_1_1 = _GEN_10847[3:0]; // @[Filter.scala 226:35 Filter.scala 228:37 Filter.scala 231:35 Filter.scala 233:35 Filter.scala 235:35 Filter.scala 237:35]
  assign io_pixelVal_out_1_2 = _GEN_10852[3:0]; // @[Filter.scala 226:35 Filter.scala 228:37 Filter.scala 231:35 Filter.scala 233:35 Filter.scala 235:35 Filter.scala 237:35]
  assign io_pixelVal_out_1_3 = _GEN_10857[3:0]; // @[Filter.scala 226:35 Filter.scala 228:37 Filter.scala 231:35 Filter.scala 233:35 Filter.scala 235:35 Filter.scala 237:35]
  assign io_pixelVal_out_1_4 = _GEN_10862[3:0]; // @[Filter.scala 226:35 Filter.scala 228:37 Filter.scala 231:35 Filter.scala 233:35 Filter.scala 235:35 Filter.scala 237:35]
  assign io_pixelVal_out_1_5 = _GEN_10867[3:0]; // @[Filter.scala 226:35 Filter.scala 228:37 Filter.scala 231:35 Filter.scala 233:35 Filter.scala 235:35 Filter.scala 237:35]
  assign io_pixelVal_out_1_6 = _GEN_10872[3:0]; // @[Filter.scala 226:35 Filter.scala 228:37 Filter.scala 231:35 Filter.scala 233:35 Filter.scala 235:35 Filter.scala 237:35]
  assign io_pixelVal_out_2_0 = _GEN_10877[3:0]; // @[Filter.scala 226:35 Filter.scala 228:37 Filter.scala 231:35 Filter.scala 233:35 Filter.scala 235:35 Filter.scala 237:35]
  assign io_pixelVal_out_2_1 = _GEN_10882[3:0]; // @[Filter.scala 226:35 Filter.scala 228:37 Filter.scala 231:35 Filter.scala 233:35 Filter.scala 235:35 Filter.scala 237:35]
  assign io_pixelVal_out_2_2 = _GEN_10887[3:0]; // @[Filter.scala 226:35 Filter.scala 228:37 Filter.scala 231:35 Filter.scala 233:35 Filter.scala 235:35 Filter.scala 237:35]
  assign io_pixelVal_out_2_3 = _GEN_10892[3:0]; // @[Filter.scala 226:35 Filter.scala 228:37 Filter.scala 231:35 Filter.scala 233:35 Filter.scala 235:35 Filter.scala 237:35]
  assign io_pixelVal_out_2_4 = _GEN_10897[3:0]; // @[Filter.scala 226:35 Filter.scala 228:37 Filter.scala 231:35 Filter.scala 233:35 Filter.scala 235:35 Filter.scala 237:35]
  assign io_pixelVal_out_2_5 = _GEN_10902[3:0]; // @[Filter.scala 226:35 Filter.scala 228:37 Filter.scala 231:35 Filter.scala 233:35 Filter.scala 235:35 Filter.scala 237:35]
  assign io_pixelVal_out_2_6 = _GEN_10907[3:0]; // @[Filter.scala 226:35 Filter.scala 228:37 Filter.scala 231:35 Filter.scala 233:35 Filter.scala 235:35 Filter.scala 237:35]
  assign io_valid_out = validOut; // @[Filter.scala 244:18]
  assign KernelConvolution_clock = clock;
  assign KernelConvolution_reset = reset;
  assign KernelConvolution_io_kernelVal_in = _GEN_10992 & _GEN_10919 ? $signed(5'sh0) : $signed(_GEN_55); // @[Filter.scala 194:41]
  assign KernelConvolution_io_pixelVal_in_0 = _GEN_1180[3:0]; // @[Filter.scala 208:53 Filter.scala 210:51 Filter.scala 212:51]
  assign KernelConvolution_io_pixelVal_in_1 = _GEN_2698[3:0]; // @[Filter.scala 208:53 Filter.scala 210:51 Filter.scala 212:51]
  assign KernelConvolution_io_pixelVal_in_2 = _GEN_4216[3:0]; // @[Filter.scala 208:53 Filter.scala 210:51 Filter.scala 212:51]
  assign KernelConvolution_io_pixelVal_in_3 = _GEN_5734[3:0]; // @[Filter.scala 208:53 Filter.scala 210:51 Filter.scala 212:51]
  assign KernelConvolution_io_pixelVal_in_4 = _GEN_7252[3:0]; // @[Filter.scala 208:53 Filter.scala 210:51 Filter.scala 212:51]
  assign KernelConvolution_io_pixelVal_in_5 = _GEN_8770[3:0]; // @[Filter.scala 208:53 Filter.scala 210:51 Filter.scala 212:51]
  assign KernelConvolution_io_pixelVal_in_6 = _GEN_10288[3:0]; // @[Filter.scala 208:53 Filter.scala 210:51 Filter.scala 212:51]
  assign KernelConvolution_1_clock = clock;
  assign KernelConvolution_1_reset = reset;
  assign KernelConvolution_1_io_kernelVal_in = _GEN_10992 & _GEN_10919 ? $signed(5'sh0) : $signed(_GEN_55); // @[Filter.scala 194:41]
  assign KernelConvolution_1_io_pixelVal_in_0 = _GEN_1434[3:0]; // @[Filter.scala 208:53 Filter.scala 210:51 Filter.scala 212:51]
  assign KernelConvolution_1_io_pixelVal_in_1 = _GEN_2952[3:0]; // @[Filter.scala 208:53 Filter.scala 210:51 Filter.scala 212:51]
  assign KernelConvolution_1_io_pixelVal_in_2 = _GEN_4470[3:0]; // @[Filter.scala 208:53 Filter.scala 210:51 Filter.scala 212:51]
  assign KernelConvolution_1_io_pixelVal_in_3 = _GEN_5988[3:0]; // @[Filter.scala 208:53 Filter.scala 210:51 Filter.scala 212:51]
  assign KernelConvolution_1_io_pixelVal_in_4 = _GEN_7506[3:0]; // @[Filter.scala 208:53 Filter.scala 210:51 Filter.scala 212:51]
  assign KernelConvolution_1_io_pixelVal_in_5 = _GEN_9024[3:0]; // @[Filter.scala 208:53 Filter.scala 210:51 Filter.scala 212:51]
  assign KernelConvolution_1_io_pixelVal_in_6 = _GEN_10542[3:0]; // @[Filter.scala 208:53 Filter.scala 210:51 Filter.scala 212:51]
  assign KernelConvolution_2_clock = clock;
  assign KernelConvolution_2_reset = reset;
  assign KernelConvolution_2_io_kernelVal_in = _GEN_10992 & _GEN_10919 ? $signed(5'sh0) : $signed(_GEN_55); // @[Filter.scala 194:41]
  assign KernelConvolution_2_io_pixelVal_in_0 = _GEN_1688[3:0]; // @[Filter.scala 208:53 Filter.scala 210:51 Filter.scala 212:51]
  assign KernelConvolution_2_io_pixelVal_in_1 = _GEN_3206[3:0]; // @[Filter.scala 208:53 Filter.scala 210:51 Filter.scala 212:51]
  assign KernelConvolution_2_io_pixelVal_in_2 = _GEN_4724[3:0]; // @[Filter.scala 208:53 Filter.scala 210:51 Filter.scala 212:51]
  assign KernelConvolution_2_io_pixelVal_in_3 = _GEN_6242[3:0]; // @[Filter.scala 208:53 Filter.scala 210:51 Filter.scala 212:51]
  assign KernelConvolution_2_io_pixelVal_in_4 = _GEN_7760[3:0]; // @[Filter.scala 208:53 Filter.scala 210:51 Filter.scala 212:51]
  assign KernelConvolution_2_io_pixelVal_in_5 = _GEN_9278[3:0]; // @[Filter.scala 208:53 Filter.scala 210:51 Filter.scala 212:51]
  assign KernelConvolution_2_io_pixelVal_in_6 = _GEN_10796[3:0]; // @[Filter.scala 208:53 Filter.scala 210:51 Filter.scala 212:51]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  kernelCounter = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  imageCounterX = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  imageCounterY = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  pixelIndex = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  pixOut_0_0 = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  pixOut_0_1 = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  pixOut_0_2 = _RAND_6[8:0];
  _RAND_7 = {1{`RANDOM}};
  pixOut_0_3 = _RAND_7[8:0];
  _RAND_8 = {1{`RANDOM}};
  pixOut_0_4 = _RAND_8[8:0];
  _RAND_9 = {1{`RANDOM}};
  pixOut_0_5 = _RAND_9[8:0];
  _RAND_10 = {1{`RANDOM}};
  pixOut_0_6 = _RAND_10[8:0];
  _RAND_11 = {1{`RANDOM}};
  pixOut_1_0 = _RAND_11[8:0];
  _RAND_12 = {1{`RANDOM}};
  pixOut_1_1 = _RAND_12[8:0];
  _RAND_13 = {1{`RANDOM}};
  pixOut_1_2 = _RAND_13[8:0];
  _RAND_14 = {1{`RANDOM}};
  pixOut_1_3 = _RAND_14[8:0];
  _RAND_15 = {1{`RANDOM}};
  pixOut_1_4 = _RAND_15[8:0];
  _RAND_16 = {1{`RANDOM}};
  pixOut_1_5 = _RAND_16[8:0];
  _RAND_17 = {1{`RANDOM}};
  pixOut_1_6 = _RAND_17[8:0];
  _RAND_18 = {1{`RANDOM}};
  pixOut_2_0 = _RAND_18[8:0];
  _RAND_19 = {1{`RANDOM}};
  pixOut_2_1 = _RAND_19[8:0];
  _RAND_20 = {1{`RANDOM}};
  pixOut_2_2 = _RAND_20[8:0];
  _RAND_21 = {1{`RANDOM}};
  pixOut_2_3 = _RAND_21[8:0];
  _RAND_22 = {1{`RANDOM}};
  pixOut_2_4 = _RAND_22[8:0];
  _RAND_23 = {1{`RANDOM}};
  pixOut_2_5 = _RAND_23[8:0];
  _RAND_24 = {1{`RANDOM}};
  pixOut_2_6 = _RAND_24[8:0];
  _RAND_25 = {1{`RANDOM}};
  validOut = _RAND_25[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      kernelCounter <= 4'h0;
    end else if (kernelCountReset) begin
      kernelCounter <= 4'h0;
    end else begin
      kernelCounter <= _T_14;
    end
    if (reset) begin
      imageCounterX <= 2'h0;
    end else if (imageCounterXReset) begin
      imageCounterX <= 2'h0;
    end else begin
      imageCounterX <= _T_20;
    end
    if (reset) begin
      imageCounterY <= 2'h0;
    end else if (imageCounterXReset) begin
      if (_T_21) begin
        imageCounterY <= 2'h0;
      end else begin
        imageCounterY <= _T_23;
      end
    end
    if (reset) begin
      pixelIndex <= 32'h0;
    end else if (kernelCountReset) begin
      if (_T_731) begin
        pixelIndex <= 32'h0;
      end else begin
        pixelIndex <= _T_729;
      end
    end
    if (reset) begin
      pixOut_0_0 <= 9'sh0;
    end else begin
      pixOut_0_0 <= _T_497[8:0];
    end
    if (reset) begin
      pixOut_0_1 <= 9'sh0;
    end else begin
      pixOut_0_1 <= _T_508[8:0];
    end
    if (reset) begin
      pixOut_0_2 <= 9'sh0;
    end else begin
      pixOut_0_2 <= _T_519[8:0];
    end
    if (reset) begin
      pixOut_0_3 <= 9'sh0;
    end else begin
      pixOut_0_3 <= _T_530[8:0];
    end
    if (reset) begin
      pixOut_0_4 <= 9'sh0;
    end else begin
      pixOut_0_4 <= _T_541[8:0];
    end
    if (reset) begin
      pixOut_0_5 <= 9'sh0;
    end else begin
      pixOut_0_5 <= _T_552[8:0];
    end
    if (reset) begin
      pixOut_0_6 <= 9'sh0;
    end else begin
      pixOut_0_6 <= _T_563[8:0];
    end
    if (reset) begin
      pixOut_1_0 <= 9'sh0;
    end else begin
      pixOut_1_0 <= _T_574[8:0];
    end
    if (reset) begin
      pixOut_1_1 <= 9'sh0;
    end else begin
      pixOut_1_1 <= _T_585[8:0];
    end
    if (reset) begin
      pixOut_1_2 <= 9'sh0;
    end else begin
      pixOut_1_2 <= _T_596[8:0];
    end
    if (reset) begin
      pixOut_1_3 <= 9'sh0;
    end else begin
      pixOut_1_3 <= _T_607[8:0];
    end
    if (reset) begin
      pixOut_1_4 <= 9'sh0;
    end else begin
      pixOut_1_4 <= _T_618[8:0];
    end
    if (reset) begin
      pixOut_1_5 <= 9'sh0;
    end else begin
      pixOut_1_5 <= _T_629[8:0];
    end
    if (reset) begin
      pixOut_1_6 <= 9'sh0;
    end else begin
      pixOut_1_6 <= _T_640[8:0];
    end
    if (reset) begin
      pixOut_2_0 <= 9'sh0;
    end else begin
      pixOut_2_0 <= _T_651[8:0];
    end
    if (reset) begin
      pixOut_2_1 <= 9'sh0;
    end else begin
      pixOut_2_1 <= _T_662[8:0];
    end
    if (reset) begin
      pixOut_2_2 <= 9'sh0;
    end else begin
      pixOut_2_2 <= _T_673[8:0];
    end
    if (reset) begin
      pixOut_2_3 <= 9'sh0;
    end else begin
      pixOut_2_3 <= _T_684[8:0];
    end
    if (reset) begin
      pixOut_2_4 <= 9'sh0;
    end else begin
      pixOut_2_4 <= _T_695[8:0];
    end
    if (reset) begin
      pixOut_2_5 <= 9'sh0;
    end else begin
      pixOut_2_5 <= _T_706[8:0];
    end
    if (reset) begin
      pixOut_2_6 <= 9'sh0;
    end else begin
      pixOut_2_6 <= _T_717[8:0];
    end
    if (reset) begin
      validOut <= 1'h0;
    end else begin
      validOut <= KernelConvolution_io_valid_out;
    end
  end
endmodule
module VideoBuffer(
  input         clock,
  input         reset,
  input  [3:0]  io_pixelVal_in_0_0,
  input  [3:0]  io_pixelVal_in_0_1,
  input  [3:0]  io_pixelVal_in_0_2,
  input  [3:0]  io_pixelVal_in_0_3,
  input  [3:0]  io_pixelVal_in_0_4,
  input  [3:0]  io_pixelVal_in_0_5,
  input  [3:0]  io_pixelVal_in_0_6,
  input  [3:0]  io_pixelVal_in_1_0,
  input  [3:0]  io_pixelVal_in_1_1,
  input  [3:0]  io_pixelVal_in_1_2,
  input  [3:0]  io_pixelVal_in_1_3,
  input  [3:0]  io_pixelVal_in_1_4,
  input  [3:0]  io_pixelVal_in_1_5,
  input  [3:0]  io_pixelVal_in_1_6,
  input  [3:0]  io_pixelVal_in_2_0,
  input  [3:0]  io_pixelVal_in_2_1,
  input  [3:0]  io_pixelVal_in_2_2,
  input  [3:0]  io_pixelVal_in_2_3,
  input  [3:0]  io_pixelVal_in_2_4,
  input  [3:0]  io_pixelVal_in_2_5,
  input  [3:0]  io_pixelVal_in_2_6,
  input         io_valid_in,
  input  [10:0] io_rowIndex,
  input  [10:0] io_colIndex,
  output [3:0]  io_pixelVal_out_0,
  output [3:0]  io_pixelVal_out_1,
  output [3:0]  io_pixelVal_out_2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] image_0_0; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_1; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_2; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_3; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_4; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_5; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_6; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_7; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_8; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_9; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_10; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_11; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_12; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_13; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_14; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_15; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_16; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_17; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_18; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_19; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_20; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_21; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_22; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_23; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_24; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_25; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_26; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_27; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_28; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_29; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_30; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_31; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_32; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_33; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_34; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_35; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_36; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_37; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_38; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_39; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_40; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_41; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_42; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_43; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_44; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_45; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_46; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_47; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_48; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_49; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_50; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_51; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_52; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_53; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_54; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_55; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_56; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_57; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_58; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_59; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_60; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_61; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_62; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_63; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_64; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_65; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_66; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_67; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_68; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_69; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_70; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_71; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_72; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_73; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_74; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_75; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_76; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_77; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_78; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_79; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_80; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_81; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_82; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_83; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_84; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_85; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_86; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_87; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_88; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_89; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_90; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_91; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_92; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_93; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_94; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_95; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_96; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_97; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_98; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_99; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_100; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_101; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_102; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_103; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_104; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_105; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_106; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_107; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_108; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_109; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_110; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_111; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_112; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_113; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_114; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_115; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_116; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_117; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_118; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_119; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_120; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_121; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_122; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_123; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_124; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_125; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_126; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_127; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_128; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_129; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_130; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_131; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_132; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_133; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_134; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_135; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_136; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_137; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_138; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_139; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_140; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_141; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_142; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_143; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_144; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_145; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_146; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_147; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_148; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_149; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_150; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_151; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_152; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_153; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_154; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_155; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_156; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_157; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_158; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_159; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_160; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_161; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_162; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_163; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_164; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_165; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_166; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_167; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_168; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_169; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_170; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_171; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_172; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_173; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_174; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_175; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_176; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_177; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_178; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_179; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_180; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_181; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_182; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_183; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_184; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_185; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_186; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_187; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_188; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_189; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_190; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_191; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_192; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_193; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_194; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_195; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_196; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_197; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_198; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_199; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_200; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_201; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_202; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_203; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_204; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_205; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_206; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_207; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_208; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_209; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_210; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_211; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_212; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_213; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_214; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_215; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_216; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_217; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_218; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_219; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_220; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_221; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_222; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_223; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_224; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_225; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_226; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_227; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_228; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_229; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_230; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_231; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_232; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_233; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_234; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_235; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_236; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_237; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_238; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_239; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_240; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_241; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_242; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_243; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_244; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_245; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_246; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_247; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_248; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_249; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_250; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_251; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_1_0; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_1; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_2; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_3; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_4; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_5; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_6; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_7; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_8; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_9; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_10; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_11; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_12; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_13; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_14; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_15; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_16; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_17; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_18; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_19; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_20; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_21; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_22; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_23; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_24; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_25; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_26; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_27; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_28; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_29; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_30; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_31; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_32; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_33; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_34; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_35; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_36; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_37; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_38; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_39; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_40; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_41; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_42; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_43; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_44; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_45; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_46; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_47; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_48; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_49; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_50; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_51; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_52; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_53; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_54; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_55; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_56; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_57; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_58; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_59; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_60; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_61; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_62; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_63; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_64; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_65; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_66; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_67; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_68; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_69; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_70; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_71; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_72; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_73; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_74; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_75; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_76; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_77; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_78; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_79; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_80; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_81; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_82; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_83; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_84; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_85; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_86; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_87; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_88; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_89; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_90; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_91; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_92; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_93; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_94; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_95; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_96; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_97; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_98; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_99; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_100; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_101; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_102; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_103; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_104; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_105; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_106; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_107; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_108; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_109; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_110; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_111; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_112; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_113; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_114; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_115; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_116; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_117; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_118; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_119; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_120; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_121; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_122; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_123; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_124; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_125; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_126; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_127; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_128; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_129; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_130; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_131; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_132; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_133; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_134; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_135; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_136; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_137; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_138; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_139; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_140; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_141; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_142; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_143; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_144; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_145; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_146; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_147; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_148; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_149; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_150; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_151; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_152; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_153; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_154; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_155; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_156; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_157; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_158; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_159; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_160; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_161; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_162; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_163; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_164; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_165; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_166; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_167; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_168; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_169; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_170; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_171; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_172; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_173; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_174; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_175; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_176; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_177; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_178; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_179; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_180; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_181; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_182; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_183; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_184; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_185; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_186; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_187; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_188; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_189; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_190; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_191; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_192; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_193; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_194; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_195; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_196; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_197; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_198; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_199; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_200; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_201; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_202; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_203; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_204; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_205; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_206; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_207; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_208; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_209; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_210; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_211; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_212; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_213; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_214; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_215; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_216; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_217; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_218; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_219; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_220; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_221; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_222; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_223; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_224; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_225; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_226; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_227; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_228; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_229; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_230; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_231; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_232; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_233; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_234; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_235; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_236; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_237; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_238; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_239; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_240; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_241; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_242; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_243; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_244; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_245; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_246; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_247; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_248; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_249; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_250; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_251; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_2_0; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_1; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_2; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_3; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_4; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_5; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_6; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_7; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_8; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_9; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_10; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_11; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_12; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_13; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_14; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_15; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_16; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_17; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_18; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_19; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_20; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_21; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_22; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_23; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_24; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_25; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_26; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_27; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_28; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_29; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_30; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_31; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_32; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_33; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_34; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_35; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_36; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_37; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_38; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_39; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_40; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_41; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_42; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_43; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_44; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_45; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_46; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_47; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_48; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_49; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_50; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_51; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_52; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_53; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_54; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_55; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_56; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_57; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_58; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_59; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_60; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_61; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_62; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_63; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_64; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_65; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_66; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_67; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_68; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_69; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_70; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_71; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_72; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_73; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_74; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_75; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_76; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_77; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_78; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_79; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_80; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_81; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_82; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_83; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_84; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_85; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_86; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_87; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_88; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_89; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_90; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_91; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_92; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_93; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_94; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_95; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_96; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_97; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_98; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_99; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_100; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_101; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_102; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_103; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_104; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_105; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_106; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_107; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_108; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_109; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_110; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_111; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_112; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_113; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_114; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_115; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_116; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_117; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_118; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_119; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_120; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_121; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_122; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_123; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_124; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_125; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_126; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_127; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_128; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_129; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_130; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_131; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_132; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_133; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_134; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_135; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_136; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_137; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_138; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_139; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_140; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_141; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_142; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_143; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_144; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_145; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_146; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_147; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_148; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_149; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_150; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_151; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_152; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_153; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_154; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_155; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_156; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_157; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_158; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_159; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_160; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_161; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_162; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_163; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_164; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_165; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_166; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_167; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_168; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_169; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_170; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_171; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_172; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_173; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_174; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_175; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_176; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_177; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_178; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_179; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_180; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_181; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_182; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_183; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_184; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_185; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_186; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_187; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_188; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_189; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_190; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_191; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_192; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_193; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_194; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_195; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_196; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_197; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_198; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_199; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_200; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_201; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_202; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_203; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_204; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_205; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_206; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_207; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_208; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_209; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_210; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_211; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_212; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_213; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_214; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_215; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_216; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_217; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_218; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_219; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_220; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_221; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_222; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_223; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_224; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_225; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_226; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_227; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_228; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_229; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_230; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_231; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_232; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_233; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_234; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_235; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_236; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_237; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_238; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_239; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_240; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_241; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_242; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_243; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_244; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_245; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_246; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_247; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_248; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_249; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_250; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_251; // @[VideoBuffer.scala 21:25]
  reg [31:0] pixelIndex; // @[VideoBuffer.scala 24:33]
  wire [15:0] _T_3 = io_rowIndex * 11'h15; // @[VideoBuffer.scala 27:54]
  wire [15:0] _GEN_6806 = {{5'd0}, io_colIndex}; // @[VideoBuffer.scala 27:69]
  wire [15:0] _T_5 = _T_3 + _GEN_6806; // @[VideoBuffer.scala 27:69]
  wire [3:0] _GEN_1 = 8'h1 == _T_5[7:0] ? image_0_1 : image_0_0; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2 = 8'h2 == _T_5[7:0] ? image_0_2 : _GEN_1; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3 = 8'h3 == _T_5[7:0] ? image_0_3 : _GEN_2; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4 = 8'h4 == _T_5[7:0] ? image_0_4 : _GEN_3; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_5 = 8'h5 == _T_5[7:0] ? image_0_5 : _GEN_4; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_6 = 8'h6 == _T_5[7:0] ? image_0_6 : _GEN_5; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_7 = 8'h7 == _T_5[7:0] ? image_0_7 : _GEN_6; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_8 = 8'h8 == _T_5[7:0] ? image_0_8 : _GEN_7; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_9 = 8'h9 == _T_5[7:0] ? image_0_9 : _GEN_8; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_10 = 8'ha == _T_5[7:0] ? image_0_10 : _GEN_9; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_11 = 8'hb == _T_5[7:0] ? image_0_11 : _GEN_10; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_12 = 8'hc == _T_5[7:0] ? image_0_12 : _GEN_11; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_13 = 8'hd == _T_5[7:0] ? image_0_13 : _GEN_12; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_14 = 8'he == _T_5[7:0] ? image_0_14 : _GEN_13; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_15 = 8'hf == _T_5[7:0] ? image_0_15 : _GEN_14; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_16 = 8'h10 == _T_5[7:0] ? image_0_16 : _GEN_15; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_17 = 8'h11 == _T_5[7:0] ? image_0_17 : _GEN_16; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_18 = 8'h12 == _T_5[7:0] ? image_0_18 : _GEN_17; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_19 = 8'h13 == _T_5[7:0] ? image_0_19 : _GEN_18; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_20 = 8'h14 == _T_5[7:0] ? image_0_20 : _GEN_19; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_21 = 8'h15 == _T_5[7:0] ? image_0_21 : _GEN_20; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_22 = 8'h16 == _T_5[7:0] ? image_0_22 : _GEN_21; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_23 = 8'h17 == _T_5[7:0] ? image_0_23 : _GEN_22; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_24 = 8'h18 == _T_5[7:0] ? image_0_24 : _GEN_23; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_25 = 8'h19 == _T_5[7:0] ? image_0_25 : _GEN_24; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_26 = 8'h1a == _T_5[7:0] ? image_0_26 : _GEN_25; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_27 = 8'h1b == _T_5[7:0] ? image_0_27 : _GEN_26; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_28 = 8'h1c == _T_5[7:0] ? image_0_28 : _GEN_27; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_29 = 8'h1d == _T_5[7:0] ? image_0_29 : _GEN_28; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_30 = 8'h1e == _T_5[7:0] ? image_0_30 : _GEN_29; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_31 = 8'h1f == _T_5[7:0] ? image_0_31 : _GEN_30; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_32 = 8'h20 == _T_5[7:0] ? image_0_32 : _GEN_31; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_33 = 8'h21 == _T_5[7:0] ? image_0_33 : _GEN_32; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_34 = 8'h22 == _T_5[7:0] ? image_0_34 : _GEN_33; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_35 = 8'h23 == _T_5[7:0] ? image_0_35 : _GEN_34; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_36 = 8'h24 == _T_5[7:0] ? image_0_36 : _GEN_35; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_37 = 8'h25 == _T_5[7:0] ? image_0_37 : _GEN_36; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_38 = 8'h26 == _T_5[7:0] ? image_0_38 : _GEN_37; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_39 = 8'h27 == _T_5[7:0] ? image_0_39 : _GEN_38; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_40 = 8'h28 == _T_5[7:0] ? image_0_40 : _GEN_39; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_41 = 8'h29 == _T_5[7:0] ? image_0_41 : _GEN_40; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_42 = 8'h2a == _T_5[7:0] ? image_0_42 : _GEN_41; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_43 = 8'h2b == _T_5[7:0] ? image_0_43 : _GEN_42; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_44 = 8'h2c == _T_5[7:0] ? image_0_44 : _GEN_43; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_45 = 8'h2d == _T_5[7:0] ? image_0_45 : _GEN_44; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_46 = 8'h2e == _T_5[7:0] ? image_0_46 : _GEN_45; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_47 = 8'h2f == _T_5[7:0] ? image_0_47 : _GEN_46; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_48 = 8'h30 == _T_5[7:0] ? image_0_48 : _GEN_47; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_49 = 8'h31 == _T_5[7:0] ? image_0_49 : _GEN_48; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_50 = 8'h32 == _T_5[7:0] ? image_0_50 : _GEN_49; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_51 = 8'h33 == _T_5[7:0] ? image_0_51 : _GEN_50; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_52 = 8'h34 == _T_5[7:0] ? image_0_52 : _GEN_51; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_53 = 8'h35 == _T_5[7:0] ? image_0_53 : _GEN_52; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_54 = 8'h36 == _T_5[7:0] ? image_0_54 : _GEN_53; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_55 = 8'h37 == _T_5[7:0] ? image_0_55 : _GEN_54; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_56 = 8'h38 == _T_5[7:0] ? image_0_56 : _GEN_55; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_57 = 8'h39 == _T_5[7:0] ? image_0_57 : _GEN_56; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_58 = 8'h3a == _T_5[7:0] ? image_0_58 : _GEN_57; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_59 = 8'h3b == _T_5[7:0] ? image_0_59 : _GEN_58; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_60 = 8'h3c == _T_5[7:0] ? image_0_60 : _GEN_59; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_61 = 8'h3d == _T_5[7:0] ? image_0_61 : _GEN_60; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_62 = 8'h3e == _T_5[7:0] ? image_0_62 : _GEN_61; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_63 = 8'h3f == _T_5[7:0] ? image_0_63 : _GEN_62; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_64 = 8'h40 == _T_5[7:0] ? image_0_64 : _GEN_63; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_65 = 8'h41 == _T_5[7:0] ? image_0_65 : _GEN_64; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_66 = 8'h42 == _T_5[7:0] ? image_0_66 : _GEN_65; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_67 = 8'h43 == _T_5[7:0] ? image_0_67 : _GEN_66; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_68 = 8'h44 == _T_5[7:0] ? image_0_68 : _GEN_67; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_69 = 8'h45 == _T_5[7:0] ? image_0_69 : _GEN_68; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_70 = 8'h46 == _T_5[7:0] ? image_0_70 : _GEN_69; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_71 = 8'h47 == _T_5[7:0] ? image_0_71 : _GEN_70; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_72 = 8'h48 == _T_5[7:0] ? image_0_72 : _GEN_71; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_73 = 8'h49 == _T_5[7:0] ? image_0_73 : _GEN_72; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_74 = 8'h4a == _T_5[7:0] ? image_0_74 : _GEN_73; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_75 = 8'h4b == _T_5[7:0] ? image_0_75 : _GEN_74; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_76 = 8'h4c == _T_5[7:0] ? image_0_76 : _GEN_75; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_77 = 8'h4d == _T_5[7:0] ? image_0_77 : _GEN_76; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_78 = 8'h4e == _T_5[7:0] ? image_0_78 : _GEN_77; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_79 = 8'h4f == _T_5[7:0] ? image_0_79 : _GEN_78; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_80 = 8'h50 == _T_5[7:0] ? image_0_80 : _GEN_79; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_81 = 8'h51 == _T_5[7:0] ? image_0_81 : _GEN_80; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_82 = 8'h52 == _T_5[7:0] ? image_0_82 : _GEN_81; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_83 = 8'h53 == _T_5[7:0] ? image_0_83 : _GEN_82; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_84 = 8'h54 == _T_5[7:0] ? image_0_84 : _GEN_83; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_85 = 8'h55 == _T_5[7:0] ? image_0_85 : _GEN_84; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_86 = 8'h56 == _T_5[7:0] ? image_0_86 : _GEN_85; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_87 = 8'h57 == _T_5[7:0] ? image_0_87 : _GEN_86; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_88 = 8'h58 == _T_5[7:0] ? image_0_88 : _GEN_87; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_89 = 8'h59 == _T_5[7:0] ? image_0_89 : _GEN_88; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_90 = 8'h5a == _T_5[7:0] ? image_0_90 : _GEN_89; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_91 = 8'h5b == _T_5[7:0] ? image_0_91 : _GEN_90; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_92 = 8'h5c == _T_5[7:0] ? image_0_92 : _GEN_91; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_93 = 8'h5d == _T_5[7:0] ? image_0_93 : _GEN_92; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_94 = 8'h5e == _T_5[7:0] ? image_0_94 : _GEN_93; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_95 = 8'h5f == _T_5[7:0] ? image_0_95 : _GEN_94; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_96 = 8'h60 == _T_5[7:0] ? image_0_96 : _GEN_95; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_97 = 8'h61 == _T_5[7:0] ? image_0_97 : _GEN_96; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_98 = 8'h62 == _T_5[7:0] ? image_0_98 : _GEN_97; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_99 = 8'h63 == _T_5[7:0] ? image_0_99 : _GEN_98; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_100 = 8'h64 == _T_5[7:0] ? image_0_100 : _GEN_99; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_101 = 8'h65 == _T_5[7:0] ? image_0_101 : _GEN_100; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_102 = 8'h66 == _T_5[7:0] ? image_0_102 : _GEN_101; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_103 = 8'h67 == _T_5[7:0] ? image_0_103 : _GEN_102; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_104 = 8'h68 == _T_5[7:0] ? image_0_104 : _GEN_103; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_105 = 8'h69 == _T_5[7:0] ? image_0_105 : _GEN_104; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_106 = 8'h6a == _T_5[7:0] ? image_0_106 : _GEN_105; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_107 = 8'h6b == _T_5[7:0] ? image_0_107 : _GEN_106; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_108 = 8'h6c == _T_5[7:0] ? image_0_108 : _GEN_107; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_109 = 8'h6d == _T_5[7:0] ? image_0_109 : _GEN_108; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_110 = 8'h6e == _T_5[7:0] ? image_0_110 : _GEN_109; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_111 = 8'h6f == _T_5[7:0] ? image_0_111 : _GEN_110; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_112 = 8'h70 == _T_5[7:0] ? image_0_112 : _GEN_111; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_113 = 8'h71 == _T_5[7:0] ? image_0_113 : _GEN_112; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_114 = 8'h72 == _T_5[7:0] ? image_0_114 : _GEN_113; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_115 = 8'h73 == _T_5[7:0] ? image_0_115 : _GEN_114; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_116 = 8'h74 == _T_5[7:0] ? image_0_116 : _GEN_115; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_117 = 8'h75 == _T_5[7:0] ? image_0_117 : _GEN_116; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_118 = 8'h76 == _T_5[7:0] ? image_0_118 : _GEN_117; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_119 = 8'h77 == _T_5[7:0] ? image_0_119 : _GEN_118; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_120 = 8'h78 == _T_5[7:0] ? image_0_120 : _GEN_119; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_121 = 8'h79 == _T_5[7:0] ? image_0_121 : _GEN_120; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_122 = 8'h7a == _T_5[7:0] ? image_0_122 : _GEN_121; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_123 = 8'h7b == _T_5[7:0] ? image_0_123 : _GEN_122; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_124 = 8'h7c == _T_5[7:0] ? image_0_124 : _GEN_123; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_125 = 8'h7d == _T_5[7:0] ? image_0_125 : _GEN_124; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_126 = 8'h7e == _T_5[7:0] ? image_0_126 : _GEN_125; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_127 = 8'h7f == _T_5[7:0] ? image_0_127 : _GEN_126; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_128 = 8'h80 == _T_5[7:0] ? image_0_128 : _GEN_127; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_129 = 8'h81 == _T_5[7:0] ? image_0_129 : _GEN_128; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_130 = 8'h82 == _T_5[7:0] ? image_0_130 : _GEN_129; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_131 = 8'h83 == _T_5[7:0] ? image_0_131 : _GEN_130; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_132 = 8'h84 == _T_5[7:0] ? image_0_132 : _GEN_131; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_133 = 8'h85 == _T_5[7:0] ? image_0_133 : _GEN_132; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_134 = 8'h86 == _T_5[7:0] ? image_0_134 : _GEN_133; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_135 = 8'h87 == _T_5[7:0] ? image_0_135 : _GEN_134; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_136 = 8'h88 == _T_5[7:0] ? image_0_136 : _GEN_135; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_137 = 8'h89 == _T_5[7:0] ? image_0_137 : _GEN_136; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_138 = 8'h8a == _T_5[7:0] ? image_0_138 : _GEN_137; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_139 = 8'h8b == _T_5[7:0] ? image_0_139 : _GEN_138; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_140 = 8'h8c == _T_5[7:0] ? image_0_140 : _GEN_139; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_141 = 8'h8d == _T_5[7:0] ? image_0_141 : _GEN_140; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_142 = 8'h8e == _T_5[7:0] ? image_0_142 : _GEN_141; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_143 = 8'h8f == _T_5[7:0] ? image_0_143 : _GEN_142; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_144 = 8'h90 == _T_5[7:0] ? image_0_144 : _GEN_143; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_145 = 8'h91 == _T_5[7:0] ? image_0_145 : _GEN_144; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_146 = 8'h92 == _T_5[7:0] ? image_0_146 : _GEN_145; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_147 = 8'h93 == _T_5[7:0] ? image_0_147 : _GEN_146; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_148 = 8'h94 == _T_5[7:0] ? image_0_148 : _GEN_147; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_149 = 8'h95 == _T_5[7:0] ? image_0_149 : _GEN_148; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_150 = 8'h96 == _T_5[7:0] ? image_0_150 : _GEN_149; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_151 = 8'h97 == _T_5[7:0] ? image_0_151 : _GEN_150; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_152 = 8'h98 == _T_5[7:0] ? image_0_152 : _GEN_151; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_153 = 8'h99 == _T_5[7:0] ? image_0_153 : _GEN_152; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_154 = 8'h9a == _T_5[7:0] ? image_0_154 : _GEN_153; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_155 = 8'h9b == _T_5[7:0] ? image_0_155 : _GEN_154; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_156 = 8'h9c == _T_5[7:0] ? image_0_156 : _GEN_155; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_157 = 8'h9d == _T_5[7:0] ? image_0_157 : _GEN_156; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_158 = 8'h9e == _T_5[7:0] ? image_0_158 : _GEN_157; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_159 = 8'h9f == _T_5[7:0] ? image_0_159 : _GEN_158; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_160 = 8'ha0 == _T_5[7:0] ? image_0_160 : _GEN_159; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_161 = 8'ha1 == _T_5[7:0] ? image_0_161 : _GEN_160; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_162 = 8'ha2 == _T_5[7:0] ? image_0_162 : _GEN_161; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_163 = 8'ha3 == _T_5[7:0] ? image_0_163 : _GEN_162; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_164 = 8'ha4 == _T_5[7:0] ? image_0_164 : _GEN_163; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_165 = 8'ha5 == _T_5[7:0] ? image_0_165 : _GEN_164; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_166 = 8'ha6 == _T_5[7:0] ? image_0_166 : _GEN_165; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_167 = 8'ha7 == _T_5[7:0] ? image_0_167 : _GEN_166; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_168 = 8'ha8 == _T_5[7:0] ? image_0_168 : _GEN_167; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_169 = 8'ha9 == _T_5[7:0] ? image_0_169 : _GEN_168; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_170 = 8'haa == _T_5[7:0] ? image_0_170 : _GEN_169; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_171 = 8'hab == _T_5[7:0] ? image_0_171 : _GEN_170; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_172 = 8'hac == _T_5[7:0] ? image_0_172 : _GEN_171; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_173 = 8'had == _T_5[7:0] ? image_0_173 : _GEN_172; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_174 = 8'hae == _T_5[7:0] ? image_0_174 : _GEN_173; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_175 = 8'haf == _T_5[7:0] ? image_0_175 : _GEN_174; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_176 = 8'hb0 == _T_5[7:0] ? image_0_176 : _GEN_175; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_177 = 8'hb1 == _T_5[7:0] ? image_0_177 : _GEN_176; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_178 = 8'hb2 == _T_5[7:0] ? image_0_178 : _GEN_177; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_179 = 8'hb3 == _T_5[7:0] ? image_0_179 : _GEN_178; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_180 = 8'hb4 == _T_5[7:0] ? image_0_180 : _GEN_179; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_181 = 8'hb5 == _T_5[7:0] ? image_0_181 : _GEN_180; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_182 = 8'hb6 == _T_5[7:0] ? image_0_182 : _GEN_181; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_183 = 8'hb7 == _T_5[7:0] ? image_0_183 : _GEN_182; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_184 = 8'hb8 == _T_5[7:0] ? image_0_184 : _GEN_183; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_185 = 8'hb9 == _T_5[7:0] ? image_0_185 : _GEN_184; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_186 = 8'hba == _T_5[7:0] ? image_0_186 : _GEN_185; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_187 = 8'hbb == _T_5[7:0] ? image_0_187 : _GEN_186; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_188 = 8'hbc == _T_5[7:0] ? image_0_188 : _GEN_187; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_189 = 8'hbd == _T_5[7:0] ? image_0_189 : _GEN_188; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_190 = 8'hbe == _T_5[7:0] ? image_0_190 : _GEN_189; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_191 = 8'hbf == _T_5[7:0] ? image_0_191 : _GEN_190; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_192 = 8'hc0 == _T_5[7:0] ? image_0_192 : _GEN_191; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_193 = 8'hc1 == _T_5[7:0] ? image_0_193 : _GEN_192; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_194 = 8'hc2 == _T_5[7:0] ? image_0_194 : _GEN_193; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_195 = 8'hc3 == _T_5[7:0] ? image_0_195 : _GEN_194; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_196 = 8'hc4 == _T_5[7:0] ? image_0_196 : _GEN_195; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_197 = 8'hc5 == _T_5[7:0] ? image_0_197 : _GEN_196; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_198 = 8'hc6 == _T_5[7:0] ? image_0_198 : _GEN_197; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_199 = 8'hc7 == _T_5[7:0] ? image_0_199 : _GEN_198; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_200 = 8'hc8 == _T_5[7:0] ? image_0_200 : _GEN_199; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_201 = 8'hc9 == _T_5[7:0] ? image_0_201 : _GEN_200; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_202 = 8'hca == _T_5[7:0] ? image_0_202 : _GEN_201; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_203 = 8'hcb == _T_5[7:0] ? image_0_203 : _GEN_202; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_204 = 8'hcc == _T_5[7:0] ? image_0_204 : _GEN_203; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_205 = 8'hcd == _T_5[7:0] ? image_0_205 : _GEN_204; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_206 = 8'hce == _T_5[7:0] ? image_0_206 : _GEN_205; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_207 = 8'hcf == _T_5[7:0] ? image_0_207 : _GEN_206; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_208 = 8'hd0 == _T_5[7:0] ? image_0_208 : _GEN_207; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_209 = 8'hd1 == _T_5[7:0] ? image_0_209 : _GEN_208; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_210 = 8'hd2 == _T_5[7:0] ? image_0_210 : _GEN_209; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_211 = 8'hd3 == _T_5[7:0] ? image_0_211 : _GEN_210; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_212 = 8'hd4 == _T_5[7:0] ? image_0_212 : _GEN_211; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_213 = 8'hd5 == _T_5[7:0] ? image_0_213 : _GEN_212; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_214 = 8'hd6 == _T_5[7:0] ? image_0_214 : _GEN_213; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_215 = 8'hd7 == _T_5[7:0] ? image_0_215 : _GEN_214; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_216 = 8'hd8 == _T_5[7:0] ? image_0_216 : _GEN_215; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_217 = 8'hd9 == _T_5[7:0] ? image_0_217 : _GEN_216; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_218 = 8'hda == _T_5[7:0] ? image_0_218 : _GEN_217; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_219 = 8'hdb == _T_5[7:0] ? image_0_219 : _GEN_218; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_220 = 8'hdc == _T_5[7:0] ? image_0_220 : _GEN_219; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_221 = 8'hdd == _T_5[7:0] ? image_0_221 : _GEN_220; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_222 = 8'hde == _T_5[7:0] ? image_0_222 : _GEN_221; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_223 = 8'hdf == _T_5[7:0] ? image_0_223 : _GEN_222; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_224 = 8'he0 == _T_5[7:0] ? image_0_224 : _GEN_223; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_225 = 8'he1 == _T_5[7:0] ? image_0_225 : _GEN_224; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_226 = 8'he2 == _T_5[7:0] ? image_0_226 : _GEN_225; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_227 = 8'he3 == _T_5[7:0] ? image_0_227 : _GEN_226; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_228 = 8'he4 == _T_5[7:0] ? image_0_228 : _GEN_227; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_229 = 8'he5 == _T_5[7:0] ? image_0_229 : _GEN_228; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_230 = 8'he6 == _T_5[7:0] ? image_0_230 : _GEN_229; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_231 = 8'he7 == _T_5[7:0] ? image_0_231 : _GEN_230; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_232 = 8'he8 == _T_5[7:0] ? image_0_232 : _GEN_231; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_233 = 8'he9 == _T_5[7:0] ? image_0_233 : _GEN_232; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_234 = 8'hea == _T_5[7:0] ? image_0_234 : _GEN_233; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_235 = 8'heb == _T_5[7:0] ? image_0_235 : _GEN_234; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_236 = 8'hec == _T_5[7:0] ? image_0_236 : _GEN_235; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_237 = 8'hed == _T_5[7:0] ? image_0_237 : _GEN_236; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_238 = 8'hee == _T_5[7:0] ? image_0_238 : _GEN_237; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_239 = 8'hef == _T_5[7:0] ? image_0_239 : _GEN_238; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_240 = 8'hf0 == _T_5[7:0] ? image_0_240 : _GEN_239; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_241 = 8'hf1 == _T_5[7:0] ? image_0_241 : _GEN_240; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_242 = 8'hf2 == _T_5[7:0] ? image_0_242 : _GEN_241; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_243 = 8'hf3 == _T_5[7:0] ? image_0_243 : _GEN_242; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_244 = 8'hf4 == _T_5[7:0] ? image_0_244 : _GEN_243; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_245 = 8'hf5 == _T_5[7:0] ? image_0_245 : _GEN_244; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_246 = 8'hf6 == _T_5[7:0] ? image_0_246 : _GEN_245; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_247 = 8'hf7 == _T_5[7:0] ? image_0_247 : _GEN_246; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_248 = 8'hf8 == _T_5[7:0] ? image_0_248 : _GEN_247; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_249 = 8'hf9 == _T_5[7:0] ? image_0_249 : _GEN_248; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_250 = 8'hfa == _T_5[7:0] ? image_0_250 : _GEN_249; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_253 = 8'h1 == _T_5[7:0] ? image_1_1 : image_1_0; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_254 = 8'h2 == _T_5[7:0] ? image_1_2 : _GEN_253; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_255 = 8'h3 == _T_5[7:0] ? image_1_3 : _GEN_254; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_256 = 8'h4 == _T_5[7:0] ? image_1_4 : _GEN_255; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_257 = 8'h5 == _T_5[7:0] ? image_1_5 : _GEN_256; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_258 = 8'h6 == _T_5[7:0] ? image_1_6 : _GEN_257; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_259 = 8'h7 == _T_5[7:0] ? image_1_7 : _GEN_258; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_260 = 8'h8 == _T_5[7:0] ? image_1_8 : _GEN_259; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_261 = 8'h9 == _T_5[7:0] ? image_1_9 : _GEN_260; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_262 = 8'ha == _T_5[7:0] ? image_1_10 : _GEN_261; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_263 = 8'hb == _T_5[7:0] ? image_1_11 : _GEN_262; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_264 = 8'hc == _T_5[7:0] ? image_1_12 : _GEN_263; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_265 = 8'hd == _T_5[7:0] ? image_1_13 : _GEN_264; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_266 = 8'he == _T_5[7:0] ? image_1_14 : _GEN_265; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_267 = 8'hf == _T_5[7:0] ? image_1_15 : _GEN_266; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_268 = 8'h10 == _T_5[7:0] ? image_1_16 : _GEN_267; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_269 = 8'h11 == _T_5[7:0] ? image_1_17 : _GEN_268; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_270 = 8'h12 == _T_5[7:0] ? image_1_18 : _GEN_269; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_271 = 8'h13 == _T_5[7:0] ? image_1_19 : _GEN_270; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_272 = 8'h14 == _T_5[7:0] ? image_1_20 : _GEN_271; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_273 = 8'h15 == _T_5[7:0] ? image_1_21 : _GEN_272; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_274 = 8'h16 == _T_5[7:0] ? image_1_22 : _GEN_273; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_275 = 8'h17 == _T_5[7:0] ? image_1_23 : _GEN_274; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_276 = 8'h18 == _T_5[7:0] ? image_1_24 : _GEN_275; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_277 = 8'h19 == _T_5[7:0] ? image_1_25 : _GEN_276; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_278 = 8'h1a == _T_5[7:0] ? image_1_26 : _GEN_277; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_279 = 8'h1b == _T_5[7:0] ? image_1_27 : _GEN_278; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_280 = 8'h1c == _T_5[7:0] ? image_1_28 : _GEN_279; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_281 = 8'h1d == _T_5[7:0] ? image_1_29 : _GEN_280; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_282 = 8'h1e == _T_5[7:0] ? image_1_30 : _GEN_281; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_283 = 8'h1f == _T_5[7:0] ? image_1_31 : _GEN_282; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_284 = 8'h20 == _T_5[7:0] ? image_1_32 : _GEN_283; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_285 = 8'h21 == _T_5[7:0] ? image_1_33 : _GEN_284; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_286 = 8'h22 == _T_5[7:0] ? image_1_34 : _GEN_285; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_287 = 8'h23 == _T_5[7:0] ? image_1_35 : _GEN_286; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_288 = 8'h24 == _T_5[7:0] ? image_1_36 : _GEN_287; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_289 = 8'h25 == _T_5[7:0] ? image_1_37 : _GEN_288; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_290 = 8'h26 == _T_5[7:0] ? image_1_38 : _GEN_289; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_291 = 8'h27 == _T_5[7:0] ? image_1_39 : _GEN_290; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_292 = 8'h28 == _T_5[7:0] ? image_1_40 : _GEN_291; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_293 = 8'h29 == _T_5[7:0] ? image_1_41 : _GEN_292; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_294 = 8'h2a == _T_5[7:0] ? image_1_42 : _GEN_293; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_295 = 8'h2b == _T_5[7:0] ? image_1_43 : _GEN_294; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_296 = 8'h2c == _T_5[7:0] ? image_1_44 : _GEN_295; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_297 = 8'h2d == _T_5[7:0] ? image_1_45 : _GEN_296; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_298 = 8'h2e == _T_5[7:0] ? image_1_46 : _GEN_297; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_299 = 8'h2f == _T_5[7:0] ? image_1_47 : _GEN_298; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_300 = 8'h30 == _T_5[7:0] ? image_1_48 : _GEN_299; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_301 = 8'h31 == _T_5[7:0] ? image_1_49 : _GEN_300; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_302 = 8'h32 == _T_5[7:0] ? image_1_50 : _GEN_301; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_303 = 8'h33 == _T_5[7:0] ? image_1_51 : _GEN_302; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_304 = 8'h34 == _T_5[7:0] ? image_1_52 : _GEN_303; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_305 = 8'h35 == _T_5[7:0] ? image_1_53 : _GEN_304; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_306 = 8'h36 == _T_5[7:0] ? image_1_54 : _GEN_305; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_307 = 8'h37 == _T_5[7:0] ? image_1_55 : _GEN_306; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_308 = 8'h38 == _T_5[7:0] ? image_1_56 : _GEN_307; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_309 = 8'h39 == _T_5[7:0] ? image_1_57 : _GEN_308; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_310 = 8'h3a == _T_5[7:0] ? image_1_58 : _GEN_309; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_311 = 8'h3b == _T_5[7:0] ? image_1_59 : _GEN_310; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_312 = 8'h3c == _T_5[7:0] ? image_1_60 : _GEN_311; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_313 = 8'h3d == _T_5[7:0] ? image_1_61 : _GEN_312; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_314 = 8'h3e == _T_5[7:0] ? image_1_62 : _GEN_313; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_315 = 8'h3f == _T_5[7:0] ? image_1_63 : _GEN_314; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_316 = 8'h40 == _T_5[7:0] ? image_1_64 : _GEN_315; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_317 = 8'h41 == _T_5[7:0] ? image_1_65 : _GEN_316; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_318 = 8'h42 == _T_5[7:0] ? image_1_66 : _GEN_317; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_319 = 8'h43 == _T_5[7:0] ? image_1_67 : _GEN_318; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_320 = 8'h44 == _T_5[7:0] ? image_1_68 : _GEN_319; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_321 = 8'h45 == _T_5[7:0] ? image_1_69 : _GEN_320; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_322 = 8'h46 == _T_5[7:0] ? image_1_70 : _GEN_321; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_323 = 8'h47 == _T_5[7:0] ? image_1_71 : _GEN_322; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_324 = 8'h48 == _T_5[7:0] ? image_1_72 : _GEN_323; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_325 = 8'h49 == _T_5[7:0] ? image_1_73 : _GEN_324; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_326 = 8'h4a == _T_5[7:0] ? image_1_74 : _GEN_325; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_327 = 8'h4b == _T_5[7:0] ? image_1_75 : _GEN_326; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_328 = 8'h4c == _T_5[7:0] ? image_1_76 : _GEN_327; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_329 = 8'h4d == _T_5[7:0] ? image_1_77 : _GEN_328; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_330 = 8'h4e == _T_5[7:0] ? image_1_78 : _GEN_329; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_331 = 8'h4f == _T_5[7:0] ? image_1_79 : _GEN_330; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_332 = 8'h50 == _T_5[7:0] ? image_1_80 : _GEN_331; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_333 = 8'h51 == _T_5[7:0] ? image_1_81 : _GEN_332; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_334 = 8'h52 == _T_5[7:0] ? image_1_82 : _GEN_333; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_335 = 8'h53 == _T_5[7:0] ? image_1_83 : _GEN_334; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_336 = 8'h54 == _T_5[7:0] ? image_1_84 : _GEN_335; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_337 = 8'h55 == _T_5[7:0] ? image_1_85 : _GEN_336; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_338 = 8'h56 == _T_5[7:0] ? image_1_86 : _GEN_337; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_339 = 8'h57 == _T_5[7:0] ? image_1_87 : _GEN_338; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_340 = 8'h58 == _T_5[7:0] ? image_1_88 : _GEN_339; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_341 = 8'h59 == _T_5[7:0] ? image_1_89 : _GEN_340; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_342 = 8'h5a == _T_5[7:0] ? image_1_90 : _GEN_341; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_343 = 8'h5b == _T_5[7:0] ? image_1_91 : _GEN_342; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_344 = 8'h5c == _T_5[7:0] ? image_1_92 : _GEN_343; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_345 = 8'h5d == _T_5[7:0] ? image_1_93 : _GEN_344; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_346 = 8'h5e == _T_5[7:0] ? image_1_94 : _GEN_345; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_347 = 8'h5f == _T_5[7:0] ? image_1_95 : _GEN_346; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_348 = 8'h60 == _T_5[7:0] ? image_1_96 : _GEN_347; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_349 = 8'h61 == _T_5[7:0] ? image_1_97 : _GEN_348; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_350 = 8'h62 == _T_5[7:0] ? image_1_98 : _GEN_349; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_351 = 8'h63 == _T_5[7:0] ? image_1_99 : _GEN_350; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_352 = 8'h64 == _T_5[7:0] ? image_1_100 : _GEN_351; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_353 = 8'h65 == _T_5[7:0] ? image_1_101 : _GEN_352; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_354 = 8'h66 == _T_5[7:0] ? image_1_102 : _GEN_353; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_355 = 8'h67 == _T_5[7:0] ? image_1_103 : _GEN_354; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_356 = 8'h68 == _T_5[7:0] ? image_1_104 : _GEN_355; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_357 = 8'h69 == _T_5[7:0] ? image_1_105 : _GEN_356; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_358 = 8'h6a == _T_5[7:0] ? image_1_106 : _GEN_357; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_359 = 8'h6b == _T_5[7:0] ? image_1_107 : _GEN_358; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_360 = 8'h6c == _T_5[7:0] ? image_1_108 : _GEN_359; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_361 = 8'h6d == _T_5[7:0] ? image_1_109 : _GEN_360; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_362 = 8'h6e == _T_5[7:0] ? image_1_110 : _GEN_361; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_363 = 8'h6f == _T_5[7:0] ? image_1_111 : _GEN_362; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_364 = 8'h70 == _T_5[7:0] ? image_1_112 : _GEN_363; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_365 = 8'h71 == _T_5[7:0] ? image_1_113 : _GEN_364; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_366 = 8'h72 == _T_5[7:0] ? image_1_114 : _GEN_365; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_367 = 8'h73 == _T_5[7:0] ? image_1_115 : _GEN_366; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_368 = 8'h74 == _T_5[7:0] ? image_1_116 : _GEN_367; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_369 = 8'h75 == _T_5[7:0] ? image_1_117 : _GEN_368; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_370 = 8'h76 == _T_5[7:0] ? image_1_118 : _GEN_369; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_371 = 8'h77 == _T_5[7:0] ? image_1_119 : _GEN_370; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_372 = 8'h78 == _T_5[7:0] ? image_1_120 : _GEN_371; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_373 = 8'h79 == _T_5[7:0] ? image_1_121 : _GEN_372; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_374 = 8'h7a == _T_5[7:0] ? image_1_122 : _GEN_373; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_375 = 8'h7b == _T_5[7:0] ? image_1_123 : _GEN_374; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_376 = 8'h7c == _T_5[7:0] ? image_1_124 : _GEN_375; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_377 = 8'h7d == _T_5[7:0] ? image_1_125 : _GEN_376; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_378 = 8'h7e == _T_5[7:0] ? image_1_126 : _GEN_377; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_379 = 8'h7f == _T_5[7:0] ? image_1_127 : _GEN_378; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_380 = 8'h80 == _T_5[7:0] ? image_1_128 : _GEN_379; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_381 = 8'h81 == _T_5[7:0] ? image_1_129 : _GEN_380; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_382 = 8'h82 == _T_5[7:0] ? image_1_130 : _GEN_381; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_383 = 8'h83 == _T_5[7:0] ? image_1_131 : _GEN_382; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_384 = 8'h84 == _T_5[7:0] ? image_1_132 : _GEN_383; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_385 = 8'h85 == _T_5[7:0] ? image_1_133 : _GEN_384; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_386 = 8'h86 == _T_5[7:0] ? image_1_134 : _GEN_385; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_387 = 8'h87 == _T_5[7:0] ? image_1_135 : _GEN_386; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_388 = 8'h88 == _T_5[7:0] ? image_1_136 : _GEN_387; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_389 = 8'h89 == _T_5[7:0] ? image_1_137 : _GEN_388; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_390 = 8'h8a == _T_5[7:0] ? image_1_138 : _GEN_389; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_391 = 8'h8b == _T_5[7:0] ? image_1_139 : _GEN_390; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_392 = 8'h8c == _T_5[7:0] ? image_1_140 : _GEN_391; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_393 = 8'h8d == _T_5[7:0] ? image_1_141 : _GEN_392; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_394 = 8'h8e == _T_5[7:0] ? image_1_142 : _GEN_393; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_395 = 8'h8f == _T_5[7:0] ? image_1_143 : _GEN_394; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_396 = 8'h90 == _T_5[7:0] ? image_1_144 : _GEN_395; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_397 = 8'h91 == _T_5[7:0] ? image_1_145 : _GEN_396; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_398 = 8'h92 == _T_5[7:0] ? image_1_146 : _GEN_397; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_399 = 8'h93 == _T_5[7:0] ? image_1_147 : _GEN_398; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_400 = 8'h94 == _T_5[7:0] ? image_1_148 : _GEN_399; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_401 = 8'h95 == _T_5[7:0] ? image_1_149 : _GEN_400; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_402 = 8'h96 == _T_5[7:0] ? image_1_150 : _GEN_401; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_403 = 8'h97 == _T_5[7:0] ? image_1_151 : _GEN_402; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_404 = 8'h98 == _T_5[7:0] ? image_1_152 : _GEN_403; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_405 = 8'h99 == _T_5[7:0] ? image_1_153 : _GEN_404; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_406 = 8'h9a == _T_5[7:0] ? image_1_154 : _GEN_405; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_407 = 8'h9b == _T_5[7:0] ? image_1_155 : _GEN_406; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_408 = 8'h9c == _T_5[7:0] ? image_1_156 : _GEN_407; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_409 = 8'h9d == _T_5[7:0] ? image_1_157 : _GEN_408; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_410 = 8'h9e == _T_5[7:0] ? image_1_158 : _GEN_409; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_411 = 8'h9f == _T_5[7:0] ? image_1_159 : _GEN_410; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_412 = 8'ha0 == _T_5[7:0] ? image_1_160 : _GEN_411; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_413 = 8'ha1 == _T_5[7:0] ? image_1_161 : _GEN_412; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_414 = 8'ha2 == _T_5[7:0] ? image_1_162 : _GEN_413; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_415 = 8'ha3 == _T_5[7:0] ? image_1_163 : _GEN_414; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_416 = 8'ha4 == _T_5[7:0] ? image_1_164 : _GEN_415; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_417 = 8'ha5 == _T_5[7:0] ? image_1_165 : _GEN_416; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_418 = 8'ha6 == _T_5[7:0] ? image_1_166 : _GEN_417; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_419 = 8'ha7 == _T_5[7:0] ? image_1_167 : _GEN_418; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_420 = 8'ha8 == _T_5[7:0] ? image_1_168 : _GEN_419; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_421 = 8'ha9 == _T_5[7:0] ? image_1_169 : _GEN_420; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_422 = 8'haa == _T_5[7:0] ? image_1_170 : _GEN_421; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_423 = 8'hab == _T_5[7:0] ? image_1_171 : _GEN_422; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_424 = 8'hac == _T_5[7:0] ? image_1_172 : _GEN_423; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_425 = 8'had == _T_5[7:0] ? image_1_173 : _GEN_424; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_426 = 8'hae == _T_5[7:0] ? image_1_174 : _GEN_425; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_427 = 8'haf == _T_5[7:0] ? image_1_175 : _GEN_426; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_428 = 8'hb0 == _T_5[7:0] ? image_1_176 : _GEN_427; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_429 = 8'hb1 == _T_5[7:0] ? image_1_177 : _GEN_428; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_430 = 8'hb2 == _T_5[7:0] ? image_1_178 : _GEN_429; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_431 = 8'hb3 == _T_5[7:0] ? image_1_179 : _GEN_430; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_432 = 8'hb4 == _T_5[7:0] ? image_1_180 : _GEN_431; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_433 = 8'hb5 == _T_5[7:0] ? image_1_181 : _GEN_432; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_434 = 8'hb6 == _T_5[7:0] ? image_1_182 : _GEN_433; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_435 = 8'hb7 == _T_5[7:0] ? image_1_183 : _GEN_434; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_436 = 8'hb8 == _T_5[7:0] ? image_1_184 : _GEN_435; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_437 = 8'hb9 == _T_5[7:0] ? image_1_185 : _GEN_436; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_438 = 8'hba == _T_5[7:0] ? image_1_186 : _GEN_437; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_439 = 8'hbb == _T_5[7:0] ? image_1_187 : _GEN_438; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_440 = 8'hbc == _T_5[7:0] ? image_1_188 : _GEN_439; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_441 = 8'hbd == _T_5[7:0] ? image_1_189 : _GEN_440; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_442 = 8'hbe == _T_5[7:0] ? image_1_190 : _GEN_441; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_443 = 8'hbf == _T_5[7:0] ? image_1_191 : _GEN_442; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_444 = 8'hc0 == _T_5[7:0] ? image_1_192 : _GEN_443; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_445 = 8'hc1 == _T_5[7:0] ? image_1_193 : _GEN_444; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_446 = 8'hc2 == _T_5[7:0] ? image_1_194 : _GEN_445; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_447 = 8'hc3 == _T_5[7:0] ? image_1_195 : _GEN_446; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_448 = 8'hc4 == _T_5[7:0] ? image_1_196 : _GEN_447; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_449 = 8'hc5 == _T_5[7:0] ? image_1_197 : _GEN_448; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_450 = 8'hc6 == _T_5[7:0] ? image_1_198 : _GEN_449; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_451 = 8'hc7 == _T_5[7:0] ? image_1_199 : _GEN_450; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_452 = 8'hc8 == _T_5[7:0] ? image_1_200 : _GEN_451; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_453 = 8'hc9 == _T_5[7:0] ? image_1_201 : _GEN_452; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_454 = 8'hca == _T_5[7:0] ? image_1_202 : _GEN_453; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_455 = 8'hcb == _T_5[7:0] ? image_1_203 : _GEN_454; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_456 = 8'hcc == _T_5[7:0] ? image_1_204 : _GEN_455; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_457 = 8'hcd == _T_5[7:0] ? image_1_205 : _GEN_456; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_458 = 8'hce == _T_5[7:0] ? image_1_206 : _GEN_457; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_459 = 8'hcf == _T_5[7:0] ? image_1_207 : _GEN_458; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_460 = 8'hd0 == _T_5[7:0] ? image_1_208 : _GEN_459; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_461 = 8'hd1 == _T_5[7:0] ? image_1_209 : _GEN_460; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_462 = 8'hd2 == _T_5[7:0] ? image_1_210 : _GEN_461; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_463 = 8'hd3 == _T_5[7:0] ? image_1_211 : _GEN_462; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_464 = 8'hd4 == _T_5[7:0] ? image_1_212 : _GEN_463; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_465 = 8'hd5 == _T_5[7:0] ? image_1_213 : _GEN_464; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_466 = 8'hd6 == _T_5[7:0] ? image_1_214 : _GEN_465; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_467 = 8'hd7 == _T_5[7:0] ? image_1_215 : _GEN_466; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_468 = 8'hd8 == _T_5[7:0] ? image_1_216 : _GEN_467; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_469 = 8'hd9 == _T_5[7:0] ? image_1_217 : _GEN_468; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_470 = 8'hda == _T_5[7:0] ? image_1_218 : _GEN_469; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_471 = 8'hdb == _T_5[7:0] ? image_1_219 : _GEN_470; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_472 = 8'hdc == _T_5[7:0] ? image_1_220 : _GEN_471; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_473 = 8'hdd == _T_5[7:0] ? image_1_221 : _GEN_472; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_474 = 8'hde == _T_5[7:0] ? image_1_222 : _GEN_473; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_475 = 8'hdf == _T_5[7:0] ? image_1_223 : _GEN_474; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_476 = 8'he0 == _T_5[7:0] ? image_1_224 : _GEN_475; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_477 = 8'he1 == _T_5[7:0] ? image_1_225 : _GEN_476; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_478 = 8'he2 == _T_5[7:0] ? image_1_226 : _GEN_477; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_479 = 8'he3 == _T_5[7:0] ? image_1_227 : _GEN_478; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_480 = 8'he4 == _T_5[7:0] ? image_1_228 : _GEN_479; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_481 = 8'he5 == _T_5[7:0] ? image_1_229 : _GEN_480; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_482 = 8'he6 == _T_5[7:0] ? image_1_230 : _GEN_481; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_483 = 8'he7 == _T_5[7:0] ? image_1_231 : _GEN_482; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_484 = 8'he8 == _T_5[7:0] ? image_1_232 : _GEN_483; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_485 = 8'he9 == _T_5[7:0] ? image_1_233 : _GEN_484; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_486 = 8'hea == _T_5[7:0] ? image_1_234 : _GEN_485; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_487 = 8'heb == _T_5[7:0] ? image_1_235 : _GEN_486; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_488 = 8'hec == _T_5[7:0] ? image_1_236 : _GEN_487; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_489 = 8'hed == _T_5[7:0] ? image_1_237 : _GEN_488; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_490 = 8'hee == _T_5[7:0] ? image_1_238 : _GEN_489; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_491 = 8'hef == _T_5[7:0] ? image_1_239 : _GEN_490; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_492 = 8'hf0 == _T_5[7:0] ? image_1_240 : _GEN_491; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_493 = 8'hf1 == _T_5[7:0] ? image_1_241 : _GEN_492; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_494 = 8'hf2 == _T_5[7:0] ? image_1_242 : _GEN_493; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_495 = 8'hf3 == _T_5[7:0] ? image_1_243 : _GEN_494; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_496 = 8'hf4 == _T_5[7:0] ? image_1_244 : _GEN_495; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_497 = 8'hf5 == _T_5[7:0] ? image_1_245 : _GEN_496; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_498 = 8'hf6 == _T_5[7:0] ? image_1_246 : _GEN_497; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_499 = 8'hf7 == _T_5[7:0] ? image_1_247 : _GEN_498; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_500 = 8'hf8 == _T_5[7:0] ? image_1_248 : _GEN_499; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_501 = 8'hf9 == _T_5[7:0] ? image_1_249 : _GEN_500; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_502 = 8'hfa == _T_5[7:0] ? image_1_250 : _GEN_501; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_505 = 8'h1 == _T_5[7:0] ? image_2_1 : image_2_0; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_506 = 8'h2 == _T_5[7:0] ? image_2_2 : _GEN_505; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_507 = 8'h3 == _T_5[7:0] ? image_2_3 : _GEN_506; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_508 = 8'h4 == _T_5[7:0] ? image_2_4 : _GEN_507; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_509 = 8'h5 == _T_5[7:0] ? image_2_5 : _GEN_508; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_510 = 8'h6 == _T_5[7:0] ? image_2_6 : _GEN_509; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_511 = 8'h7 == _T_5[7:0] ? image_2_7 : _GEN_510; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_512 = 8'h8 == _T_5[7:0] ? image_2_8 : _GEN_511; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_513 = 8'h9 == _T_5[7:0] ? image_2_9 : _GEN_512; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_514 = 8'ha == _T_5[7:0] ? image_2_10 : _GEN_513; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_515 = 8'hb == _T_5[7:0] ? image_2_11 : _GEN_514; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_516 = 8'hc == _T_5[7:0] ? image_2_12 : _GEN_515; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_517 = 8'hd == _T_5[7:0] ? image_2_13 : _GEN_516; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_518 = 8'he == _T_5[7:0] ? image_2_14 : _GEN_517; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_519 = 8'hf == _T_5[7:0] ? image_2_15 : _GEN_518; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_520 = 8'h10 == _T_5[7:0] ? image_2_16 : _GEN_519; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_521 = 8'h11 == _T_5[7:0] ? image_2_17 : _GEN_520; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_522 = 8'h12 == _T_5[7:0] ? image_2_18 : _GEN_521; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_523 = 8'h13 == _T_5[7:0] ? image_2_19 : _GEN_522; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_524 = 8'h14 == _T_5[7:0] ? image_2_20 : _GEN_523; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_525 = 8'h15 == _T_5[7:0] ? image_2_21 : _GEN_524; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_526 = 8'h16 == _T_5[7:0] ? image_2_22 : _GEN_525; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_527 = 8'h17 == _T_5[7:0] ? image_2_23 : _GEN_526; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_528 = 8'h18 == _T_5[7:0] ? image_2_24 : _GEN_527; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_529 = 8'h19 == _T_5[7:0] ? image_2_25 : _GEN_528; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_530 = 8'h1a == _T_5[7:0] ? image_2_26 : _GEN_529; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_531 = 8'h1b == _T_5[7:0] ? image_2_27 : _GEN_530; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_532 = 8'h1c == _T_5[7:0] ? image_2_28 : _GEN_531; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_533 = 8'h1d == _T_5[7:0] ? image_2_29 : _GEN_532; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_534 = 8'h1e == _T_5[7:0] ? image_2_30 : _GEN_533; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_535 = 8'h1f == _T_5[7:0] ? image_2_31 : _GEN_534; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_536 = 8'h20 == _T_5[7:0] ? image_2_32 : _GEN_535; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_537 = 8'h21 == _T_5[7:0] ? image_2_33 : _GEN_536; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_538 = 8'h22 == _T_5[7:0] ? image_2_34 : _GEN_537; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_539 = 8'h23 == _T_5[7:0] ? image_2_35 : _GEN_538; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_540 = 8'h24 == _T_5[7:0] ? image_2_36 : _GEN_539; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_541 = 8'h25 == _T_5[7:0] ? image_2_37 : _GEN_540; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_542 = 8'h26 == _T_5[7:0] ? image_2_38 : _GEN_541; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_543 = 8'h27 == _T_5[7:0] ? image_2_39 : _GEN_542; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_544 = 8'h28 == _T_5[7:0] ? image_2_40 : _GEN_543; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_545 = 8'h29 == _T_5[7:0] ? image_2_41 : _GEN_544; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_546 = 8'h2a == _T_5[7:0] ? image_2_42 : _GEN_545; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_547 = 8'h2b == _T_5[7:0] ? image_2_43 : _GEN_546; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_548 = 8'h2c == _T_5[7:0] ? image_2_44 : _GEN_547; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_549 = 8'h2d == _T_5[7:0] ? image_2_45 : _GEN_548; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_550 = 8'h2e == _T_5[7:0] ? image_2_46 : _GEN_549; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_551 = 8'h2f == _T_5[7:0] ? image_2_47 : _GEN_550; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_552 = 8'h30 == _T_5[7:0] ? image_2_48 : _GEN_551; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_553 = 8'h31 == _T_5[7:0] ? image_2_49 : _GEN_552; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_554 = 8'h32 == _T_5[7:0] ? image_2_50 : _GEN_553; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_555 = 8'h33 == _T_5[7:0] ? image_2_51 : _GEN_554; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_556 = 8'h34 == _T_5[7:0] ? image_2_52 : _GEN_555; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_557 = 8'h35 == _T_5[7:0] ? image_2_53 : _GEN_556; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_558 = 8'h36 == _T_5[7:0] ? image_2_54 : _GEN_557; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_559 = 8'h37 == _T_5[7:0] ? image_2_55 : _GEN_558; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_560 = 8'h38 == _T_5[7:0] ? image_2_56 : _GEN_559; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_561 = 8'h39 == _T_5[7:0] ? image_2_57 : _GEN_560; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_562 = 8'h3a == _T_5[7:0] ? image_2_58 : _GEN_561; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_563 = 8'h3b == _T_5[7:0] ? image_2_59 : _GEN_562; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_564 = 8'h3c == _T_5[7:0] ? image_2_60 : _GEN_563; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_565 = 8'h3d == _T_5[7:0] ? image_2_61 : _GEN_564; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_566 = 8'h3e == _T_5[7:0] ? image_2_62 : _GEN_565; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_567 = 8'h3f == _T_5[7:0] ? image_2_63 : _GEN_566; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_568 = 8'h40 == _T_5[7:0] ? image_2_64 : _GEN_567; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_569 = 8'h41 == _T_5[7:0] ? image_2_65 : _GEN_568; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_570 = 8'h42 == _T_5[7:0] ? image_2_66 : _GEN_569; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_571 = 8'h43 == _T_5[7:0] ? image_2_67 : _GEN_570; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_572 = 8'h44 == _T_5[7:0] ? image_2_68 : _GEN_571; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_573 = 8'h45 == _T_5[7:0] ? image_2_69 : _GEN_572; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_574 = 8'h46 == _T_5[7:0] ? image_2_70 : _GEN_573; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_575 = 8'h47 == _T_5[7:0] ? image_2_71 : _GEN_574; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_576 = 8'h48 == _T_5[7:0] ? image_2_72 : _GEN_575; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_577 = 8'h49 == _T_5[7:0] ? image_2_73 : _GEN_576; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_578 = 8'h4a == _T_5[7:0] ? image_2_74 : _GEN_577; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_579 = 8'h4b == _T_5[7:0] ? image_2_75 : _GEN_578; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_580 = 8'h4c == _T_5[7:0] ? image_2_76 : _GEN_579; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_581 = 8'h4d == _T_5[7:0] ? image_2_77 : _GEN_580; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_582 = 8'h4e == _T_5[7:0] ? image_2_78 : _GEN_581; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_583 = 8'h4f == _T_5[7:0] ? image_2_79 : _GEN_582; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_584 = 8'h50 == _T_5[7:0] ? image_2_80 : _GEN_583; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_585 = 8'h51 == _T_5[7:0] ? image_2_81 : _GEN_584; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_586 = 8'h52 == _T_5[7:0] ? image_2_82 : _GEN_585; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_587 = 8'h53 == _T_5[7:0] ? image_2_83 : _GEN_586; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_588 = 8'h54 == _T_5[7:0] ? image_2_84 : _GEN_587; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_589 = 8'h55 == _T_5[7:0] ? image_2_85 : _GEN_588; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_590 = 8'h56 == _T_5[7:0] ? image_2_86 : _GEN_589; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_591 = 8'h57 == _T_5[7:0] ? image_2_87 : _GEN_590; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_592 = 8'h58 == _T_5[7:0] ? image_2_88 : _GEN_591; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_593 = 8'h59 == _T_5[7:0] ? image_2_89 : _GEN_592; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_594 = 8'h5a == _T_5[7:0] ? image_2_90 : _GEN_593; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_595 = 8'h5b == _T_5[7:0] ? image_2_91 : _GEN_594; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_596 = 8'h5c == _T_5[7:0] ? image_2_92 : _GEN_595; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_597 = 8'h5d == _T_5[7:0] ? image_2_93 : _GEN_596; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_598 = 8'h5e == _T_5[7:0] ? image_2_94 : _GEN_597; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_599 = 8'h5f == _T_5[7:0] ? image_2_95 : _GEN_598; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_600 = 8'h60 == _T_5[7:0] ? image_2_96 : _GEN_599; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_601 = 8'h61 == _T_5[7:0] ? image_2_97 : _GEN_600; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_602 = 8'h62 == _T_5[7:0] ? image_2_98 : _GEN_601; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_603 = 8'h63 == _T_5[7:0] ? image_2_99 : _GEN_602; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_604 = 8'h64 == _T_5[7:0] ? image_2_100 : _GEN_603; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_605 = 8'h65 == _T_5[7:0] ? image_2_101 : _GEN_604; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_606 = 8'h66 == _T_5[7:0] ? image_2_102 : _GEN_605; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_607 = 8'h67 == _T_5[7:0] ? image_2_103 : _GEN_606; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_608 = 8'h68 == _T_5[7:0] ? image_2_104 : _GEN_607; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_609 = 8'h69 == _T_5[7:0] ? image_2_105 : _GEN_608; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_610 = 8'h6a == _T_5[7:0] ? image_2_106 : _GEN_609; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_611 = 8'h6b == _T_5[7:0] ? image_2_107 : _GEN_610; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_612 = 8'h6c == _T_5[7:0] ? image_2_108 : _GEN_611; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_613 = 8'h6d == _T_5[7:0] ? image_2_109 : _GEN_612; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_614 = 8'h6e == _T_5[7:0] ? image_2_110 : _GEN_613; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_615 = 8'h6f == _T_5[7:0] ? image_2_111 : _GEN_614; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_616 = 8'h70 == _T_5[7:0] ? image_2_112 : _GEN_615; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_617 = 8'h71 == _T_5[7:0] ? image_2_113 : _GEN_616; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_618 = 8'h72 == _T_5[7:0] ? image_2_114 : _GEN_617; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_619 = 8'h73 == _T_5[7:0] ? image_2_115 : _GEN_618; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_620 = 8'h74 == _T_5[7:0] ? image_2_116 : _GEN_619; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_621 = 8'h75 == _T_5[7:0] ? image_2_117 : _GEN_620; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_622 = 8'h76 == _T_5[7:0] ? image_2_118 : _GEN_621; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_623 = 8'h77 == _T_5[7:0] ? image_2_119 : _GEN_622; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_624 = 8'h78 == _T_5[7:0] ? image_2_120 : _GEN_623; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_625 = 8'h79 == _T_5[7:0] ? image_2_121 : _GEN_624; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_626 = 8'h7a == _T_5[7:0] ? image_2_122 : _GEN_625; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_627 = 8'h7b == _T_5[7:0] ? image_2_123 : _GEN_626; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_628 = 8'h7c == _T_5[7:0] ? image_2_124 : _GEN_627; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_629 = 8'h7d == _T_5[7:0] ? image_2_125 : _GEN_628; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_630 = 8'h7e == _T_5[7:0] ? image_2_126 : _GEN_629; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_631 = 8'h7f == _T_5[7:0] ? image_2_127 : _GEN_630; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_632 = 8'h80 == _T_5[7:0] ? image_2_128 : _GEN_631; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_633 = 8'h81 == _T_5[7:0] ? image_2_129 : _GEN_632; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_634 = 8'h82 == _T_5[7:0] ? image_2_130 : _GEN_633; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_635 = 8'h83 == _T_5[7:0] ? image_2_131 : _GEN_634; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_636 = 8'h84 == _T_5[7:0] ? image_2_132 : _GEN_635; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_637 = 8'h85 == _T_5[7:0] ? image_2_133 : _GEN_636; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_638 = 8'h86 == _T_5[7:0] ? image_2_134 : _GEN_637; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_639 = 8'h87 == _T_5[7:0] ? image_2_135 : _GEN_638; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_640 = 8'h88 == _T_5[7:0] ? image_2_136 : _GEN_639; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_641 = 8'h89 == _T_5[7:0] ? image_2_137 : _GEN_640; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_642 = 8'h8a == _T_5[7:0] ? image_2_138 : _GEN_641; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_643 = 8'h8b == _T_5[7:0] ? image_2_139 : _GEN_642; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_644 = 8'h8c == _T_5[7:0] ? image_2_140 : _GEN_643; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_645 = 8'h8d == _T_5[7:0] ? image_2_141 : _GEN_644; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_646 = 8'h8e == _T_5[7:0] ? image_2_142 : _GEN_645; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_647 = 8'h8f == _T_5[7:0] ? image_2_143 : _GEN_646; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_648 = 8'h90 == _T_5[7:0] ? image_2_144 : _GEN_647; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_649 = 8'h91 == _T_5[7:0] ? image_2_145 : _GEN_648; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_650 = 8'h92 == _T_5[7:0] ? image_2_146 : _GEN_649; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_651 = 8'h93 == _T_5[7:0] ? image_2_147 : _GEN_650; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_652 = 8'h94 == _T_5[7:0] ? image_2_148 : _GEN_651; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_653 = 8'h95 == _T_5[7:0] ? image_2_149 : _GEN_652; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_654 = 8'h96 == _T_5[7:0] ? image_2_150 : _GEN_653; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_655 = 8'h97 == _T_5[7:0] ? image_2_151 : _GEN_654; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_656 = 8'h98 == _T_5[7:0] ? image_2_152 : _GEN_655; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_657 = 8'h99 == _T_5[7:0] ? image_2_153 : _GEN_656; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_658 = 8'h9a == _T_5[7:0] ? image_2_154 : _GEN_657; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_659 = 8'h9b == _T_5[7:0] ? image_2_155 : _GEN_658; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_660 = 8'h9c == _T_5[7:0] ? image_2_156 : _GEN_659; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_661 = 8'h9d == _T_5[7:0] ? image_2_157 : _GEN_660; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_662 = 8'h9e == _T_5[7:0] ? image_2_158 : _GEN_661; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_663 = 8'h9f == _T_5[7:0] ? image_2_159 : _GEN_662; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_664 = 8'ha0 == _T_5[7:0] ? image_2_160 : _GEN_663; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_665 = 8'ha1 == _T_5[7:0] ? image_2_161 : _GEN_664; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_666 = 8'ha2 == _T_5[7:0] ? image_2_162 : _GEN_665; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_667 = 8'ha3 == _T_5[7:0] ? image_2_163 : _GEN_666; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_668 = 8'ha4 == _T_5[7:0] ? image_2_164 : _GEN_667; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_669 = 8'ha5 == _T_5[7:0] ? image_2_165 : _GEN_668; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_670 = 8'ha6 == _T_5[7:0] ? image_2_166 : _GEN_669; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_671 = 8'ha7 == _T_5[7:0] ? image_2_167 : _GEN_670; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_672 = 8'ha8 == _T_5[7:0] ? image_2_168 : _GEN_671; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_673 = 8'ha9 == _T_5[7:0] ? image_2_169 : _GEN_672; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_674 = 8'haa == _T_5[7:0] ? image_2_170 : _GEN_673; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_675 = 8'hab == _T_5[7:0] ? image_2_171 : _GEN_674; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_676 = 8'hac == _T_5[7:0] ? image_2_172 : _GEN_675; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_677 = 8'had == _T_5[7:0] ? image_2_173 : _GEN_676; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_678 = 8'hae == _T_5[7:0] ? image_2_174 : _GEN_677; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_679 = 8'haf == _T_5[7:0] ? image_2_175 : _GEN_678; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_680 = 8'hb0 == _T_5[7:0] ? image_2_176 : _GEN_679; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_681 = 8'hb1 == _T_5[7:0] ? image_2_177 : _GEN_680; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_682 = 8'hb2 == _T_5[7:0] ? image_2_178 : _GEN_681; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_683 = 8'hb3 == _T_5[7:0] ? image_2_179 : _GEN_682; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_684 = 8'hb4 == _T_5[7:0] ? image_2_180 : _GEN_683; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_685 = 8'hb5 == _T_5[7:0] ? image_2_181 : _GEN_684; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_686 = 8'hb6 == _T_5[7:0] ? image_2_182 : _GEN_685; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_687 = 8'hb7 == _T_5[7:0] ? image_2_183 : _GEN_686; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_688 = 8'hb8 == _T_5[7:0] ? image_2_184 : _GEN_687; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_689 = 8'hb9 == _T_5[7:0] ? image_2_185 : _GEN_688; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_690 = 8'hba == _T_5[7:0] ? image_2_186 : _GEN_689; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_691 = 8'hbb == _T_5[7:0] ? image_2_187 : _GEN_690; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_692 = 8'hbc == _T_5[7:0] ? image_2_188 : _GEN_691; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_693 = 8'hbd == _T_5[7:0] ? image_2_189 : _GEN_692; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_694 = 8'hbe == _T_5[7:0] ? image_2_190 : _GEN_693; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_695 = 8'hbf == _T_5[7:0] ? image_2_191 : _GEN_694; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_696 = 8'hc0 == _T_5[7:0] ? image_2_192 : _GEN_695; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_697 = 8'hc1 == _T_5[7:0] ? image_2_193 : _GEN_696; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_698 = 8'hc2 == _T_5[7:0] ? image_2_194 : _GEN_697; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_699 = 8'hc3 == _T_5[7:0] ? image_2_195 : _GEN_698; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_700 = 8'hc4 == _T_5[7:0] ? image_2_196 : _GEN_699; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_701 = 8'hc5 == _T_5[7:0] ? image_2_197 : _GEN_700; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_702 = 8'hc6 == _T_5[7:0] ? image_2_198 : _GEN_701; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_703 = 8'hc7 == _T_5[7:0] ? image_2_199 : _GEN_702; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_704 = 8'hc8 == _T_5[7:0] ? image_2_200 : _GEN_703; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_705 = 8'hc9 == _T_5[7:0] ? image_2_201 : _GEN_704; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_706 = 8'hca == _T_5[7:0] ? image_2_202 : _GEN_705; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_707 = 8'hcb == _T_5[7:0] ? image_2_203 : _GEN_706; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_708 = 8'hcc == _T_5[7:0] ? image_2_204 : _GEN_707; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_709 = 8'hcd == _T_5[7:0] ? image_2_205 : _GEN_708; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_710 = 8'hce == _T_5[7:0] ? image_2_206 : _GEN_709; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_711 = 8'hcf == _T_5[7:0] ? image_2_207 : _GEN_710; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_712 = 8'hd0 == _T_5[7:0] ? image_2_208 : _GEN_711; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_713 = 8'hd1 == _T_5[7:0] ? image_2_209 : _GEN_712; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_714 = 8'hd2 == _T_5[7:0] ? image_2_210 : _GEN_713; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_715 = 8'hd3 == _T_5[7:0] ? image_2_211 : _GEN_714; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_716 = 8'hd4 == _T_5[7:0] ? image_2_212 : _GEN_715; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_717 = 8'hd5 == _T_5[7:0] ? image_2_213 : _GEN_716; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_718 = 8'hd6 == _T_5[7:0] ? image_2_214 : _GEN_717; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_719 = 8'hd7 == _T_5[7:0] ? image_2_215 : _GEN_718; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_720 = 8'hd8 == _T_5[7:0] ? image_2_216 : _GEN_719; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_721 = 8'hd9 == _T_5[7:0] ? image_2_217 : _GEN_720; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_722 = 8'hda == _T_5[7:0] ? image_2_218 : _GEN_721; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_723 = 8'hdb == _T_5[7:0] ? image_2_219 : _GEN_722; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_724 = 8'hdc == _T_5[7:0] ? image_2_220 : _GEN_723; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_725 = 8'hdd == _T_5[7:0] ? image_2_221 : _GEN_724; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_726 = 8'hde == _T_5[7:0] ? image_2_222 : _GEN_725; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_727 = 8'hdf == _T_5[7:0] ? image_2_223 : _GEN_726; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_728 = 8'he0 == _T_5[7:0] ? image_2_224 : _GEN_727; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_729 = 8'he1 == _T_5[7:0] ? image_2_225 : _GEN_728; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_730 = 8'he2 == _T_5[7:0] ? image_2_226 : _GEN_729; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_731 = 8'he3 == _T_5[7:0] ? image_2_227 : _GEN_730; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_732 = 8'he4 == _T_5[7:0] ? image_2_228 : _GEN_731; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_733 = 8'he5 == _T_5[7:0] ? image_2_229 : _GEN_732; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_734 = 8'he6 == _T_5[7:0] ? image_2_230 : _GEN_733; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_735 = 8'he7 == _T_5[7:0] ? image_2_231 : _GEN_734; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_736 = 8'he8 == _T_5[7:0] ? image_2_232 : _GEN_735; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_737 = 8'he9 == _T_5[7:0] ? image_2_233 : _GEN_736; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_738 = 8'hea == _T_5[7:0] ? image_2_234 : _GEN_737; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_739 = 8'heb == _T_5[7:0] ? image_2_235 : _GEN_738; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_740 = 8'hec == _T_5[7:0] ? image_2_236 : _GEN_739; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_741 = 8'hed == _T_5[7:0] ? image_2_237 : _GEN_740; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_742 = 8'hee == _T_5[7:0] ? image_2_238 : _GEN_741; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_743 = 8'hef == _T_5[7:0] ? image_2_239 : _GEN_742; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_744 = 8'hf0 == _T_5[7:0] ? image_2_240 : _GEN_743; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_745 = 8'hf1 == _T_5[7:0] ? image_2_241 : _GEN_744; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_746 = 8'hf2 == _T_5[7:0] ? image_2_242 : _GEN_745; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_747 = 8'hf3 == _T_5[7:0] ? image_2_243 : _GEN_746; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_748 = 8'hf4 == _T_5[7:0] ? image_2_244 : _GEN_747; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_749 = 8'hf5 == _T_5[7:0] ? image_2_245 : _GEN_748; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_750 = 8'hf6 == _T_5[7:0] ? image_2_246 : _GEN_749; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_751 = 8'hf7 == _T_5[7:0] ? image_2_247 : _GEN_750; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_752 = 8'hf8 == _T_5[7:0] ? image_2_248 : _GEN_751; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_753 = 8'hf9 == _T_5[7:0] ? image_2_249 : _GEN_752; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_754 = 8'hfa == _T_5[7:0] ? image_2_250 : _GEN_753; // @[VideoBuffer.scala 27:30]
  wire [32:0] _T_15 = {{1'd0}, pixelIndex}; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_19 = pixelIndex + 32'h1; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_22 = pixelIndex + 32'h2; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_25 = pixelIndex + 32'h3; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_28 = pixelIndex + 32'h4; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_31 = pixelIndex + 32'h5; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_34 = pixelIndex + 32'h6; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_79 = pixelIndex + 32'h7; // @[VideoBuffer.scala 36:34]
  wire [8:0] _T_80 = 5'h15 * 5'hc; // @[VideoBuffer.scala 37:42]
  wire [31:0] _GEN_6809 = {{23'd0}, _T_80}; // @[VideoBuffer.scala 37:25]
  wire  _T_81 = pixelIndex == _GEN_6809; // @[VideoBuffer.scala 37:25]
  assign io_pixelVal_out_0 = 8'hfb == _T_5[7:0] ? image_0_251 : _GEN_250; // @[VideoBuffer.scala 27:30]
  assign io_pixelVal_out_1 = 8'hfb == _T_5[7:0] ? image_1_251 : _GEN_502; // @[VideoBuffer.scala 27:30]
  assign io_pixelVal_out_2 = 8'hfb == _T_5[7:0] ? image_2_251 : _GEN_754; // @[VideoBuffer.scala 27:30]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  image_0_0 = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  image_0_1 = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  image_0_2 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  image_0_3 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  image_0_4 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  image_0_5 = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  image_0_6 = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  image_0_7 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  image_0_8 = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  image_0_9 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  image_0_10 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  image_0_11 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  image_0_12 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  image_0_13 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  image_0_14 = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  image_0_15 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  image_0_16 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  image_0_17 = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  image_0_18 = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  image_0_19 = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  image_0_20 = _RAND_20[3:0];
  _RAND_21 = {1{`RANDOM}};
  image_0_21 = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  image_0_22 = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  image_0_23 = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  image_0_24 = _RAND_24[3:0];
  _RAND_25 = {1{`RANDOM}};
  image_0_25 = _RAND_25[3:0];
  _RAND_26 = {1{`RANDOM}};
  image_0_26 = _RAND_26[3:0];
  _RAND_27 = {1{`RANDOM}};
  image_0_27 = _RAND_27[3:0];
  _RAND_28 = {1{`RANDOM}};
  image_0_28 = _RAND_28[3:0];
  _RAND_29 = {1{`RANDOM}};
  image_0_29 = _RAND_29[3:0];
  _RAND_30 = {1{`RANDOM}};
  image_0_30 = _RAND_30[3:0];
  _RAND_31 = {1{`RANDOM}};
  image_0_31 = _RAND_31[3:0];
  _RAND_32 = {1{`RANDOM}};
  image_0_32 = _RAND_32[3:0];
  _RAND_33 = {1{`RANDOM}};
  image_0_33 = _RAND_33[3:0];
  _RAND_34 = {1{`RANDOM}};
  image_0_34 = _RAND_34[3:0];
  _RAND_35 = {1{`RANDOM}};
  image_0_35 = _RAND_35[3:0];
  _RAND_36 = {1{`RANDOM}};
  image_0_36 = _RAND_36[3:0];
  _RAND_37 = {1{`RANDOM}};
  image_0_37 = _RAND_37[3:0];
  _RAND_38 = {1{`RANDOM}};
  image_0_38 = _RAND_38[3:0];
  _RAND_39 = {1{`RANDOM}};
  image_0_39 = _RAND_39[3:0];
  _RAND_40 = {1{`RANDOM}};
  image_0_40 = _RAND_40[3:0];
  _RAND_41 = {1{`RANDOM}};
  image_0_41 = _RAND_41[3:0];
  _RAND_42 = {1{`RANDOM}};
  image_0_42 = _RAND_42[3:0];
  _RAND_43 = {1{`RANDOM}};
  image_0_43 = _RAND_43[3:0];
  _RAND_44 = {1{`RANDOM}};
  image_0_44 = _RAND_44[3:0];
  _RAND_45 = {1{`RANDOM}};
  image_0_45 = _RAND_45[3:0];
  _RAND_46 = {1{`RANDOM}};
  image_0_46 = _RAND_46[3:0];
  _RAND_47 = {1{`RANDOM}};
  image_0_47 = _RAND_47[3:0];
  _RAND_48 = {1{`RANDOM}};
  image_0_48 = _RAND_48[3:0];
  _RAND_49 = {1{`RANDOM}};
  image_0_49 = _RAND_49[3:0];
  _RAND_50 = {1{`RANDOM}};
  image_0_50 = _RAND_50[3:0];
  _RAND_51 = {1{`RANDOM}};
  image_0_51 = _RAND_51[3:0];
  _RAND_52 = {1{`RANDOM}};
  image_0_52 = _RAND_52[3:0];
  _RAND_53 = {1{`RANDOM}};
  image_0_53 = _RAND_53[3:0];
  _RAND_54 = {1{`RANDOM}};
  image_0_54 = _RAND_54[3:0];
  _RAND_55 = {1{`RANDOM}};
  image_0_55 = _RAND_55[3:0];
  _RAND_56 = {1{`RANDOM}};
  image_0_56 = _RAND_56[3:0];
  _RAND_57 = {1{`RANDOM}};
  image_0_57 = _RAND_57[3:0];
  _RAND_58 = {1{`RANDOM}};
  image_0_58 = _RAND_58[3:0];
  _RAND_59 = {1{`RANDOM}};
  image_0_59 = _RAND_59[3:0];
  _RAND_60 = {1{`RANDOM}};
  image_0_60 = _RAND_60[3:0];
  _RAND_61 = {1{`RANDOM}};
  image_0_61 = _RAND_61[3:0];
  _RAND_62 = {1{`RANDOM}};
  image_0_62 = _RAND_62[3:0];
  _RAND_63 = {1{`RANDOM}};
  image_0_63 = _RAND_63[3:0];
  _RAND_64 = {1{`RANDOM}};
  image_0_64 = _RAND_64[3:0];
  _RAND_65 = {1{`RANDOM}};
  image_0_65 = _RAND_65[3:0];
  _RAND_66 = {1{`RANDOM}};
  image_0_66 = _RAND_66[3:0];
  _RAND_67 = {1{`RANDOM}};
  image_0_67 = _RAND_67[3:0];
  _RAND_68 = {1{`RANDOM}};
  image_0_68 = _RAND_68[3:0];
  _RAND_69 = {1{`RANDOM}};
  image_0_69 = _RAND_69[3:0];
  _RAND_70 = {1{`RANDOM}};
  image_0_70 = _RAND_70[3:0];
  _RAND_71 = {1{`RANDOM}};
  image_0_71 = _RAND_71[3:0];
  _RAND_72 = {1{`RANDOM}};
  image_0_72 = _RAND_72[3:0];
  _RAND_73 = {1{`RANDOM}};
  image_0_73 = _RAND_73[3:0];
  _RAND_74 = {1{`RANDOM}};
  image_0_74 = _RAND_74[3:0];
  _RAND_75 = {1{`RANDOM}};
  image_0_75 = _RAND_75[3:0];
  _RAND_76 = {1{`RANDOM}};
  image_0_76 = _RAND_76[3:0];
  _RAND_77 = {1{`RANDOM}};
  image_0_77 = _RAND_77[3:0];
  _RAND_78 = {1{`RANDOM}};
  image_0_78 = _RAND_78[3:0];
  _RAND_79 = {1{`RANDOM}};
  image_0_79 = _RAND_79[3:0];
  _RAND_80 = {1{`RANDOM}};
  image_0_80 = _RAND_80[3:0];
  _RAND_81 = {1{`RANDOM}};
  image_0_81 = _RAND_81[3:0];
  _RAND_82 = {1{`RANDOM}};
  image_0_82 = _RAND_82[3:0];
  _RAND_83 = {1{`RANDOM}};
  image_0_83 = _RAND_83[3:0];
  _RAND_84 = {1{`RANDOM}};
  image_0_84 = _RAND_84[3:0];
  _RAND_85 = {1{`RANDOM}};
  image_0_85 = _RAND_85[3:0];
  _RAND_86 = {1{`RANDOM}};
  image_0_86 = _RAND_86[3:0];
  _RAND_87 = {1{`RANDOM}};
  image_0_87 = _RAND_87[3:0];
  _RAND_88 = {1{`RANDOM}};
  image_0_88 = _RAND_88[3:0];
  _RAND_89 = {1{`RANDOM}};
  image_0_89 = _RAND_89[3:0];
  _RAND_90 = {1{`RANDOM}};
  image_0_90 = _RAND_90[3:0];
  _RAND_91 = {1{`RANDOM}};
  image_0_91 = _RAND_91[3:0];
  _RAND_92 = {1{`RANDOM}};
  image_0_92 = _RAND_92[3:0];
  _RAND_93 = {1{`RANDOM}};
  image_0_93 = _RAND_93[3:0];
  _RAND_94 = {1{`RANDOM}};
  image_0_94 = _RAND_94[3:0];
  _RAND_95 = {1{`RANDOM}};
  image_0_95 = _RAND_95[3:0];
  _RAND_96 = {1{`RANDOM}};
  image_0_96 = _RAND_96[3:0];
  _RAND_97 = {1{`RANDOM}};
  image_0_97 = _RAND_97[3:0];
  _RAND_98 = {1{`RANDOM}};
  image_0_98 = _RAND_98[3:0];
  _RAND_99 = {1{`RANDOM}};
  image_0_99 = _RAND_99[3:0];
  _RAND_100 = {1{`RANDOM}};
  image_0_100 = _RAND_100[3:0];
  _RAND_101 = {1{`RANDOM}};
  image_0_101 = _RAND_101[3:0];
  _RAND_102 = {1{`RANDOM}};
  image_0_102 = _RAND_102[3:0];
  _RAND_103 = {1{`RANDOM}};
  image_0_103 = _RAND_103[3:0];
  _RAND_104 = {1{`RANDOM}};
  image_0_104 = _RAND_104[3:0];
  _RAND_105 = {1{`RANDOM}};
  image_0_105 = _RAND_105[3:0];
  _RAND_106 = {1{`RANDOM}};
  image_0_106 = _RAND_106[3:0];
  _RAND_107 = {1{`RANDOM}};
  image_0_107 = _RAND_107[3:0];
  _RAND_108 = {1{`RANDOM}};
  image_0_108 = _RAND_108[3:0];
  _RAND_109 = {1{`RANDOM}};
  image_0_109 = _RAND_109[3:0];
  _RAND_110 = {1{`RANDOM}};
  image_0_110 = _RAND_110[3:0];
  _RAND_111 = {1{`RANDOM}};
  image_0_111 = _RAND_111[3:0];
  _RAND_112 = {1{`RANDOM}};
  image_0_112 = _RAND_112[3:0];
  _RAND_113 = {1{`RANDOM}};
  image_0_113 = _RAND_113[3:0];
  _RAND_114 = {1{`RANDOM}};
  image_0_114 = _RAND_114[3:0];
  _RAND_115 = {1{`RANDOM}};
  image_0_115 = _RAND_115[3:0];
  _RAND_116 = {1{`RANDOM}};
  image_0_116 = _RAND_116[3:0];
  _RAND_117 = {1{`RANDOM}};
  image_0_117 = _RAND_117[3:0];
  _RAND_118 = {1{`RANDOM}};
  image_0_118 = _RAND_118[3:0];
  _RAND_119 = {1{`RANDOM}};
  image_0_119 = _RAND_119[3:0];
  _RAND_120 = {1{`RANDOM}};
  image_0_120 = _RAND_120[3:0];
  _RAND_121 = {1{`RANDOM}};
  image_0_121 = _RAND_121[3:0];
  _RAND_122 = {1{`RANDOM}};
  image_0_122 = _RAND_122[3:0];
  _RAND_123 = {1{`RANDOM}};
  image_0_123 = _RAND_123[3:0];
  _RAND_124 = {1{`RANDOM}};
  image_0_124 = _RAND_124[3:0];
  _RAND_125 = {1{`RANDOM}};
  image_0_125 = _RAND_125[3:0];
  _RAND_126 = {1{`RANDOM}};
  image_0_126 = _RAND_126[3:0];
  _RAND_127 = {1{`RANDOM}};
  image_0_127 = _RAND_127[3:0];
  _RAND_128 = {1{`RANDOM}};
  image_0_128 = _RAND_128[3:0];
  _RAND_129 = {1{`RANDOM}};
  image_0_129 = _RAND_129[3:0];
  _RAND_130 = {1{`RANDOM}};
  image_0_130 = _RAND_130[3:0];
  _RAND_131 = {1{`RANDOM}};
  image_0_131 = _RAND_131[3:0];
  _RAND_132 = {1{`RANDOM}};
  image_0_132 = _RAND_132[3:0];
  _RAND_133 = {1{`RANDOM}};
  image_0_133 = _RAND_133[3:0];
  _RAND_134 = {1{`RANDOM}};
  image_0_134 = _RAND_134[3:0];
  _RAND_135 = {1{`RANDOM}};
  image_0_135 = _RAND_135[3:0];
  _RAND_136 = {1{`RANDOM}};
  image_0_136 = _RAND_136[3:0];
  _RAND_137 = {1{`RANDOM}};
  image_0_137 = _RAND_137[3:0];
  _RAND_138 = {1{`RANDOM}};
  image_0_138 = _RAND_138[3:0];
  _RAND_139 = {1{`RANDOM}};
  image_0_139 = _RAND_139[3:0];
  _RAND_140 = {1{`RANDOM}};
  image_0_140 = _RAND_140[3:0];
  _RAND_141 = {1{`RANDOM}};
  image_0_141 = _RAND_141[3:0];
  _RAND_142 = {1{`RANDOM}};
  image_0_142 = _RAND_142[3:0];
  _RAND_143 = {1{`RANDOM}};
  image_0_143 = _RAND_143[3:0];
  _RAND_144 = {1{`RANDOM}};
  image_0_144 = _RAND_144[3:0];
  _RAND_145 = {1{`RANDOM}};
  image_0_145 = _RAND_145[3:0];
  _RAND_146 = {1{`RANDOM}};
  image_0_146 = _RAND_146[3:0];
  _RAND_147 = {1{`RANDOM}};
  image_0_147 = _RAND_147[3:0];
  _RAND_148 = {1{`RANDOM}};
  image_0_148 = _RAND_148[3:0];
  _RAND_149 = {1{`RANDOM}};
  image_0_149 = _RAND_149[3:0];
  _RAND_150 = {1{`RANDOM}};
  image_0_150 = _RAND_150[3:0];
  _RAND_151 = {1{`RANDOM}};
  image_0_151 = _RAND_151[3:0];
  _RAND_152 = {1{`RANDOM}};
  image_0_152 = _RAND_152[3:0];
  _RAND_153 = {1{`RANDOM}};
  image_0_153 = _RAND_153[3:0];
  _RAND_154 = {1{`RANDOM}};
  image_0_154 = _RAND_154[3:0];
  _RAND_155 = {1{`RANDOM}};
  image_0_155 = _RAND_155[3:0];
  _RAND_156 = {1{`RANDOM}};
  image_0_156 = _RAND_156[3:0];
  _RAND_157 = {1{`RANDOM}};
  image_0_157 = _RAND_157[3:0];
  _RAND_158 = {1{`RANDOM}};
  image_0_158 = _RAND_158[3:0];
  _RAND_159 = {1{`RANDOM}};
  image_0_159 = _RAND_159[3:0];
  _RAND_160 = {1{`RANDOM}};
  image_0_160 = _RAND_160[3:0];
  _RAND_161 = {1{`RANDOM}};
  image_0_161 = _RAND_161[3:0];
  _RAND_162 = {1{`RANDOM}};
  image_0_162 = _RAND_162[3:0];
  _RAND_163 = {1{`RANDOM}};
  image_0_163 = _RAND_163[3:0];
  _RAND_164 = {1{`RANDOM}};
  image_0_164 = _RAND_164[3:0];
  _RAND_165 = {1{`RANDOM}};
  image_0_165 = _RAND_165[3:0];
  _RAND_166 = {1{`RANDOM}};
  image_0_166 = _RAND_166[3:0];
  _RAND_167 = {1{`RANDOM}};
  image_0_167 = _RAND_167[3:0];
  _RAND_168 = {1{`RANDOM}};
  image_0_168 = _RAND_168[3:0];
  _RAND_169 = {1{`RANDOM}};
  image_0_169 = _RAND_169[3:0];
  _RAND_170 = {1{`RANDOM}};
  image_0_170 = _RAND_170[3:0];
  _RAND_171 = {1{`RANDOM}};
  image_0_171 = _RAND_171[3:0];
  _RAND_172 = {1{`RANDOM}};
  image_0_172 = _RAND_172[3:0];
  _RAND_173 = {1{`RANDOM}};
  image_0_173 = _RAND_173[3:0];
  _RAND_174 = {1{`RANDOM}};
  image_0_174 = _RAND_174[3:0];
  _RAND_175 = {1{`RANDOM}};
  image_0_175 = _RAND_175[3:0];
  _RAND_176 = {1{`RANDOM}};
  image_0_176 = _RAND_176[3:0];
  _RAND_177 = {1{`RANDOM}};
  image_0_177 = _RAND_177[3:0];
  _RAND_178 = {1{`RANDOM}};
  image_0_178 = _RAND_178[3:0];
  _RAND_179 = {1{`RANDOM}};
  image_0_179 = _RAND_179[3:0];
  _RAND_180 = {1{`RANDOM}};
  image_0_180 = _RAND_180[3:0];
  _RAND_181 = {1{`RANDOM}};
  image_0_181 = _RAND_181[3:0];
  _RAND_182 = {1{`RANDOM}};
  image_0_182 = _RAND_182[3:0];
  _RAND_183 = {1{`RANDOM}};
  image_0_183 = _RAND_183[3:0];
  _RAND_184 = {1{`RANDOM}};
  image_0_184 = _RAND_184[3:0];
  _RAND_185 = {1{`RANDOM}};
  image_0_185 = _RAND_185[3:0];
  _RAND_186 = {1{`RANDOM}};
  image_0_186 = _RAND_186[3:0];
  _RAND_187 = {1{`RANDOM}};
  image_0_187 = _RAND_187[3:0];
  _RAND_188 = {1{`RANDOM}};
  image_0_188 = _RAND_188[3:0];
  _RAND_189 = {1{`RANDOM}};
  image_0_189 = _RAND_189[3:0];
  _RAND_190 = {1{`RANDOM}};
  image_0_190 = _RAND_190[3:0];
  _RAND_191 = {1{`RANDOM}};
  image_0_191 = _RAND_191[3:0];
  _RAND_192 = {1{`RANDOM}};
  image_0_192 = _RAND_192[3:0];
  _RAND_193 = {1{`RANDOM}};
  image_0_193 = _RAND_193[3:0];
  _RAND_194 = {1{`RANDOM}};
  image_0_194 = _RAND_194[3:0];
  _RAND_195 = {1{`RANDOM}};
  image_0_195 = _RAND_195[3:0];
  _RAND_196 = {1{`RANDOM}};
  image_0_196 = _RAND_196[3:0];
  _RAND_197 = {1{`RANDOM}};
  image_0_197 = _RAND_197[3:0];
  _RAND_198 = {1{`RANDOM}};
  image_0_198 = _RAND_198[3:0];
  _RAND_199 = {1{`RANDOM}};
  image_0_199 = _RAND_199[3:0];
  _RAND_200 = {1{`RANDOM}};
  image_0_200 = _RAND_200[3:0];
  _RAND_201 = {1{`RANDOM}};
  image_0_201 = _RAND_201[3:0];
  _RAND_202 = {1{`RANDOM}};
  image_0_202 = _RAND_202[3:0];
  _RAND_203 = {1{`RANDOM}};
  image_0_203 = _RAND_203[3:0];
  _RAND_204 = {1{`RANDOM}};
  image_0_204 = _RAND_204[3:0];
  _RAND_205 = {1{`RANDOM}};
  image_0_205 = _RAND_205[3:0];
  _RAND_206 = {1{`RANDOM}};
  image_0_206 = _RAND_206[3:0];
  _RAND_207 = {1{`RANDOM}};
  image_0_207 = _RAND_207[3:0];
  _RAND_208 = {1{`RANDOM}};
  image_0_208 = _RAND_208[3:0];
  _RAND_209 = {1{`RANDOM}};
  image_0_209 = _RAND_209[3:0];
  _RAND_210 = {1{`RANDOM}};
  image_0_210 = _RAND_210[3:0];
  _RAND_211 = {1{`RANDOM}};
  image_0_211 = _RAND_211[3:0];
  _RAND_212 = {1{`RANDOM}};
  image_0_212 = _RAND_212[3:0];
  _RAND_213 = {1{`RANDOM}};
  image_0_213 = _RAND_213[3:0];
  _RAND_214 = {1{`RANDOM}};
  image_0_214 = _RAND_214[3:0];
  _RAND_215 = {1{`RANDOM}};
  image_0_215 = _RAND_215[3:0];
  _RAND_216 = {1{`RANDOM}};
  image_0_216 = _RAND_216[3:0];
  _RAND_217 = {1{`RANDOM}};
  image_0_217 = _RAND_217[3:0];
  _RAND_218 = {1{`RANDOM}};
  image_0_218 = _RAND_218[3:0];
  _RAND_219 = {1{`RANDOM}};
  image_0_219 = _RAND_219[3:0];
  _RAND_220 = {1{`RANDOM}};
  image_0_220 = _RAND_220[3:0];
  _RAND_221 = {1{`RANDOM}};
  image_0_221 = _RAND_221[3:0];
  _RAND_222 = {1{`RANDOM}};
  image_0_222 = _RAND_222[3:0];
  _RAND_223 = {1{`RANDOM}};
  image_0_223 = _RAND_223[3:0];
  _RAND_224 = {1{`RANDOM}};
  image_0_224 = _RAND_224[3:0];
  _RAND_225 = {1{`RANDOM}};
  image_0_225 = _RAND_225[3:0];
  _RAND_226 = {1{`RANDOM}};
  image_0_226 = _RAND_226[3:0];
  _RAND_227 = {1{`RANDOM}};
  image_0_227 = _RAND_227[3:0];
  _RAND_228 = {1{`RANDOM}};
  image_0_228 = _RAND_228[3:0];
  _RAND_229 = {1{`RANDOM}};
  image_0_229 = _RAND_229[3:0];
  _RAND_230 = {1{`RANDOM}};
  image_0_230 = _RAND_230[3:0];
  _RAND_231 = {1{`RANDOM}};
  image_0_231 = _RAND_231[3:0];
  _RAND_232 = {1{`RANDOM}};
  image_0_232 = _RAND_232[3:0];
  _RAND_233 = {1{`RANDOM}};
  image_0_233 = _RAND_233[3:0];
  _RAND_234 = {1{`RANDOM}};
  image_0_234 = _RAND_234[3:0];
  _RAND_235 = {1{`RANDOM}};
  image_0_235 = _RAND_235[3:0];
  _RAND_236 = {1{`RANDOM}};
  image_0_236 = _RAND_236[3:0];
  _RAND_237 = {1{`RANDOM}};
  image_0_237 = _RAND_237[3:0];
  _RAND_238 = {1{`RANDOM}};
  image_0_238 = _RAND_238[3:0];
  _RAND_239 = {1{`RANDOM}};
  image_0_239 = _RAND_239[3:0];
  _RAND_240 = {1{`RANDOM}};
  image_0_240 = _RAND_240[3:0];
  _RAND_241 = {1{`RANDOM}};
  image_0_241 = _RAND_241[3:0];
  _RAND_242 = {1{`RANDOM}};
  image_0_242 = _RAND_242[3:0];
  _RAND_243 = {1{`RANDOM}};
  image_0_243 = _RAND_243[3:0];
  _RAND_244 = {1{`RANDOM}};
  image_0_244 = _RAND_244[3:0];
  _RAND_245 = {1{`RANDOM}};
  image_0_245 = _RAND_245[3:0];
  _RAND_246 = {1{`RANDOM}};
  image_0_246 = _RAND_246[3:0];
  _RAND_247 = {1{`RANDOM}};
  image_0_247 = _RAND_247[3:0];
  _RAND_248 = {1{`RANDOM}};
  image_0_248 = _RAND_248[3:0];
  _RAND_249 = {1{`RANDOM}};
  image_0_249 = _RAND_249[3:0];
  _RAND_250 = {1{`RANDOM}};
  image_0_250 = _RAND_250[3:0];
  _RAND_251 = {1{`RANDOM}};
  image_0_251 = _RAND_251[3:0];
  _RAND_252 = {1{`RANDOM}};
  image_1_0 = _RAND_252[3:0];
  _RAND_253 = {1{`RANDOM}};
  image_1_1 = _RAND_253[3:0];
  _RAND_254 = {1{`RANDOM}};
  image_1_2 = _RAND_254[3:0];
  _RAND_255 = {1{`RANDOM}};
  image_1_3 = _RAND_255[3:0];
  _RAND_256 = {1{`RANDOM}};
  image_1_4 = _RAND_256[3:0];
  _RAND_257 = {1{`RANDOM}};
  image_1_5 = _RAND_257[3:0];
  _RAND_258 = {1{`RANDOM}};
  image_1_6 = _RAND_258[3:0];
  _RAND_259 = {1{`RANDOM}};
  image_1_7 = _RAND_259[3:0];
  _RAND_260 = {1{`RANDOM}};
  image_1_8 = _RAND_260[3:0];
  _RAND_261 = {1{`RANDOM}};
  image_1_9 = _RAND_261[3:0];
  _RAND_262 = {1{`RANDOM}};
  image_1_10 = _RAND_262[3:0];
  _RAND_263 = {1{`RANDOM}};
  image_1_11 = _RAND_263[3:0];
  _RAND_264 = {1{`RANDOM}};
  image_1_12 = _RAND_264[3:0];
  _RAND_265 = {1{`RANDOM}};
  image_1_13 = _RAND_265[3:0];
  _RAND_266 = {1{`RANDOM}};
  image_1_14 = _RAND_266[3:0];
  _RAND_267 = {1{`RANDOM}};
  image_1_15 = _RAND_267[3:0];
  _RAND_268 = {1{`RANDOM}};
  image_1_16 = _RAND_268[3:0];
  _RAND_269 = {1{`RANDOM}};
  image_1_17 = _RAND_269[3:0];
  _RAND_270 = {1{`RANDOM}};
  image_1_18 = _RAND_270[3:0];
  _RAND_271 = {1{`RANDOM}};
  image_1_19 = _RAND_271[3:0];
  _RAND_272 = {1{`RANDOM}};
  image_1_20 = _RAND_272[3:0];
  _RAND_273 = {1{`RANDOM}};
  image_1_21 = _RAND_273[3:0];
  _RAND_274 = {1{`RANDOM}};
  image_1_22 = _RAND_274[3:0];
  _RAND_275 = {1{`RANDOM}};
  image_1_23 = _RAND_275[3:0];
  _RAND_276 = {1{`RANDOM}};
  image_1_24 = _RAND_276[3:0];
  _RAND_277 = {1{`RANDOM}};
  image_1_25 = _RAND_277[3:0];
  _RAND_278 = {1{`RANDOM}};
  image_1_26 = _RAND_278[3:0];
  _RAND_279 = {1{`RANDOM}};
  image_1_27 = _RAND_279[3:0];
  _RAND_280 = {1{`RANDOM}};
  image_1_28 = _RAND_280[3:0];
  _RAND_281 = {1{`RANDOM}};
  image_1_29 = _RAND_281[3:0];
  _RAND_282 = {1{`RANDOM}};
  image_1_30 = _RAND_282[3:0];
  _RAND_283 = {1{`RANDOM}};
  image_1_31 = _RAND_283[3:0];
  _RAND_284 = {1{`RANDOM}};
  image_1_32 = _RAND_284[3:0];
  _RAND_285 = {1{`RANDOM}};
  image_1_33 = _RAND_285[3:0];
  _RAND_286 = {1{`RANDOM}};
  image_1_34 = _RAND_286[3:0];
  _RAND_287 = {1{`RANDOM}};
  image_1_35 = _RAND_287[3:0];
  _RAND_288 = {1{`RANDOM}};
  image_1_36 = _RAND_288[3:0];
  _RAND_289 = {1{`RANDOM}};
  image_1_37 = _RAND_289[3:0];
  _RAND_290 = {1{`RANDOM}};
  image_1_38 = _RAND_290[3:0];
  _RAND_291 = {1{`RANDOM}};
  image_1_39 = _RAND_291[3:0];
  _RAND_292 = {1{`RANDOM}};
  image_1_40 = _RAND_292[3:0];
  _RAND_293 = {1{`RANDOM}};
  image_1_41 = _RAND_293[3:0];
  _RAND_294 = {1{`RANDOM}};
  image_1_42 = _RAND_294[3:0];
  _RAND_295 = {1{`RANDOM}};
  image_1_43 = _RAND_295[3:0];
  _RAND_296 = {1{`RANDOM}};
  image_1_44 = _RAND_296[3:0];
  _RAND_297 = {1{`RANDOM}};
  image_1_45 = _RAND_297[3:0];
  _RAND_298 = {1{`RANDOM}};
  image_1_46 = _RAND_298[3:0];
  _RAND_299 = {1{`RANDOM}};
  image_1_47 = _RAND_299[3:0];
  _RAND_300 = {1{`RANDOM}};
  image_1_48 = _RAND_300[3:0];
  _RAND_301 = {1{`RANDOM}};
  image_1_49 = _RAND_301[3:0];
  _RAND_302 = {1{`RANDOM}};
  image_1_50 = _RAND_302[3:0];
  _RAND_303 = {1{`RANDOM}};
  image_1_51 = _RAND_303[3:0];
  _RAND_304 = {1{`RANDOM}};
  image_1_52 = _RAND_304[3:0];
  _RAND_305 = {1{`RANDOM}};
  image_1_53 = _RAND_305[3:0];
  _RAND_306 = {1{`RANDOM}};
  image_1_54 = _RAND_306[3:0];
  _RAND_307 = {1{`RANDOM}};
  image_1_55 = _RAND_307[3:0];
  _RAND_308 = {1{`RANDOM}};
  image_1_56 = _RAND_308[3:0];
  _RAND_309 = {1{`RANDOM}};
  image_1_57 = _RAND_309[3:0];
  _RAND_310 = {1{`RANDOM}};
  image_1_58 = _RAND_310[3:0];
  _RAND_311 = {1{`RANDOM}};
  image_1_59 = _RAND_311[3:0];
  _RAND_312 = {1{`RANDOM}};
  image_1_60 = _RAND_312[3:0];
  _RAND_313 = {1{`RANDOM}};
  image_1_61 = _RAND_313[3:0];
  _RAND_314 = {1{`RANDOM}};
  image_1_62 = _RAND_314[3:0];
  _RAND_315 = {1{`RANDOM}};
  image_1_63 = _RAND_315[3:0];
  _RAND_316 = {1{`RANDOM}};
  image_1_64 = _RAND_316[3:0];
  _RAND_317 = {1{`RANDOM}};
  image_1_65 = _RAND_317[3:0];
  _RAND_318 = {1{`RANDOM}};
  image_1_66 = _RAND_318[3:0];
  _RAND_319 = {1{`RANDOM}};
  image_1_67 = _RAND_319[3:0];
  _RAND_320 = {1{`RANDOM}};
  image_1_68 = _RAND_320[3:0];
  _RAND_321 = {1{`RANDOM}};
  image_1_69 = _RAND_321[3:0];
  _RAND_322 = {1{`RANDOM}};
  image_1_70 = _RAND_322[3:0];
  _RAND_323 = {1{`RANDOM}};
  image_1_71 = _RAND_323[3:0];
  _RAND_324 = {1{`RANDOM}};
  image_1_72 = _RAND_324[3:0];
  _RAND_325 = {1{`RANDOM}};
  image_1_73 = _RAND_325[3:0];
  _RAND_326 = {1{`RANDOM}};
  image_1_74 = _RAND_326[3:0];
  _RAND_327 = {1{`RANDOM}};
  image_1_75 = _RAND_327[3:0];
  _RAND_328 = {1{`RANDOM}};
  image_1_76 = _RAND_328[3:0];
  _RAND_329 = {1{`RANDOM}};
  image_1_77 = _RAND_329[3:0];
  _RAND_330 = {1{`RANDOM}};
  image_1_78 = _RAND_330[3:0];
  _RAND_331 = {1{`RANDOM}};
  image_1_79 = _RAND_331[3:0];
  _RAND_332 = {1{`RANDOM}};
  image_1_80 = _RAND_332[3:0];
  _RAND_333 = {1{`RANDOM}};
  image_1_81 = _RAND_333[3:0];
  _RAND_334 = {1{`RANDOM}};
  image_1_82 = _RAND_334[3:0];
  _RAND_335 = {1{`RANDOM}};
  image_1_83 = _RAND_335[3:0];
  _RAND_336 = {1{`RANDOM}};
  image_1_84 = _RAND_336[3:0];
  _RAND_337 = {1{`RANDOM}};
  image_1_85 = _RAND_337[3:0];
  _RAND_338 = {1{`RANDOM}};
  image_1_86 = _RAND_338[3:0];
  _RAND_339 = {1{`RANDOM}};
  image_1_87 = _RAND_339[3:0];
  _RAND_340 = {1{`RANDOM}};
  image_1_88 = _RAND_340[3:0];
  _RAND_341 = {1{`RANDOM}};
  image_1_89 = _RAND_341[3:0];
  _RAND_342 = {1{`RANDOM}};
  image_1_90 = _RAND_342[3:0];
  _RAND_343 = {1{`RANDOM}};
  image_1_91 = _RAND_343[3:0];
  _RAND_344 = {1{`RANDOM}};
  image_1_92 = _RAND_344[3:0];
  _RAND_345 = {1{`RANDOM}};
  image_1_93 = _RAND_345[3:0];
  _RAND_346 = {1{`RANDOM}};
  image_1_94 = _RAND_346[3:0];
  _RAND_347 = {1{`RANDOM}};
  image_1_95 = _RAND_347[3:0];
  _RAND_348 = {1{`RANDOM}};
  image_1_96 = _RAND_348[3:0];
  _RAND_349 = {1{`RANDOM}};
  image_1_97 = _RAND_349[3:0];
  _RAND_350 = {1{`RANDOM}};
  image_1_98 = _RAND_350[3:0];
  _RAND_351 = {1{`RANDOM}};
  image_1_99 = _RAND_351[3:0];
  _RAND_352 = {1{`RANDOM}};
  image_1_100 = _RAND_352[3:0];
  _RAND_353 = {1{`RANDOM}};
  image_1_101 = _RAND_353[3:0];
  _RAND_354 = {1{`RANDOM}};
  image_1_102 = _RAND_354[3:0];
  _RAND_355 = {1{`RANDOM}};
  image_1_103 = _RAND_355[3:0];
  _RAND_356 = {1{`RANDOM}};
  image_1_104 = _RAND_356[3:0];
  _RAND_357 = {1{`RANDOM}};
  image_1_105 = _RAND_357[3:0];
  _RAND_358 = {1{`RANDOM}};
  image_1_106 = _RAND_358[3:0];
  _RAND_359 = {1{`RANDOM}};
  image_1_107 = _RAND_359[3:0];
  _RAND_360 = {1{`RANDOM}};
  image_1_108 = _RAND_360[3:0];
  _RAND_361 = {1{`RANDOM}};
  image_1_109 = _RAND_361[3:0];
  _RAND_362 = {1{`RANDOM}};
  image_1_110 = _RAND_362[3:0];
  _RAND_363 = {1{`RANDOM}};
  image_1_111 = _RAND_363[3:0];
  _RAND_364 = {1{`RANDOM}};
  image_1_112 = _RAND_364[3:0];
  _RAND_365 = {1{`RANDOM}};
  image_1_113 = _RAND_365[3:0];
  _RAND_366 = {1{`RANDOM}};
  image_1_114 = _RAND_366[3:0];
  _RAND_367 = {1{`RANDOM}};
  image_1_115 = _RAND_367[3:0];
  _RAND_368 = {1{`RANDOM}};
  image_1_116 = _RAND_368[3:0];
  _RAND_369 = {1{`RANDOM}};
  image_1_117 = _RAND_369[3:0];
  _RAND_370 = {1{`RANDOM}};
  image_1_118 = _RAND_370[3:0];
  _RAND_371 = {1{`RANDOM}};
  image_1_119 = _RAND_371[3:0];
  _RAND_372 = {1{`RANDOM}};
  image_1_120 = _RAND_372[3:0];
  _RAND_373 = {1{`RANDOM}};
  image_1_121 = _RAND_373[3:0];
  _RAND_374 = {1{`RANDOM}};
  image_1_122 = _RAND_374[3:0];
  _RAND_375 = {1{`RANDOM}};
  image_1_123 = _RAND_375[3:0];
  _RAND_376 = {1{`RANDOM}};
  image_1_124 = _RAND_376[3:0];
  _RAND_377 = {1{`RANDOM}};
  image_1_125 = _RAND_377[3:0];
  _RAND_378 = {1{`RANDOM}};
  image_1_126 = _RAND_378[3:0];
  _RAND_379 = {1{`RANDOM}};
  image_1_127 = _RAND_379[3:0];
  _RAND_380 = {1{`RANDOM}};
  image_1_128 = _RAND_380[3:0];
  _RAND_381 = {1{`RANDOM}};
  image_1_129 = _RAND_381[3:0];
  _RAND_382 = {1{`RANDOM}};
  image_1_130 = _RAND_382[3:0];
  _RAND_383 = {1{`RANDOM}};
  image_1_131 = _RAND_383[3:0];
  _RAND_384 = {1{`RANDOM}};
  image_1_132 = _RAND_384[3:0];
  _RAND_385 = {1{`RANDOM}};
  image_1_133 = _RAND_385[3:0];
  _RAND_386 = {1{`RANDOM}};
  image_1_134 = _RAND_386[3:0];
  _RAND_387 = {1{`RANDOM}};
  image_1_135 = _RAND_387[3:0];
  _RAND_388 = {1{`RANDOM}};
  image_1_136 = _RAND_388[3:0];
  _RAND_389 = {1{`RANDOM}};
  image_1_137 = _RAND_389[3:0];
  _RAND_390 = {1{`RANDOM}};
  image_1_138 = _RAND_390[3:0];
  _RAND_391 = {1{`RANDOM}};
  image_1_139 = _RAND_391[3:0];
  _RAND_392 = {1{`RANDOM}};
  image_1_140 = _RAND_392[3:0];
  _RAND_393 = {1{`RANDOM}};
  image_1_141 = _RAND_393[3:0];
  _RAND_394 = {1{`RANDOM}};
  image_1_142 = _RAND_394[3:0];
  _RAND_395 = {1{`RANDOM}};
  image_1_143 = _RAND_395[3:0];
  _RAND_396 = {1{`RANDOM}};
  image_1_144 = _RAND_396[3:0];
  _RAND_397 = {1{`RANDOM}};
  image_1_145 = _RAND_397[3:0];
  _RAND_398 = {1{`RANDOM}};
  image_1_146 = _RAND_398[3:0];
  _RAND_399 = {1{`RANDOM}};
  image_1_147 = _RAND_399[3:0];
  _RAND_400 = {1{`RANDOM}};
  image_1_148 = _RAND_400[3:0];
  _RAND_401 = {1{`RANDOM}};
  image_1_149 = _RAND_401[3:0];
  _RAND_402 = {1{`RANDOM}};
  image_1_150 = _RAND_402[3:0];
  _RAND_403 = {1{`RANDOM}};
  image_1_151 = _RAND_403[3:0];
  _RAND_404 = {1{`RANDOM}};
  image_1_152 = _RAND_404[3:0];
  _RAND_405 = {1{`RANDOM}};
  image_1_153 = _RAND_405[3:0];
  _RAND_406 = {1{`RANDOM}};
  image_1_154 = _RAND_406[3:0];
  _RAND_407 = {1{`RANDOM}};
  image_1_155 = _RAND_407[3:0];
  _RAND_408 = {1{`RANDOM}};
  image_1_156 = _RAND_408[3:0];
  _RAND_409 = {1{`RANDOM}};
  image_1_157 = _RAND_409[3:0];
  _RAND_410 = {1{`RANDOM}};
  image_1_158 = _RAND_410[3:0];
  _RAND_411 = {1{`RANDOM}};
  image_1_159 = _RAND_411[3:0];
  _RAND_412 = {1{`RANDOM}};
  image_1_160 = _RAND_412[3:0];
  _RAND_413 = {1{`RANDOM}};
  image_1_161 = _RAND_413[3:0];
  _RAND_414 = {1{`RANDOM}};
  image_1_162 = _RAND_414[3:0];
  _RAND_415 = {1{`RANDOM}};
  image_1_163 = _RAND_415[3:0];
  _RAND_416 = {1{`RANDOM}};
  image_1_164 = _RAND_416[3:0];
  _RAND_417 = {1{`RANDOM}};
  image_1_165 = _RAND_417[3:0];
  _RAND_418 = {1{`RANDOM}};
  image_1_166 = _RAND_418[3:0];
  _RAND_419 = {1{`RANDOM}};
  image_1_167 = _RAND_419[3:0];
  _RAND_420 = {1{`RANDOM}};
  image_1_168 = _RAND_420[3:0];
  _RAND_421 = {1{`RANDOM}};
  image_1_169 = _RAND_421[3:0];
  _RAND_422 = {1{`RANDOM}};
  image_1_170 = _RAND_422[3:0];
  _RAND_423 = {1{`RANDOM}};
  image_1_171 = _RAND_423[3:0];
  _RAND_424 = {1{`RANDOM}};
  image_1_172 = _RAND_424[3:0];
  _RAND_425 = {1{`RANDOM}};
  image_1_173 = _RAND_425[3:0];
  _RAND_426 = {1{`RANDOM}};
  image_1_174 = _RAND_426[3:0];
  _RAND_427 = {1{`RANDOM}};
  image_1_175 = _RAND_427[3:0];
  _RAND_428 = {1{`RANDOM}};
  image_1_176 = _RAND_428[3:0];
  _RAND_429 = {1{`RANDOM}};
  image_1_177 = _RAND_429[3:0];
  _RAND_430 = {1{`RANDOM}};
  image_1_178 = _RAND_430[3:0];
  _RAND_431 = {1{`RANDOM}};
  image_1_179 = _RAND_431[3:0];
  _RAND_432 = {1{`RANDOM}};
  image_1_180 = _RAND_432[3:0];
  _RAND_433 = {1{`RANDOM}};
  image_1_181 = _RAND_433[3:0];
  _RAND_434 = {1{`RANDOM}};
  image_1_182 = _RAND_434[3:0];
  _RAND_435 = {1{`RANDOM}};
  image_1_183 = _RAND_435[3:0];
  _RAND_436 = {1{`RANDOM}};
  image_1_184 = _RAND_436[3:0];
  _RAND_437 = {1{`RANDOM}};
  image_1_185 = _RAND_437[3:0];
  _RAND_438 = {1{`RANDOM}};
  image_1_186 = _RAND_438[3:0];
  _RAND_439 = {1{`RANDOM}};
  image_1_187 = _RAND_439[3:0];
  _RAND_440 = {1{`RANDOM}};
  image_1_188 = _RAND_440[3:0];
  _RAND_441 = {1{`RANDOM}};
  image_1_189 = _RAND_441[3:0];
  _RAND_442 = {1{`RANDOM}};
  image_1_190 = _RAND_442[3:0];
  _RAND_443 = {1{`RANDOM}};
  image_1_191 = _RAND_443[3:0];
  _RAND_444 = {1{`RANDOM}};
  image_1_192 = _RAND_444[3:0];
  _RAND_445 = {1{`RANDOM}};
  image_1_193 = _RAND_445[3:0];
  _RAND_446 = {1{`RANDOM}};
  image_1_194 = _RAND_446[3:0];
  _RAND_447 = {1{`RANDOM}};
  image_1_195 = _RAND_447[3:0];
  _RAND_448 = {1{`RANDOM}};
  image_1_196 = _RAND_448[3:0];
  _RAND_449 = {1{`RANDOM}};
  image_1_197 = _RAND_449[3:0];
  _RAND_450 = {1{`RANDOM}};
  image_1_198 = _RAND_450[3:0];
  _RAND_451 = {1{`RANDOM}};
  image_1_199 = _RAND_451[3:0];
  _RAND_452 = {1{`RANDOM}};
  image_1_200 = _RAND_452[3:0];
  _RAND_453 = {1{`RANDOM}};
  image_1_201 = _RAND_453[3:0];
  _RAND_454 = {1{`RANDOM}};
  image_1_202 = _RAND_454[3:0];
  _RAND_455 = {1{`RANDOM}};
  image_1_203 = _RAND_455[3:0];
  _RAND_456 = {1{`RANDOM}};
  image_1_204 = _RAND_456[3:0];
  _RAND_457 = {1{`RANDOM}};
  image_1_205 = _RAND_457[3:0];
  _RAND_458 = {1{`RANDOM}};
  image_1_206 = _RAND_458[3:0];
  _RAND_459 = {1{`RANDOM}};
  image_1_207 = _RAND_459[3:0];
  _RAND_460 = {1{`RANDOM}};
  image_1_208 = _RAND_460[3:0];
  _RAND_461 = {1{`RANDOM}};
  image_1_209 = _RAND_461[3:0];
  _RAND_462 = {1{`RANDOM}};
  image_1_210 = _RAND_462[3:0];
  _RAND_463 = {1{`RANDOM}};
  image_1_211 = _RAND_463[3:0];
  _RAND_464 = {1{`RANDOM}};
  image_1_212 = _RAND_464[3:0];
  _RAND_465 = {1{`RANDOM}};
  image_1_213 = _RAND_465[3:0];
  _RAND_466 = {1{`RANDOM}};
  image_1_214 = _RAND_466[3:0];
  _RAND_467 = {1{`RANDOM}};
  image_1_215 = _RAND_467[3:0];
  _RAND_468 = {1{`RANDOM}};
  image_1_216 = _RAND_468[3:0];
  _RAND_469 = {1{`RANDOM}};
  image_1_217 = _RAND_469[3:0];
  _RAND_470 = {1{`RANDOM}};
  image_1_218 = _RAND_470[3:0];
  _RAND_471 = {1{`RANDOM}};
  image_1_219 = _RAND_471[3:0];
  _RAND_472 = {1{`RANDOM}};
  image_1_220 = _RAND_472[3:0];
  _RAND_473 = {1{`RANDOM}};
  image_1_221 = _RAND_473[3:0];
  _RAND_474 = {1{`RANDOM}};
  image_1_222 = _RAND_474[3:0];
  _RAND_475 = {1{`RANDOM}};
  image_1_223 = _RAND_475[3:0];
  _RAND_476 = {1{`RANDOM}};
  image_1_224 = _RAND_476[3:0];
  _RAND_477 = {1{`RANDOM}};
  image_1_225 = _RAND_477[3:0];
  _RAND_478 = {1{`RANDOM}};
  image_1_226 = _RAND_478[3:0];
  _RAND_479 = {1{`RANDOM}};
  image_1_227 = _RAND_479[3:0];
  _RAND_480 = {1{`RANDOM}};
  image_1_228 = _RAND_480[3:0];
  _RAND_481 = {1{`RANDOM}};
  image_1_229 = _RAND_481[3:0];
  _RAND_482 = {1{`RANDOM}};
  image_1_230 = _RAND_482[3:0];
  _RAND_483 = {1{`RANDOM}};
  image_1_231 = _RAND_483[3:0];
  _RAND_484 = {1{`RANDOM}};
  image_1_232 = _RAND_484[3:0];
  _RAND_485 = {1{`RANDOM}};
  image_1_233 = _RAND_485[3:0];
  _RAND_486 = {1{`RANDOM}};
  image_1_234 = _RAND_486[3:0];
  _RAND_487 = {1{`RANDOM}};
  image_1_235 = _RAND_487[3:0];
  _RAND_488 = {1{`RANDOM}};
  image_1_236 = _RAND_488[3:0];
  _RAND_489 = {1{`RANDOM}};
  image_1_237 = _RAND_489[3:0];
  _RAND_490 = {1{`RANDOM}};
  image_1_238 = _RAND_490[3:0];
  _RAND_491 = {1{`RANDOM}};
  image_1_239 = _RAND_491[3:0];
  _RAND_492 = {1{`RANDOM}};
  image_1_240 = _RAND_492[3:0];
  _RAND_493 = {1{`RANDOM}};
  image_1_241 = _RAND_493[3:0];
  _RAND_494 = {1{`RANDOM}};
  image_1_242 = _RAND_494[3:0];
  _RAND_495 = {1{`RANDOM}};
  image_1_243 = _RAND_495[3:0];
  _RAND_496 = {1{`RANDOM}};
  image_1_244 = _RAND_496[3:0];
  _RAND_497 = {1{`RANDOM}};
  image_1_245 = _RAND_497[3:0];
  _RAND_498 = {1{`RANDOM}};
  image_1_246 = _RAND_498[3:0];
  _RAND_499 = {1{`RANDOM}};
  image_1_247 = _RAND_499[3:0];
  _RAND_500 = {1{`RANDOM}};
  image_1_248 = _RAND_500[3:0];
  _RAND_501 = {1{`RANDOM}};
  image_1_249 = _RAND_501[3:0];
  _RAND_502 = {1{`RANDOM}};
  image_1_250 = _RAND_502[3:0];
  _RAND_503 = {1{`RANDOM}};
  image_1_251 = _RAND_503[3:0];
  _RAND_504 = {1{`RANDOM}};
  image_2_0 = _RAND_504[3:0];
  _RAND_505 = {1{`RANDOM}};
  image_2_1 = _RAND_505[3:0];
  _RAND_506 = {1{`RANDOM}};
  image_2_2 = _RAND_506[3:0];
  _RAND_507 = {1{`RANDOM}};
  image_2_3 = _RAND_507[3:0];
  _RAND_508 = {1{`RANDOM}};
  image_2_4 = _RAND_508[3:0];
  _RAND_509 = {1{`RANDOM}};
  image_2_5 = _RAND_509[3:0];
  _RAND_510 = {1{`RANDOM}};
  image_2_6 = _RAND_510[3:0];
  _RAND_511 = {1{`RANDOM}};
  image_2_7 = _RAND_511[3:0];
  _RAND_512 = {1{`RANDOM}};
  image_2_8 = _RAND_512[3:0];
  _RAND_513 = {1{`RANDOM}};
  image_2_9 = _RAND_513[3:0];
  _RAND_514 = {1{`RANDOM}};
  image_2_10 = _RAND_514[3:0];
  _RAND_515 = {1{`RANDOM}};
  image_2_11 = _RAND_515[3:0];
  _RAND_516 = {1{`RANDOM}};
  image_2_12 = _RAND_516[3:0];
  _RAND_517 = {1{`RANDOM}};
  image_2_13 = _RAND_517[3:0];
  _RAND_518 = {1{`RANDOM}};
  image_2_14 = _RAND_518[3:0];
  _RAND_519 = {1{`RANDOM}};
  image_2_15 = _RAND_519[3:0];
  _RAND_520 = {1{`RANDOM}};
  image_2_16 = _RAND_520[3:0];
  _RAND_521 = {1{`RANDOM}};
  image_2_17 = _RAND_521[3:0];
  _RAND_522 = {1{`RANDOM}};
  image_2_18 = _RAND_522[3:0];
  _RAND_523 = {1{`RANDOM}};
  image_2_19 = _RAND_523[3:0];
  _RAND_524 = {1{`RANDOM}};
  image_2_20 = _RAND_524[3:0];
  _RAND_525 = {1{`RANDOM}};
  image_2_21 = _RAND_525[3:0];
  _RAND_526 = {1{`RANDOM}};
  image_2_22 = _RAND_526[3:0];
  _RAND_527 = {1{`RANDOM}};
  image_2_23 = _RAND_527[3:0];
  _RAND_528 = {1{`RANDOM}};
  image_2_24 = _RAND_528[3:0];
  _RAND_529 = {1{`RANDOM}};
  image_2_25 = _RAND_529[3:0];
  _RAND_530 = {1{`RANDOM}};
  image_2_26 = _RAND_530[3:0];
  _RAND_531 = {1{`RANDOM}};
  image_2_27 = _RAND_531[3:0];
  _RAND_532 = {1{`RANDOM}};
  image_2_28 = _RAND_532[3:0];
  _RAND_533 = {1{`RANDOM}};
  image_2_29 = _RAND_533[3:0];
  _RAND_534 = {1{`RANDOM}};
  image_2_30 = _RAND_534[3:0];
  _RAND_535 = {1{`RANDOM}};
  image_2_31 = _RAND_535[3:0];
  _RAND_536 = {1{`RANDOM}};
  image_2_32 = _RAND_536[3:0];
  _RAND_537 = {1{`RANDOM}};
  image_2_33 = _RAND_537[3:0];
  _RAND_538 = {1{`RANDOM}};
  image_2_34 = _RAND_538[3:0];
  _RAND_539 = {1{`RANDOM}};
  image_2_35 = _RAND_539[3:0];
  _RAND_540 = {1{`RANDOM}};
  image_2_36 = _RAND_540[3:0];
  _RAND_541 = {1{`RANDOM}};
  image_2_37 = _RAND_541[3:0];
  _RAND_542 = {1{`RANDOM}};
  image_2_38 = _RAND_542[3:0];
  _RAND_543 = {1{`RANDOM}};
  image_2_39 = _RAND_543[3:0];
  _RAND_544 = {1{`RANDOM}};
  image_2_40 = _RAND_544[3:0];
  _RAND_545 = {1{`RANDOM}};
  image_2_41 = _RAND_545[3:0];
  _RAND_546 = {1{`RANDOM}};
  image_2_42 = _RAND_546[3:0];
  _RAND_547 = {1{`RANDOM}};
  image_2_43 = _RAND_547[3:0];
  _RAND_548 = {1{`RANDOM}};
  image_2_44 = _RAND_548[3:0];
  _RAND_549 = {1{`RANDOM}};
  image_2_45 = _RAND_549[3:0];
  _RAND_550 = {1{`RANDOM}};
  image_2_46 = _RAND_550[3:0];
  _RAND_551 = {1{`RANDOM}};
  image_2_47 = _RAND_551[3:0];
  _RAND_552 = {1{`RANDOM}};
  image_2_48 = _RAND_552[3:0];
  _RAND_553 = {1{`RANDOM}};
  image_2_49 = _RAND_553[3:0];
  _RAND_554 = {1{`RANDOM}};
  image_2_50 = _RAND_554[3:0];
  _RAND_555 = {1{`RANDOM}};
  image_2_51 = _RAND_555[3:0];
  _RAND_556 = {1{`RANDOM}};
  image_2_52 = _RAND_556[3:0];
  _RAND_557 = {1{`RANDOM}};
  image_2_53 = _RAND_557[3:0];
  _RAND_558 = {1{`RANDOM}};
  image_2_54 = _RAND_558[3:0];
  _RAND_559 = {1{`RANDOM}};
  image_2_55 = _RAND_559[3:0];
  _RAND_560 = {1{`RANDOM}};
  image_2_56 = _RAND_560[3:0];
  _RAND_561 = {1{`RANDOM}};
  image_2_57 = _RAND_561[3:0];
  _RAND_562 = {1{`RANDOM}};
  image_2_58 = _RAND_562[3:0];
  _RAND_563 = {1{`RANDOM}};
  image_2_59 = _RAND_563[3:0];
  _RAND_564 = {1{`RANDOM}};
  image_2_60 = _RAND_564[3:0];
  _RAND_565 = {1{`RANDOM}};
  image_2_61 = _RAND_565[3:0];
  _RAND_566 = {1{`RANDOM}};
  image_2_62 = _RAND_566[3:0];
  _RAND_567 = {1{`RANDOM}};
  image_2_63 = _RAND_567[3:0];
  _RAND_568 = {1{`RANDOM}};
  image_2_64 = _RAND_568[3:0];
  _RAND_569 = {1{`RANDOM}};
  image_2_65 = _RAND_569[3:0];
  _RAND_570 = {1{`RANDOM}};
  image_2_66 = _RAND_570[3:0];
  _RAND_571 = {1{`RANDOM}};
  image_2_67 = _RAND_571[3:0];
  _RAND_572 = {1{`RANDOM}};
  image_2_68 = _RAND_572[3:0];
  _RAND_573 = {1{`RANDOM}};
  image_2_69 = _RAND_573[3:0];
  _RAND_574 = {1{`RANDOM}};
  image_2_70 = _RAND_574[3:0];
  _RAND_575 = {1{`RANDOM}};
  image_2_71 = _RAND_575[3:0];
  _RAND_576 = {1{`RANDOM}};
  image_2_72 = _RAND_576[3:0];
  _RAND_577 = {1{`RANDOM}};
  image_2_73 = _RAND_577[3:0];
  _RAND_578 = {1{`RANDOM}};
  image_2_74 = _RAND_578[3:0];
  _RAND_579 = {1{`RANDOM}};
  image_2_75 = _RAND_579[3:0];
  _RAND_580 = {1{`RANDOM}};
  image_2_76 = _RAND_580[3:0];
  _RAND_581 = {1{`RANDOM}};
  image_2_77 = _RAND_581[3:0];
  _RAND_582 = {1{`RANDOM}};
  image_2_78 = _RAND_582[3:0];
  _RAND_583 = {1{`RANDOM}};
  image_2_79 = _RAND_583[3:0];
  _RAND_584 = {1{`RANDOM}};
  image_2_80 = _RAND_584[3:0];
  _RAND_585 = {1{`RANDOM}};
  image_2_81 = _RAND_585[3:0];
  _RAND_586 = {1{`RANDOM}};
  image_2_82 = _RAND_586[3:0];
  _RAND_587 = {1{`RANDOM}};
  image_2_83 = _RAND_587[3:0];
  _RAND_588 = {1{`RANDOM}};
  image_2_84 = _RAND_588[3:0];
  _RAND_589 = {1{`RANDOM}};
  image_2_85 = _RAND_589[3:0];
  _RAND_590 = {1{`RANDOM}};
  image_2_86 = _RAND_590[3:0];
  _RAND_591 = {1{`RANDOM}};
  image_2_87 = _RAND_591[3:0];
  _RAND_592 = {1{`RANDOM}};
  image_2_88 = _RAND_592[3:0];
  _RAND_593 = {1{`RANDOM}};
  image_2_89 = _RAND_593[3:0];
  _RAND_594 = {1{`RANDOM}};
  image_2_90 = _RAND_594[3:0];
  _RAND_595 = {1{`RANDOM}};
  image_2_91 = _RAND_595[3:0];
  _RAND_596 = {1{`RANDOM}};
  image_2_92 = _RAND_596[3:0];
  _RAND_597 = {1{`RANDOM}};
  image_2_93 = _RAND_597[3:0];
  _RAND_598 = {1{`RANDOM}};
  image_2_94 = _RAND_598[3:0];
  _RAND_599 = {1{`RANDOM}};
  image_2_95 = _RAND_599[3:0];
  _RAND_600 = {1{`RANDOM}};
  image_2_96 = _RAND_600[3:0];
  _RAND_601 = {1{`RANDOM}};
  image_2_97 = _RAND_601[3:0];
  _RAND_602 = {1{`RANDOM}};
  image_2_98 = _RAND_602[3:0];
  _RAND_603 = {1{`RANDOM}};
  image_2_99 = _RAND_603[3:0];
  _RAND_604 = {1{`RANDOM}};
  image_2_100 = _RAND_604[3:0];
  _RAND_605 = {1{`RANDOM}};
  image_2_101 = _RAND_605[3:0];
  _RAND_606 = {1{`RANDOM}};
  image_2_102 = _RAND_606[3:0];
  _RAND_607 = {1{`RANDOM}};
  image_2_103 = _RAND_607[3:0];
  _RAND_608 = {1{`RANDOM}};
  image_2_104 = _RAND_608[3:0];
  _RAND_609 = {1{`RANDOM}};
  image_2_105 = _RAND_609[3:0];
  _RAND_610 = {1{`RANDOM}};
  image_2_106 = _RAND_610[3:0];
  _RAND_611 = {1{`RANDOM}};
  image_2_107 = _RAND_611[3:0];
  _RAND_612 = {1{`RANDOM}};
  image_2_108 = _RAND_612[3:0];
  _RAND_613 = {1{`RANDOM}};
  image_2_109 = _RAND_613[3:0];
  _RAND_614 = {1{`RANDOM}};
  image_2_110 = _RAND_614[3:0];
  _RAND_615 = {1{`RANDOM}};
  image_2_111 = _RAND_615[3:0];
  _RAND_616 = {1{`RANDOM}};
  image_2_112 = _RAND_616[3:0];
  _RAND_617 = {1{`RANDOM}};
  image_2_113 = _RAND_617[3:0];
  _RAND_618 = {1{`RANDOM}};
  image_2_114 = _RAND_618[3:0];
  _RAND_619 = {1{`RANDOM}};
  image_2_115 = _RAND_619[3:0];
  _RAND_620 = {1{`RANDOM}};
  image_2_116 = _RAND_620[3:0];
  _RAND_621 = {1{`RANDOM}};
  image_2_117 = _RAND_621[3:0];
  _RAND_622 = {1{`RANDOM}};
  image_2_118 = _RAND_622[3:0];
  _RAND_623 = {1{`RANDOM}};
  image_2_119 = _RAND_623[3:0];
  _RAND_624 = {1{`RANDOM}};
  image_2_120 = _RAND_624[3:0];
  _RAND_625 = {1{`RANDOM}};
  image_2_121 = _RAND_625[3:0];
  _RAND_626 = {1{`RANDOM}};
  image_2_122 = _RAND_626[3:0];
  _RAND_627 = {1{`RANDOM}};
  image_2_123 = _RAND_627[3:0];
  _RAND_628 = {1{`RANDOM}};
  image_2_124 = _RAND_628[3:0];
  _RAND_629 = {1{`RANDOM}};
  image_2_125 = _RAND_629[3:0];
  _RAND_630 = {1{`RANDOM}};
  image_2_126 = _RAND_630[3:0];
  _RAND_631 = {1{`RANDOM}};
  image_2_127 = _RAND_631[3:0];
  _RAND_632 = {1{`RANDOM}};
  image_2_128 = _RAND_632[3:0];
  _RAND_633 = {1{`RANDOM}};
  image_2_129 = _RAND_633[3:0];
  _RAND_634 = {1{`RANDOM}};
  image_2_130 = _RAND_634[3:0];
  _RAND_635 = {1{`RANDOM}};
  image_2_131 = _RAND_635[3:0];
  _RAND_636 = {1{`RANDOM}};
  image_2_132 = _RAND_636[3:0];
  _RAND_637 = {1{`RANDOM}};
  image_2_133 = _RAND_637[3:0];
  _RAND_638 = {1{`RANDOM}};
  image_2_134 = _RAND_638[3:0];
  _RAND_639 = {1{`RANDOM}};
  image_2_135 = _RAND_639[3:0];
  _RAND_640 = {1{`RANDOM}};
  image_2_136 = _RAND_640[3:0];
  _RAND_641 = {1{`RANDOM}};
  image_2_137 = _RAND_641[3:0];
  _RAND_642 = {1{`RANDOM}};
  image_2_138 = _RAND_642[3:0];
  _RAND_643 = {1{`RANDOM}};
  image_2_139 = _RAND_643[3:0];
  _RAND_644 = {1{`RANDOM}};
  image_2_140 = _RAND_644[3:0];
  _RAND_645 = {1{`RANDOM}};
  image_2_141 = _RAND_645[3:0];
  _RAND_646 = {1{`RANDOM}};
  image_2_142 = _RAND_646[3:0];
  _RAND_647 = {1{`RANDOM}};
  image_2_143 = _RAND_647[3:0];
  _RAND_648 = {1{`RANDOM}};
  image_2_144 = _RAND_648[3:0];
  _RAND_649 = {1{`RANDOM}};
  image_2_145 = _RAND_649[3:0];
  _RAND_650 = {1{`RANDOM}};
  image_2_146 = _RAND_650[3:0];
  _RAND_651 = {1{`RANDOM}};
  image_2_147 = _RAND_651[3:0];
  _RAND_652 = {1{`RANDOM}};
  image_2_148 = _RAND_652[3:0];
  _RAND_653 = {1{`RANDOM}};
  image_2_149 = _RAND_653[3:0];
  _RAND_654 = {1{`RANDOM}};
  image_2_150 = _RAND_654[3:0];
  _RAND_655 = {1{`RANDOM}};
  image_2_151 = _RAND_655[3:0];
  _RAND_656 = {1{`RANDOM}};
  image_2_152 = _RAND_656[3:0];
  _RAND_657 = {1{`RANDOM}};
  image_2_153 = _RAND_657[3:0];
  _RAND_658 = {1{`RANDOM}};
  image_2_154 = _RAND_658[3:0];
  _RAND_659 = {1{`RANDOM}};
  image_2_155 = _RAND_659[3:0];
  _RAND_660 = {1{`RANDOM}};
  image_2_156 = _RAND_660[3:0];
  _RAND_661 = {1{`RANDOM}};
  image_2_157 = _RAND_661[3:0];
  _RAND_662 = {1{`RANDOM}};
  image_2_158 = _RAND_662[3:0];
  _RAND_663 = {1{`RANDOM}};
  image_2_159 = _RAND_663[3:0];
  _RAND_664 = {1{`RANDOM}};
  image_2_160 = _RAND_664[3:0];
  _RAND_665 = {1{`RANDOM}};
  image_2_161 = _RAND_665[3:0];
  _RAND_666 = {1{`RANDOM}};
  image_2_162 = _RAND_666[3:0];
  _RAND_667 = {1{`RANDOM}};
  image_2_163 = _RAND_667[3:0];
  _RAND_668 = {1{`RANDOM}};
  image_2_164 = _RAND_668[3:0];
  _RAND_669 = {1{`RANDOM}};
  image_2_165 = _RAND_669[3:0];
  _RAND_670 = {1{`RANDOM}};
  image_2_166 = _RAND_670[3:0];
  _RAND_671 = {1{`RANDOM}};
  image_2_167 = _RAND_671[3:0];
  _RAND_672 = {1{`RANDOM}};
  image_2_168 = _RAND_672[3:0];
  _RAND_673 = {1{`RANDOM}};
  image_2_169 = _RAND_673[3:0];
  _RAND_674 = {1{`RANDOM}};
  image_2_170 = _RAND_674[3:0];
  _RAND_675 = {1{`RANDOM}};
  image_2_171 = _RAND_675[3:0];
  _RAND_676 = {1{`RANDOM}};
  image_2_172 = _RAND_676[3:0];
  _RAND_677 = {1{`RANDOM}};
  image_2_173 = _RAND_677[3:0];
  _RAND_678 = {1{`RANDOM}};
  image_2_174 = _RAND_678[3:0];
  _RAND_679 = {1{`RANDOM}};
  image_2_175 = _RAND_679[3:0];
  _RAND_680 = {1{`RANDOM}};
  image_2_176 = _RAND_680[3:0];
  _RAND_681 = {1{`RANDOM}};
  image_2_177 = _RAND_681[3:0];
  _RAND_682 = {1{`RANDOM}};
  image_2_178 = _RAND_682[3:0];
  _RAND_683 = {1{`RANDOM}};
  image_2_179 = _RAND_683[3:0];
  _RAND_684 = {1{`RANDOM}};
  image_2_180 = _RAND_684[3:0];
  _RAND_685 = {1{`RANDOM}};
  image_2_181 = _RAND_685[3:0];
  _RAND_686 = {1{`RANDOM}};
  image_2_182 = _RAND_686[3:0];
  _RAND_687 = {1{`RANDOM}};
  image_2_183 = _RAND_687[3:0];
  _RAND_688 = {1{`RANDOM}};
  image_2_184 = _RAND_688[3:0];
  _RAND_689 = {1{`RANDOM}};
  image_2_185 = _RAND_689[3:0];
  _RAND_690 = {1{`RANDOM}};
  image_2_186 = _RAND_690[3:0];
  _RAND_691 = {1{`RANDOM}};
  image_2_187 = _RAND_691[3:0];
  _RAND_692 = {1{`RANDOM}};
  image_2_188 = _RAND_692[3:0];
  _RAND_693 = {1{`RANDOM}};
  image_2_189 = _RAND_693[3:0];
  _RAND_694 = {1{`RANDOM}};
  image_2_190 = _RAND_694[3:0];
  _RAND_695 = {1{`RANDOM}};
  image_2_191 = _RAND_695[3:0];
  _RAND_696 = {1{`RANDOM}};
  image_2_192 = _RAND_696[3:0];
  _RAND_697 = {1{`RANDOM}};
  image_2_193 = _RAND_697[3:0];
  _RAND_698 = {1{`RANDOM}};
  image_2_194 = _RAND_698[3:0];
  _RAND_699 = {1{`RANDOM}};
  image_2_195 = _RAND_699[3:0];
  _RAND_700 = {1{`RANDOM}};
  image_2_196 = _RAND_700[3:0];
  _RAND_701 = {1{`RANDOM}};
  image_2_197 = _RAND_701[3:0];
  _RAND_702 = {1{`RANDOM}};
  image_2_198 = _RAND_702[3:0];
  _RAND_703 = {1{`RANDOM}};
  image_2_199 = _RAND_703[3:0];
  _RAND_704 = {1{`RANDOM}};
  image_2_200 = _RAND_704[3:0];
  _RAND_705 = {1{`RANDOM}};
  image_2_201 = _RAND_705[3:0];
  _RAND_706 = {1{`RANDOM}};
  image_2_202 = _RAND_706[3:0];
  _RAND_707 = {1{`RANDOM}};
  image_2_203 = _RAND_707[3:0];
  _RAND_708 = {1{`RANDOM}};
  image_2_204 = _RAND_708[3:0];
  _RAND_709 = {1{`RANDOM}};
  image_2_205 = _RAND_709[3:0];
  _RAND_710 = {1{`RANDOM}};
  image_2_206 = _RAND_710[3:0];
  _RAND_711 = {1{`RANDOM}};
  image_2_207 = _RAND_711[3:0];
  _RAND_712 = {1{`RANDOM}};
  image_2_208 = _RAND_712[3:0];
  _RAND_713 = {1{`RANDOM}};
  image_2_209 = _RAND_713[3:0];
  _RAND_714 = {1{`RANDOM}};
  image_2_210 = _RAND_714[3:0];
  _RAND_715 = {1{`RANDOM}};
  image_2_211 = _RAND_715[3:0];
  _RAND_716 = {1{`RANDOM}};
  image_2_212 = _RAND_716[3:0];
  _RAND_717 = {1{`RANDOM}};
  image_2_213 = _RAND_717[3:0];
  _RAND_718 = {1{`RANDOM}};
  image_2_214 = _RAND_718[3:0];
  _RAND_719 = {1{`RANDOM}};
  image_2_215 = _RAND_719[3:0];
  _RAND_720 = {1{`RANDOM}};
  image_2_216 = _RAND_720[3:0];
  _RAND_721 = {1{`RANDOM}};
  image_2_217 = _RAND_721[3:0];
  _RAND_722 = {1{`RANDOM}};
  image_2_218 = _RAND_722[3:0];
  _RAND_723 = {1{`RANDOM}};
  image_2_219 = _RAND_723[3:0];
  _RAND_724 = {1{`RANDOM}};
  image_2_220 = _RAND_724[3:0];
  _RAND_725 = {1{`RANDOM}};
  image_2_221 = _RAND_725[3:0];
  _RAND_726 = {1{`RANDOM}};
  image_2_222 = _RAND_726[3:0];
  _RAND_727 = {1{`RANDOM}};
  image_2_223 = _RAND_727[3:0];
  _RAND_728 = {1{`RANDOM}};
  image_2_224 = _RAND_728[3:0];
  _RAND_729 = {1{`RANDOM}};
  image_2_225 = _RAND_729[3:0];
  _RAND_730 = {1{`RANDOM}};
  image_2_226 = _RAND_730[3:0];
  _RAND_731 = {1{`RANDOM}};
  image_2_227 = _RAND_731[3:0];
  _RAND_732 = {1{`RANDOM}};
  image_2_228 = _RAND_732[3:0];
  _RAND_733 = {1{`RANDOM}};
  image_2_229 = _RAND_733[3:0];
  _RAND_734 = {1{`RANDOM}};
  image_2_230 = _RAND_734[3:0];
  _RAND_735 = {1{`RANDOM}};
  image_2_231 = _RAND_735[3:0];
  _RAND_736 = {1{`RANDOM}};
  image_2_232 = _RAND_736[3:0];
  _RAND_737 = {1{`RANDOM}};
  image_2_233 = _RAND_737[3:0];
  _RAND_738 = {1{`RANDOM}};
  image_2_234 = _RAND_738[3:0];
  _RAND_739 = {1{`RANDOM}};
  image_2_235 = _RAND_739[3:0];
  _RAND_740 = {1{`RANDOM}};
  image_2_236 = _RAND_740[3:0];
  _RAND_741 = {1{`RANDOM}};
  image_2_237 = _RAND_741[3:0];
  _RAND_742 = {1{`RANDOM}};
  image_2_238 = _RAND_742[3:0];
  _RAND_743 = {1{`RANDOM}};
  image_2_239 = _RAND_743[3:0];
  _RAND_744 = {1{`RANDOM}};
  image_2_240 = _RAND_744[3:0];
  _RAND_745 = {1{`RANDOM}};
  image_2_241 = _RAND_745[3:0];
  _RAND_746 = {1{`RANDOM}};
  image_2_242 = _RAND_746[3:0];
  _RAND_747 = {1{`RANDOM}};
  image_2_243 = _RAND_747[3:0];
  _RAND_748 = {1{`RANDOM}};
  image_2_244 = _RAND_748[3:0];
  _RAND_749 = {1{`RANDOM}};
  image_2_245 = _RAND_749[3:0];
  _RAND_750 = {1{`RANDOM}};
  image_2_246 = _RAND_750[3:0];
  _RAND_751 = {1{`RANDOM}};
  image_2_247 = _RAND_751[3:0];
  _RAND_752 = {1{`RANDOM}};
  image_2_248 = _RAND_752[3:0];
  _RAND_753 = {1{`RANDOM}};
  image_2_249 = _RAND_753[3:0];
  _RAND_754 = {1{`RANDOM}};
  image_2_250 = _RAND_754[3:0];
  _RAND_755 = {1{`RANDOM}};
  image_2_251 = _RAND_755[3:0];
  _RAND_756 = {1{`RANDOM}};
  pixelIndex = _RAND_756[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      image_0_0 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h0 == _T_34[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_6;
      end else if (8'h0 == _T_31[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_5;
      end else if (8'h0 == _T_28[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_4;
      end else if (8'h0 == _T_25[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_3;
      end else if (8'h0 == _T_22[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_2;
      end else if (8'h0 == _T_19[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_1;
      end else if (8'h0 == _T_15[7:0]) begin
        image_0_0 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_1 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1 == _T_34[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_6;
      end else if (8'h1 == _T_31[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_5;
      end else if (8'h1 == _T_28[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_4;
      end else if (8'h1 == _T_25[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_3;
      end else if (8'h1 == _T_22[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_2;
      end else if (8'h1 == _T_19[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_1;
      end else if (8'h1 == _T_15[7:0]) begin
        image_0_1 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_2 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2 == _T_34[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_6;
      end else if (8'h2 == _T_31[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_5;
      end else if (8'h2 == _T_28[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_4;
      end else if (8'h2 == _T_25[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_3;
      end else if (8'h2 == _T_22[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_2;
      end else if (8'h2 == _T_19[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_1;
      end else if (8'h2 == _T_15[7:0]) begin
        image_0_2 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_3 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3 == _T_34[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_6;
      end else if (8'h3 == _T_31[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_5;
      end else if (8'h3 == _T_28[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_4;
      end else if (8'h3 == _T_25[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_3;
      end else if (8'h3 == _T_22[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_2;
      end else if (8'h3 == _T_19[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_1;
      end else if (8'h3 == _T_15[7:0]) begin
        image_0_3 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_4 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4 == _T_34[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_6;
      end else if (8'h4 == _T_31[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_5;
      end else if (8'h4 == _T_28[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_4;
      end else if (8'h4 == _T_25[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_3;
      end else if (8'h4 == _T_22[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_2;
      end else if (8'h4 == _T_19[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_1;
      end else if (8'h4 == _T_15[7:0]) begin
        image_0_4 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_5 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5 == _T_34[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_6;
      end else if (8'h5 == _T_31[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_5;
      end else if (8'h5 == _T_28[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_4;
      end else if (8'h5 == _T_25[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_3;
      end else if (8'h5 == _T_22[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_2;
      end else if (8'h5 == _T_19[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_1;
      end else if (8'h5 == _T_15[7:0]) begin
        image_0_5 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_6 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6 == _T_34[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_6;
      end else if (8'h6 == _T_31[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_5;
      end else if (8'h6 == _T_28[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_4;
      end else if (8'h6 == _T_25[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_3;
      end else if (8'h6 == _T_22[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_2;
      end else if (8'h6 == _T_19[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_1;
      end else if (8'h6 == _T_15[7:0]) begin
        image_0_6 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_7 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7 == _T_34[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_6;
      end else if (8'h7 == _T_31[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_5;
      end else if (8'h7 == _T_28[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_4;
      end else if (8'h7 == _T_25[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_3;
      end else if (8'h7 == _T_22[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_2;
      end else if (8'h7 == _T_19[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_1;
      end else if (8'h7 == _T_15[7:0]) begin
        image_0_7 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_8 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8 == _T_34[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_6;
      end else if (8'h8 == _T_31[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_5;
      end else if (8'h8 == _T_28[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_4;
      end else if (8'h8 == _T_25[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_3;
      end else if (8'h8 == _T_22[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_2;
      end else if (8'h8 == _T_19[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_1;
      end else if (8'h8 == _T_15[7:0]) begin
        image_0_8 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_9 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h9 == _T_34[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_6;
      end else if (8'h9 == _T_31[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_5;
      end else if (8'h9 == _T_28[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_4;
      end else if (8'h9 == _T_25[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_3;
      end else if (8'h9 == _T_22[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_2;
      end else if (8'h9 == _T_19[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_1;
      end else if (8'h9 == _T_15[7:0]) begin
        image_0_9 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_10 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha == _T_34[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_6;
      end else if (8'ha == _T_31[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_5;
      end else if (8'ha == _T_28[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_4;
      end else if (8'ha == _T_25[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_3;
      end else if (8'ha == _T_22[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_2;
      end else if (8'ha == _T_19[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_1;
      end else if (8'ha == _T_15[7:0]) begin
        image_0_10 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_11 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb == _T_34[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_6;
      end else if (8'hb == _T_31[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_5;
      end else if (8'hb == _T_28[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_4;
      end else if (8'hb == _T_25[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_3;
      end else if (8'hb == _T_22[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_2;
      end else if (8'hb == _T_19[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_1;
      end else if (8'hb == _T_15[7:0]) begin
        image_0_11 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_12 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hc == _T_34[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_6;
      end else if (8'hc == _T_31[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_5;
      end else if (8'hc == _T_28[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_4;
      end else if (8'hc == _T_25[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_3;
      end else if (8'hc == _T_22[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_2;
      end else if (8'hc == _T_19[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_1;
      end else if (8'hc == _T_15[7:0]) begin
        image_0_12 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_13 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hd == _T_34[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_6;
      end else if (8'hd == _T_31[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_5;
      end else if (8'hd == _T_28[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_4;
      end else if (8'hd == _T_25[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_3;
      end else if (8'hd == _T_22[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_2;
      end else if (8'hd == _T_19[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_1;
      end else if (8'hd == _T_15[7:0]) begin
        image_0_13 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_14 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'he == _T_34[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_6;
      end else if (8'he == _T_31[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_5;
      end else if (8'he == _T_28[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_4;
      end else if (8'he == _T_25[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_3;
      end else if (8'he == _T_22[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_2;
      end else if (8'he == _T_19[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_1;
      end else if (8'he == _T_15[7:0]) begin
        image_0_14 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_15 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hf == _T_34[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_6;
      end else if (8'hf == _T_31[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_5;
      end else if (8'hf == _T_28[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_4;
      end else if (8'hf == _T_25[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_3;
      end else if (8'hf == _T_22[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_2;
      end else if (8'hf == _T_19[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_1;
      end else if (8'hf == _T_15[7:0]) begin
        image_0_15 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_16 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h10 == _T_34[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_6;
      end else if (8'h10 == _T_31[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_5;
      end else if (8'h10 == _T_28[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_4;
      end else if (8'h10 == _T_25[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_3;
      end else if (8'h10 == _T_22[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_2;
      end else if (8'h10 == _T_19[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_1;
      end else if (8'h10 == _T_15[7:0]) begin
        image_0_16 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_17 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h11 == _T_34[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_6;
      end else if (8'h11 == _T_31[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_5;
      end else if (8'h11 == _T_28[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_4;
      end else if (8'h11 == _T_25[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_3;
      end else if (8'h11 == _T_22[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_2;
      end else if (8'h11 == _T_19[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_1;
      end else if (8'h11 == _T_15[7:0]) begin
        image_0_17 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_18 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h12 == _T_34[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_6;
      end else if (8'h12 == _T_31[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_5;
      end else if (8'h12 == _T_28[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_4;
      end else if (8'h12 == _T_25[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_3;
      end else if (8'h12 == _T_22[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_2;
      end else if (8'h12 == _T_19[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_1;
      end else if (8'h12 == _T_15[7:0]) begin
        image_0_18 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_19 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h13 == _T_34[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_6;
      end else if (8'h13 == _T_31[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_5;
      end else if (8'h13 == _T_28[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_4;
      end else if (8'h13 == _T_25[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_3;
      end else if (8'h13 == _T_22[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_2;
      end else if (8'h13 == _T_19[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_1;
      end else if (8'h13 == _T_15[7:0]) begin
        image_0_19 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_20 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h14 == _T_34[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_6;
      end else if (8'h14 == _T_31[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_5;
      end else if (8'h14 == _T_28[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_4;
      end else if (8'h14 == _T_25[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_3;
      end else if (8'h14 == _T_22[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_2;
      end else if (8'h14 == _T_19[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_1;
      end else if (8'h14 == _T_15[7:0]) begin
        image_0_20 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_21 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h15 == _T_34[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_6;
      end else if (8'h15 == _T_31[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_5;
      end else if (8'h15 == _T_28[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_4;
      end else if (8'h15 == _T_25[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_3;
      end else if (8'h15 == _T_22[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_2;
      end else if (8'h15 == _T_19[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_1;
      end else if (8'h15 == _T_15[7:0]) begin
        image_0_21 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_22 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h16 == _T_34[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_6;
      end else if (8'h16 == _T_31[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_5;
      end else if (8'h16 == _T_28[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_4;
      end else if (8'h16 == _T_25[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_3;
      end else if (8'h16 == _T_22[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_2;
      end else if (8'h16 == _T_19[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_1;
      end else if (8'h16 == _T_15[7:0]) begin
        image_0_22 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_23 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h17 == _T_34[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_6;
      end else if (8'h17 == _T_31[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_5;
      end else if (8'h17 == _T_28[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_4;
      end else if (8'h17 == _T_25[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_3;
      end else if (8'h17 == _T_22[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_2;
      end else if (8'h17 == _T_19[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_1;
      end else if (8'h17 == _T_15[7:0]) begin
        image_0_23 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_24 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h18 == _T_34[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_6;
      end else if (8'h18 == _T_31[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_5;
      end else if (8'h18 == _T_28[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_4;
      end else if (8'h18 == _T_25[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_3;
      end else if (8'h18 == _T_22[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_2;
      end else if (8'h18 == _T_19[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_1;
      end else if (8'h18 == _T_15[7:0]) begin
        image_0_24 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_25 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h19 == _T_34[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_6;
      end else if (8'h19 == _T_31[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_5;
      end else if (8'h19 == _T_28[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_4;
      end else if (8'h19 == _T_25[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_3;
      end else if (8'h19 == _T_22[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_2;
      end else if (8'h19 == _T_19[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_1;
      end else if (8'h19 == _T_15[7:0]) begin
        image_0_25 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_26 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1a == _T_34[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_6;
      end else if (8'h1a == _T_31[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_5;
      end else if (8'h1a == _T_28[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_4;
      end else if (8'h1a == _T_25[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_3;
      end else if (8'h1a == _T_22[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_2;
      end else if (8'h1a == _T_19[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_1;
      end else if (8'h1a == _T_15[7:0]) begin
        image_0_26 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_27 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1b == _T_34[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_6;
      end else if (8'h1b == _T_31[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_5;
      end else if (8'h1b == _T_28[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_4;
      end else if (8'h1b == _T_25[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_3;
      end else if (8'h1b == _T_22[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_2;
      end else if (8'h1b == _T_19[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_1;
      end else if (8'h1b == _T_15[7:0]) begin
        image_0_27 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_28 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1c == _T_34[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_6;
      end else if (8'h1c == _T_31[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_5;
      end else if (8'h1c == _T_28[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_4;
      end else if (8'h1c == _T_25[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_3;
      end else if (8'h1c == _T_22[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_2;
      end else if (8'h1c == _T_19[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_1;
      end else if (8'h1c == _T_15[7:0]) begin
        image_0_28 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_29 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1d == _T_34[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_6;
      end else if (8'h1d == _T_31[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_5;
      end else if (8'h1d == _T_28[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_4;
      end else if (8'h1d == _T_25[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_3;
      end else if (8'h1d == _T_22[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_2;
      end else if (8'h1d == _T_19[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_1;
      end else if (8'h1d == _T_15[7:0]) begin
        image_0_29 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_30 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1e == _T_34[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_6;
      end else if (8'h1e == _T_31[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_5;
      end else if (8'h1e == _T_28[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_4;
      end else if (8'h1e == _T_25[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_3;
      end else if (8'h1e == _T_22[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_2;
      end else if (8'h1e == _T_19[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_1;
      end else if (8'h1e == _T_15[7:0]) begin
        image_0_30 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_31 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h1f == _T_34[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_6;
      end else if (8'h1f == _T_31[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_5;
      end else if (8'h1f == _T_28[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_4;
      end else if (8'h1f == _T_25[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_3;
      end else if (8'h1f == _T_22[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_2;
      end else if (8'h1f == _T_19[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_1;
      end else if (8'h1f == _T_15[7:0]) begin
        image_0_31 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_32 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h20 == _T_34[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_6;
      end else if (8'h20 == _T_31[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_5;
      end else if (8'h20 == _T_28[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_4;
      end else if (8'h20 == _T_25[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_3;
      end else if (8'h20 == _T_22[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_2;
      end else if (8'h20 == _T_19[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_1;
      end else if (8'h20 == _T_15[7:0]) begin
        image_0_32 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_33 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h21 == _T_34[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_6;
      end else if (8'h21 == _T_31[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_5;
      end else if (8'h21 == _T_28[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_4;
      end else if (8'h21 == _T_25[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_3;
      end else if (8'h21 == _T_22[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_2;
      end else if (8'h21 == _T_19[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_1;
      end else if (8'h21 == _T_15[7:0]) begin
        image_0_33 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_34 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h22 == _T_34[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_6;
      end else if (8'h22 == _T_31[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_5;
      end else if (8'h22 == _T_28[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_4;
      end else if (8'h22 == _T_25[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_3;
      end else if (8'h22 == _T_22[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_2;
      end else if (8'h22 == _T_19[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_1;
      end else if (8'h22 == _T_15[7:0]) begin
        image_0_34 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_35 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h23 == _T_34[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_6;
      end else if (8'h23 == _T_31[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_5;
      end else if (8'h23 == _T_28[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_4;
      end else if (8'h23 == _T_25[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_3;
      end else if (8'h23 == _T_22[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_2;
      end else if (8'h23 == _T_19[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_1;
      end else if (8'h23 == _T_15[7:0]) begin
        image_0_35 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_36 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h24 == _T_34[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_6;
      end else if (8'h24 == _T_31[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_5;
      end else if (8'h24 == _T_28[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_4;
      end else if (8'h24 == _T_25[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_3;
      end else if (8'h24 == _T_22[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_2;
      end else if (8'h24 == _T_19[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_1;
      end else if (8'h24 == _T_15[7:0]) begin
        image_0_36 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_37 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h25 == _T_34[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_6;
      end else if (8'h25 == _T_31[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_5;
      end else if (8'h25 == _T_28[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_4;
      end else if (8'h25 == _T_25[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_3;
      end else if (8'h25 == _T_22[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_2;
      end else if (8'h25 == _T_19[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_1;
      end else if (8'h25 == _T_15[7:0]) begin
        image_0_37 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_38 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h26 == _T_34[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_6;
      end else if (8'h26 == _T_31[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_5;
      end else if (8'h26 == _T_28[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_4;
      end else if (8'h26 == _T_25[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_3;
      end else if (8'h26 == _T_22[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_2;
      end else if (8'h26 == _T_19[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_1;
      end else if (8'h26 == _T_15[7:0]) begin
        image_0_38 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_39 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h27 == _T_34[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_6;
      end else if (8'h27 == _T_31[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_5;
      end else if (8'h27 == _T_28[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_4;
      end else if (8'h27 == _T_25[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_3;
      end else if (8'h27 == _T_22[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_2;
      end else if (8'h27 == _T_19[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_1;
      end else if (8'h27 == _T_15[7:0]) begin
        image_0_39 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_40 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h28 == _T_34[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_6;
      end else if (8'h28 == _T_31[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_5;
      end else if (8'h28 == _T_28[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_4;
      end else if (8'h28 == _T_25[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_3;
      end else if (8'h28 == _T_22[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_2;
      end else if (8'h28 == _T_19[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_1;
      end else if (8'h28 == _T_15[7:0]) begin
        image_0_40 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_41 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h29 == _T_34[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_6;
      end else if (8'h29 == _T_31[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_5;
      end else if (8'h29 == _T_28[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_4;
      end else if (8'h29 == _T_25[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_3;
      end else if (8'h29 == _T_22[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_2;
      end else if (8'h29 == _T_19[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_1;
      end else if (8'h29 == _T_15[7:0]) begin
        image_0_41 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_42 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2a == _T_34[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_6;
      end else if (8'h2a == _T_31[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_5;
      end else if (8'h2a == _T_28[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_4;
      end else if (8'h2a == _T_25[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_3;
      end else if (8'h2a == _T_22[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_2;
      end else if (8'h2a == _T_19[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_1;
      end else if (8'h2a == _T_15[7:0]) begin
        image_0_42 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_43 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2b == _T_34[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_6;
      end else if (8'h2b == _T_31[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_5;
      end else if (8'h2b == _T_28[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_4;
      end else if (8'h2b == _T_25[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_3;
      end else if (8'h2b == _T_22[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_2;
      end else if (8'h2b == _T_19[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_1;
      end else if (8'h2b == _T_15[7:0]) begin
        image_0_43 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_44 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2c == _T_34[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_6;
      end else if (8'h2c == _T_31[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_5;
      end else if (8'h2c == _T_28[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_4;
      end else if (8'h2c == _T_25[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_3;
      end else if (8'h2c == _T_22[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_2;
      end else if (8'h2c == _T_19[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_1;
      end else if (8'h2c == _T_15[7:0]) begin
        image_0_44 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_45 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2d == _T_34[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_6;
      end else if (8'h2d == _T_31[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_5;
      end else if (8'h2d == _T_28[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_4;
      end else if (8'h2d == _T_25[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_3;
      end else if (8'h2d == _T_22[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_2;
      end else if (8'h2d == _T_19[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_1;
      end else if (8'h2d == _T_15[7:0]) begin
        image_0_45 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_46 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2e == _T_34[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_6;
      end else if (8'h2e == _T_31[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_5;
      end else if (8'h2e == _T_28[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_4;
      end else if (8'h2e == _T_25[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_3;
      end else if (8'h2e == _T_22[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_2;
      end else if (8'h2e == _T_19[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_1;
      end else if (8'h2e == _T_15[7:0]) begin
        image_0_46 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_47 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h2f == _T_34[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_6;
      end else if (8'h2f == _T_31[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_5;
      end else if (8'h2f == _T_28[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_4;
      end else if (8'h2f == _T_25[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_3;
      end else if (8'h2f == _T_22[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_2;
      end else if (8'h2f == _T_19[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_1;
      end else if (8'h2f == _T_15[7:0]) begin
        image_0_47 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_48 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h30 == _T_34[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_6;
      end else if (8'h30 == _T_31[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_5;
      end else if (8'h30 == _T_28[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_4;
      end else if (8'h30 == _T_25[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_3;
      end else if (8'h30 == _T_22[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_2;
      end else if (8'h30 == _T_19[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_1;
      end else if (8'h30 == _T_15[7:0]) begin
        image_0_48 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_49 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h31 == _T_34[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_6;
      end else if (8'h31 == _T_31[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_5;
      end else if (8'h31 == _T_28[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_4;
      end else if (8'h31 == _T_25[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_3;
      end else if (8'h31 == _T_22[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_2;
      end else if (8'h31 == _T_19[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_1;
      end else if (8'h31 == _T_15[7:0]) begin
        image_0_49 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_50 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h32 == _T_34[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_6;
      end else if (8'h32 == _T_31[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_5;
      end else if (8'h32 == _T_28[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_4;
      end else if (8'h32 == _T_25[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_3;
      end else if (8'h32 == _T_22[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_2;
      end else if (8'h32 == _T_19[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_1;
      end else if (8'h32 == _T_15[7:0]) begin
        image_0_50 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_51 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h33 == _T_34[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_6;
      end else if (8'h33 == _T_31[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_5;
      end else if (8'h33 == _T_28[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_4;
      end else if (8'h33 == _T_25[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_3;
      end else if (8'h33 == _T_22[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_2;
      end else if (8'h33 == _T_19[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_1;
      end else if (8'h33 == _T_15[7:0]) begin
        image_0_51 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_52 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h34 == _T_34[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_6;
      end else if (8'h34 == _T_31[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_5;
      end else if (8'h34 == _T_28[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_4;
      end else if (8'h34 == _T_25[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_3;
      end else if (8'h34 == _T_22[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_2;
      end else if (8'h34 == _T_19[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_1;
      end else if (8'h34 == _T_15[7:0]) begin
        image_0_52 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_53 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h35 == _T_34[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_6;
      end else if (8'h35 == _T_31[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_5;
      end else if (8'h35 == _T_28[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_4;
      end else if (8'h35 == _T_25[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_3;
      end else if (8'h35 == _T_22[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_2;
      end else if (8'h35 == _T_19[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_1;
      end else if (8'h35 == _T_15[7:0]) begin
        image_0_53 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_54 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h36 == _T_34[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_6;
      end else if (8'h36 == _T_31[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_5;
      end else if (8'h36 == _T_28[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_4;
      end else if (8'h36 == _T_25[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_3;
      end else if (8'h36 == _T_22[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_2;
      end else if (8'h36 == _T_19[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_1;
      end else if (8'h36 == _T_15[7:0]) begin
        image_0_54 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_55 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h37 == _T_34[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_6;
      end else if (8'h37 == _T_31[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_5;
      end else if (8'h37 == _T_28[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_4;
      end else if (8'h37 == _T_25[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_3;
      end else if (8'h37 == _T_22[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_2;
      end else if (8'h37 == _T_19[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_1;
      end else if (8'h37 == _T_15[7:0]) begin
        image_0_55 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_56 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h38 == _T_34[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_6;
      end else if (8'h38 == _T_31[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_5;
      end else if (8'h38 == _T_28[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_4;
      end else if (8'h38 == _T_25[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_3;
      end else if (8'h38 == _T_22[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_2;
      end else if (8'h38 == _T_19[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_1;
      end else if (8'h38 == _T_15[7:0]) begin
        image_0_56 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_57 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h39 == _T_34[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_6;
      end else if (8'h39 == _T_31[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_5;
      end else if (8'h39 == _T_28[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_4;
      end else if (8'h39 == _T_25[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_3;
      end else if (8'h39 == _T_22[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_2;
      end else if (8'h39 == _T_19[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_1;
      end else if (8'h39 == _T_15[7:0]) begin
        image_0_57 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_58 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3a == _T_34[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_6;
      end else if (8'h3a == _T_31[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_5;
      end else if (8'h3a == _T_28[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_4;
      end else if (8'h3a == _T_25[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_3;
      end else if (8'h3a == _T_22[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_2;
      end else if (8'h3a == _T_19[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_1;
      end else if (8'h3a == _T_15[7:0]) begin
        image_0_58 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_59 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3b == _T_34[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_6;
      end else if (8'h3b == _T_31[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_5;
      end else if (8'h3b == _T_28[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_4;
      end else if (8'h3b == _T_25[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_3;
      end else if (8'h3b == _T_22[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_2;
      end else if (8'h3b == _T_19[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_1;
      end else if (8'h3b == _T_15[7:0]) begin
        image_0_59 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_60 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3c == _T_34[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_6;
      end else if (8'h3c == _T_31[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_5;
      end else if (8'h3c == _T_28[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_4;
      end else if (8'h3c == _T_25[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_3;
      end else if (8'h3c == _T_22[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_2;
      end else if (8'h3c == _T_19[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_1;
      end else if (8'h3c == _T_15[7:0]) begin
        image_0_60 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_61 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3d == _T_34[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_6;
      end else if (8'h3d == _T_31[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_5;
      end else if (8'h3d == _T_28[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_4;
      end else if (8'h3d == _T_25[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_3;
      end else if (8'h3d == _T_22[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_2;
      end else if (8'h3d == _T_19[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_1;
      end else if (8'h3d == _T_15[7:0]) begin
        image_0_61 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_62 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3e == _T_34[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_6;
      end else if (8'h3e == _T_31[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_5;
      end else if (8'h3e == _T_28[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_4;
      end else if (8'h3e == _T_25[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_3;
      end else if (8'h3e == _T_22[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_2;
      end else if (8'h3e == _T_19[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_1;
      end else if (8'h3e == _T_15[7:0]) begin
        image_0_62 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_63 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h3f == _T_34[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_6;
      end else if (8'h3f == _T_31[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_5;
      end else if (8'h3f == _T_28[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_4;
      end else if (8'h3f == _T_25[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_3;
      end else if (8'h3f == _T_22[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_2;
      end else if (8'h3f == _T_19[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_1;
      end else if (8'h3f == _T_15[7:0]) begin
        image_0_63 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_64 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h40 == _T_34[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_6;
      end else if (8'h40 == _T_31[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_5;
      end else if (8'h40 == _T_28[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_4;
      end else if (8'h40 == _T_25[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_3;
      end else if (8'h40 == _T_22[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_2;
      end else if (8'h40 == _T_19[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_1;
      end else if (8'h40 == _T_15[7:0]) begin
        image_0_64 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_65 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h41 == _T_34[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_6;
      end else if (8'h41 == _T_31[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_5;
      end else if (8'h41 == _T_28[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_4;
      end else if (8'h41 == _T_25[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_3;
      end else if (8'h41 == _T_22[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_2;
      end else if (8'h41 == _T_19[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_1;
      end else if (8'h41 == _T_15[7:0]) begin
        image_0_65 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_66 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h42 == _T_34[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_6;
      end else if (8'h42 == _T_31[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_5;
      end else if (8'h42 == _T_28[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_4;
      end else if (8'h42 == _T_25[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_3;
      end else if (8'h42 == _T_22[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_2;
      end else if (8'h42 == _T_19[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_1;
      end else if (8'h42 == _T_15[7:0]) begin
        image_0_66 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_67 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h43 == _T_34[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_6;
      end else if (8'h43 == _T_31[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_5;
      end else if (8'h43 == _T_28[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_4;
      end else if (8'h43 == _T_25[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_3;
      end else if (8'h43 == _T_22[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_2;
      end else if (8'h43 == _T_19[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_1;
      end else if (8'h43 == _T_15[7:0]) begin
        image_0_67 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_68 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h44 == _T_34[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_6;
      end else if (8'h44 == _T_31[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_5;
      end else if (8'h44 == _T_28[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_4;
      end else if (8'h44 == _T_25[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_3;
      end else if (8'h44 == _T_22[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_2;
      end else if (8'h44 == _T_19[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_1;
      end else if (8'h44 == _T_15[7:0]) begin
        image_0_68 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_69 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h45 == _T_34[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_6;
      end else if (8'h45 == _T_31[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_5;
      end else if (8'h45 == _T_28[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_4;
      end else if (8'h45 == _T_25[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_3;
      end else if (8'h45 == _T_22[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_2;
      end else if (8'h45 == _T_19[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_1;
      end else if (8'h45 == _T_15[7:0]) begin
        image_0_69 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_70 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h46 == _T_34[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_6;
      end else if (8'h46 == _T_31[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_5;
      end else if (8'h46 == _T_28[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_4;
      end else if (8'h46 == _T_25[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_3;
      end else if (8'h46 == _T_22[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_2;
      end else if (8'h46 == _T_19[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_1;
      end else if (8'h46 == _T_15[7:0]) begin
        image_0_70 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_71 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h47 == _T_34[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_6;
      end else if (8'h47 == _T_31[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_5;
      end else if (8'h47 == _T_28[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_4;
      end else if (8'h47 == _T_25[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_3;
      end else if (8'h47 == _T_22[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_2;
      end else if (8'h47 == _T_19[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_1;
      end else if (8'h47 == _T_15[7:0]) begin
        image_0_71 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_72 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h48 == _T_34[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_6;
      end else if (8'h48 == _T_31[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_5;
      end else if (8'h48 == _T_28[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_4;
      end else if (8'h48 == _T_25[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_3;
      end else if (8'h48 == _T_22[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_2;
      end else if (8'h48 == _T_19[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_1;
      end else if (8'h48 == _T_15[7:0]) begin
        image_0_72 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_73 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h49 == _T_34[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_6;
      end else if (8'h49 == _T_31[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_5;
      end else if (8'h49 == _T_28[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_4;
      end else if (8'h49 == _T_25[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_3;
      end else if (8'h49 == _T_22[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_2;
      end else if (8'h49 == _T_19[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_1;
      end else if (8'h49 == _T_15[7:0]) begin
        image_0_73 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_74 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4a == _T_34[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_6;
      end else if (8'h4a == _T_31[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_5;
      end else if (8'h4a == _T_28[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_4;
      end else if (8'h4a == _T_25[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_3;
      end else if (8'h4a == _T_22[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_2;
      end else if (8'h4a == _T_19[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_1;
      end else if (8'h4a == _T_15[7:0]) begin
        image_0_74 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_75 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4b == _T_34[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_6;
      end else if (8'h4b == _T_31[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_5;
      end else if (8'h4b == _T_28[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_4;
      end else if (8'h4b == _T_25[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_3;
      end else if (8'h4b == _T_22[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_2;
      end else if (8'h4b == _T_19[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_1;
      end else if (8'h4b == _T_15[7:0]) begin
        image_0_75 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_76 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4c == _T_34[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_6;
      end else if (8'h4c == _T_31[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_5;
      end else if (8'h4c == _T_28[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_4;
      end else if (8'h4c == _T_25[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_3;
      end else if (8'h4c == _T_22[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_2;
      end else if (8'h4c == _T_19[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_1;
      end else if (8'h4c == _T_15[7:0]) begin
        image_0_76 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_77 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4d == _T_34[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_6;
      end else if (8'h4d == _T_31[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_5;
      end else if (8'h4d == _T_28[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_4;
      end else if (8'h4d == _T_25[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_3;
      end else if (8'h4d == _T_22[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_2;
      end else if (8'h4d == _T_19[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_1;
      end else if (8'h4d == _T_15[7:0]) begin
        image_0_77 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_78 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4e == _T_34[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_6;
      end else if (8'h4e == _T_31[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_5;
      end else if (8'h4e == _T_28[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_4;
      end else if (8'h4e == _T_25[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_3;
      end else if (8'h4e == _T_22[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_2;
      end else if (8'h4e == _T_19[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_1;
      end else if (8'h4e == _T_15[7:0]) begin
        image_0_78 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_79 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h4f == _T_34[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_6;
      end else if (8'h4f == _T_31[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_5;
      end else if (8'h4f == _T_28[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_4;
      end else if (8'h4f == _T_25[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_3;
      end else if (8'h4f == _T_22[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_2;
      end else if (8'h4f == _T_19[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_1;
      end else if (8'h4f == _T_15[7:0]) begin
        image_0_79 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_80 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h50 == _T_34[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_6;
      end else if (8'h50 == _T_31[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_5;
      end else if (8'h50 == _T_28[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_4;
      end else if (8'h50 == _T_25[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_3;
      end else if (8'h50 == _T_22[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_2;
      end else if (8'h50 == _T_19[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_1;
      end else if (8'h50 == _T_15[7:0]) begin
        image_0_80 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_81 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h51 == _T_34[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_6;
      end else if (8'h51 == _T_31[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_5;
      end else if (8'h51 == _T_28[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_4;
      end else if (8'h51 == _T_25[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_3;
      end else if (8'h51 == _T_22[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_2;
      end else if (8'h51 == _T_19[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_1;
      end else if (8'h51 == _T_15[7:0]) begin
        image_0_81 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_82 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h52 == _T_34[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_6;
      end else if (8'h52 == _T_31[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_5;
      end else if (8'h52 == _T_28[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_4;
      end else if (8'h52 == _T_25[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_3;
      end else if (8'h52 == _T_22[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_2;
      end else if (8'h52 == _T_19[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_1;
      end else if (8'h52 == _T_15[7:0]) begin
        image_0_82 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_83 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h53 == _T_34[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_6;
      end else if (8'h53 == _T_31[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_5;
      end else if (8'h53 == _T_28[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_4;
      end else if (8'h53 == _T_25[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_3;
      end else if (8'h53 == _T_22[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_2;
      end else if (8'h53 == _T_19[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_1;
      end else if (8'h53 == _T_15[7:0]) begin
        image_0_83 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_84 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h54 == _T_34[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_6;
      end else if (8'h54 == _T_31[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_5;
      end else if (8'h54 == _T_28[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_4;
      end else if (8'h54 == _T_25[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_3;
      end else if (8'h54 == _T_22[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_2;
      end else if (8'h54 == _T_19[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_1;
      end else if (8'h54 == _T_15[7:0]) begin
        image_0_84 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_85 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h55 == _T_34[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_6;
      end else if (8'h55 == _T_31[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_5;
      end else if (8'h55 == _T_28[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_4;
      end else if (8'h55 == _T_25[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_3;
      end else if (8'h55 == _T_22[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_2;
      end else if (8'h55 == _T_19[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_1;
      end else if (8'h55 == _T_15[7:0]) begin
        image_0_85 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_86 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h56 == _T_34[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_6;
      end else if (8'h56 == _T_31[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_5;
      end else if (8'h56 == _T_28[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_4;
      end else if (8'h56 == _T_25[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_3;
      end else if (8'h56 == _T_22[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_2;
      end else if (8'h56 == _T_19[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_1;
      end else if (8'h56 == _T_15[7:0]) begin
        image_0_86 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_87 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h57 == _T_34[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_6;
      end else if (8'h57 == _T_31[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_5;
      end else if (8'h57 == _T_28[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_4;
      end else if (8'h57 == _T_25[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_3;
      end else if (8'h57 == _T_22[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_2;
      end else if (8'h57 == _T_19[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_1;
      end else if (8'h57 == _T_15[7:0]) begin
        image_0_87 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_88 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h58 == _T_34[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_6;
      end else if (8'h58 == _T_31[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_5;
      end else if (8'h58 == _T_28[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_4;
      end else if (8'h58 == _T_25[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_3;
      end else if (8'h58 == _T_22[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_2;
      end else if (8'h58 == _T_19[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_1;
      end else if (8'h58 == _T_15[7:0]) begin
        image_0_88 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_89 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h59 == _T_34[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_6;
      end else if (8'h59 == _T_31[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_5;
      end else if (8'h59 == _T_28[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_4;
      end else if (8'h59 == _T_25[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_3;
      end else if (8'h59 == _T_22[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_2;
      end else if (8'h59 == _T_19[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_1;
      end else if (8'h59 == _T_15[7:0]) begin
        image_0_89 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_90 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5a == _T_34[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_6;
      end else if (8'h5a == _T_31[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_5;
      end else if (8'h5a == _T_28[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_4;
      end else if (8'h5a == _T_25[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_3;
      end else if (8'h5a == _T_22[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_2;
      end else if (8'h5a == _T_19[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_1;
      end else if (8'h5a == _T_15[7:0]) begin
        image_0_90 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_91 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5b == _T_34[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_6;
      end else if (8'h5b == _T_31[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_5;
      end else if (8'h5b == _T_28[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_4;
      end else if (8'h5b == _T_25[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_3;
      end else if (8'h5b == _T_22[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_2;
      end else if (8'h5b == _T_19[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_1;
      end else if (8'h5b == _T_15[7:0]) begin
        image_0_91 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_92 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5c == _T_34[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_6;
      end else if (8'h5c == _T_31[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_5;
      end else if (8'h5c == _T_28[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_4;
      end else if (8'h5c == _T_25[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_3;
      end else if (8'h5c == _T_22[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_2;
      end else if (8'h5c == _T_19[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_1;
      end else if (8'h5c == _T_15[7:0]) begin
        image_0_92 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_93 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5d == _T_34[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_6;
      end else if (8'h5d == _T_31[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_5;
      end else if (8'h5d == _T_28[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_4;
      end else if (8'h5d == _T_25[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_3;
      end else if (8'h5d == _T_22[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_2;
      end else if (8'h5d == _T_19[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_1;
      end else if (8'h5d == _T_15[7:0]) begin
        image_0_93 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_94 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5e == _T_34[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_6;
      end else if (8'h5e == _T_31[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_5;
      end else if (8'h5e == _T_28[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_4;
      end else if (8'h5e == _T_25[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_3;
      end else if (8'h5e == _T_22[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_2;
      end else if (8'h5e == _T_19[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_1;
      end else if (8'h5e == _T_15[7:0]) begin
        image_0_94 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_95 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h5f == _T_34[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_6;
      end else if (8'h5f == _T_31[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_5;
      end else if (8'h5f == _T_28[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_4;
      end else if (8'h5f == _T_25[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_3;
      end else if (8'h5f == _T_22[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_2;
      end else if (8'h5f == _T_19[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_1;
      end else if (8'h5f == _T_15[7:0]) begin
        image_0_95 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_96 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h60 == _T_34[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_6;
      end else if (8'h60 == _T_31[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_5;
      end else if (8'h60 == _T_28[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_4;
      end else if (8'h60 == _T_25[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_3;
      end else if (8'h60 == _T_22[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_2;
      end else if (8'h60 == _T_19[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_1;
      end else if (8'h60 == _T_15[7:0]) begin
        image_0_96 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_97 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h61 == _T_34[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_6;
      end else if (8'h61 == _T_31[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_5;
      end else if (8'h61 == _T_28[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_4;
      end else if (8'h61 == _T_25[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_3;
      end else if (8'h61 == _T_22[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_2;
      end else if (8'h61 == _T_19[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_1;
      end else if (8'h61 == _T_15[7:0]) begin
        image_0_97 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_98 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h62 == _T_34[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_6;
      end else if (8'h62 == _T_31[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_5;
      end else if (8'h62 == _T_28[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_4;
      end else if (8'h62 == _T_25[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_3;
      end else if (8'h62 == _T_22[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_2;
      end else if (8'h62 == _T_19[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_1;
      end else if (8'h62 == _T_15[7:0]) begin
        image_0_98 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_99 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h63 == _T_34[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_6;
      end else if (8'h63 == _T_31[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_5;
      end else if (8'h63 == _T_28[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_4;
      end else if (8'h63 == _T_25[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_3;
      end else if (8'h63 == _T_22[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_2;
      end else if (8'h63 == _T_19[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_1;
      end else if (8'h63 == _T_15[7:0]) begin
        image_0_99 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_100 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h64 == _T_34[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_6;
      end else if (8'h64 == _T_31[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_5;
      end else if (8'h64 == _T_28[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_4;
      end else if (8'h64 == _T_25[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_3;
      end else if (8'h64 == _T_22[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_2;
      end else if (8'h64 == _T_19[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_1;
      end else if (8'h64 == _T_15[7:0]) begin
        image_0_100 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_101 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h65 == _T_34[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_6;
      end else if (8'h65 == _T_31[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_5;
      end else if (8'h65 == _T_28[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_4;
      end else if (8'h65 == _T_25[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_3;
      end else if (8'h65 == _T_22[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_2;
      end else if (8'h65 == _T_19[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_1;
      end else if (8'h65 == _T_15[7:0]) begin
        image_0_101 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_102 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h66 == _T_34[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_6;
      end else if (8'h66 == _T_31[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_5;
      end else if (8'h66 == _T_28[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_4;
      end else if (8'h66 == _T_25[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_3;
      end else if (8'h66 == _T_22[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_2;
      end else if (8'h66 == _T_19[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_1;
      end else if (8'h66 == _T_15[7:0]) begin
        image_0_102 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_103 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h67 == _T_34[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_6;
      end else if (8'h67 == _T_31[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_5;
      end else if (8'h67 == _T_28[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_4;
      end else if (8'h67 == _T_25[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_3;
      end else if (8'h67 == _T_22[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_2;
      end else if (8'h67 == _T_19[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_1;
      end else if (8'h67 == _T_15[7:0]) begin
        image_0_103 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_104 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h68 == _T_34[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_6;
      end else if (8'h68 == _T_31[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_5;
      end else if (8'h68 == _T_28[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_4;
      end else if (8'h68 == _T_25[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_3;
      end else if (8'h68 == _T_22[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_2;
      end else if (8'h68 == _T_19[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_1;
      end else if (8'h68 == _T_15[7:0]) begin
        image_0_104 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_105 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h69 == _T_34[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_6;
      end else if (8'h69 == _T_31[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_5;
      end else if (8'h69 == _T_28[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_4;
      end else if (8'h69 == _T_25[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_3;
      end else if (8'h69 == _T_22[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_2;
      end else if (8'h69 == _T_19[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_1;
      end else if (8'h69 == _T_15[7:0]) begin
        image_0_105 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_106 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6a == _T_34[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_6;
      end else if (8'h6a == _T_31[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_5;
      end else if (8'h6a == _T_28[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_4;
      end else if (8'h6a == _T_25[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_3;
      end else if (8'h6a == _T_22[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_2;
      end else if (8'h6a == _T_19[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_1;
      end else if (8'h6a == _T_15[7:0]) begin
        image_0_106 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_107 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6b == _T_34[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_6;
      end else if (8'h6b == _T_31[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_5;
      end else if (8'h6b == _T_28[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_4;
      end else if (8'h6b == _T_25[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_3;
      end else if (8'h6b == _T_22[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_2;
      end else if (8'h6b == _T_19[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_1;
      end else if (8'h6b == _T_15[7:0]) begin
        image_0_107 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_108 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6c == _T_34[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_6;
      end else if (8'h6c == _T_31[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_5;
      end else if (8'h6c == _T_28[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_4;
      end else if (8'h6c == _T_25[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_3;
      end else if (8'h6c == _T_22[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_2;
      end else if (8'h6c == _T_19[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_1;
      end else if (8'h6c == _T_15[7:0]) begin
        image_0_108 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_109 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6d == _T_34[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_6;
      end else if (8'h6d == _T_31[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_5;
      end else if (8'h6d == _T_28[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_4;
      end else if (8'h6d == _T_25[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_3;
      end else if (8'h6d == _T_22[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_2;
      end else if (8'h6d == _T_19[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_1;
      end else if (8'h6d == _T_15[7:0]) begin
        image_0_109 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_110 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6e == _T_34[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_6;
      end else if (8'h6e == _T_31[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_5;
      end else if (8'h6e == _T_28[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_4;
      end else if (8'h6e == _T_25[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_3;
      end else if (8'h6e == _T_22[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_2;
      end else if (8'h6e == _T_19[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_1;
      end else if (8'h6e == _T_15[7:0]) begin
        image_0_110 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_111 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h6f == _T_34[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_6;
      end else if (8'h6f == _T_31[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_5;
      end else if (8'h6f == _T_28[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_4;
      end else if (8'h6f == _T_25[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_3;
      end else if (8'h6f == _T_22[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_2;
      end else if (8'h6f == _T_19[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_1;
      end else if (8'h6f == _T_15[7:0]) begin
        image_0_111 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_112 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h70 == _T_34[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_6;
      end else if (8'h70 == _T_31[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_5;
      end else if (8'h70 == _T_28[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_4;
      end else if (8'h70 == _T_25[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_3;
      end else if (8'h70 == _T_22[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_2;
      end else if (8'h70 == _T_19[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_1;
      end else if (8'h70 == _T_15[7:0]) begin
        image_0_112 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_113 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h71 == _T_34[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_6;
      end else if (8'h71 == _T_31[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_5;
      end else if (8'h71 == _T_28[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_4;
      end else if (8'h71 == _T_25[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_3;
      end else if (8'h71 == _T_22[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_2;
      end else if (8'h71 == _T_19[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_1;
      end else if (8'h71 == _T_15[7:0]) begin
        image_0_113 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_114 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h72 == _T_34[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_6;
      end else if (8'h72 == _T_31[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_5;
      end else if (8'h72 == _T_28[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_4;
      end else if (8'h72 == _T_25[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_3;
      end else if (8'h72 == _T_22[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_2;
      end else if (8'h72 == _T_19[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_1;
      end else if (8'h72 == _T_15[7:0]) begin
        image_0_114 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_115 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h73 == _T_34[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_6;
      end else if (8'h73 == _T_31[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_5;
      end else if (8'h73 == _T_28[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_4;
      end else if (8'h73 == _T_25[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_3;
      end else if (8'h73 == _T_22[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_2;
      end else if (8'h73 == _T_19[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_1;
      end else if (8'h73 == _T_15[7:0]) begin
        image_0_115 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_116 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h74 == _T_34[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_6;
      end else if (8'h74 == _T_31[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_5;
      end else if (8'h74 == _T_28[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_4;
      end else if (8'h74 == _T_25[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_3;
      end else if (8'h74 == _T_22[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_2;
      end else if (8'h74 == _T_19[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_1;
      end else if (8'h74 == _T_15[7:0]) begin
        image_0_116 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_117 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h75 == _T_34[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_6;
      end else if (8'h75 == _T_31[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_5;
      end else if (8'h75 == _T_28[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_4;
      end else if (8'h75 == _T_25[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_3;
      end else if (8'h75 == _T_22[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_2;
      end else if (8'h75 == _T_19[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_1;
      end else if (8'h75 == _T_15[7:0]) begin
        image_0_117 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_118 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h76 == _T_34[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_6;
      end else if (8'h76 == _T_31[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_5;
      end else if (8'h76 == _T_28[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_4;
      end else if (8'h76 == _T_25[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_3;
      end else if (8'h76 == _T_22[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_2;
      end else if (8'h76 == _T_19[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_1;
      end else if (8'h76 == _T_15[7:0]) begin
        image_0_118 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_119 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h77 == _T_34[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_6;
      end else if (8'h77 == _T_31[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_5;
      end else if (8'h77 == _T_28[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_4;
      end else if (8'h77 == _T_25[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_3;
      end else if (8'h77 == _T_22[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_2;
      end else if (8'h77 == _T_19[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_1;
      end else if (8'h77 == _T_15[7:0]) begin
        image_0_119 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_120 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h78 == _T_34[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_6;
      end else if (8'h78 == _T_31[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_5;
      end else if (8'h78 == _T_28[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_4;
      end else if (8'h78 == _T_25[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_3;
      end else if (8'h78 == _T_22[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_2;
      end else if (8'h78 == _T_19[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_1;
      end else if (8'h78 == _T_15[7:0]) begin
        image_0_120 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_121 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h79 == _T_34[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_6;
      end else if (8'h79 == _T_31[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_5;
      end else if (8'h79 == _T_28[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_4;
      end else if (8'h79 == _T_25[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_3;
      end else if (8'h79 == _T_22[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_2;
      end else if (8'h79 == _T_19[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_1;
      end else if (8'h79 == _T_15[7:0]) begin
        image_0_121 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_122 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7a == _T_34[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_6;
      end else if (8'h7a == _T_31[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_5;
      end else if (8'h7a == _T_28[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_4;
      end else if (8'h7a == _T_25[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_3;
      end else if (8'h7a == _T_22[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_2;
      end else if (8'h7a == _T_19[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_1;
      end else if (8'h7a == _T_15[7:0]) begin
        image_0_122 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_123 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7b == _T_34[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_6;
      end else if (8'h7b == _T_31[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_5;
      end else if (8'h7b == _T_28[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_4;
      end else if (8'h7b == _T_25[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_3;
      end else if (8'h7b == _T_22[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_2;
      end else if (8'h7b == _T_19[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_1;
      end else if (8'h7b == _T_15[7:0]) begin
        image_0_123 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_124 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7c == _T_34[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_6;
      end else if (8'h7c == _T_31[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_5;
      end else if (8'h7c == _T_28[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_4;
      end else if (8'h7c == _T_25[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_3;
      end else if (8'h7c == _T_22[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_2;
      end else if (8'h7c == _T_19[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_1;
      end else if (8'h7c == _T_15[7:0]) begin
        image_0_124 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_125 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7d == _T_34[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_6;
      end else if (8'h7d == _T_31[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_5;
      end else if (8'h7d == _T_28[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_4;
      end else if (8'h7d == _T_25[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_3;
      end else if (8'h7d == _T_22[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_2;
      end else if (8'h7d == _T_19[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_1;
      end else if (8'h7d == _T_15[7:0]) begin
        image_0_125 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_126 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7e == _T_34[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_6;
      end else if (8'h7e == _T_31[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_5;
      end else if (8'h7e == _T_28[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_4;
      end else if (8'h7e == _T_25[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_3;
      end else if (8'h7e == _T_22[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_2;
      end else if (8'h7e == _T_19[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_1;
      end else if (8'h7e == _T_15[7:0]) begin
        image_0_126 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_127 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h7f == _T_34[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_6;
      end else if (8'h7f == _T_31[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_5;
      end else if (8'h7f == _T_28[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_4;
      end else if (8'h7f == _T_25[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_3;
      end else if (8'h7f == _T_22[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_2;
      end else if (8'h7f == _T_19[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_1;
      end else if (8'h7f == _T_15[7:0]) begin
        image_0_127 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_128 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h80 == _T_34[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_6;
      end else if (8'h80 == _T_31[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_5;
      end else if (8'h80 == _T_28[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_4;
      end else if (8'h80 == _T_25[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_3;
      end else if (8'h80 == _T_22[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_2;
      end else if (8'h80 == _T_19[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_1;
      end else if (8'h80 == _T_15[7:0]) begin
        image_0_128 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_129 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h81 == _T_34[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_6;
      end else if (8'h81 == _T_31[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_5;
      end else if (8'h81 == _T_28[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_4;
      end else if (8'h81 == _T_25[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_3;
      end else if (8'h81 == _T_22[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_2;
      end else if (8'h81 == _T_19[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_1;
      end else if (8'h81 == _T_15[7:0]) begin
        image_0_129 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_130 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h82 == _T_34[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_6;
      end else if (8'h82 == _T_31[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_5;
      end else if (8'h82 == _T_28[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_4;
      end else if (8'h82 == _T_25[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_3;
      end else if (8'h82 == _T_22[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_2;
      end else if (8'h82 == _T_19[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_1;
      end else if (8'h82 == _T_15[7:0]) begin
        image_0_130 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_131 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h83 == _T_34[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_6;
      end else if (8'h83 == _T_31[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_5;
      end else if (8'h83 == _T_28[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_4;
      end else if (8'h83 == _T_25[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_3;
      end else if (8'h83 == _T_22[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_2;
      end else if (8'h83 == _T_19[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_1;
      end else if (8'h83 == _T_15[7:0]) begin
        image_0_131 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_132 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h84 == _T_34[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_6;
      end else if (8'h84 == _T_31[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_5;
      end else if (8'h84 == _T_28[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_4;
      end else if (8'h84 == _T_25[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_3;
      end else if (8'h84 == _T_22[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_2;
      end else if (8'h84 == _T_19[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_1;
      end else if (8'h84 == _T_15[7:0]) begin
        image_0_132 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_133 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h85 == _T_34[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_6;
      end else if (8'h85 == _T_31[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_5;
      end else if (8'h85 == _T_28[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_4;
      end else if (8'h85 == _T_25[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_3;
      end else if (8'h85 == _T_22[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_2;
      end else if (8'h85 == _T_19[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_1;
      end else if (8'h85 == _T_15[7:0]) begin
        image_0_133 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_134 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h86 == _T_34[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_6;
      end else if (8'h86 == _T_31[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_5;
      end else if (8'h86 == _T_28[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_4;
      end else if (8'h86 == _T_25[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_3;
      end else if (8'h86 == _T_22[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_2;
      end else if (8'h86 == _T_19[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_1;
      end else if (8'h86 == _T_15[7:0]) begin
        image_0_134 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_135 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h87 == _T_34[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_6;
      end else if (8'h87 == _T_31[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_5;
      end else if (8'h87 == _T_28[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_4;
      end else if (8'h87 == _T_25[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_3;
      end else if (8'h87 == _T_22[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_2;
      end else if (8'h87 == _T_19[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_1;
      end else if (8'h87 == _T_15[7:0]) begin
        image_0_135 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_136 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h88 == _T_34[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_6;
      end else if (8'h88 == _T_31[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_5;
      end else if (8'h88 == _T_28[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_4;
      end else if (8'h88 == _T_25[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_3;
      end else if (8'h88 == _T_22[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_2;
      end else if (8'h88 == _T_19[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_1;
      end else if (8'h88 == _T_15[7:0]) begin
        image_0_136 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_137 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h89 == _T_34[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_6;
      end else if (8'h89 == _T_31[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_5;
      end else if (8'h89 == _T_28[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_4;
      end else if (8'h89 == _T_25[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_3;
      end else if (8'h89 == _T_22[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_2;
      end else if (8'h89 == _T_19[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_1;
      end else if (8'h89 == _T_15[7:0]) begin
        image_0_137 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_138 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8a == _T_34[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_6;
      end else if (8'h8a == _T_31[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_5;
      end else if (8'h8a == _T_28[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_4;
      end else if (8'h8a == _T_25[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_3;
      end else if (8'h8a == _T_22[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_2;
      end else if (8'h8a == _T_19[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_1;
      end else if (8'h8a == _T_15[7:0]) begin
        image_0_138 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_139 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8b == _T_34[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_6;
      end else if (8'h8b == _T_31[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_5;
      end else if (8'h8b == _T_28[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_4;
      end else if (8'h8b == _T_25[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_3;
      end else if (8'h8b == _T_22[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_2;
      end else if (8'h8b == _T_19[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_1;
      end else if (8'h8b == _T_15[7:0]) begin
        image_0_139 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_140 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8c == _T_34[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_6;
      end else if (8'h8c == _T_31[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_5;
      end else if (8'h8c == _T_28[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_4;
      end else if (8'h8c == _T_25[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_3;
      end else if (8'h8c == _T_22[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_2;
      end else if (8'h8c == _T_19[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_1;
      end else if (8'h8c == _T_15[7:0]) begin
        image_0_140 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_141 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8d == _T_34[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_6;
      end else if (8'h8d == _T_31[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_5;
      end else if (8'h8d == _T_28[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_4;
      end else if (8'h8d == _T_25[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_3;
      end else if (8'h8d == _T_22[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_2;
      end else if (8'h8d == _T_19[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_1;
      end else if (8'h8d == _T_15[7:0]) begin
        image_0_141 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_142 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8e == _T_34[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_6;
      end else if (8'h8e == _T_31[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_5;
      end else if (8'h8e == _T_28[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_4;
      end else if (8'h8e == _T_25[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_3;
      end else if (8'h8e == _T_22[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_2;
      end else if (8'h8e == _T_19[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_1;
      end else if (8'h8e == _T_15[7:0]) begin
        image_0_142 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_143 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h8f == _T_34[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_6;
      end else if (8'h8f == _T_31[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_5;
      end else if (8'h8f == _T_28[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_4;
      end else if (8'h8f == _T_25[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_3;
      end else if (8'h8f == _T_22[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_2;
      end else if (8'h8f == _T_19[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_1;
      end else if (8'h8f == _T_15[7:0]) begin
        image_0_143 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_144 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h90 == _T_34[7:0]) begin
        image_0_144 <= io_pixelVal_in_0_6;
      end else if (8'h90 == _T_31[7:0]) begin
        image_0_144 <= io_pixelVal_in_0_5;
      end else if (8'h90 == _T_28[7:0]) begin
        image_0_144 <= io_pixelVal_in_0_4;
      end else if (8'h90 == _T_25[7:0]) begin
        image_0_144 <= io_pixelVal_in_0_3;
      end else if (8'h90 == _T_22[7:0]) begin
        image_0_144 <= io_pixelVal_in_0_2;
      end else if (8'h90 == _T_19[7:0]) begin
        image_0_144 <= io_pixelVal_in_0_1;
      end else if (8'h90 == _T_15[7:0]) begin
        image_0_144 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_145 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h91 == _T_34[7:0]) begin
        image_0_145 <= io_pixelVal_in_0_6;
      end else if (8'h91 == _T_31[7:0]) begin
        image_0_145 <= io_pixelVal_in_0_5;
      end else if (8'h91 == _T_28[7:0]) begin
        image_0_145 <= io_pixelVal_in_0_4;
      end else if (8'h91 == _T_25[7:0]) begin
        image_0_145 <= io_pixelVal_in_0_3;
      end else if (8'h91 == _T_22[7:0]) begin
        image_0_145 <= io_pixelVal_in_0_2;
      end else if (8'h91 == _T_19[7:0]) begin
        image_0_145 <= io_pixelVal_in_0_1;
      end else if (8'h91 == _T_15[7:0]) begin
        image_0_145 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_146 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h92 == _T_34[7:0]) begin
        image_0_146 <= io_pixelVal_in_0_6;
      end else if (8'h92 == _T_31[7:0]) begin
        image_0_146 <= io_pixelVal_in_0_5;
      end else if (8'h92 == _T_28[7:0]) begin
        image_0_146 <= io_pixelVal_in_0_4;
      end else if (8'h92 == _T_25[7:0]) begin
        image_0_146 <= io_pixelVal_in_0_3;
      end else if (8'h92 == _T_22[7:0]) begin
        image_0_146 <= io_pixelVal_in_0_2;
      end else if (8'h92 == _T_19[7:0]) begin
        image_0_146 <= io_pixelVal_in_0_1;
      end else if (8'h92 == _T_15[7:0]) begin
        image_0_146 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_147 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h93 == _T_34[7:0]) begin
        image_0_147 <= io_pixelVal_in_0_6;
      end else if (8'h93 == _T_31[7:0]) begin
        image_0_147 <= io_pixelVal_in_0_5;
      end else if (8'h93 == _T_28[7:0]) begin
        image_0_147 <= io_pixelVal_in_0_4;
      end else if (8'h93 == _T_25[7:0]) begin
        image_0_147 <= io_pixelVal_in_0_3;
      end else if (8'h93 == _T_22[7:0]) begin
        image_0_147 <= io_pixelVal_in_0_2;
      end else if (8'h93 == _T_19[7:0]) begin
        image_0_147 <= io_pixelVal_in_0_1;
      end else if (8'h93 == _T_15[7:0]) begin
        image_0_147 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_148 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h94 == _T_34[7:0]) begin
        image_0_148 <= io_pixelVal_in_0_6;
      end else if (8'h94 == _T_31[7:0]) begin
        image_0_148 <= io_pixelVal_in_0_5;
      end else if (8'h94 == _T_28[7:0]) begin
        image_0_148 <= io_pixelVal_in_0_4;
      end else if (8'h94 == _T_25[7:0]) begin
        image_0_148 <= io_pixelVal_in_0_3;
      end else if (8'h94 == _T_22[7:0]) begin
        image_0_148 <= io_pixelVal_in_0_2;
      end else if (8'h94 == _T_19[7:0]) begin
        image_0_148 <= io_pixelVal_in_0_1;
      end else if (8'h94 == _T_15[7:0]) begin
        image_0_148 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_149 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h95 == _T_34[7:0]) begin
        image_0_149 <= io_pixelVal_in_0_6;
      end else if (8'h95 == _T_31[7:0]) begin
        image_0_149 <= io_pixelVal_in_0_5;
      end else if (8'h95 == _T_28[7:0]) begin
        image_0_149 <= io_pixelVal_in_0_4;
      end else if (8'h95 == _T_25[7:0]) begin
        image_0_149 <= io_pixelVal_in_0_3;
      end else if (8'h95 == _T_22[7:0]) begin
        image_0_149 <= io_pixelVal_in_0_2;
      end else if (8'h95 == _T_19[7:0]) begin
        image_0_149 <= io_pixelVal_in_0_1;
      end else if (8'h95 == _T_15[7:0]) begin
        image_0_149 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_150 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h96 == _T_34[7:0]) begin
        image_0_150 <= io_pixelVal_in_0_6;
      end else if (8'h96 == _T_31[7:0]) begin
        image_0_150 <= io_pixelVal_in_0_5;
      end else if (8'h96 == _T_28[7:0]) begin
        image_0_150 <= io_pixelVal_in_0_4;
      end else if (8'h96 == _T_25[7:0]) begin
        image_0_150 <= io_pixelVal_in_0_3;
      end else if (8'h96 == _T_22[7:0]) begin
        image_0_150 <= io_pixelVal_in_0_2;
      end else if (8'h96 == _T_19[7:0]) begin
        image_0_150 <= io_pixelVal_in_0_1;
      end else if (8'h96 == _T_15[7:0]) begin
        image_0_150 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_151 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h97 == _T_34[7:0]) begin
        image_0_151 <= io_pixelVal_in_0_6;
      end else if (8'h97 == _T_31[7:0]) begin
        image_0_151 <= io_pixelVal_in_0_5;
      end else if (8'h97 == _T_28[7:0]) begin
        image_0_151 <= io_pixelVal_in_0_4;
      end else if (8'h97 == _T_25[7:0]) begin
        image_0_151 <= io_pixelVal_in_0_3;
      end else if (8'h97 == _T_22[7:0]) begin
        image_0_151 <= io_pixelVal_in_0_2;
      end else if (8'h97 == _T_19[7:0]) begin
        image_0_151 <= io_pixelVal_in_0_1;
      end else if (8'h97 == _T_15[7:0]) begin
        image_0_151 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_152 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h98 == _T_34[7:0]) begin
        image_0_152 <= io_pixelVal_in_0_6;
      end else if (8'h98 == _T_31[7:0]) begin
        image_0_152 <= io_pixelVal_in_0_5;
      end else if (8'h98 == _T_28[7:0]) begin
        image_0_152 <= io_pixelVal_in_0_4;
      end else if (8'h98 == _T_25[7:0]) begin
        image_0_152 <= io_pixelVal_in_0_3;
      end else if (8'h98 == _T_22[7:0]) begin
        image_0_152 <= io_pixelVal_in_0_2;
      end else if (8'h98 == _T_19[7:0]) begin
        image_0_152 <= io_pixelVal_in_0_1;
      end else if (8'h98 == _T_15[7:0]) begin
        image_0_152 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_153 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h99 == _T_34[7:0]) begin
        image_0_153 <= io_pixelVal_in_0_6;
      end else if (8'h99 == _T_31[7:0]) begin
        image_0_153 <= io_pixelVal_in_0_5;
      end else if (8'h99 == _T_28[7:0]) begin
        image_0_153 <= io_pixelVal_in_0_4;
      end else if (8'h99 == _T_25[7:0]) begin
        image_0_153 <= io_pixelVal_in_0_3;
      end else if (8'h99 == _T_22[7:0]) begin
        image_0_153 <= io_pixelVal_in_0_2;
      end else if (8'h99 == _T_19[7:0]) begin
        image_0_153 <= io_pixelVal_in_0_1;
      end else if (8'h99 == _T_15[7:0]) begin
        image_0_153 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_154 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h9a == _T_34[7:0]) begin
        image_0_154 <= io_pixelVal_in_0_6;
      end else if (8'h9a == _T_31[7:0]) begin
        image_0_154 <= io_pixelVal_in_0_5;
      end else if (8'h9a == _T_28[7:0]) begin
        image_0_154 <= io_pixelVal_in_0_4;
      end else if (8'h9a == _T_25[7:0]) begin
        image_0_154 <= io_pixelVal_in_0_3;
      end else if (8'h9a == _T_22[7:0]) begin
        image_0_154 <= io_pixelVal_in_0_2;
      end else if (8'h9a == _T_19[7:0]) begin
        image_0_154 <= io_pixelVal_in_0_1;
      end else if (8'h9a == _T_15[7:0]) begin
        image_0_154 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_155 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h9b == _T_34[7:0]) begin
        image_0_155 <= io_pixelVal_in_0_6;
      end else if (8'h9b == _T_31[7:0]) begin
        image_0_155 <= io_pixelVal_in_0_5;
      end else if (8'h9b == _T_28[7:0]) begin
        image_0_155 <= io_pixelVal_in_0_4;
      end else if (8'h9b == _T_25[7:0]) begin
        image_0_155 <= io_pixelVal_in_0_3;
      end else if (8'h9b == _T_22[7:0]) begin
        image_0_155 <= io_pixelVal_in_0_2;
      end else if (8'h9b == _T_19[7:0]) begin
        image_0_155 <= io_pixelVal_in_0_1;
      end else if (8'h9b == _T_15[7:0]) begin
        image_0_155 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_156 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h9c == _T_34[7:0]) begin
        image_0_156 <= io_pixelVal_in_0_6;
      end else if (8'h9c == _T_31[7:0]) begin
        image_0_156 <= io_pixelVal_in_0_5;
      end else if (8'h9c == _T_28[7:0]) begin
        image_0_156 <= io_pixelVal_in_0_4;
      end else if (8'h9c == _T_25[7:0]) begin
        image_0_156 <= io_pixelVal_in_0_3;
      end else if (8'h9c == _T_22[7:0]) begin
        image_0_156 <= io_pixelVal_in_0_2;
      end else if (8'h9c == _T_19[7:0]) begin
        image_0_156 <= io_pixelVal_in_0_1;
      end else if (8'h9c == _T_15[7:0]) begin
        image_0_156 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_157 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h9d == _T_34[7:0]) begin
        image_0_157 <= io_pixelVal_in_0_6;
      end else if (8'h9d == _T_31[7:0]) begin
        image_0_157 <= io_pixelVal_in_0_5;
      end else if (8'h9d == _T_28[7:0]) begin
        image_0_157 <= io_pixelVal_in_0_4;
      end else if (8'h9d == _T_25[7:0]) begin
        image_0_157 <= io_pixelVal_in_0_3;
      end else if (8'h9d == _T_22[7:0]) begin
        image_0_157 <= io_pixelVal_in_0_2;
      end else if (8'h9d == _T_19[7:0]) begin
        image_0_157 <= io_pixelVal_in_0_1;
      end else if (8'h9d == _T_15[7:0]) begin
        image_0_157 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_158 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h9e == _T_34[7:0]) begin
        image_0_158 <= io_pixelVal_in_0_6;
      end else if (8'h9e == _T_31[7:0]) begin
        image_0_158 <= io_pixelVal_in_0_5;
      end else if (8'h9e == _T_28[7:0]) begin
        image_0_158 <= io_pixelVal_in_0_4;
      end else if (8'h9e == _T_25[7:0]) begin
        image_0_158 <= io_pixelVal_in_0_3;
      end else if (8'h9e == _T_22[7:0]) begin
        image_0_158 <= io_pixelVal_in_0_2;
      end else if (8'h9e == _T_19[7:0]) begin
        image_0_158 <= io_pixelVal_in_0_1;
      end else if (8'h9e == _T_15[7:0]) begin
        image_0_158 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_159 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'h9f == _T_34[7:0]) begin
        image_0_159 <= io_pixelVal_in_0_6;
      end else if (8'h9f == _T_31[7:0]) begin
        image_0_159 <= io_pixelVal_in_0_5;
      end else if (8'h9f == _T_28[7:0]) begin
        image_0_159 <= io_pixelVal_in_0_4;
      end else if (8'h9f == _T_25[7:0]) begin
        image_0_159 <= io_pixelVal_in_0_3;
      end else if (8'h9f == _T_22[7:0]) begin
        image_0_159 <= io_pixelVal_in_0_2;
      end else if (8'h9f == _T_19[7:0]) begin
        image_0_159 <= io_pixelVal_in_0_1;
      end else if (8'h9f == _T_15[7:0]) begin
        image_0_159 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_160 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha0 == _T_34[7:0]) begin
        image_0_160 <= io_pixelVal_in_0_6;
      end else if (8'ha0 == _T_31[7:0]) begin
        image_0_160 <= io_pixelVal_in_0_5;
      end else if (8'ha0 == _T_28[7:0]) begin
        image_0_160 <= io_pixelVal_in_0_4;
      end else if (8'ha0 == _T_25[7:0]) begin
        image_0_160 <= io_pixelVal_in_0_3;
      end else if (8'ha0 == _T_22[7:0]) begin
        image_0_160 <= io_pixelVal_in_0_2;
      end else if (8'ha0 == _T_19[7:0]) begin
        image_0_160 <= io_pixelVal_in_0_1;
      end else if (8'ha0 == _T_15[7:0]) begin
        image_0_160 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_161 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha1 == _T_34[7:0]) begin
        image_0_161 <= io_pixelVal_in_0_6;
      end else if (8'ha1 == _T_31[7:0]) begin
        image_0_161 <= io_pixelVal_in_0_5;
      end else if (8'ha1 == _T_28[7:0]) begin
        image_0_161 <= io_pixelVal_in_0_4;
      end else if (8'ha1 == _T_25[7:0]) begin
        image_0_161 <= io_pixelVal_in_0_3;
      end else if (8'ha1 == _T_22[7:0]) begin
        image_0_161 <= io_pixelVal_in_0_2;
      end else if (8'ha1 == _T_19[7:0]) begin
        image_0_161 <= io_pixelVal_in_0_1;
      end else if (8'ha1 == _T_15[7:0]) begin
        image_0_161 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_162 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha2 == _T_34[7:0]) begin
        image_0_162 <= io_pixelVal_in_0_6;
      end else if (8'ha2 == _T_31[7:0]) begin
        image_0_162 <= io_pixelVal_in_0_5;
      end else if (8'ha2 == _T_28[7:0]) begin
        image_0_162 <= io_pixelVal_in_0_4;
      end else if (8'ha2 == _T_25[7:0]) begin
        image_0_162 <= io_pixelVal_in_0_3;
      end else if (8'ha2 == _T_22[7:0]) begin
        image_0_162 <= io_pixelVal_in_0_2;
      end else if (8'ha2 == _T_19[7:0]) begin
        image_0_162 <= io_pixelVal_in_0_1;
      end else if (8'ha2 == _T_15[7:0]) begin
        image_0_162 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_163 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha3 == _T_34[7:0]) begin
        image_0_163 <= io_pixelVal_in_0_6;
      end else if (8'ha3 == _T_31[7:0]) begin
        image_0_163 <= io_pixelVal_in_0_5;
      end else if (8'ha3 == _T_28[7:0]) begin
        image_0_163 <= io_pixelVal_in_0_4;
      end else if (8'ha3 == _T_25[7:0]) begin
        image_0_163 <= io_pixelVal_in_0_3;
      end else if (8'ha3 == _T_22[7:0]) begin
        image_0_163 <= io_pixelVal_in_0_2;
      end else if (8'ha3 == _T_19[7:0]) begin
        image_0_163 <= io_pixelVal_in_0_1;
      end else if (8'ha3 == _T_15[7:0]) begin
        image_0_163 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_164 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha4 == _T_34[7:0]) begin
        image_0_164 <= io_pixelVal_in_0_6;
      end else if (8'ha4 == _T_31[7:0]) begin
        image_0_164 <= io_pixelVal_in_0_5;
      end else if (8'ha4 == _T_28[7:0]) begin
        image_0_164 <= io_pixelVal_in_0_4;
      end else if (8'ha4 == _T_25[7:0]) begin
        image_0_164 <= io_pixelVal_in_0_3;
      end else if (8'ha4 == _T_22[7:0]) begin
        image_0_164 <= io_pixelVal_in_0_2;
      end else if (8'ha4 == _T_19[7:0]) begin
        image_0_164 <= io_pixelVal_in_0_1;
      end else if (8'ha4 == _T_15[7:0]) begin
        image_0_164 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_165 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha5 == _T_34[7:0]) begin
        image_0_165 <= io_pixelVal_in_0_6;
      end else if (8'ha5 == _T_31[7:0]) begin
        image_0_165 <= io_pixelVal_in_0_5;
      end else if (8'ha5 == _T_28[7:0]) begin
        image_0_165 <= io_pixelVal_in_0_4;
      end else if (8'ha5 == _T_25[7:0]) begin
        image_0_165 <= io_pixelVal_in_0_3;
      end else if (8'ha5 == _T_22[7:0]) begin
        image_0_165 <= io_pixelVal_in_0_2;
      end else if (8'ha5 == _T_19[7:0]) begin
        image_0_165 <= io_pixelVal_in_0_1;
      end else if (8'ha5 == _T_15[7:0]) begin
        image_0_165 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_166 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha6 == _T_34[7:0]) begin
        image_0_166 <= io_pixelVal_in_0_6;
      end else if (8'ha6 == _T_31[7:0]) begin
        image_0_166 <= io_pixelVal_in_0_5;
      end else if (8'ha6 == _T_28[7:0]) begin
        image_0_166 <= io_pixelVal_in_0_4;
      end else if (8'ha6 == _T_25[7:0]) begin
        image_0_166 <= io_pixelVal_in_0_3;
      end else if (8'ha6 == _T_22[7:0]) begin
        image_0_166 <= io_pixelVal_in_0_2;
      end else if (8'ha6 == _T_19[7:0]) begin
        image_0_166 <= io_pixelVal_in_0_1;
      end else if (8'ha6 == _T_15[7:0]) begin
        image_0_166 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_167 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha7 == _T_34[7:0]) begin
        image_0_167 <= io_pixelVal_in_0_6;
      end else if (8'ha7 == _T_31[7:0]) begin
        image_0_167 <= io_pixelVal_in_0_5;
      end else if (8'ha7 == _T_28[7:0]) begin
        image_0_167 <= io_pixelVal_in_0_4;
      end else if (8'ha7 == _T_25[7:0]) begin
        image_0_167 <= io_pixelVal_in_0_3;
      end else if (8'ha7 == _T_22[7:0]) begin
        image_0_167 <= io_pixelVal_in_0_2;
      end else if (8'ha7 == _T_19[7:0]) begin
        image_0_167 <= io_pixelVal_in_0_1;
      end else if (8'ha7 == _T_15[7:0]) begin
        image_0_167 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_168 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha8 == _T_34[7:0]) begin
        image_0_168 <= io_pixelVal_in_0_6;
      end else if (8'ha8 == _T_31[7:0]) begin
        image_0_168 <= io_pixelVal_in_0_5;
      end else if (8'ha8 == _T_28[7:0]) begin
        image_0_168 <= io_pixelVal_in_0_4;
      end else if (8'ha8 == _T_25[7:0]) begin
        image_0_168 <= io_pixelVal_in_0_3;
      end else if (8'ha8 == _T_22[7:0]) begin
        image_0_168 <= io_pixelVal_in_0_2;
      end else if (8'ha8 == _T_19[7:0]) begin
        image_0_168 <= io_pixelVal_in_0_1;
      end else if (8'ha8 == _T_15[7:0]) begin
        image_0_168 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_169 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'ha9 == _T_34[7:0]) begin
        image_0_169 <= io_pixelVal_in_0_6;
      end else if (8'ha9 == _T_31[7:0]) begin
        image_0_169 <= io_pixelVal_in_0_5;
      end else if (8'ha9 == _T_28[7:0]) begin
        image_0_169 <= io_pixelVal_in_0_4;
      end else if (8'ha9 == _T_25[7:0]) begin
        image_0_169 <= io_pixelVal_in_0_3;
      end else if (8'ha9 == _T_22[7:0]) begin
        image_0_169 <= io_pixelVal_in_0_2;
      end else if (8'ha9 == _T_19[7:0]) begin
        image_0_169 <= io_pixelVal_in_0_1;
      end else if (8'ha9 == _T_15[7:0]) begin
        image_0_169 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_170 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'haa == _T_34[7:0]) begin
        image_0_170 <= io_pixelVal_in_0_6;
      end else if (8'haa == _T_31[7:0]) begin
        image_0_170 <= io_pixelVal_in_0_5;
      end else if (8'haa == _T_28[7:0]) begin
        image_0_170 <= io_pixelVal_in_0_4;
      end else if (8'haa == _T_25[7:0]) begin
        image_0_170 <= io_pixelVal_in_0_3;
      end else if (8'haa == _T_22[7:0]) begin
        image_0_170 <= io_pixelVal_in_0_2;
      end else if (8'haa == _T_19[7:0]) begin
        image_0_170 <= io_pixelVal_in_0_1;
      end else if (8'haa == _T_15[7:0]) begin
        image_0_170 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_171 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hab == _T_34[7:0]) begin
        image_0_171 <= io_pixelVal_in_0_6;
      end else if (8'hab == _T_31[7:0]) begin
        image_0_171 <= io_pixelVal_in_0_5;
      end else if (8'hab == _T_28[7:0]) begin
        image_0_171 <= io_pixelVal_in_0_4;
      end else if (8'hab == _T_25[7:0]) begin
        image_0_171 <= io_pixelVal_in_0_3;
      end else if (8'hab == _T_22[7:0]) begin
        image_0_171 <= io_pixelVal_in_0_2;
      end else if (8'hab == _T_19[7:0]) begin
        image_0_171 <= io_pixelVal_in_0_1;
      end else if (8'hab == _T_15[7:0]) begin
        image_0_171 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_172 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hac == _T_34[7:0]) begin
        image_0_172 <= io_pixelVal_in_0_6;
      end else if (8'hac == _T_31[7:0]) begin
        image_0_172 <= io_pixelVal_in_0_5;
      end else if (8'hac == _T_28[7:0]) begin
        image_0_172 <= io_pixelVal_in_0_4;
      end else if (8'hac == _T_25[7:0]) begin
        image_0_172 <= io_pixelVal_in_0_3;
      end else if (8'hac == _T_22[7:0]) begin
        image_0_172 <= io_pixelVal_in_0_2;
      end else if (8'hac == _T_19[7:0]) begin
        image_0_172 <= io_pixelVal_in_0_1;
      end else if (8'hac == _T_15[7:0]) begin
        image_0_172 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_173 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'had == _T_34[7:0]) begin
        image_0_173 <= io_pixelVal_in_0_6;
      end else if (8'had == _T_31[7:0]) begin
        image_0_173 <= io_pixelVal_in_0_5;
      end else if (8'had == _T_28[7:0]) begin
        image_0_173 <= io_pixelVal_in_0_4;
      end else if (8'had == _T_25[7:0]) begin
        image_0_173 <= io_pixelVal_in_0_3;
      end else if (8'had == _T_22[7:0]) begin
        image_0_173 <= io_pixelVal_in_0_2;
      end else if (8'had == _T_19[7:0]) begin
        image_0_173 <= io_pixelVal_in_0_1;
      end else if (8'had == _T_15[7:0]) begin
        image_0_173 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_174 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hae == _T_34[7:0]) begin
        image_0_174 <= io_pixelVal_in_0_6;
      end else if (8'hae == _T_31[7:0]) begin
        image_0_174 <= io_pixelVal_in_0_5;
      end else if (8'hae == _T_28[7:0]) begin
        image_0_174 <= io_pixelVal_in_0_4;
      end else if (8'hae == _T_25[7:0]) begin
        image_0_174 <= io_pixelVal_in_0_3;
      end else if (8'hae == _T_22[7:0]) begin
        image_0_174 <= io_pixelVal_in_0_2;
      end else if (8'hae == _T_19[7:0]) begin
        image_0_174 <= io_pixelVal_in_0_1;
      end else if (8'hae == _T_15[7:0]) begin
        image_0_174 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_175 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'haf == _T_34[7:0]) begin
        image_0_175 <= io_pixelVal_in_0_6;
      end else if (8'haf == _T_31[7:0]) begin
        image_0_175 <= io_pixelVal_in_0_5;
      end else if (8'haf == _T_28[7:0]) begin
        image_0_175 <= io_pixelVal_in_0_4;
      end else if (8'haf == _T_25[7:0]) begin
        image_0_175 <= io_pixelVal_in_0_3;
      end else if (8'haf == _T_22[7:0]) begin
        image_0_175 <= io_pixelVal_in_0_2;
      end else if (8'haf == _T_19[7:0]) begin
        image_0_175 <= io_pixelVal_in_0_1;
      end else if (8'haf == _T_15[7:0]) begin
        image_0_175 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_176 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb0 == _T_34[7:0]) begin
        image_0_176 <= io_pixelVal_in_0_6;
      end else if (8'hb0 == _T_31[7:0]) begin
        image_0_176 <= io_pixelVal_in_0_5;
      end else if (8'hb0 == _T_28[7:0]) begin
        image_0_176 <= io_pixelVal_in_0_4;
      end else if (8'hb0 == _T_25[7:0]) begin
        image_0_176 <= io_pixelVal_in_0_3;
      end else if (8'hb0 == _T_22[7:0]) begin
        image_0_176 <= io_pixelVal_in_0_2;
      end else if (8'hb0 == _T_19[7:0]) begin
        image_0_176 <= io_pixelVal_in_0_1;
      end else if (8'hb0 == _T_15[7:0]) begin
        image_0_176 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_177 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb1 == _T_34[7:0]) begin
        image_0_177 <= io_pixelVal_in_0_6;
      end else if (8'hb1 == _T_31[7:0]) begin
        image_0_177 <= io_pixelVal_in_0_5;
      end else if (8'hb1 == _T_28[7:0]) begin
        image_0_177 <= io_pixelVal_in_0_4;
      end else if (8'hb1 == _T_25[7:0]) begin
        image_0_177 <= io_pixelVal_in_0_3;
      end else if (8'hb1 == _T_22[7:0]) begin
        image_0_177 <= io_pixelVal_in_0_2;
      end else if (8'hb1 == _T_19[7:0]) begin
        image_0_177 <= io_pixelVal_in_0_1;
      end else if (8'hb1 == _T_15[7:0]) begin
        image_0_177 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_178 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb2 == _T_34[7:0]) begin
        image_0_178 <= io_pixelVal_in_0_6;
      end else if (8'hb2 == _T_31[7:0]) begin
        image_0_178 <= io_pixelVal_in_0_5;
      end else if (8'hb2 == _T_28[7:0]) begin
        image_0_178 <= io_pixelVal_in_0_4;
      end else if (8'hb2 == _T_25[7:0]) begin
        image_0_178 <= io_pixelVal_in_0_3;
      end else if (8'hb2 == _T_22[7:0]) begin
        image_0_178 <= io_pixelVal_in_0_2;
      end else if (8'hb2 == _T_19[7:0]) begin
        image_0_178 <= io_pixelVal_in_0_1;
      end else if (8'hb2 == _T_15[7:0]) begin
        image_0_178 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_179 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb3 == _T_34[7:0]) begin
        image_0_179 <= io_pixelVal_in_0_6;
      end else if (8'hb3 == _T_31[7:0]) begin
        image_0_179 <= io_pixelVal_in_0_5;
      end else if (8'hb3 == _T_28[7:0]) begin
        image_0_179 <= io_pixelVal_in_0_4;
      end else if (8'hb3 == _T_25[7:0]) begin
        image_0_179 <= io_pixelVal_in_0_3;
      end else if (8'hb3 == _T_22[7:0]) begin
        image_0_179 <= io_pixelVal_in_0_2;
      end else if (8'hb3 == _T_19[7:0]) begin
        image_0_179 <= io_pixelVal_in_0_1;
      end else if (8'hb3 == _T_15[7:0]) begin
        image_0_179 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_180 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb4 == _T_34[7:0]) begin
        image_0_180 <= io_pixelVal_in_0_6;
      end else if (8'hb4 == _T_31[7:0]) begin
        image_0_180 <= io_pixelVal_in_0_5;
      end else if (8'hb4 == _T_28[7:0]) begin
        image_0_180 <= io_pixelVal_in_0_4;
      end else if (8'hb4 == _T_25[7:0]) begin
        image_0_180 <= io_pixelVal_in_0_3;
      end else if (8'hb4 == _T_22[7:0]) begin
        image_0_180 <= io_pixelVal_in_0_2;
      end else if (8'hb4 == _T_19[7:0]) begin
        image_0_180 <= io_pixelVal_in_0_1;
      end else if (8'hb4 == _T_15[7:0]) begin
        image_0_180 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_181 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb5 == _T_34[7:0]) begin
        image_0_181 <= io_pixelVal_in_0_6;
      end else if (8'hb5 == _T_31[7:0]) begin
        image_0_181 <= io_pixelVal_in_0_5;
      end else if (8'hb5 == _T_28[7:0]) begin
        image_0_181 <= io_pixelVal_in_0_4;
      end else if (8'hb5 == _T_25[7:0]) begin
        image_0_181 <= io_pixelVal_in_0_3;
      end else if (8'hb5 == _T_22[7:0]) begin
        image_0_181 <= io_pixelVal_in_0_2;
      end else if (8'hb5 == _T_19[7:0]) begin
        image_0_181 <= io_pixelVal_in_0_1;
      end else if (8'hb5 == _T_15[7:0]) begin
        image_0_181 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_182 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb6 == _T_34[7:0]) begin
        image_0_182 <= io_pixelVal_in_0_6;
      end else if (8'hb6 == _T_31[7:0]) begin
        image_0_182 <= io_pixelVal_in_0_5;
      end else if (8'hb6 == _T_28[7:0]) begin
        image_0_182 <= io_pixelVal_in_0_4;
      end else if (8'hb6 == _T_25[7:0]) begin
        image_0_182 <= io_pixelVal_in_0_3;
      end else if (8'hb6 == _T_22[7:0]) begin
        image_0_182 <= io_pixelVal_in_0_2;
      end else if (8'hb6 == _T_19[7:0]) begin
        image_0_182 <= io_pixelVal_in_0_1;
      end else if (8'hb6 == _T_15[7:0]) begin
        image_0_182 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_183 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb7 == _T_34[7:0]) begin
        image_0_183 <= io_pixelVal_in_0_6;
      end else if (8'hb7 == _T_31[7:0]) begin
        image_0_183 <= io_pixelVal_in_0_5;
      end else if (8'hb7 == _T_28[7:0]) begin
        image_0_183 <= io_pixelVal_in_0_4;
      end else if (8'hb7 == _T_25[7:0]) begin
        image_0_183 <= io_pixelVal_in_0_3;
      end else if (8'hb7 == _T_22[7:0]) begin
        image_0_183 <= io_pixelVal_in_0_2;
      end else if (8'hb7 == _T_19[7:0]) begin
        image_0_183 <= io_pixelVal_in_0_1;
      end else if (8'hb7 == _T_15[7:0]) begin
        image_0_183 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_184 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb8 == _T_34[7:0]) begin
        image_0_184 <= io_pixelVal_in_0_6;
      end else if (8'hb8 == _T_31[7:0]) begin
        image_0_184 <= io_pixelVal_in_0_5;
      end else if (8'hb8 == _T_28[7:0]) begin
        image_0_184 <= io_pixelVal_in_0_4;
      end else if (8'hb8 == _T_25[7:0]) begin
        image_0_184 <= io_pixelVal_in_0_3;
      end else if (8'hb8 == _T_22[7:0]) begin
        image_0_184 <= io_pixelVal_in_0_2;
      end else if (8'hb8 == _T_19[7:0]) begin
        image_0_184 <= io_pixelVal_in_0_1;
      end else if (8'hb8 == _T_15[7:0]) begin
        image_0_184 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_185 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hb9 == _T_34[7:0]) begin
        image_0_185 <= io_pixelVal_in_0_6;
      end else if (8'hb9 == _T_31[7:0]) begin
        image_0_185 <= io_pixelVal_in_0_5;
      end else if (8'hb9 == _T_28[7:0]) begin
        image_0_185 <= io_pixelVal_in_0_4;
      end else if (8'hb9 == _T_25[7:0]) begin
        image_0_185 <= io_pixelVal_in_0_3;
      end else if (8'hb9 == _T_22[7:0]) begin
        image_0_185 <= io_pixelVal_in_0_2;
      end else if (8'hb9 == _T_19[7:0]) begin
        image_0_185 <= io_pixelVal_in_0_1;
      end else if (8'hb9 == _T_15[7:0]) begin
        image_0_185 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_186 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hba == _T_34[7:0]) begin
        image_0_186 <= io_pixelVal_in_0_6;
      end else if (8'hba == _T_31[7:0]) begin
        image_0_186 <= io_pixelVal_in_0_5;
      end else if (8'hba == _T_28[7:0]) begin
        image_0_186 <= io_pixelVal_in_0_4;
      end else if (8'hba == _T_25[7:0]) begin
        image_0_186 <= io_pixelVal_in_0_3;
      end else if (8'hba == _T_22[7:0]) begin
        image_0_186 <= io_pixelVal_in_0_2;
      end else if (8'hba == _T_19[7:0]) begin
        image_0_186 <= io_pixelVal_in_0_1;
      end else if (8'hba == _T_15[7:0]) begin
        image_0_186 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_187 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hbb == _T_34[7:0]) begin
        image_0_187 <= io_pixelVal_in_0_6;
      end else if (8'hbb == _T_31[7:0]) begin
        image_0_187 <= io_pixelVal_in_0_5;
      end else if (8'hbb == _T_28[7:0]) begin
        image_0_187 <= io_pixelVal_in_0_4;
      end else if (8'hbb == _T_25[7:0]) begin
        image_0_187 <= io_pixelVal_in_0_3;
      end else if (8'hbb == _T_22[7:0]) begin
        image_0_187 <= io_pixelVal_in_0_2;
      end else if (8'hbb == _T_19[7:0]) begin
        image_0_187 <= io_pixelVal_in_0_1;
      end else if (8'hbb == _T_15[7:0]) begin
        image_0_187 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_188 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hbc == _T_34[7:0]) begin
        image_0_188 <= io_pixelVal_in_0_6;
      end else if (8'hbc == _T_31[7:0]) begin
        image_0_188 <= io_pixelVal_in_0_5;
      end else if (8'hbc == _T_28[7:0]) begin
        image_0_188 <= io_pixelVal_in_0_4;
      end else if (8'hbc == _T_25[7:0]) begin
        image_0_188 <= io_pixelVal_in_0_3;
      end else if (8'hbc == _T_22[7:0]) begin
        image_0_188 <= io_pixelVal_in_0_2;
      end else if (8'hbc == _T_19[7:0]) begin
        image_0_188 <= io_pixelVal_in_0_1;
      end else if (8'hbc == _T_15[7:0]) begin
        image_0_188 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_189 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hbd == _T_34[7:0]) begin
        image_0_189 <= io_pixelVal_in_0_6;
      end else if (8'hbd == _T_31[7:0]) begin
        image_0_189 <= io_pixelVal_in_0_5;
      end else if (8'hbd == _T_28[7:0]) begin
        image_0_189 <= io_pixelVal_in_0_4;
      end else if (8'hbd == _T_25[7:0]) begin
        image_0_189 <= io_pixelVal_in_0_3;
      end else if (8'hbd == _T_22[7:0]) begin
        image_0_189 <= io_pixelVal_in_0_2;
      end else if (8'hbd == _T_19[7:0]) begin
        image_0_189 <= io_pixelVal_in_0_1;
      end else if (8'hbd == _T_15[7:0]) begin
        image_0_189 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_190 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hbe == _T_34[7:0]) begin
        image_0_190 <= io_pixelVal_in_0_6;
      end else if (8'hbe == _T_31[7:0]) begin
        image_0_190 <= io_pixelVal_in_0_5;
      end else if (8'hbe == _T_28[7:0]) begin
        image_0_190 <= io_pixelVal_in_0_4;
      end else if (8'hbe == _T_25[7:0]) begin
        image_0_190 <= io_pixelVal_in_0_3;
      end else if (8'hbe == _T_22[7:0]) begin
        image_0_190 <= io_pixelVal_in_0_2;
      end else if (8'hbe == _T_19[7:0]) begin
        image_0_190 <= io_pixelVal_in_0_1;
      end else if (8'hbe == _T_15[7:0]) begin
        image_0_190 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_191 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hbf == _T_34[7:0]) begin
        image_0_191 <= io_pixelVal_in_0_6;
      end else if (8'hbf == _T_31[7:0]) begin
        image_0_191 <= io_pixelVal_in_0_5;
      end else if (8'hbf == _T_28[7:0]) begin
        image_0_191 <= io_pixelVal_in_0_4;
      end else if (8'hbf == _T_25[7:0]) begin
        image_0_191 <= io_pixelVal_in_0_3;
      end else if (8'hbf == _T_22[7:0]) begin
        image_0_191 <= io_pixelVal_in_0_2;
      end else if (8'hbf == _T_19[7:0]) begin
        image_0_191 <= io_pixelVal_in_0_1;
      end else if (8'hbf == _T_15[7:0]) begin
        image_0_191 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_192 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hc0 == _T_34[7:0]) begin
        image_0_192 <= io_pixelVal_in_0_6;
      end else if (8'hc0 == _T_31[7:0]) begin
        image_0_192 <= io_pixelVal_in_0_5;
      end else if (8'hc0 == _T_28[7:0]) begin
        image_0_192 <= io_pixelVal_in_0_4;
      end else if (8'hc0 == _T_25[7:0]) begin
        image_0_192 <= io_pixelVal_in_0_3;
      end else if (8'hc0 == _T_22[7:0]) begin
        image_0_192 <= io_pixelVal_in_0_2;
      end else if (8'hc0 == _T_19[7:0]) begin
        image_0_192 <= io_pixelVal_in_0_1;
      end else if (8'hc0 == _T_15[7:0]) begin
        image_0_192 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_193 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hc1 == _T_34[7:0]) begin
        image_0_193 <= io_pixelVal_in_0_6;
      end else if (8'hc1 == _T_31[7:0]) begin
        image_0_193 <= io_pixelVal_in_0_5;
      end else if (8'hc1 == _T_28[7:0]) begin
        image_0_193 <= io_pixelVal_in_0_4;
      end else if (8'hc1 == _T_25[7:0]) begin
        image_0_193 <= io_pixelVal_in_0_3;
      end else if (8'hc1 == _T_22[7:0]) begin
        image_0_193 <= io_pixelVal_in_0_2;
      end else if (8'hc1 == _T_19[7:0]) begin
        image_0_193 <= io_pixelVal_in_0_1;
      end else if (8'hc1 == _T_15[7:0]) begin
        image_0_193 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_194 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hc2 == _T_34[7:0]) begin
        image_0_194 <= io_pixelVal_in_0_6;
      end else if (8'hc2 == _T_31[7:0]) begin
        image_0_194 <= io_pixelVal_in_0_5;
      end else if (8'hc2 == _T_28[7:0]) begin
        image_0_194 <= io_pixelVal_in_0_4;
      end else if (8'hc2 == _T_25[7:0]) begin
        image_0_194 <= io_pixelVal_in_0_3;
      end else if (8'hc2 == _T_22[7:0]) begin
        image_0_194 <= io_pixelVal_in_0_2;
      end else if (8'hc2 == _T_19[7:0]) begin
        image_0_194 <= io_pixelVal_in_0_1;
      end else if (8'hc2 == _T_15[7:0]) begin
        image_0_194 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_195 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hc3 == _T_34[7:0]) begin
        image_0_195 <= io_pixelVal_in_0_6;
      end else if (8'hc3 == _T_31[7:0]) begin
        image_0_195 <= io_pixelVal_in_0_5;
      end else if (8'hc3 == _T_28[7:0]) begin
        image_0_195 <= io_pixelVal_in_0_4;
      end else if (8'hc3 == _T_25[7:0]) begin
        image_0_195 <= io_pixelVal_in_0_3;
      end else if (8'hc3 == _T_22[7:0]) begin
        image_0_195 <= io_pixelVal_in_0_2;
      end else if (8'hc3 == _T_19[7:0]) begin
        image_0_195 <= io_pixelVal_in_0_1;
      end else if (8'hc3 == _T_15[7:0]) begin
        image_0_195 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_196 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hc4 == _T_34[7:0]) begin
        image_0_196 <= io_pixelVal_in_0_6;
      end else if (8'hc4 == _T_31[7:0]) begin
        image_0_196 <= io_pixelVal_in_0_5;
      end else if (8'hc4 == _T_28[7:0]) begin
        image_0_196 <= io_pixelVal_in_0_4;
      end else if (8'hc4 == _T_25[7:0]) begin
        image_0_196 <= io_pixelVal_in_0_3;
      end else if (8'hc4 == _T_22[7:0]) begin
        image_0_196 <= io_pixelVal_in_0_2;
      end else if (8'hc4 == _T_19[7:0]) begin
        image_0_196 <= io_pixelVal_in_0_1;
      end else if (8'hc4 == _T_15[7:0]) begin
        image_0_196 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_197 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hc5 == _T_34[7:0]) begin
        image_0_197 <= io_pixelVal_in_0_6;
      end else if (8'hc5 == _T_31[7:0]) begin
        image_0_197 <= io_pixelVal_in_0_5;
      end else if (8'hc5 == _T_28[7:0]) begin
        image_0_197 <= io_pixelVal_in_0_4;
      end else if (8'hc5 == _T_25[7:0]) begin
        image_0_197 <= io_pixelVal_in_0_3;
      end else if (8'hc5 == _T_22[7:0]) begin
        image_0_197 <= io_pixelVal_in_0_2;
      end else if (8'hc5 == _T_19[7:0]) begin
        image_0_197 <= io_pixelVal_in_0_1;
      end else if (8'hc5 == _T_15[7:0]) begin
        image_0_197 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_198 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hc6 == _T_34[7:0]) begin
        image_0_198 <= io_pixelVal_in_0_6;
      end else if (8'hc6 == _T_31[7:0]) begin
        image_0_198 <= io_pixelVal_in_0_5;
      end else if (8'hc6 == _T_28[7:0]) begin
        image_0_198 <= io_pixelVal_in_0_4;
      end else if (8'hc6 == _T_25[7:0]) begin
        image_0_198 <= io_pixelVal_in_0_3;
      end else if (8'hc6 == _T_22[7:0]) begin
        image_0_198 <= io_pixelVal_in_0_2;
      end else if (8'hc6 == _T_19[7:0]) begin
        image_0_198 <= io_pixelVal_in_0_1;
      end else if (8'hc6 == _T_15[7:0]) begin
        image_0_198 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_199 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hc7 == _T_34[7:0]) begin
        image_0_199 <= io_pixelVal_in_0_6;
      end else if (8'hc7 == _T_31[7:0]) begin
        image_0_199 <= io_pixelVal_in_0_5;
      end else if (8'hc7 == _T_28[7:0]) begin
        image_0_199 <= io_pixelVal_in_0_4;
      end else if (8'hc7 == _T_25[7:0]) begin
        image_0_199 <= io_pixelVal_in_0_3;
      end else if (8'hc7 == _T_22[7:0]) begin
        image_0_199 <= io_pixelVal_in_0_2;
      end else if (8'hc7 == _T_19[7:0]) begin
        image_0_199 <= io_pixelVal_in_0_1;
      end else if (8'hc7 == _T_15[7:0]) begin
        image_0_199 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_200 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hc8 == _T_34[7:0]) begin
        image_0_200 <= io_pixelVal_in_0_6;
      end else if (8'hc8 == _T_31[7:0]) begin
        image_0_200 <= io_pixelVal_in_0_5;
      end else if (8'hc8 == _T_28[7:0]) begin
        image_0_200 <= io_pixelVal_in_0_4;
      end else if (8'hc8 == _T_25[7:0]) begin
        image_0_200 <= io_pixelVal_in_0_3;
      end else if (8'hc8 == _T_22[7:0]) begin
        image_0_200 <= io_pixelVal_in_0_2;
      end else if (8'hc8 == _T_19[7:0]) begin
        image_0_200 <= io_pixelVal_in_0_1;
      end else if (8'hc8 == _T_15[7:0]) begin
        image_0_200 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_201 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hc9 == _T_34[7:0]) begin
        image_0_201 <= io_pixelVal_in_0_6;
      end else if (8'hc9 == _T_31[7:0]) begin
        image_0_201 <= io_pixelVal_in_0_5;
      end else if (8'hc9 == _T_28[7:0]) begin
        image_0_201 <= io_pixelVal_in_0_4;
      end else if (8'hc9 == _T_25[7:0]) begin
        image_0_201 <= io_pixelVal_in_0_3;
      end else if (8'hc9 == _T_22[7:0]) begin
        image_0_201 <= io_pixelVal_in_0_2;
      end else if (8'hc9 == _T_19[7:0]) begin
        image_0_201 <= io_pixelVal_in_0_1;
      end else if (8'hc9 == _T_15[7:0]) begin
        image_0_201 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_202 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hca == _T_34[7:0]) begin
        image_0_202 <= io_pixelVal_in_0_6;
      end else if (8'hca == _T_31[7:0]) begin
        image_0_202 <= io_pixelVal_in_0_5;
      end else if (8'hca == _T_28[7:0]) begin
        image_0_202 <= io_pixelVal_in_0_4;
      end else if (8'hca == _T_25[7:0]) begin
        image_0_202 <= io_pixelVal_in_0_3;
      end else if (8'hca == _T_22[7:0]) begin
        image_0_202 <= io_pixelVal_in_0_2;
      end else if (8'hca == _T_19[7:0]) begin
        image_0_202 <= io_pixelVal_in_0_1;
      end else if (8'hca == _T_15[7:0]) begin
        image_0_202 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_203 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hcb == _T_34[7:0]) begin
        image_0_203 <= io_pixelVal_in_0_6;
      end else if (8'hcb == _T_31[7:0]) begin
        image_0_203 <= io_pixelVal_in_0_5;
      end else if (8'hcb == _T_28[7:0]) begin
        image_0_203 <= io_pixelVal_in_0_4;
      end else if (8'hcb == _T_25[7:0]) begin
        image_0_203 <= io_pixelVal_in_0_3;
      end else if (8'hcb == _T_22[7:0]) begin
        image_0_203 <= io_pixelVal_in_0_2;
      end else if (8'hcb == _T_19[7:0]) begin
        image_0_203 <= io_pixelVal_in_0_1;
      end else if (8'hcb == _T_15[7:0]) begin
        image_0_203 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_204 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hcc == _T_34[7:0]) begin
        image_0_204 <= io_pixelVal_in_0_6;
      end else if (8'hcc == _T_31[7:0]) begin
        image_0_204 <= io_pixelVal_in_0_5;
      end else if (8'hcc == _T_28[7:0]) begin
        image_0_204 <= io_pixelVal_in_0_4;
      end else if (8'hcc == _T_25[7:0]) begin
        image_0_204 <= io_pixelVal_in_0_3;
      end else if (8'hcc == _T_22[7:0]) begin
        image_0_204 <= io_pixelVal_in_0_2;
      end else if (8'hcc == _T_19[7:0]) begin
        image_0_204 <= io_pixelVal_in_0_1;
      end else if (8'hcc == _T_15[7:0]) begin
        image_0_204 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_205 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hcd == _T_34[7:0]) begin
        image_0_205 <= io_pixelVal_in_0_6;
      end else if (8'hcd == _T_31[7:0]) begin
        image_0_205 <= io_pixelVal_in_0_5;
      end else if (8'hcd == _T_28[7:0]) begin
        image_0_205 <= io_pixelVal_in_0_4;
      end else if (8'hcd == _T_25[7:0]) begin
        image_0_205 <= io_pixelVal_in_0_3;
      end else if (8'hcd == _T_22[7:0]) begin
        image_0_205 <= io_pixelVal_in_0_2;
      end else if (8'hcd == _T_19[7:0]) begin
        image_0_205 <= io_pixelVal_in_0_1;
      end else if (8'hcd == _T_15[7:0]) begin
        image_0_205 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_206 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hce == _T_34[7:0]) begin
        image_0_206 <= io_pixelVal_in_0_6;
      end else if (8'hce == _T_31[7:0]) begin
        image_0_206 <= io_pixelVal_in_0_5;
      end else if (8'hce == _T_28[7:0]) begin
        image_0_206 <= io_pixelVal_in_0_4;
      end else if (8'hce == _T_25[7:0]) begin
        image_0_206 <= io_pixelVal_in_0_3;
      end else if (8'hce == _T_22[7:0]) begin
        image_0_206 <= io_pixelVal_in_0_2;
      end else if (8'hce == _T_19[7:0]) begin
        image_0_206 <= io_pixelVal_in_0_1;
      end else if (8'hce == _T_15[7:0]) begin
        image_0_206 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_207 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hcf == _T_34[7:0]) begin
        image_0_207 <= io_pixelVal_in_0_6;
      end else if (8'hcf == _T_31[7:0]) begin
        image_0_207 <= io_pixelVal_in_0_5;
      end else if (8'hcf == _T_28[7:0]) begin
        image_0_207 <= io_pixelVal_in_0_4;
      end else if (8'hcf == _T_25[7:0]) begin
        image_0_207 <= io_pixelVal_in_0_3;
      end else if (8'hcf == _T_22[7:0]) begin
        image_0_207 <= io_pixelVal_in_0_2;
      end else if (8'hcf == _T_19[7:0]) begin
        image_0_207 <= io_pixelVal_in_0_1;
      end else if (8'hcf == _T_15[7:0]) begin
        image_0_207 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_208 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hd0 == _T_34[7:0]) begin
        image_0_208 <= io_pixelVal_in_0_6;
      end else if (8'hd0 == _T_31[7:0]) begin
        image_0_208 <= io_pixelVal_in_0_5;
      end else if (8'hd0 == _T_28[7:0]) begin
        image_0_208 <= io_pixelVal_in_0_4;
      end else if (8'hd0 == _T_25[7:0]) begin
        image_0_208 <= io_pixelVal_in_0_3;
      end else if (8'hd0 == _T_22[7:0]) begin
        image_0_208 <= io_pixelVal_in_0_2;
      end else if (8'hd0 == _T_19[7:0]) begin
        image_0_208 <= io_pixelVal_in_0_1;
      end else if (8'hd0 == _T_15[7:0]) begin
        image_0_208 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_209 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hd1 == _T_34[7:0]) begin
        image_0_209 <= io_pixelVal_in_0_6;
      end else if (8'hd1 == _T_31[7:0]) begin
        image_0_209 <= io_pixelVal_in_0_5;
      end else if (8'hd1 == _T_28[7:0]) begin
        image_0_209 <= io_pixelVal_in_0_4;
      end else if (8'hd1 == _T_25[7:0]) begin
        image_0_209 <= io_pixelVal_in_0_3;
      end else if (8'hd1 == _T_22[7:0]) begin
        image_0_209 <= io_pixelVal_in_0_2;
      end else if (8'hd1 == _T_19[7:0]) begin
        image_0_209 <= io_pixelVal_in_0_1;
      end else if (8'hd1 == _T_15[7:0]) begin
        image_0_209 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_210 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hd2 == _T_34[7:0]) begin
        image_0_210 <= io_pixelVal_in_0_6;
      end else if (8'hd2 == _T_31[7:0]) begin
        image_0_210 <= io_pixelVal_in_0_5;
      end else if (8'hd2 == _T_28[7:0]) begin
        image_0_210 <= io_pixelVal_in_0_4;
      end else if (8'hd2 == _T_25[7:0]) begin
        image_0_210 <= io_pixelVal_in_0_3;
      end else if (8'hd2 == _T_22[7:0]) begin
        image_0_210 <= io_pixelVal_in_0_2;
      end else if (8'hd2 == _T_19[7:0]) begin
        image_0_210 <= io_pixelVal_in_0_1;
      end else if (8'hd2 == _T_15[7:0]) begin
        image_0_210 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_211 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hd3 == _T_34[7:0]) begin
        image_0_211 <= io_pixelVal_in_0_6;
      end else if (8'hd3 == _T_31[7:0]) begin
        image_0_211 <= io_pixelVal_in_0_5;
      end else if (8'hd3 == _T_28[7:0]) begin
        image_0_211 <= io_pixelVal_in_0_4;
      end else if (8'hd3 == _T_25[7:0]) begin
        image_0_211 <= io_pixelVal_in_0_3;
      end else if (8'hd3 == _T_22[7:0]) begin
        image_0_211 <= io_pixelVal_in_0_2;
      end else if (8'hd3 == _T_19[7:0]) begin
        image_0_211 <= io_pixelVal_in_0_1;
      end else if (8'hd3 == _T_15[7:0]) begin
        image_0_211 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_212 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hd4 == _T_34[7:0]) begin
        image_0_212 <= io_pixelVal_in_0_6;
      end else if (8'hd4 == _T_31[7:0]) begin
        image_0_212 <= io_pixelVal_in_0_5;
      end else if (8'hd4 == _T_28[7:0]) begin
        image_0_212 <= io_pixelVal_in_0_4;
      end else if (8'hd4 == _T_25[7:0]) begin
        image_0_212 <= io_pixelVal_in_0_3;
      end else if (8'hd4 == _T_22[7:0]) begin
        image_0_212 <= io_pixelVal_in_0_2;
      end else if (8'hd4 == _T_19[7:0]) begin
        image_0_212 <= io_pixelVal_in_0_1;
      end else if (8'hd4 == _T_15[7:0]) begin
        image_0_212 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_213 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hd5 == _T_34[7:0]) begin
        image_0_213 <= io_pixelVal_in_0_6;
      end else if (8'hd5 == _T_31[7:0]) begin
        image_0_213 <= io_pixelVal_in_0_5;
      end else if (8'hd5 == _T_28[7:0]) begin
        image_0_213 <= io_pixelVal_in_0_4;
      end else if (8'hd5 == _T_25[7:0]) begin
        image_0_213 <= io_pixelVal_in_0_3;
      end else if (8'hd5 == _T_22[7:0]) begin
        image_0_213 <= io_pixelVal_in_0_2;
      end else if (8'hd5 == _T_19[7:0]) begin
        image_0_213 <= io_pixelVal_in_0_1;
      end else if (8'hd5 == _T_15[7:0]) begin
        image_0_213 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_214 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hd6 == _T_34[7:0]) begin
        image_0_214 <= io_pixelVal_in_0_6;
      end else if (8'hd6 == _T_31[7:0]) begin
        image_0_214 <= io_pixelVal_in_0_5;
      end else if (8'hd6 == _T_28[7:0]) begin
        image_0_214 <= io_pixelVal_in_0_4;
      end else if (8'hd6 == _T_25[7:0]) begin
        image_0_214 <= io_pixelVal_in_0_3;
      end else if (8'hd6 == _T_22[7:0]) begin
        image_0_214 <= io_pixelVal_in_0_2;
      end else if (8'hd6 == _T_19[7:0]) begin
        image_0_214 <= io_pixelVal_in_0_1;
      end else if (8'hd6 == _T_15[7:0]) begin
        image_0_214 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_215 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hd7 == _T_34[7:0]) begin
        image_0_215 <= io_pixelVal_in_0_6;
      end else if (8'hd7 == _T_31[7:0]) begin
        image_0_215 <= io_pixelVal_in_0_5;
      end else if (8'hd7 == _T_28[7:0]) begin
        image_0_215 <= io_pixelVal_in_0_4;
      end else if (8'hd7 == _T_25[7:0]) begin
        image_0_215 <= io_pixelVal_in_0_3;
      end else if (8'hd7 == _T_22[7:0]) begin
        image_0_215 <= io_pixelVal_in_0_2;
      end else if (8'hd7 == _T_19[7:0]) begin
        image_0_215 <= io_pixelVal_in_0_1;
      end else if (8'hd7 == _T_15[7:0]) begin
        image_0_215 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_216 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hd8 == _T_34[7:0]) begin
        image_0_216 <= io_pixelVal_in_0_6;
      end else if (8'hd8 == _T_31[7:0]) begin
        image_0_216 <= io_pixelVal_in_0_5;
      end else if (8'hd8 == _T_28[7:0]) begin
        image_0_216 <= io_pixelVal_in_0_4;
      end else if (8'hd8 == _T_25[7:0]) begin
        image_0_216 <= io_pixelVal_in_0_3;
      end else if (8'hd8 == _T_22[7:0]) begin
        image_0_216 <= io_pixelVal_in_0_2;
      end else if (8'hd8 == _T_19[7:0]) begin
        image_0_216 <= io_pixelVal_in_0_1;
      end else if (8'hd8 == _T_15[7:0]) begin
        image_0_216 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_217 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hd9 == _T_34[7:0]) begin
        image_0_217 <= io_pixelVal_in_0_6;
      end else if (8'hd9 == _T_31[7:0]) begin
        image_0_217 <= io_pixelVal_in_0_5;
      end else if (8'hd9 == _T_28[7:0]) begin
        image_0_217 <= io_pixelVal_in_0_4;
      end else if (8'hd9 == _T_25[7:0]) begin
        image_0_217 <= io_pixelVal_in_0_3;
      end else if (8'hd9 == _T_22[7:0]) begin
        image_0_217 <= io_pixelVal_in_0_2;
      end else if (8'hd9 == _T_19[7:0]) begin
        image_0_217 <= io_pixelVal_in_0_1;
      end else if (8'hd9 == _T_15[7:0]) begin
        image_0_217 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_218 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hda == _T_34[7:0]) begin
        image_0_218 <= io_pixelVal_in_0_6;
      end else if (8'hda == _T_31[7:0]) begin
        image_0_218 <= io_pixelVal_in_0_5;
      end else if (8'hda == _T_28[7:0]) begin
        image_0_218 <= io_pixelVal_in_0_4;
      end else if (8'hda == _T_25[7:0]) begin
        image_0_218 <= io_pixelVal_in_0_3;
      end else if (8'hda == _T_22[7:0]) begin
        image_0_218 <= io_pixelVal_in_0_2;
      end else if (8'hda == _T_19[7:0]) begin
        image_0_218 <= io_pixelVal_in_0_1;
      end else if (8'hda == _T_15[7:0]) begin
        image_0_218 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_219 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hdb == _T_34[7:0]) begin
        image_0_219 <= io_pixelVal_in_0_6;
      end else if (8'hdb == _T_31[7:0]) begin
        image_0_219 <= io_pixelVal_in_0_5;
      end else if (8'hdb == _T_28[7:0]) begin
        image_0_219 <= io_pixelVal_in_0_4;
      end else if (8'hdb == _T_25[7:0]) begin
        image_0_219 <= io_pixelVal_in_0_3;
      end else if (8'hdb == _T_22[7:0]) begin
        image_0_219 <= io_pixelVal_in_0_2;
      end else if (8'hdb == _T_19[7:0]) begin
        image_0_219 <= io_pixelVal_in_0_1;
      end else if (8'hdb == _T_15[7:0]) begin
        image_0_219 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_220 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hdc == _T_34[7:0]) begin
        image_0_220 <= io_pixelVal_in_0_6;
      end else if (8'hdc == _T_31[7:0]) begin
        image_0_220 <= io_pixelVal_in_0_5;
      end else if (8'hdc == _T_28[7:0]) begin
        image_0_220 <= io_pixelVal_in_0_4;
      end else if (8'hdc == _T_25[7:0]) begin
        image_0_220 <= io_pixelVal_in_0_3;
      end else if (8'hdc == _T_22[7:0]) begin
        image_0_220 <= io_pixelVal_in_0_2;
      end else if (8'hdc == _T_19[7:0]) begin
        image_0_220 <= io_pixelVal_in_0_1;
      end else if (8'hdc == _T_15[7:0]) begin
        image_0_220 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_221 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hdd == _T_34[7:0]) begin
        image_0_221 <= io_pixelVal_in_0_6;
      end else if (8'hdd == _T_31[7:0]) begin
        image_0_221 <= io_pixelVal_in_0_5;
      end else if (8'hdd == _T_28[7:0]) begin
        image_0_221 <= io_pixelVal_in_0_4;
      end else if (8'hdd == _T_25[7:0]) begin
        image_0_221 <= io_pixelVal_in_0_3;
      end else if (8'hdd == _T_22[7:0]) begin
        image_0_221 <= io_pixelVal_in_0_2;
      end else if (8'hdd == _T_19[7:0]) begin
        image_0_221 <= io_pixelVal_in_0_1;
      end else if (8'hdd == _T_15[7:0]) begin
        image_0_221 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_222 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hde == _T_34[7:0]) begin
        image_0_222 <= io_pixelVal_in_0_6;
      end else if (8'hde == _T_31[7:0]) begin
        image_0_222 <= io_pixelVal_in_0_5;
      end else if (8'hde == _T_28[7:0]) begin
        image_0_222 <= io_pixelVal_in_0_4;
      end else if (8'hde == _T_25[7:0]) begin
        image_0_222 <= io_pixelVal_in_0_3;
      end else if (8'hde == _T_22[7:0]) begin
        image_0_222 <= io_pixelVal_in_0_2;
      end else if (8'hde == _T_19[7:0]) begin
        image_0_222 <= io_pixelVal_in_0_1;
      end else if (8'hde == _T_15[7:0]) begin
        image_0_222 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_223 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hdf == _T_34[7:0]) begin
        image_0_223 <= io_pixelVal_in_0_6;
      end else if (8'hdf == _T_31[7:0]) begin
        image_0_223 <= io_pixelVal_in_0_5;
      end else if (8'hdf == _T_28[7:0]) begin
        image_0_223 <= io_pixelVal_in_0_4;
      end else if (8'hdf == _T_25[7:0]) begin
        image_0_223 <= io_pixelVal_in_0_3;
      end else if (8'hdf == _T_22[7:0]) begin
        image_0_223 <= io_pixelVal_in_0_2;
      end else if (8'hdf == _T_19[7:0]) begin
        image_0_223 <= io_pixelVal_in_0_1;
      end else if (8'hdf == _T_15[7:0]) begin
        image_0_223 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_224 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'he0 == _T_34[7:0]) begin
        image_0_224 <= io_pixelVal_in_0_6;
      end else if (8'he0 == _T_31[7:0]) begin
        image_0_224 <= io_pixelVal_in_0_5;
      end else if (8'he0 == _T_28[7:0]) begin
        image_0_224 <= io_pixelVal_in_0_4;
      end else if (8'he0 == _T_25[7:0]) begin
        image_0_224 <= io_pixelVal_in_0_3;
      end else if (8'he0 == _T_22[7:0]) begin
        image_0_224 <= io_pixelVal_in_0_2;
      end else if (8'he0 == _T_19[7:0]) begin
        image_0_224 <= io_pixelVal_in_0_1;
      end else if (8'he0 == _T_15[7:0]) begin
        image_0_224 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_225 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'he1 == _T_34[7:0]) begin
        image_0_225 <= io_pixelVal_in_0_6;
      end else if (8'he1 == _T_31[7:0]) begin
        image_0_225 <= io_pixelVal_in_0_5;
      end else if (8'he1 == _T_28[7:0]) begin
        image_0_225 <= io_pixelVal_in_0_4;
      end else if (8'he1 == _T_25[7:0]) begin
        image_0_225 <= io_pixelVal_in_0_3;
      end else if (8'he1 == _T_22[7:0]) begin
        image_0_225 <= io_pixelVal_in_0_2;
      end else if (8'he1 == _T_19[7:0]) begin
        image_0_225 <= io_pixelVal_in_0_1;
      end else if (8'he1 == _T_15[7:0]) begin
        image_0_225 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_226 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'he2 == _T_34[7:0]) begin
        image_0_226 <= io_pixelVal_in_0_6;
      end else if (8'he2 == _T_31[7:0]) begin
        image_0_226 <= io_pixelVal_in_0_5;
      end else if (8'he2 == _T_28[7:0]) begin
        image_0_226 <= io_pixelVal_in_0_4;
      end else if (8'he2 == _T_25[7:0]) begin
        image_0_226 <= io_pixelVal_in_0_3;
      end else if (8'he2 == _T_22[7:0]) begin
        image_0_226 <= io_pixelVal_in_0_2;
      end else if (8'he2 == _T_19[7:0]) begin
        image_0_226 <= io_pixelVal_in_0_1;
      end else if (8'he2 == _T_15[7:0]) begin
        image_0_226 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_227 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'he3 == _T_34[7:0]) begin
        image_0_227 <= io_pixelVal_in_0_6;
      end else if (8'he3 == _T_31[7:0]) begin
        image_0_227 <= io_pixelVal_in_0_5;
      end else if (8'he3 == _T_28[7:0]) begin
        image_0_227 <= io_pixelVal_in_0_4;
      end else if (8'he3 == _T_25[7:0]) begin
        image_0_227 <= io_pixelVal_in_0_3;
      end else if (8'he3 == _T_22[7:0]) begin
        image_0_227 <= io_pixelVal_in_0_2;
      end else if (8'he3 == _T_19[7:0]) begin
        image_0_227 <= io_pixelVal_in_0_1;
      end else if (8'he3 == _T_15[7:0]) begin
        image_0_227 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_228 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'he4 == _T_34[7:0]) begin
        image_0_228 <= io_pixelVal_in_0_6;
      end else if (8'he4 == _T_31[7:0]) begin
        image_0_228 <= io_pixelVal_in_0_5;
      end else if (8'he4 == _T_28[7:0]) begin
        image_0_228 <= io_pixelVal_in_0_4;
      end else if (8'he4 == _T_25[7:0]) begin
        image_0_228 <= io_pixelVal_in_0_3;
      end else if (8'he4 == _T_22[7:0]) begin
        image_0_228 <= io_pixelVal_in_0_2;
      end else if (8'he4 == _T_19[7:0]) begin
        image_0_228 <= io_pixelVal_in_0_1;
      end else if (8'he4 == _T_15[7:0]) begin
        image_0_228 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_229 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'he5 == _T_34[7:0]) begin
        image_0_229 <= io_pixelVal_in_0_6;
      end else if (8'he5 == _T_31[7:0]) begin
        image_0_229 <= io_pixelVal_in_0_5;
      end else if (8'he5 == _T_28[7:0]) begin
        image_0_229 <= io_pixelVal_in_0_4;
      end else if (8'he5 == _T_25[7:0]) begin
        image_0_229 <= io_pixelVal_in_0_3;
      end else if (8'he5 == _T_22[7:0]) begin
        image_0_229 <= io_pixelVal_in_0_2;
      end else if (8'he5 == _T_19[7:0]) begin
        image_0_229 <= io_pixelVal_in_0_1;
      end else if (8'he5 == _T_15[7:0]) begin
        image_0_229 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_230 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'he6 == _T_34[7:0]) begin
        image_0_230 <= io_pixelVal_in_0_6;
      end else if (8'he6 == _T_31[7:0]) begin
        image_0_230 <= io_pixelVal_in_0_5;
      end else if (8'he6 == _T_28[7:0]) begin
        image_0_230 <= io_pixelVal_in_0_4;
      end else if (8'he6 == _T_25[7:0]) begin
        image_0_230 <= io_pixelVal_in_0_3;
      end else if (8'he6 == _T_22[7:0]) begin
        image_0_230 <= io_pixelVal_in_0_2;
      end else if (8'he6 == _T_19[7:0]) begin
        image_0_230 <= io_pixelVal_in_0_1;
      end else if (8'he6 == _T_15[7:0]) begin
        image_0_230 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_231 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'he7 == _T_34[7:0]) begin
        image_0_231 <= io_pixelVal_in_0_6;
      end else if (8'he7 == _T_31[7:0]) begin
        image_0_231 <= io_pixelVal_in_0_5;
      end else if (8'he7 == _T_28[7:0]) begin
        image_0_231 <= io_pixelVal_in_0_4;
      end else if (8'he7 == _T_25[7:0]) begin
        image_0_231 <= io_pixelVal_in_0_3;
      end else if (8'he7 == _T_22[7:0]) begin
        image_0_231 <= io_pixelVal_in_0_2;
      end else if (8'he7 == _T_19[7:0]) begin
        image_0_231 <= io_pixelVal_in_0_1;
      end else if (8'he7 == _T_15[7:0]) begin
        image_0_231 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_232 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'he8 == _T_34[7:0]) begin
        image_0_232 <= io_pixelVal_in_0_6;
      end else if (8'he8 == _T_31[7:0]) begin
        image_0_232 <= io_pixelVal_in_0_5;
      end else if (8'he8 == _T_28[7:0]) begin
        image_0_232 <= io_pixelVal_in_0_4;
      end else if (8'he8 == _T_25[7:0]) begin
        image_0_232 <= io_pixelVal_in_0_3;
      end else if (8'he8 == _T_22[7:0]) begin
        image_0_232 <= io_pixelVal_in_0_2;
      end else if (8'he8 == _T_19[7:0]) begin
        image_0_232 <= io_pixelVal_in_0_1;
      end else if (8'he8 == _T_15[7:0]) begin
        image_0_232 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_233 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'he9 == _T_34[7:0]) begin
        image_0_233 <= io_pixelVal_in_0_6;
      end else if (8'he9 == _T_31[7:0]) begin
        image_0_233 <= io_pixelVal_in_0_5;
      end else if (8'he9 == _T_28[7:0]) begin
        image_0_233 <= io_pixelVal_in_0_4;
      end else if (8'he9 == _T_25[7:0]) begin
        image_0_233 <= io_pixelVal_in_0_3;
      end else if (8'he9 == _T_22[7:0]) begin
        image_0_233 <= io_pixelVal_in_0_2;
      end else if (8'he9 == _T_19[7:0]) begin
        image_0_233 <= io_pixelVal_in_0_1;
      end else if (8'he9 == _T_15[7:0]) begin
        image_0_233 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_234 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hea == _T_34[7:0]) begin
        image_0_234 <= io_pixelVal_in_0_6;
      end else if (8'hea == _T_31[7:0]) begin
        image_0_234 <= io_pixelVal_in_0_5;
      end else if (8'hea == _T_28[7:0]) begin
        image_0_234 <= io_pixelVal_in_0_4;
      end else if (8'hea == _T_25[7:0]) begin
        image_0_234 <= io_pixelVal_in_0_3;
      end else if (8'hea == _T_22[7:0]) begin
        image_0_234 <= io_pixelVal_in_0_2;
      end else if (8'hea == _T_19[7:0]) begin
        image_0_234 <= io_pixelVal_in_0_1;
      end else if (8'hea == _T_15[7:0]) begin
        image_0_234 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_235 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'heb == _T_34[7:0]) begin
        image_0_235 <= io_pixelVal_in_0_6;
      end else if (8'heb == _T_31[7:0]) begin
        image_0_235 <= io_pixelVal_in_0_5;
      end else if (8'heb == _T_28[7:0]) begin
        image_0_235 <= io_pixelVal_in_0_4;
      end else if (8'heb == _T_25[7:0]) begin
        image_0_235 <= io_pixelVal_in_0_3;
      end else if (8'heb == _T_22[7:0]) begin
        image_0_235 <= io_pixelVal_in_0_2;
      end else if (8'heb == _T_19[7:0]) begin
        image_0_235 <= io_pixelVal_in_0_1;
      end else if (8'heb == _T_15[7:0]) begin
        image_0_235 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_236 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hec == _T_34[7:0]) begin
        image_0_236 <= io_pixelVal_in_0_6;
      end else if (8'hec == _T_31[7:0]) begin
        image_0_236 <= io_pixelVal_in_0_5;
      end else if (8'hec == _T_28[7:0]) begin
        image_0_236 <= io_pixelVal_in_0_4;
      end else if (8'hec == _T_25[7:0]) begin
        image_0_236 <= io_pixelVal_in_0_3;
      end else if (8'hec == _T_22[7:0]) begin
        image_0_236 <= io_pixelVal_in_0_2;
      end else if (8'hec == _T_19[7:0]) begin
        image_0_236 <= io_pixelVal_in_0_1;
      end else if (8'hec == _T_15[7:0]) begin
        image_0_236 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_237 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hed == _T_34[7:0]) begin
        image_0_237 <= io_pixelVal_in_0_6;
      end else if (8'hed == _T_31[7:0]) begin
        image_0_237 <= io_pixelVal_in_0_5;
      end else if (8'hed == _T_28[7:0]) begin
        image_0_237 <= io_pixelVal_in_0_4;
      end else if (8'hed == _T_25[7:0]) begin
        image_0_237 <= io_pixelVal_in_0_3;
      end else if (8'hed == _T_22[7:0]) begin
        image_0_237 <= io_pixelVal_in_0_2;
      end else if (8'hed == _T_19[7:0]) begin
        image_0_237 <= io_pixelVal_in_0_1;
      end else if (8'hed == _T_15[7:0]) begin
        image_0_237 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_238 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hee == _T_34[7:0]) begin
        image_0_238 <= io_pixelVal_in_0_6;
      end else if (8'hee == _T_31[7:0]) begin
        image_0_238 <= io_pixelVal_in_0_5;
      end else if (8'hee == _T_28[7:0]) begin
        image_0_238 <= io_pixelVal_in_0_4;
      end else if (8'hee == _T_25[7:0]) begin
        image_0_238 <= io_pixelVal_in_0_3;
      end else if (8'hee == _T_22[7:0]) begin
        image_0_238 <= io_pixelVal_in_0_2;
      end else if (8'hee == _T_19[7:0]) begin
        image_0_238 <= io_pixelVal_in_0_1;
      end else if (8'hee == _T_15[7:0]) begin
        image_0_238 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_239 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hef == _T_34[7:0]) begin
        image_0_239 <= io_pixelVal_in_0_6;
      end else if (8'hef == _T_31[7:0]) begin
        image_0_239 <= io_pixelVal_in_0_5;
      end else if (8'hef == _T_28[7:0]) begin
        image_0_239 <= io_pixelVal_in_0_4;
      end else if (8'hef == _T_25[7:0]) begin
        image_0_239 <= io_pixelVal_in_0_3;
      end else if (8'hef == _T_22[7:0]) begin
        image_0_239 <= io_pixelVal_in_0_2;
      end else if (8'hef == _T_19[7:0]) begin
        image_0_239 <= io_pixelVal_in_0_1;
      end else if (8'hef == _T_15[7:0]) begin
        image_0_239 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_240 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hf0 == _T_34[7:0]) begin
        image_0_240 <= io_pixelVal_in_0_6;
      end else if (8'hf0 == _T_31[7:0]) begin
        image_0_240 <= io_pixelVal_in_0_5;
      end else if (8'hf0 == _T_28[7:0]) begin
        image_0_240 <= io_pixelVal_in_0_4;
      end else if (8'hf0 == _T_25[7:0]) begin
        image_0_240 <= io_pixelVal_in_0_3;
      end else if (8'hf0 == _T_22[7:0]) begin
        image_0_240 <= io_pixelVal_in_0_2;
      end else if (8'hf0 == _T_19[7:0]) begin
        image_0_240 <= io_pixelVal_in_0_1;
      end else if (8'hf0 == _T_15[7:0]) begin
        image_0_240 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_241 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hf1 == _T_34[7:0]) begin
        image_0_241 <= io_pixelVal_in_0_6;
      end else if (8'hf1 == _T_31[7:0]) begin
        image_0_241 <= io_pixelVal_in_0_5;
      end else if (8'hf1 == _T_28[7:0]) begin
        image_0_241 <= io_pixelVal_in_0_4;
      end else if (8'hf1 == _T_25[7:0]) begin
        image_0_241 <= io_pixelVal_in_0_3;
      end else if (8'hf1 == _T_22[7:0]) begin
        image_0_241 <= io_pixelVal_in_0_2;
      end else if (8'hf1 == _T_19[7:0]) begin
        image_0_241 <= io_pixelVal_in_0_1;
      end else if (8'hf1 == _T_15[7:0]) begin
        image_0_241 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_242 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hf2 == _T_34[7:0]) begin
        image_0_242 <= io_pixelVal_in_0_6;
      end else if (8'hf2 == _T_31[7:0]) begin
        image_0_242 <= io_pixelVal_in_0_5;
      end else if (8'hf2 == _T_28[7:0]) begin
        image_0_242 <= io_pixelVal_in_0_4;
      end else if (8'hf2 == _T_25[7:0]) begin
        image_0_242 <= io_pixelVal_in_0_3;
      end else if (8'hf2 == _T_22[7:0]) begin
        image_0_242 <= io_pixelVal_in_0_2;
      end else if (8'hf2 == _T_19[7:0]) begin
        image_0_242 <= io_pixelVal_in_0_1;
      end else if (8'hf2 == _T_15[7:0]) begin
        image_0_242 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_243 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hf3 == _T_34[7:0]) begin
        image_0_243 <= io_pixelVal_in_0_6;
      end else if (8'hf3 == _T_31[7:0]) begin
        image_0_243 <= io_pixelVal_in_0_5;
      end else if (8'hf3 == _T_28[7:0]) begin
        image_0_243 <= io_pixelVal_in_0_4;
      end else if (8'hf3 == _T_25[7:0]) begin
        image_0_243 <= io_pixelVal_in_0_3;
      end else if (8'hf3 == _T_22[7:0]) begin
        image_0_243 <= io_pixelVal_in_0_2;
      end else if (8'hf3 == _T_19[7:0]) begin
        image_0_243 <= io_pixelVal_in_0_1;
      end else if (8'hf3 == _T_15[7:0]) begin
        image_0_243 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_244 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hf4 == _T_34[7:0]) begin
        image_0_244 <= io_pixelVal_in_0_6;
      end else if (8'hf4 == _T_31[7:0]) begin
        image_0_244 <= io_pixelVal_in_0_5;
      end else if (8'hf4 == _T_28[7:0]) begin
        image_0_244 <= io_pixelVal_in_0_4;
      end else if (8'hf4 == _T_25[7:0]) begin
        image_0_244 <= io_pixelVal_in_0_3;
      end else if (8'hf4 == _T_22[7:0]) begin
        image_0_244 <= io_pixelVal_in_0_2;
      end else if (8'hf4 == _T_19[7:0]) begin
        image_0_244 <= io_pixelVal_in_0_1;
      end else if (8'hf4 == _T_15[7:0]) begin
        image_0_244 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_245 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hf5 == _T_34[7:0]) begin
        image_0_245 <= io_pixelVal_in_0_6;
      end else if (8'hf5 == _T_31[7:0]) begin
        image_0_245 <= io_pixelVal_in_0_5;
      end else if (8'hf5 == _T_28[7:0]) begin
        image_0_245 <= io_pixelVal_in_0_4;
      end else if (8'hf5 == _T_25[7:0]) begin
        image_0_245 <= io_pixelVal_in_0_3;
      end else if (8'hf5 == _T_22[7:0]) begin
        image_0_245 <= io_pixelVal_in_0_2;
      end else if (8'hf5 == _T_19[7:0]) begin
        image_0_245 <= io_pixelVal_in_0_1;
      end else if (8'hf5 == _T_15[7:0]) begin
        image_0_245 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_246 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hf6 == _T_34[7:0]) begin
        image_0_246 <= io_pixelVal_in_0_6;
      end else if (8'hf6 == _T_31[7:0]) begin
        image_0_246 <= io_pixelVal_in_0_5;
      end else if (8'hf6 == _T_28[7:0]) begin
        image_0_246 <= io_pixelVal_in_0_4;
      end else if (8'hf6 == _T_25[7:0]) begin
        image_0_246 <= io_pixelVal_in_0_3;
      end else if (8'hf6 == _T_22[7:0]) begin
        image_0_246 <= io_pixelVal_in_0_2;
      end else if (8'hf6 == _T_19[7:0]) begin
        image_0_246 <= io_pixelVal_in_0_1;
      end else if (8'hf6 == _T_15[7:0]) begin
        image_0_246 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_247 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hf7 == _T_34[7:0]) begin
        image_0_247 <= io_pixelVal_in_0_6;
      end else if (8'hf7 == _T_31[7:0]) begin
        image_0_247 <= io_pixelVal_in_0_5;
      end else if (8'hf7 == _T_28[7:0]) begin
        image_0_247 <= io_pixelVal_in_0_4;
      end else if (8'hf7 == _T_25[7:0]) begin
        image_0_247 <= io_pixelVal_in_0_3;
      end else if (8'hf7 == _T_22[7:0]) begin
        image_0_247 <= io_pixelVal_in_0_2;
      end else if (8'hf7 == _T_19[7:0]) begin
        image_0_247 <= io_pixelVal_in_0_1;
      end else if (8'hf7 == _T_15[7:0]) begin
        image_0_247 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_248 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hf8 == _T_34[7:0]) begin
        image_0_248 <= io_pixelVal_in_0_6;
      end else if (8'hf8 == _T_31[7:0]) begin
        image_0_248 <= io_pixelVal_in_0_5;
      end else if (8'hf8 == _T_28[7:0]) begin
        image_0_248 <= io_pixelVal_in_0_4;
      end else if (8'hf8 == _T_25[7:0]) begin
        image_0_248 <= io_pixelVal_in_0_3;
      end else if (8'hf8 == _T_22[7:0]) begin
        image_0_248 <= io_pixelVal_in_0_2;
      end else if (8'hf8 == _T_19[7:0]) begin
        image_0_248 <= io_pixelVal_in_0_1;
      end else if (8'hf8 == _T_15[7:0]) begin
        image_0_248 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_249 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hf9 == _T_34[7:0]) begin
        image_0_249 <= io_pixelVal_in_0_6;
      end else if (8'hf9 == _T_31[7:0]) begin
        image_0_249 <= io_pixelVal_in_0_5;
      end else if (8'hf9 == _T_28[7:0]) begin
        image_0_249 <= io_pixelVal_in_0_4;
      end else if (8'hf9 == _T_25[7:0]) begin
        image_0_249 <= io_pixelVal_in_0_3;
      end else if (8'hf9 == _T_22[7:0]) begin
        image_0_249 <= io_pixelVal_in_0_2;
      end else if (8'hf9 == _T_19[7:0]) begin
        image_0_249 <= io_pixelVal_in_0_1;
      end else if (8'hf9 == _T_15[7:0]) begin
        image_0_249 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_250 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hfa == _T_34[7:0]) begin
        image_0_250 <= io_pixelVal_in_0_6;
      end else if (8'hfa == _T_31[7:0]) begin
        image_0_250 <= io_pixelVal_in_0_5;
      end else if (8'hfa == _T_28[7:0]) begin
        image_0_250 <= io_pixelVal_in_0_4;
      end else if (8'hfa == _T_25[7:0]) begin
        image_0_250 <= io_pixelVal_in_0_3;
      end else if (8'hfa == _T_22[7:0]) begin
        image_0_250 <= io_pixelVal_in_0_2;
      end else if (8'hfa == _T_19[7:0]) begin
        image_0_250 <= io_pixelVal_in_0_1;
      end else if (8'hfa == _T_15[7:0]) begin
        image_0_250 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_251 <= 4'hf;
    end else if (io_valid_in) begin
      if (8'hfb == _T_34[7:0]) begin
        image_0_251 <= io_pixelVal_in_0_6;
      end else if (8'hfb == _T_31[7:0]) begin
        image_0_251 <= io_pixelVal_in_0_5;
      end else if (8'hfb == _T_28[7:0]) begin
        image_0_251 <= io_pixelVal_in_0_4;
      end else if (8'hfb == _T_25[7:0]) begin
        image_0_251 <= io_pixelVal_in_0_3;
      end else if (8'hfb == _T_22[7:0]) begin
        image_0_251 <= io_pixelVal_in_0_2;
      end else if (8'hfb == _T_19[7:0]) begin
        image_0_251 <= io_pixelVal_in_0_1;
      end else if (8'hfb == _T_15[7:0]) begin
        image_0_251 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_1_0 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h0 == _T_34[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_6;
      end else if (8'h0 == _T_31[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_5;
      end else if (8'h0 == _T_28[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_4;
      end else if (8'h0 == _T_25[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_3;
      end else if (8'h0 == _T_22[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_2;
      end else if (8'h0 == _T_19[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_1;
      end else if (8'h0 == _T_15[7:0]) begin
        image_1_0 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_1 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1 == _T_34[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_6;
      end else if (8'h1 == _T_31[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_5;
      end else if (8'h1 == _T_28[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_4;
      end else if (8'h1 == _T_25[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_3;
      end else if (8'h1 == _T_22[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_2;
      end else if (8'h1 == _T_19[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_1;
      end else if (8'h1 == _T_15[7:0]) begin
        image_1_1 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_2 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2 == _T_34[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_6;
      end else if (8'h2 == _T_31[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_5;
      end else if (8'h2 == _T_28[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_4;
      end else if (8'h2 == _T_25[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_3;
      end else if (8'h2 == _T_22[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_2;
      end else if (8'h2 == _T_19[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_1;
      end else if (8'h2 == _T_15[7:0]) begin
        image_1_2 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_3 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3 == _T_34[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_6;
      end else if (8'h3 == _T_31[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_5;
      end else if (8'h3 == _T_28[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_4;
      end else if (8'h3 == _T_25[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_3;
      end else if (8'h3 == _T_22[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_2;
      end else if (8'h3 == _T_19[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_1;
      end else if (8'h3 == _T_15[7:0]) begin
        image_1_3 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_4 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4 == _T_34[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_6;
      end else if (8'h4 == _T_31[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_5;
      end else if (8'h4 == _T_28[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_4;
      end else if (8'h4 == _T_25[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_3;
      end else if (8'h4 == _T_22[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_2;
      end else if (8'h4 == _T_19[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_1;
      end else if (8'h4 == _T_15[7:0]) begin
        image_1_4 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_5 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5 == _T_34[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_6;
      end else if (8'h5 == _T_31[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_5;
      end else if (8'h5 == _T_28[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_4;
      end else if (8'h5 == _T_25[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_3;
      end else if (8'h5 == _T_22[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_2;
      end else if (8'h5 == _T_19[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_1;
      end else if (8'h5 == _T_15[7:0]) begin
        image_1_5 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_6 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6 == _T_34[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_6;
      end else if (8'h6 == _T_31[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_5;
      end else if (8'h6 == _T_28[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_4;
      end else if (8'h6 == _T_25[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_3;
      end else if (8'h6 == _T_22[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_2;
      end else if (8'h6 == _T_19[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_1;
      end else if (8'h6 == _T_15[7:0]) begin
        image_1_6 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_7 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7 == _T_34[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_6;
      end else if (8'h7 == _T_31[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_5;
      end else if (8'h7 == _T_28[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_4;
      end else if (8'h7 == _T_25[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_3;
      end else if (8'h7 == _T_22[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_2;
      end else if (8'h7 == _T_19[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_1;
      end else if (8'h7 == _T_15[7:0]) begin
        image_1_7 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_8 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8 == _T_34[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_6;
      end else if (8'h8 == _T_31[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_5;
      end else if (8'h8 == _T_28[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_4;
      end else if (8'h8 == _T_25[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_3;
      end else if (8'h8 == _T_22[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_2;
      end else if (8'h8 == _T_19[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_1;
      end else if (8'h8 == _T_15[7:0]) begin
        image_1_8 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_9 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9 == _T_34[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_6;
      end else if (8'h9 == _T_31[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_5;
      end else if (8'h9 == _T_28[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_4;
      end else if (8'h9 == _T_25[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_3;
      end else if (8'h9 == _T_22[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_2;
      end else if (8'h9 == _T_19[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_1;
      end else if (8'h9 == _T_15[7:0]) begin
        image_1_9 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_10 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha == _T_34[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_6;
      end else if (8'ha == _T_31[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_5;
      end else if (8'ha == _T_28[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_4;
      end else if (8'ha == _T_25[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_3;
      end else if (8'ha == _T_22[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_2;
      end else if (8'ha == _T_19[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_1;
      end else if (8'ha == _T_15[7:0]) begin
        image_1_10 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_11 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb == _T_34[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_6;
      end else if (8'hb == _T_31[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_5;
      end else if (8'hb == _T_28[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_4;
      end else if (8'hb == _T_25[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_3;
      end else if (8'hb == _T_22[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_2;
      end else if (8'hb == _T_19[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_1;
      end else if (8'hb == _T_15[7:0]) begin
        image_1_11 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_12 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc == _T_34[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_6;
      end else if (8'hc == _T_31[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_5;
      end else if (8'hc == _T_28[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_4;
      end else if (8'hc == _T_25[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_3;
      end else if (8'hc == _T_22[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_2;
      end else if (8'hc == _T_19[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_1;
      end else if (8'hc == _T_15[7:0]) begin
        image_1_12 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_13 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd == _T_34[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_6;
      end else if (8'hd == _T_31[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_5;
      end else if (8'hd == _T_28[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_4;
      end else if (8'hd == _T_25[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_3;
      end else if (8'hd == _T_22[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_2;
      end else if (8'hd == _T_19[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_1;
      end else if (8'hd == _T_15[7:0]) begin
        image_1_13 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_14 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he == _T_34[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_6;
      end else if (8'he == _T_31[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_5;
      end else if (8'he == _T_28[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_4;
      end else if (8'he == _T_25[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_3;
      end else if (8'he == _T_22[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_2;
      end else if (8'he == _T_19[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_1;
      end else if (8'he == _T_15[7:0]) begin
        image_1_14 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_15 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf == _T_34[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_6;
      end else if (8'hf == _T_31[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_5;
      end else if (8'hf == _T_28[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_4;
      end else if (8'hf == _T_25[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_3;
      end else if (8'hf == _T_22[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_2;
      end else if (8'hf == _T_19[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_1;
      end else if (8'hf == _T_15[7:0]) begin
        image_1_15 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_16 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h10 == _T_34[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_6;
      end else if (8'h10 == _T_31[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_5;
      end else if (8'h10 == _T_28[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_4;
      end else if (8'h10 == _T_25[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_3;
      end else if (8'h10 == _T_22[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_2;
      end else if (8'h10 == _T_19[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_1;
      end else if (8'h10 == _T_15[7:0]) begin
        image_1_16 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_17 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h11 == _T_34[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_6;
      end else if (8'h11 == _T_31[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_5;
      end else if (8'h11 == _T_28[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_4;
      end else if (8'h11 == _T_25[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_3;
      end else if (8'h11 == _T_22[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_2;
      end else if (8'h11 == _T_19[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_1;
      end else if (8'h11 == _T_15[7:0]) begin
        image_1_17 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_18 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h12 == _T_34[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_6;
      end else if (8'h12 == _T_31[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_5;
      end else if (8'h12 == _T_28[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_4;
      end else if (8'h12 == _T_25[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_3;
      end else if (8'h12 == _T_22[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_2;
      end else if (8'h12 == _T_19[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_1;
      end else if (8'h12 == _T_15[7:0]) begin
        image_1_18 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_19 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h13 == _T_34[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_6;
      end else if (8'h13 == _T_31[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_5;
      end else if (8'h13 == _T_28[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_4;
      end else if (8'h13 == _T_25[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_3;
      end else if (8'h13 == _T_22[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_2;
      end else if (8'h13 == _T_19[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_1;
      end else if (8'h13 == _T_15[7:0]) begin
        image_1_19 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_20 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h14 == _T_34[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_6;
      end else if (8'h14 == _T_31[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_5;
      end else if (8'h14 == _T_28[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_4;
      end else if (8'h14 == _T_25[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_3;
      end else if (8'h14 == _T_22[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_2;
      end else if (8'h14 == _T_19[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_1;
      end else if (8'h14 == _T_15[7:0]) begin
        image_1_20 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_21 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h15 == _T_34[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_6;
      end else if (8'h15 == _T_31[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_5;
      end else if (8'h15 == _T_28[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_4;
      end else if (8'h15 == _T_25[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_3;
      end else if (8'h15 == _T_22[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_2;
      end else if (8'h15 == _T_19[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_1;
      end else if (8'h15 == _T_15[7:0]) begin
        image_1_21 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_22 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h16 == _T_34[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_6;
      end else if (8'h16 == _T_31[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_5;
      end else if (8'h16 == _T_28[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_4;
      end else if (8'h16 == _T_25[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_3;
      end else if (8'h16 == _T_22[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_2;
      end else if (8'h16 == _T_19[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_1;
      end else if (8'h16 == _T_15[7:0]) begin
        image_1_22 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_23 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h17 == _T_34[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_6;
      end else if (8'h17 == _T_31[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_5;
      end else if (8'h17 == _T_28[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_4;
      end else if (8'h17 == _T_25[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_3;
      end else if (8'h17 == _T_22[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_2;
      end else if (8'h17 == _T_19[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_1;
      end else if (8'h17 == _T_15[7:0]) begin
        image_1_23 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_24 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h18 == _T_34[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_6;
      end else if (8'h18 == _T_31[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_5;
      end else if (8'h18 == _T_28[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_4;
      end else if (8'h18 == _T_25[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_3;
      end else if (8'h18 == _T_22[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_2;
      end else if (8'h18 == _T_19[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_1;
      end else if (8'h18 == _T_15[7:0]) begin
        image_1_24 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_25 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h19 == _T_34[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_6;
      end else if (8'h19 == _T_31[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_5;
      end else if (8'h19 == _T_28[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_4;
      end else if (8'h19 == _T_25[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_3;
      end else if (8'h19 == _T_22[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_2;
      end else if (8'h19 == _T_19[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_1;
      end else if (8'h19 == _T_15[7:0]) begin
        image_1_25 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_26 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1a == _T_34[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_6;
      end else if (8'h1a == _T_31[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_5;
      end else if (8'h1a == _T_28[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_4;
      end else if (8'h1a == _T_25[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_3;
      end else if (8'h1a == _T_22[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_2;
      end else if (8'h1a == _T_19[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_1;
      end else if (8'h1a == _T_15[7:0]) begin
        image_1_26 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_27 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1b == _T_34[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_6;
      end else if (8'h1b == _T_31[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_5;
      end else if (8'h1b == _T_28[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_4;
      end else if (8'h1b == _T_25[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_3;
      end else if (8'h1b == _T_22[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_2;
      end else if (8'h1b == _T_19[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_1;
      end else if (8'h1b == _T_15[7:0]) begin
        image_1_27 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_28 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1c == _T_34[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_6;
      end else if (8'h1c == _T_31[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_5;
      end else if (8'h1c == _T_28[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_4;
      end else if (8'h1c == _T_25[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_3;
      end else if (8'h1c == _T_22[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_2;
      end else if (8'h1c == _T_19[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_1;
      end else if (8'h1c == _T_15[7:0]) begin
        image_1_28 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_29 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1d == _T_34[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_6;
      end else if (8'h1d == _T_31[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_5;
      end else if (8'h1d == _T_28[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_4;
      end else if (8'h1d == _T_25[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_3;
      end else if (8'h1d == _T_22[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_2;
      end else if (8'h1d == _T_19[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_1;
      end else if (8'h1d == _T_15[7:0]) begin
        image_1_29 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_30 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1e == _T_34[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_6;
      end else if (8'h1e == _T_31[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_5;
      end else if (8'h1e == _T_28[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_4;
      end else if (8'h1e == _T_25[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_3;
      end else if (8'h1e == _T_22[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_2;
      end else if (8'h1e == _T_19[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_1;
      end else if (8'h1e == _T_15[7:0]) begin
        image_1_30 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_31 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1f == _T_34[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_6;
      end else if (8'h1f == _T_31[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_5;
      end else if (8'h1f == _T_28[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_4;
      end else if (8'h1f == _T_25[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_3;
      end else if (8'h1f == _T_22[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_2;
      end else if (8'h1f == _T_19[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_1;
      end else if (8'h1f == _T_15[7:0]) begin
        image_1_31 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_32 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h20 == _T_34[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_6;
      end else if (8'h20 == _T_31[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_5;
      end else if (8'h20 == _T_28[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_4;
      end else if (8'h20 == _T_25[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_3;
      end else if (8'h20 == _T_22[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_2;
      end else if (8'h20 == _T_19[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_1;
      end else if (8'h20 == _T_15[7:0]) begin
        image_1_32 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_33 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h21 == _T_34[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_6;
      end else if (8'h21 == _T_31[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_5;
      end else if (8'h21 == _T_28[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_4;
      end else if (8'h21 == _T_25[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_3;
      end else if (8'h21 == _T_22[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_2;
      end else if (8'h21 == _T_19[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_1;
      end else if (8'h21 == _T_15[7:0]) begin
        image_1_33 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_34 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h22 == _T_34[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_6;
      end else if (8'h22 == _T_31[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_5;
      end else if (8'h22 == _T_28[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_4;
      end else if (8'h22 == _T_25[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_3;
      end else if (8'h22 == _T_22[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_2;
      end else if (8'h22 == _T_19[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_1;
      end else if (8'h22 == _T_15[7:0]) begin
        image_1_34 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_35 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h23 == _T_34[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_6;
      end else if (8'h23 == _T_31[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_5;
      end else if (8'h23 == _T_28[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_4;
      end else if (8'h23 == _T_25[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_3;
      end else if (8'h23 == _T_22[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_2;
      end else if (8'h23 == _T_19[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_1;
      end else if (8'h23 == _T_15[7:0]) begin
        image_1_35 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_36 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h24 == _T_34[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_6;
      end else if (8'h24 == _T_31[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_5;
      end else if (8'h24 == _T_28[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_4;
      end else if (8'h24 == _T_25[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_3;
      end else if (8'h24 == _T_22[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_2;
      end else if (8'h24 == _T_19[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_1;
      end else if (8'h24 == _T_15[7:0]) begin
        image_1_36 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_37 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h25 == _T_34[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_6;
      end else if (8'h25 == _T_31[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_5;
      end else if (8'h25 == _T_28[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_4;
      end else if (8'h25 == _T_25[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_3;
      end else if (8'h25 == _T_22[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_2;
      end else if (8'h25 == _T_19[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_1;
      end else if (8'h25 == _T_15[7:0]) begin
        image_1_37 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_38 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h26 == _T_34[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_6;
      end else if (8'h26 == _T_31[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_5;
      end else if (8'h26 == _T_28[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_4;
      end else if (8'h26 == _T_25[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_3;
      end else if (8'h26 == _T_22[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_2;
      end else if (8'h26 == _T_19[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_1;
      end else if (8'h26 == _T_15[7:0]) begin
        image_1_38 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_39 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h27 == _T_34[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_6;
      end else if (8'h27 == _T_31[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_5;
      end else if (8'h27 == _T_28[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_4;
      end else if (8'h27 == _T_25[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_3;
      end else if (8'h27 == _T_22[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_2;
      end else if (8'h27 == _T_19[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_1;
      end else if (8'h27 == _T_15[7:0]) begin
        image_1_39 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_40 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h28 == _T_34[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_6;
      end else if (8'h28 == _T_31[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_5;
      end else if (8'h28 == _T_28[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_4;
      end else if (8'h28 == _T_25[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_3;
      end else if (8'h28 == _T_22[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_2;
      end else if (8'h28 == _T_19[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_1;
      end else if (8'h28 == _T_15[7:0]) begin
        image_1_40 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_41 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h29 == _T_34[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_6;
      end else if (8'h29 == _T_31[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_5;
      end else if (8'h29 == _T_28[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_4;
      end else if (8'h29 == _T_25[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_3;
      end else if (8'h29 == _T_22[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_2;
      end else if (8'h29 == _T_19[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_1;
      end else if (8'h29 == _T_15[7:0]) begin
        image_1_41 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_42 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2a == _T_34[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_6;
      end else if (8'h2a == _T_31[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_5;
      end else if (8'h2a == _T_28[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_4;
      end else if (8'h2a == _T_25[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_3;
      end else if (8'h2a == _T_22[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_2;
      end else if (8'h2a == _T_19[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_1;
      end else if (8'h2a == _T_15[7:0]) begin
        image_1_42 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_43 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2b == _T_34[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_6;
      end else if (8'h2b == _T_31[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_5;
      end else if (8'h2b == _T_28[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_4;
      end else if (8'h2b == _T_25[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_3;
      end else if (8'h2b == _T_22[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_2;
      end else if (8'h2b == _T_19[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_1;
      end else if (8'h2b == _T_15[7:0]) begin
        image_1_43 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_44 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2c == _T_34[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_6;
      end else if (8'h2c == _T_31[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_5;
      end else if (8'h2c == _T_28[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_4;
      end else if (8'h2c == _T_25[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_3;
      end else if (8'h2c == _T_22[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_2;
      end else if (8'h2c == _T_19[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_1;
      end else if (8'h2c == _T_15[7:0]) begin
        image_1_44 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_45 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2d == _T_34[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_6;
      end else if (8'h2d == _T_31[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_5;
      end else if (8'h2d == _T_28[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_4;
      end else if (8'h2d == _T_25[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_3;
      end else if (8'h2d == _T_22[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_2;
      end else if (8'h2d == _T_19[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_1;
      end else if (8'h2d == _T_15[7:0]) begin
        image_1_45 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_46 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2e == _T_34[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_6;
      end else if (8'h2e == _T_31[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_5;
      end else if (8'h2e == _T_28[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_4;
      end else if (8'h2e == _T_25[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_3;
      end else if (8'h2e == _T_22[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_2;
      end else if (8'h2e == _T_19[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_1;
      end else if (8'h2e == _T_15[7:0]) begin
        image_1_46 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_47 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2f == _T_34[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_6;
      end else if (8'h2f == _T_31[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_5;
      end else if (8'h2f == _T_28[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_4;
      end else if (8'h2f == _T_25[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_3;
      end else if (8'h2f == _T_22[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_2;
      end else if (8'h2f == _T_19[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_1;
      end else if (8'h2f == _T_15[7:0]) begin
        image_1_47 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_48 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h30 == _T_34[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_6;
      end else if (8'h30 == _T_31[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_5;
      end else if (8'h30 == _T_28[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_4;
      end else if (8'h30 == _T_25[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_3;
      end else if (8'h30 == _T_22[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_2;
      end else if (8'h30 == _T_19[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_1;
      end else if (8'h30 == _T_15[7:0]) begin
        image_1_48 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_49 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h31 == _T_34[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_6;
      end else if (8'h31 == _T_31[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_5;
      end else if (8'h31 == _T_28[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_4;
      end else if (8'h31 == _T_25[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_3;
      end else if (8'h31 == _T_22[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_2;
      end else if (8'h31 == _T_19[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_1;
      end else if (8'h31 == _T_15[7:0]) begin
        image_1_49 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_50 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h32 == _T_34[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_6;
      end else if (8'h32 == _T_31[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_5;
      end else if (8'h32 == _T_28[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_4;
      end else if (8'h32 == _T_25[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_3;
      end else if (8'h32 == _T_22[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_2;
      end else if (8'h32 == _T_19[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_1;
      end else if (8'h32 == _T_15[7:0]) begin
        image_1_50 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_51 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h33 == _T_34[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_6;
      end else if (8'h33 == _T_31[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_5;
      end else if (8'h33 == _T_28[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_4;
      end else if (8'h33 == _T_25[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_3;
      end else if (8'h33 == _T_22[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_2;
      end else if (8'h33 == _T_19[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_1;
      end else if (8'h33 == _T_15[7:0]) begin
        image_1_51 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_52 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h34 == _T_34[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_6;
      end else if (8'h34 == _T_31[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_5;
      end else if (8'h34 == _T_28[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_4;
      end else if (8'h34 == _T_25[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_3;
      end else if (8'h34 == _T_22[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_2;
      end else if (8'h34 == _T_19[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_1;
      end else if (8'h34 == _T_15[7:0]) begin
        image_1_52 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_53 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h35 == _T_34[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_6;
      end else if (8'h35 == _T_31[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_5;
      end else if (8'h35 == _T_28[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_4;
      end else if (8'h35 == _T_25[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_3;
      end else if (8'h35 == _T_22[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_2;
      end else if (8'h35 == _T_19[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_1;
      end else if (8'h35 == _T_15[7:0]) begin
        image_1_53 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_54 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h36 == _T_34[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_6;
      end else if (8'h36 == _T_31[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_5;
      end else if (8'h36 == _T_28[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_4;
      end else if (8'h36 == _T_25[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_3;
      end else if (8'h36 == _T_22[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_2;
      end else if (8'h36 == _T_19[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_1;
      end else if (8'h36 == _T_15[7:0]) begin
        image_1_54 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_55 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h37 == _T_34[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_6;
      end else if (8'h37 == _T_31[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_5;
      end else if (8'h37 == _T_28[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_4;
      end else if (8'h37 == _T_25[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_3;
      end else if (8'h37 == _T_22[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_2;
      end else if (8'h37 == _T_19[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_1;
      end else if (8'h37 == _T_15[7:0]) begin
        image_1_55 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_56 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h38 == _T_34[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_6;
      end else if (8'h38 == _T_31[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_5;
      end else if (8'h38 == _T_28[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_4;
      end else if (8'h38 == _T_25[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_3;
      end else if (8'h38 == _T_22[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_2;
      end else if (8'h38 == _T_19[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_1;
      end else if (8'h38 == _T_15[7:0]) begin
        image_1_56 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_57 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h39 == _T_34[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_6;
      end else if (8'h39 == _T_31[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_5;
      end else if (8'h39 == _T_28[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_4;
      end else if (8'h39 == _T_25[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_3;
      end else if (8'h39 == _T_22[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_2;
      end else if (8'h39 == _T_19[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_1;
      end else if (8'h39 == _T_15[7:0]) begin
        image_1_57 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_58 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3a == _T_34[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_6;
      end else if (8'h3a == _T_31[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_5;
      end else if (8'h3a == _T_28[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_4;
      end else if (8'h3a == _T_25[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_3;
      end else if (8'h3a == _T_22[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_2;
      end else if (8'h3a == _T_19[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_1;
      end else if (8'h3a == _T_15[7:0]) begin
        image_1_58 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_59 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3b == _T_34[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_6;
      end else if (8'h3b == _T_31[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_5;
      end else if (8'h3b == _T_28[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_4;
      end else if (8'h3b == _T_25[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_3;
      end else if (8'h3b == _T_22[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_2;
      end else if (8'h3b == _T_19[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_1;
      end else if (8'h3b == _T_15[7:0]) begin
        image_1_59 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_60 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3c == _T_34[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_6;
      end else if (8'h3c == _T_31[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_5;
      end else if (8'h3c == _T_28[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_4;
      end else if (8'h3c == _T_25[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_3;
      end else if (8'h3c == _T_22[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_2;
      end else if (8'h3c == _T_19[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_1;
      end else if (8'h3c == _T_15[7:0]) begin
        image_1_60 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_61 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3d == _T_34[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_6;
      end else if (8'h3d == _T_31[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_5;
      end else if (8'h3d == _T_28[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_4;
      end else if (8'h3d == _T_25[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_3;
      end else if (8'h3d == _T_22[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_2;
      end else if (8'h3d == _T_19[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_1;
      end else if (8'h3d == _T_15[7:0]) begin
        image_1_61 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_62 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3e == _T_34[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_6;
      end else if (8'h3e == _T_31[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_5;
      end else if (8'h3e == _T_28[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_4;
      end else if (8'h3e == _T_25[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_3;
      end else if (8'h3e == _T_22[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_2;
      end else if (8'h3e == _T_19[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_1;
      end else if (8'h3e == _T_15[7:0]) begin
        image_1_62 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_63 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3f == _T_34[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_6;
      end else if (8'h3f == _T_31[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_5;
      end else if (8'h3f == _T_28[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_4;
      end else if (8'h3f == _T_25[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_3;
      end else if (8'h3f == _T_22[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_2;
      end else if (8'h3f == _T_19[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_1;
      end else if (8'h3f == _T_15[7:0]) begin
        image_1_63 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_64 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h40 == _T_34[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_6;
      end else if (8'h40 == _T_31[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_5;
      end else if (8'h40 == _T_28[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_4;
      end else if (8'h40 == _T_25[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_3;
      end else if (8'h40 == _T_22[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_2;
      end else if (8'h40 == _T_19[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_1;
      end else if (8'h40 == _T_15[7:0]) begin
        image_1_64 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_65 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h41 == _T_34[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_6;
      end else if (8'h41 == _T_31[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_5;
      end else if (8'h41 == _T_28[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_4;
      end else if (8'h41 == _T_25[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_3;
      end else if (8'h41 == _T_22[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_2;
      end else if (8'h41 == _T_19[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_1;
      end else if (8'h41 == _T_15[7:0]) begin
        image_1_65 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_66 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h42 == _T_34[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_6;
      end else if (8'h42 == _T_31[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_5;
      end else if (8'h42 == _T_28[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_4;
      end else if (8'h42 == _T_25[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_3;
      end else if (8'h42 == _T_22[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_2;
      end else if (8'h42 == _T_19[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_1;
      end else if (8'h42 == _T_15[7:0]) begin
        image_1_66 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_67 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h43 == _T_34[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_6;
      end else if (8'h43 == _T_31[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_5;
      end else if (8'h43 == _T_28[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_4;
      end else if (8'h43 == _T_25[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_3;
      end else if (8'h43 == _T_22[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_2;
      end else if (8'h43 == _T_19[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_1;
      end else if (8'h43 == _T_15[7:0]) begin
        image_1_67 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_68 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h44 == _T_34[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_6;
      end else if (8'h44 == _T_31[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_5;
      end else if (8'h44 == _T_28[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_4;
      end else if (8'h44 == _T_25[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_3;
      end else if (8'h44 == _T_22[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_2;
      end else if (8'h44 == _T_19[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_1;
      end else if (8'h44 == _T_15[7:0]) begin
        image_1_68 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_69 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h45 == _T_34[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_6;
      end else if (8'h45 == _T_31[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_5;
      end else if (8'h45 == _T_28[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_4;
      end else if (8'h45 == _T_25[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_3;
      end else if (8'h45 == _T_22[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_2;
      end else if (8'h45 == _T_19[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_1;
      end else if (8'h45 == _T_15[7:0]) begin
        image_1_69 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_70 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h46 == _T_34[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_6;
      end else if (8'h46 == _T_31[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_5;
      end else if (8'h46 == _T_28[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_4;
      end else if (8'h46 == _T_25[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_3;
      end else if (8'h46 == _T_22[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_2;
      end else if (8'h46 == _T_19[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_1;
      end else if (8'h46 == _T_15[7:0]) begin
        image_1_70 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_71 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h47 == _T_34[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_6;
      end else if (8'h47 == _T_31[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_5;
      end else if (8'h47 == _T_28[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_4;
      end else if (8'h47 == _T_25[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_3;
      end else if (8'h47 == _T_22[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_2;
      end else if (8'h47 == _T_19[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_1;
      end else if (8'h47 == _T_15[7:0]) begin
        image_1_71 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_72 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h48 == _T_34[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_6;
      end else if (8'h48 == _T_31[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_5;
      end else if (8'h48 == _T_28[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_4;
      end else if (8'h48 == _T_25[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_3;
      end else if (8'h48 == _T_22[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_2;
      end else if (8'h48 == _T_19[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_1;
      end else if (8'h48 == _T_15[7:0]) begin
        image_1_72 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_73 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h49 == _T_34[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_6;
      end else if (8'h49 == _T_31[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_5;
      end else if (8'h49 == _T_28[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_4;
      end else if (8'h49 == _T_25[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_3;
      end else if (8'h49 == _T_22[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_2;
      end else if (8'h49 == _T_19[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_1;
      end else if (8'h49 == _T_15[7:0]) begin
        image_1_73 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_74 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4a == _T_34[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_6;
      end else if (8'h4a == _T_31[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_5;
      end else if (8'h4a == _T_28[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_4;
      end else if (8'h4a == _T_25[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_3;
      end else if (8'h4a == _T_22[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_2;
      end else if (8'h4a == _T_19[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_1;
      end else if (8'h4a == _T_15[7:0]) begin
        image_1_74 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_75 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4b == _T_34[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_6;
      end else if (8'h4b == _T_31[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_5;
      end else if (8'h4b == _T_28[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_4;
      end else if (8'h4b == _T_25[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_3;
      end else if (8'h4b == _T_22[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_2;
      end else if (8'h4b == _T_19[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_1;
      end else if (8'h4b == _T_15[7:0]) begin
        image_1_75 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_76 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4c == _T_34[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_6;
      end else if (8'h4c == _T_31[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_5;
      end else if (8'h4c == _T_28[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_4;
      end else if (8'h4c == _T_25[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_3;
      end else if (8'h4c == _T_22[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_2;
      end else if (8'h4c == _T_19[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_1;
      end else if (8'h4c == _T_15[7:0]) begin
        image_1_76 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_77 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4d == _T_34[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_6;
      end else if (8'h4d == _T_31[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_5;
      end else if (8'h4d == _T_28[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_4;
      end else if (8'h4d == _T_25[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_3;
      end else if (8'h4d == _T_22[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_2;
      end else if (8'h4d == _T_19[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_1;
      end else if (8'h4d == _T_15[7:0]) begin
        image_1_77 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_78 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4e == _T_34[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_6;
      end else if (8'h4e == _T_31[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_5;
      end else if (8'h4e == _T_28[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_4;
      end else if (8'h4e == _T_25[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_3;
      end else if (8'h4e == _T_22[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_2;
      end else if (8'h4e == _T_19[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_1;
      end else if (8'h4e == _T_15[7:0]) begin
        image_1_78 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_79 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4f == _T_34[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_6;
      end else if (8'h4f == _T_31[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_5;
      end else if (8'h4f == _T_28[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_4;
      end else if (8'h4f == _T_25[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_3;
      end else if (8'h4f == _T_22[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_2;
      end else if (8'h4f == _T_19[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_1;
      end else if (8'h4f == _T_15[7:0]) begin
        image_1_79 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_80 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h50 == _T_34[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_6;
      end else if (8'h50 == _T_31[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_5;
      end else if (8'h50 == _T_28[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_4;
      end else if (8'h50 == _T_25[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_3;
      end else if (8'h50 == _T_22[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_2;
      end else if (8'h50 == _T_19[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_1;
      end else if (8'h50 == _T_15[7:0]) begin
        image_1_80 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_81 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h51 == _T_34[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_6;
      end else if (8'h51 == _T_31[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_5;
      end else if (8'h51 == _T_28[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_4;
      end else if (8'h51 == _T_25[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_3;
      end else if (8'h51 == _T_22[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_2;
      end else if (8'h51 == _T_19[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_1;
      end else if (8'h51 == _T_15[7:0]) begin
        image_1_81 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_82 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h52 == _T_34[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_6;
      end else if (8'h52 == _T_31[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_5;
      end else if (8'h52 == _T_28[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_4;
      end else if (8'h52 == _T_25[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_3;
      end else if (8'h52 == _T_22[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_2;
      end else if (8'h52 == _T_19[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_1;
      end else if (8'h52 == _T_15[7:0]) begin
        image_1_82 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_83 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h53 == _T_34[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_6;
      end else if (8'h53 == _T_31[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_5;
      end else if (8'h53 == _T_28[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_4;
      end else if (8'h53 == _T_25[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_3;
      end else if (8'h53 == _T_22[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_2;
      end else if (8'h53 == _T_19[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_1;
      end else if (8'h53 == _T_15[7:0]) begin
        image_1_83 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_84 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h54 == _T_34[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_6;
      end else if (8'h54 == _T_31[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_5;
      end else if (8'h54 == _T_28[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_4;
      end else if (8'h54 == _T_25[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_3;
      end else if (8'h54 == _T_22[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_2;
      end else if (8'h54 == _T_19[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_1;
      end else if (8'h54 == _T_15[7:0]) begin
        image_1_84 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_85 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h55 == _T_34[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_6;
      end else if (8'h55 == _T_31[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_5;
      end else if (8'h55 == _T_28[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_4;
      end else if (8'h55 == _T_25[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_3;
      end else if (8'h55 == _T_22[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_2;
      end else if (8'h55 == _T_19[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_1;
      end else if (8'h55 == _T_15[7:0]) begin
        image_1_85 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_86 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h56 == _T_34[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_6;
      end else if (8'h56 == _T_31[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_5;
      end else if (8'h56 == _T_28[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_4;
      end else if (8'h56 == _T_25[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_3;
      end else if (8'h56 == _T_22[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_2;
      end else if (8'h56 == _T_19[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_1;
      end else if (8'h56 == _T_15[7:0]) begin
        image_1_86 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_87 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h57 == _T_34[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_6;
      end else if (8'h57 == _T_31[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_5;
      end else if (8'h57 == _T_28[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_4;
      end else if (8'h57 == _T_25[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_3;
      end else if (8'h57 == _T_22[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_2;
      end else if (8'h57 == _T_19[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_1;
      end else if (8'h57 == _T_15[7:0]) begin
        image_1_87 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_88 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h58 == _T_34[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_6;
      end else if (8'h58 == _T_31[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_5;
      end else if (8'h58 == _T_28[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_4;
      end else if (8'h58 == _T_25[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_3;
      end else if (8'h58 == _T_22[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_2;
      end else if (8'h58 == _T_19[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_1;
      end else if (8'h58 == _T_15[7:0]) begin
        image_1_88 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_89 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h59 == _T_34[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_6;
      end else if (8'h59 == _T_31[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_5;
      end else if (8'h59 == _T_28[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_4;
      end else if (8'h59 == _T_25[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_3;
      end else if (8'h59 == _T_22[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_2;
      end else if (8'h59 == _T_19[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_1;
      end else if (8'h59 == _T_15[7:0]) begin
        image_1_89 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_90 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5a == _T_34[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_6;
      end else if (8'h5a == _T_31[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_5;
      end else if (8'h5a == _T_28[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_4;
      end else if (8'h5a == _T_25[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_3;
      end else if (8'h5a == _T_22[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_2;
      end else if (8'h5a == _T_19[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_1;
      end else if (8'h5a == _T_15[7:0]) begin
        image_1_90 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_91 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5b == _T_34[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_6;
      end else if (8'h5b == _T_31[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_5;
      end else if (8'h5b == _T_28[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_4;
      end else if (8'h5b == _T_25[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_3;
      end else if (8'h5b == _T_22[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_2;
      end else if (8'h5b == _T_19[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_1;
      end else if (8'h5b == _T_15[7:0]) begin
        image_1_91 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_92 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5c == _T_34[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_6;
      end else if (8'h5c == _T_31[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_5;
      end else if (8'h5c == _T_28[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_4;
      end else if (8'h5c == _T_25[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_3;
      end else if (8'h5c == _T_22[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_2;
      end else if (8'h5c == _T_19[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_1;
      end else if (8'h5c == _T_15[7:0]) begin
        image_1_92 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_93 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5d == _T_34[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_6;
      end else if (8'h5d == _T_31[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_5;
      end else if (8'h5d == _T_28[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_4;
      end else if (8'h5d == _T_25[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_3;
      end else if (8'h5d == _T_22[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_2;
      end else if (8'h5d == _T_19[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_1;
      end else if (8'h5d == _T_15[7:0]) begin
        image_1_93 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_94 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5e == _T_34[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_6;
      end else if (8'h5e == _T_31[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_5;
      end else if (8'h5e == _T_28[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_4;
      end else if (8'h5e == _T_25[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_3;
      end else if (8'h5e == _T_22[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_2;
      end else if (8'h5e == _T_19[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_1;
      end else if (8'h5e == _T_15[7:0]) begin
        image_1_94 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_95 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5f == _T_34[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_6;
      end else if (8'h5f == _T_31[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_5;
      end else if (8'h5f == _T_28[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_4;
      end else if (8'h5f == _T_25[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_3;
      end else if (8'h5f == _T_22[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_2;
      end else if (8'h5f == _T_19[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_1;
      end else if (8'h5f == _T_15[7:0]) begin
        image_1_95 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_96 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h60 == _T_34[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_6;
      end else if (8'h60 == _T_31[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_5;
      end else if (8'h60 == _T_28[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_4;
      end else if (8'h60 == _T_25[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_3;
      end else if (8'h60 == _T_22[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_2;
      end else if (8'h60 == _T_19[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_1;
      end else if (8'h60 == _T_15[7:0]) begin
        image_1_96 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_97 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h61 == _T_34[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_6;
      end else if (8'h61 == _T_31[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_5;
      end else if (8'h61 == _T_28[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_4;
      end else if (8'h61 == _T_25[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_3;
      end else if (8'h61 == _T_22[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_2;
      end else if (8'h61 == _T_19[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_1;
      end else if (8'h61 == _T_15[7:0]) begin
        image_1_97 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_98 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h62 == _T_34[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_6;
      end else if (8'h62 == _T_31[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_5;
      end else if (8'h62 == _T_28[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_4;
      end else if (8'h62 == _T_25[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_3;
      end else if (8'h62 == _T_22[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_2;
      end else if (8'h62 == _T_19[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_1;
      end else if (8'h62 == _T_15[7:0]) begin
        image_1_98 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_99 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h63 == _T_34[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_6;
      end else if (8'h63 == _T_31[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_5;
      end else if (8'h63 == _T_28[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_4;
      end else if (8'h63 == _T_25[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_3;
      end else if (8'h63 == _T_22[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_2;
      end else if (8'h63 == _T_19[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_1;
      end else if (8'h63 == _T_15[7:0]) begin
        image_1_99 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_100 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h64 == _T_34[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_6;
      end else if (8'h64 == _T_31[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_5;
      end else if (8'h64 == _T_28[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_4;
      end else if (8'h64 == _T_25[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_3;
      end else if (8'h64 == _T_22[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_2;
      end else if (8'h64 == _T_19[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_1;
      end else if (8'h64 == _T_15[7:0]) begin
        image_1_100 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_101 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h65 == _T_34[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_6;
      end else if (8'h65 == _T_31[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_5;
      end else if (8'h65 == _T_28[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_4;
      end else if (8'h65 == _T_25[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_3;
      end else if (8'h65 == _T_22[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_2;
      end else if (8'h65 == _T_19[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_1;
      end else if (8'h65 == _T_15[7:0]) begin
        image_1_101 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_102 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h66 == _T_34[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_6;
      end else if (8'h66 == _T_31[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_5;
      end else if (8'h66 == _T_28[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_4;
      end else if (8'h66 == _T_25[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_3;
      end else if (8'h66 == _T_22[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_2;
      end else if (8'h66 == _T_19[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_1;
      end else if (8'h66 == _T_15[7:0]) begin
        image_1_102 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_103 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h67 == _T_34[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_6;
      end else if (8'h67 == _T_31[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_5;
      end else if (8'h67 == _T_28[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_4;
      end else if (8'h67 == _T_25[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_3;
      end else if (8'h67 == _T_22[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_2;
      end else if (8'h67 == _T_19[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_1;
      end else if (8'h67 == _T_15[7:0]) begin
        image_1_103 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_104 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h68 == _T_34[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_6;
      end else if (8'h68 == _T_31[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_5;
      end else if (8'h68 == _T_28[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_4;
      end else if (8'h68 == _T_25[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_3;
      end else if (8'h68 == _T_22[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_2;
      end else if (8'h68 == _T_19[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_1;
      end else if (8'h68 == _T_15[7:0]) begin
        image_1_104 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_105 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h69 == _T_34[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_6;
      end else if (8'h69 == _T_31[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_5;
      end else if (8'h69 == _T_28[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_4;
      end else if (8'h69 == _T_25[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_3;
      end else if (8'h69 == _T_22[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_2;
      end else if (8'h69 == _T_19[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_1;
      end else if (8'h69 == _T_15[7:0]) begin
        image_1_105 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_106 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6a == _T_34[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_6;
      end else if (8'h6a == _T_31[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_5;
      end else if (8'h6a == _T_28[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_4;
      end else if (8'h6a == _T_25[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_3;
      end else if (8'h6a == _T_22[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_2;
      end else if (8'h6a == _T_19[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_1;
      end else if (8'h6a == _T_15[7:0]) begin
        image_1_106 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_107 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6b == _T_34[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_6;
      end else if (8'h6b == _T_31[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_5;
      end else if (8'h6b == _T_28[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_4;
      end else if (8'h6b == _T_25[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_3;
      end else if (8'h6b == _T_22[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_2;
      end else if (8'h6b == _T_19[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_1;
      end else if (8'h6b == _T_15[7:0]) begin
        image_1_107 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_108 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6c == _T_34[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_6;
      end else if (8'h6c == _T_31[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_5;
      end else if (8'h6c == _T_28[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_4;
      end else if (8'h6c == _T_25[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_3;
      end else if (8'h6c == _T_22[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_2;
      end else if (8'h6c == _T_19[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_1;
      end else if (8'h6c == _T_15[7:0]) begin
        image_1_108 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_109 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6d == _T_34[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_6;
      end else if (8'h6d == _T_31[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_5;
      end else if (8'h6d == _T_28[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_4;
      end else if (8'h6d == _T_25[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_3;
      end else if (8'h6d == _T_22[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_2;
      end else if (8'h6d == _T_19[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_1;
      end else if (8'h6d == _T_15[7:0]) begin
        image_1_109 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_110 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6e == _T_34[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_6;
      end else if (8'h6e == _T_31[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_5;
      end else if (8'h6e == _T_28[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_4;
      end else if (8'h6e == _T_25[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_3;
      end else if (8'h6e == _T_22[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_2;
      end else if (8'h6e == _T_19[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_1;
      end else if (8'h6e == _T_15[7:0]) begin
        image_1_110 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_111 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6f == _T_34[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_6;
      end else if (8'h6f == _T_31[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_5;
      end else if (8'h6f == _T_28[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_4;
      end else if (8'h6f == _T_25[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_3;
      end else if (8'h6f == _T_22[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_2;
      end else if (8'h6f == _T_19[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_1;
      end else if (8'h6f == _T_15[7:0]) begin
        image_1_111 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_112 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h70 == _T_34[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_6;
      end else if (8'h70 == _T_31[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_5;
      end else if (8'h70 == _T_28[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_4;
      end else if (8'h70 == _T_25[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_3;
      end else if (8'h70 == _T_22[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_2;
      end else if (8'h70 == _T_19[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_1;
      end else if (8'h70 == _T_15[7:0]) begin
        image_1_112 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_113 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h71 == _T_34[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_6;
      end else if (8'h71 == _T_31[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_5;
      end else if (8'h71 == _T_28[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_4;
      end else if (8'h71 == _T_25[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_3;
      end else if (8'h71 == _T_22[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_2;
      end else if (8'h71 == _T_19[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_1;
      end else if (8'h71 == _T_15[7:0]) begin
        image_1_113 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_114 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h72 == _T_34[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_6;
      end else if (8'h72 == _T_31[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_5;
      end else if (8'h72 == _T_28[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_4;
      end else if (8'h72 == _T_25[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_3;
      end else if (8'h72 == _T_22[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_2;
      end else if (8'h72 == _T_19[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_1;
      end else if (8'h72 == _T_15[7:0]) begin
        image_1_114 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_115 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h73 == _T_34[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_6;
      end else if (8'h73 == _T_31[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_5;
      end else if (8'h73 == _T_28[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_4;
      end else if (8'h73 == _T_25[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_3;
      end else if (8'h73 == _T_22[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_2;
      end else if (8'h73 == _T_19[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_1;
      end else if (8'h73 == _T_15[7:0]) begin
        image_1_115 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_116 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h74 == _T_34[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_6;
      end else if (8'h74 == _T_31[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_5;
      end else if (8'h74 == _T_28[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_4;
      end else if (8'h74 == _T_25[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_3;
      end else if (8'h74 == _T_22[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_2;
      end else if (8'h74 == _T_19[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_1;
      end else if (8'h74 == _T_15[7:0]) begin
        image_1_116 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_117 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h75 == _T_34[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_6;
      end else if (8'h75 == _T_31[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_5;
      end else if (8'h75 == _T_28[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_4;
      end else if (8'h75 == _T_25[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_3;
      end else if (8'h75 == _T_22[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_2;
      end else if (8'h75 == _T_19[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_1;
      end else if (8'h75 == _T_15[7:0]) begin
        image_1_117 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_118 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h76 == _T_34[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_6;
      end else if (8'h76 == _T_31[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_5;
      end else if (8'h76 == _T_28[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_4;
      end else if (8'h76 == _T_25[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_3;
      end else if (8'h76 == _T_22[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_2;
      end else if (8'h76 == _T_19[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_1;
      end else if (8'h76 == _T_15[7:0]) begin
        image_1_118 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_119 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h77 == _T_34[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_6;
      end else if (8'h77 == _T_31[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_5;
      end else if (8'h77 == _T_28[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_4;
      end else if (8'h77 == _T_25[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_3;
      end else if (8'h77 == _T_22[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_2;
      end else if (8'h77 == _T_19[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_1;
      end else if (8'h77 == _T_15[7:0]) begin
        image_1_119 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_120 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h78 == _T_34[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_6;
      end else if (8'h78 == _T_31[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_5;
      end else if (8'h78 == _T_28[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_4;
      end else if (8'h78 == _T_25[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_3;
      end else if (8'h78 == _T_22[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_2;
      end else if (8'h78 == _T_19[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_1;
      end else if (8'h78 == _T_15[7:0]) begin
        image_1_120 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_121 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h79 == _T_34[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_6;
      end else if (8'h79 == _T_31[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_5;
      end else if (8'h79 == _T_28[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_4;
      end else if (8'h79 == _T_25[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_3;
      end else if (8'h79 == _T_22[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_2;
      end else if (8'h79 == _T_19[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_1;
      end else if (8'h79 == _T_15[7:0]) begin
        image_1_121 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_122 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7a == _T_34[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_6;
      end else if (8'h7a == _T_31[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_5;
      end else if (8'h7a == _T_28[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_4;
      end else if (8'h7a == _T_25[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_3;
      end else if (8'h7a == _T_22[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_2;
      end else if (8'h7a == _T_19[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_1;
      end else if (8'h7a == _T_15[7:0]) begin
        image_1_122 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_123 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7b == _T_34[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_6;
      end else if (8'h7b == _T_31[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_5;
      end else if (8'h7b == _T_28[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_4;
      end else if (8'h7b == _T_25[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_3;
      end else if (8'h7b == _T_22[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_2;
      end else if (8'h7b == _T_19[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_1;
      end else if (8'h7b == _T_15[7:0]) begin
        image_1_123 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_124 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7c == _T_34[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_6;
      end else if (8'h7c == _T_31[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_5;
      end else if (8'h7c == _T_28[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_4;
      end else if (8'h7c == _T_25[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_3;
      end else if (8'h7c == _T_22[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_2;
      end else if (8'h7c == _T_19[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_1;
      end else if (8'h7c == _T_15[7:0]) begin
        image_1_124 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_125 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7d == _T_34[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_6;
      end else if (8'h7d == _T_31[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_5;
      end else if (8'h7d == _T_28[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_4;
      end else if (8'h7d == _T_25[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_3;
      end else if (8'h7d == _T_22[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_2;
      end else if (8'h7d == _T_19[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_1;
      end else if (8'h7d == _T_15[7:0]) begin
        image_1_125 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_126 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7e == _T_34[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_6;
      end else if (8'h7e == _T_31[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_5;
      end else if (8'h7e == _T_28[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_4;
      end else if (8'h7e == _T_25[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_3;
      end else if (8'h7e == _T_22[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_2;
      end else if (8'h7e == _T_19[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_1;
      end else if (8'h7e == _T_15[7:0]) begin
        image_1_126 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_127 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7f == _T_34[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_6;
      end else if (8'h7f == _T_31[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_5;
      end else if (8'h7f == _T_28[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_4;
      end else if (8'h7f == _T_25[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_3;
      end else if (8'h7f == _T_22[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_2;
      end else if (8'h7f == _T_19[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_1;
      end else if (8'h7f == _T_15[7:0]) begin
        image_1_127 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_128 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h80 == _T_34[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_6;
      end else if (8'h80 == _T_31[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_5;
      end else if (8'h80 == _T_28[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_4;
      end else if (8'h80 == _T_25[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_3;
      end else if (8'h80 == _T_22[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_2;
      end else if (8'h80 == _T_19[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_1;
      end else if (8'h80 == _T_15[7:0]) begin
        image_1_128 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_129 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h81 == _T_34[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_6;
      end else if (8'h81 == _T_31[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_5;
      end else if (8'h81 == _T_28[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_4;
      end else if (8'h81 == _T_25[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_3;
      end else if (8'h81 == _T_22[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_2;
      end else if (8'h81 == _T_19[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_1;
      end else if (8'h81 == _T_15[7:0]) begin
        image_1_129 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_130 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h82 == _T_34[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_6;
      end else if (8'h82 == _T_31[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_5;
      end else if (8'h82 == _T_28[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_4;
      end else if (8'h82 == _T_25[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_3;
      end else if (8'h82 == _T_22[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_2;
      end else if (8'h82 == _T_19[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_1;
      end else if (8'h82 == _T_15[7:0]) begin
        image_1_130 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_131 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h83 == _T_34[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_6;
      end else if (8'h83 == _T_31[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_5;
      end else if (8'h83 == _T_28[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_4;
      end else if (8'h83 == _T_25[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_3;
      end else if (8'h83 == _T_22[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_2;
      end else if (8'h83 == _T_19[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_1;
      end else if (8'h83 == _T_15[7:0]) begin
        image_1_131 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_132 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h84 == _T_34[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_6;
      end else if (8'h84 == _T_31[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_5;
      end else if (8'h84 == _T_28[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_4;
      end else if (8'h84 == _T_25[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_3;
      end else if (8'h84 == _T_22[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_2;
      end else if (8'h84 == _T_19[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_1;
      end else if (8'h84 == _T_15[7:0]) begin
        image_1_132 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_133 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h85 == _T_34[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_6;
      end else if (8'h85 == _T_31[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_5;
      end else if (8'h85 == _T_28[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_4;
      end else if (8'h85 == _T_25[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_3;
      end else if (8'h85 == _T_22[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_2;
      end else if (8'h85 == _T_19[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_1;
      end else if (8'h85 == _T_15[7:0]) begin
        image_1_133 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_134 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h86 == _T_34[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_6;
      end else if (8'h86 == _T_31[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_5;
      end else if (8'h86 == _T_28[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_4;
      end else if (8'h86 == _T_25[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_3;
      end else if (8'h86 == _T_22[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_2;
      end else if (8'h86 == _T_19[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_1;
      end else if (8'h86 == _T_15[7:0]) begin
        image_1_134 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_135 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h87 == _T_34[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_6;
      end else if (8'h87 == _T_31[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_5;
      end else if (8'h87 == _T_28[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_4;
      end else if (8'h87 == _T_25[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_3;
      end else if (8'h87 == _T_22[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_2;
      end else if (8'h87 == _T_19[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_1;
      end else if (8'h87 == _T_15[7:0]) begin
        image_1_135 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_136 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h88 == _T_34[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_6;
      end else if (8'h88 == _T_31[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_5;
      end else if (8'h88 == _T_28[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_4;
      end else if (8'h88 == _T_25[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_3;
      end else if (8'h88 == _T_22[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_2;
      end else if (8'h88 == _T_19[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_1;
      end else if (8'h88 == _T_15[7:0]) begin
        image_1_136 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_137 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h89 == _T_34[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_6;
      end else if (8'h89 == _T_31[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_5;
      end else if (8'h89 == _T_28[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_4;
      end else if (8'h89 == _T_25[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_3;
      end else if (8'h89 == _T_22[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_2;
      end else if (8'h89 == _T_19[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_1;
      end else if (8'h89 == _T_15[7:0]) begin
        image_1_137 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_138 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8a == _T_34[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_6;
      end else if (8'h8a == _T_31[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_5;
      end else if (8'h8a == _T_28[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_4;
      end else if (8'h8a == _T_25[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_3;
      end else if (8'h8a == _T_22[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_2;
      end else if (8'h8a == _T_19[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_1;
      end else if (8'h8a == _T_15[7:0]) begin
        image_1_138 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_139 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8b == _T_34[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_6;
      end else if (8'h8b == _T_31[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_5;
      end else if (8'h8b == _T_28[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_4;
      end else if (8'h8b == _T_25[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_3;
      end else if (8'h8b == _T_22[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_2;
      end else if (8'h8b == _T_19[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_1;
      end else if (8'h8b == _T_15[7:0]) begin
        image_1_139 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_140 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8c == _T_34[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_6;
      end else if (8'h8c == _T_31[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_5;
      end else if (8'h8c == _T_28[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_4;
      end else if (8'h8c == _T_25[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_3;
      end else if (8'h8c == _T_22[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_2;
      end else if (8'h8c == _T_19[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_1;
      end else if (8'h8c == _T_15[7:0]) begin
        image_1_140 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_141 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8d == _T_34[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_6;
      end else if (8'h8d == _T_31[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_5;
      end else if (8'h8d == _T_28[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_4;
      end else if (8'h8d == _T_25[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_3;
      end else if (8'h8d == _T_22[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_2;
      end else if (8'h8d == _T_19[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_1;
      end else if (8'h8d == _T_15[7:0]) begin
        image_1_141 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_142 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8e == _T_34[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_6;
      end else if (8'h8e == _T_31[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_5;
      end else if (8'h8e == _T_28[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_4;
      end else if (8'h8e == _T_25[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_3;
      end else if (8'h8e == _T_22[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_2;
      end else if (8'h8e == _T_19[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_1;
      end else if (8'h8e == _T_15[7:0]) begin
        image_1_142 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_143 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8f == _T_34[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_6;
      end else if (8'h8f == _T_31[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_5;
      end else if (8'h8f == _T_28[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_4;
      end else if (8'h8f == _T_25[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_3;
      end else if (8'h8f == _T_22[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_2;
      end else if (8'h8f == _T_19[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_1;
      end else if (8'h8f == _T_15[7:0]) begin
        image_1_143 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_144 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h90 == _T_34[7:0]) begin
        image_1_144 <= io_pixelVal_in_1_6;
      end else if (8'h90 == _T_31[7:0]) begin
        image_1_144 <= io_pixelVal_in_1_5;
      end else if (8'h90 == _T_28[7:0]) begin
        image_1_144 <= io_pixelVal_in_1_4;
      end else if (8'h90 == _T_25[7:0]) begin
        image_1_144 <= io_pixelVal_in_1_3;
      end else if (8'h90 == _T_22[7:0]) begin
        image_1_144 <= io_pixelVal_in_1_2;
      end else if (8'h90 == _T_19[7:0]) begin
        image_1_144 <= io_pixelVal_in_1_1;
      end else if (8'h90 == _T_15[7:0]) begin
        image_1_144 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_145 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h91 == _T_34[7:0]) begin
        image_1_145 <= io_pixelVal_in_1_6;
      end else if (8'h91 == _T_31[7:0]) begin
        image_1_145 <= io_pixelVal_in_1_5;
      end else if (8'h91 == _T_28[7:0]) begin
        image_1_145 <= io_pixelVal_in_1_4;
      end else if (8'h91 == _T_25[7:0]) begin
        image_1_145 <= io_pixelVal_in_1_3;
      end else if (8'h91 == _T_22[7:0]) begin
        image_1_145 <= io_pixelVal_in_1_2;
      end else if (8'h91 == _T_19[7:0]) begin
        image_1_145 <= io_pixelVal_in_1_1;
      end else if (8'h91 == _T_15[7:0]) begin
        image_1_145 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_146 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h92 == _T_34[7:0]) begin
        image_1_146 <= io_pixelVal_in_1_6;
      end else if (8'h92 == _T_31[7:0]) begin
        image_1_146 <= io_pixelVal_in_1_5;
      end else if (8'h92 == _T_28[7:0]) begin
        image_1_146 <= io_pixelVal_in_1_4;
      end else if (8'h92 == _T_25[7:0]) begin
        image_1_146 <= io_pixelVal_in_1_3;
      end else if (8'h92 == _T_22[7:0]) begin
        image_1_146 <= io_pixelVal_in_1_2;
      end else if (8'h92 == _T_19[7:0]) begin
        image_1_146 <= io_pixelVal_in_1_1;
      end else if (8'h92 == _T_15[7:0]) begin
        image_1_146 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_147 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h93 == _T_34[7:0]) begin
        image_1_147 <= io_pixelVal_in_1_6;
      end else if (8'h93 == _T_31[7:0]) begin
        image_1_147 <= io_pixelVal_in_1_5;
      end else if (8'h93 == _T_28[7:0]) begin
        image_1_147 <= io_pixelVal_in_1_4;
      end else if (8'h93 == _T_25[7:0]) begin
        image_1_147 <= io_pixelVal_in_1_3;
      end else if (8'h93 == _T_22[7:0]) begin
        image_1_147 <= io_pixelVal_in_1_2;
      end else if (8'h93 == _T_19[7:0]) begin
        image_1_147 <= io_pixelVal_in_1_1;
      end else if (8'h93 == _T_15[7:0]) begin
        image_1_147 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_148 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h94 == _T_34[7:0]) begin
        image_1_148 <= io_pixelVal_in_1_6;
      end else if (8'h94 == _T_31[7:0]) begin
        image_1_148 <= io_pixelVal_in_1_5;
      end else if (8'h94 == _T_28[7:0]) begin
        image_1_148 <= io_pixelVal_in_1_4;
      end else if (8'h94 == _T_25[7:0]) begin
        image_1_148 <= io_pixelVal_in_1_3;
      end else if (8'h94 == _T_22[7:0]) begin
        image_1_148 <= io_pixelVal_in_1_2;
      end else if (8'h94 == _T_19[7:0]) begin
        image_1_148 <= io_pixelVal_in_1_1;
      end else if (8'h94 == _T_15[7:0]) begin
        image_1_148 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_149 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h95 == _T_34[7:0]) begin
        image_1_149 <= io_pixelVal_in_1_6;
      end else if (8'h95 == _T_31[7:0]) begin
        image_1_149 <= io_pixelVal_in_1_5;
      end else if (8'h95 == _T_28[7:0]) begin
        image_1_149 <= io_pixelVal_in_1_4;
      end else if (8'h95 == _T_25[7:0]) begin
        image_1_149 <= io_pixelVal_in_1_3;
      end else if (8'h95 == _T_22[7:0]) begin
        image_1_149 <= io_pixelVal_in_1_2;
      end else if (8'h95 == _T_19[7:0]) begin
        image_1_149 <= io_pixelVal_in_1_1;
      end else if (8'h95 == _T_15[7:0]) begin
        image_1_149 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_150 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h96 == _T_34[7:0]) begin
        image_1_150 <= io_pixelVal_in_1_6;
      end else if (8'h96 == _T_31[7:0]) begin
        image_1_150 <= io_pixelVal_in_1_5;
      end else if (8'h96 == _T_28[7:0]) begin
        image_1_150 <= io_pixelVal_in_1_4;
      end else if (8'h96 == _T_25[7:0]) begin
        image_1_150 <= io_pixelVal_in_1_3;
      end else if (8'h96 == _T_22[7:0]) begin
        image_1_150 <= io_pixelVal_in_1_2;
      end else if (8'h96 == _T_19[7:0]) begin
        image_1_150 <= io_pixelVal_in_1_1;
      end else if (8'h96 == _T_15[7:0]) begin
        image_1_150 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_151 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h97 == _T_34[7:0]) begin
        image_1_151 <= io_pixelVal_in_1_6;
      end else if (8'h97 == _T_31[7:0]) begin
        image_1_151 <= io_pixelVal_in_1_5;
      end else if (8'h97 == _T_28[7:0]) begin
        image_1_151 <= io_pixelVal_in_1_4;
      end else if (8'h97 == _T_25[7:0]) begin
        image_1_151 <= io_pixelVal_in_1_3;
      end else if (8'h97 == _T_22[7:0]) begin
        image_1_151 <= io_pixelVal_in_1_2;
      end else if (8'h97 == _T_19[7:0]) begin
        image_1_151 <= io_pixelVal_in_1_1;
      end else if (8'h97 == _T_15[7:0]) begin
        image_1_151 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_152 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h98 == _T_34[7:0]) begin
        image_1_152 <= io_pixelVal_in_1_6;
      end else if (8'h98 == _T_31[7:0]) begin
        image_1_152 <= io_pixelVal_in_1_5;
      end else if (8'h98 == _T_28[7:0]) begin
        image_1_152 <= io_pixelVal_in_1_4;
      end else if (8'h98 == _T_25[7:0]) begin
        image_1_152 <= io_pixelVal_in_1_3;
      end else if (8'h98 == _T_22[7:0]) begin
        image_1_152 <= io_pixelVal_in_1_2;
      end else if (8'h98 == _T_19[7:0]) begin
        image_1_152 <= io_pixelVal_in_1_1;
      end else if (8'h98 == _T_15[7:0]) begin
        image_1_152 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_153 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h99 == _T_34[7:0]) begin
        image_1_153 <= io_pixelVal_in_1_6;
      end else if (8'h99 == _T_31[7:0]) begin
        image_1_153 <= io_pixelVal_in_1_5;
      end else if (8'h99 == _T_28[7:0]) begin
        image_1_153 <= io_pixelVal_in_1_4;
      end else if (8'h99 == _T_25[7:0]) begin
        image_1_153 <= io_pixelVal_in_1_3;
      end else if (8'h99 == _T_22[7:0]) begin
        image_1_153 <= io_pixelVal_in_1_2;
      end else if (8'h99 == _T_19[7:0]) begin
        image_1_153 <= io_pixelVal_in_1_1;
      end else if (8'h99 == _T_15[7:0]) begin
        image_1_153 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_154 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9a == _T_34[7:0]) begin
        image_1_154 <= io_pixelVal_in_1_6;
      end else if (8'h9a == _T_31[7:0]) begin
        image_1_154 <= io_pixelVal_in_1_5;
      end else if (8'h9a == _T_28[7:0]) begin
        image_1_154 <= io_pixelVal_in_1_4;
      end else if (8'h9a == _T_25[7:0]) begin
        image_1_154 <= io_pixelVal_in_1_3;
      end else if (8'h9a == _T_22[7:0]) begin
        image_1_154 <= io_pixelVal_in_1_2;
      end else if (8'h9a == _T_19[7:0]) begin
        image_1_154 <= io_pixelVal_in_1_1;
      end else if (8'h9a == _T_15[7:0]) begin
        image_1_154 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_155 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9b == _T_34[7:0]) begin
        image_1_155 <= io_pixelVal_in_1_6;
      end else if (8'h9b == _T_31[7:0]) begin
        image_1_155 <= io_pixelVal_in_1_5;
      end else if (8'h9b == _T_28[7:0]) begin
        image_1_155 <= io_pixelVal_in_1_4;
      end else if (8'h9b == _T_25[7:0]) begin
        image_1_155 <= io_pixelVal_in_1_3;
      end else if (8'h9b == _T_22[7:0]) begin
        image_1_155 <= io_pixelVal_in_1_2;
      end else if (8'h9b == _T_19[7:0]) begin
        image_1_155 <= io_pixelVal_in_1_1;
      end else if (8'h9b == _T_15[7:0]) begin
        image_1_155 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_156 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9c == _T_34[7:0]) begin
        image_1_156 <= io_pixelVal_in_1_6;
      end else if (8'h9c == _T_31[7:0]) begin
        image_1_156 <= io_pixelVal_in_1_5;
      end else if (8'h9c == _T_28[7:0]) begin
        image_1_156 <= io_pixelVal_in_1_4;
      end else if (8'h9c == _T_25[7:0]) begin
        image_1_156 <= io_pixelVal_in_1_3;
      end else if (8'h9c == _T_22[7:0]) begin
        image_1_156 <= io_pixelVal_in_1_2;
      end else if (8'h9c == _T_19[7:0]) begin
        image_1_156 <= io_pixelVal_in_1_1;
      end else if (8'h9c == _T_15[7:0]) begin
        image_1_156 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_157 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9d == _T_34[7:0]) begin
        image_1_157 <= io_pixelVal_in_1_6;
      end else if (8'h9d == _T_31[7:0]) begin
        image_1_157 <= io_pixelVal_in_1_5;
      end else if (8'h9d == _T_28[7:0]) begin
        image_1_157 <= io_pixelVal_in_1_4;
      end else if (8'h9d == _T_25[7:0]) begin
        image_1_157 <= io_pixelVal_in_1_3;
      end else if (8'h9d == _T_22[7:0]) begin
        image_1_157 <= io_pixelVal_in_1_2;
      end else if (8'h9d == _T_19[7:0]) begin
        image_1_157 <= io_pixelVal_in_1_1;
      end else if (8'h9d == _T_15[7:0]) begin
        image_1_157 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_158 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9e == _T_34[7:0]) begin
        image_1_158 <= io_pixelVal_in_1_6;
      end else if (8'h9e == _T_31[7:0]) begin
        image_1_158 <= io_pixelVal_in_1_5;
      end else if (8'h9e == _T_28[7:0]) begin
        image_1_158 <= io_pixelVal_in_1_4;
      end else if (8'h9e == _T_25[7:0]) begin
        image_1_158 <= io_pixelVal_in_1_3;
      end else if (8'h9e == _T_22[7:0]) begin
        image_1_158 <= io_pixelVal_in_1_2;
      end else if (8'h9e == _T_19[7:0]) begin
        image_1_158 <= io_pixelVal_in_1_1;
      end else if (8'h9e == _T_15[7:0]) begin
        image_1_158 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_159 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9f == _T_34[7:0]) begin
        image_1_159 <= io_pixelVal_in_1_6;
      end else if (8'h9f == _T_31[7:0]) begin
        image_1_159 <= io_pixelVal_in_1_5;
      end else if (8'h9f == _T_28[7:0]) begin
        image_1_159 <= io_pixelVal_in_1_4;
      end else if (8'h9f == _T_25[7:0]) begin
        image_1_159 <= io_pixelVal_in_1_3;
      end else if (8'h9f == _T_22[7:0]) begin
        image_1_159 <= io_pixelVal_in_1_2;
      end else if (8'h9f == _T_19[7:0]) begin
        image_1_159 <= io_pixelVal_in_1_1;
      end else if (8'h9f == _T_15[7:0]) begin
        image_1_159 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_160 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha0 == _T_34[7:0]) begin
        image_1_160 <= io_pixelVal_in_1_6;
      end else if (8'ha0 == _T_31[7:0]) begin
        image_1_160 <= io_pixelVal_in_1_5;
      end else if (8'ha0 == _T_28[7:0]) begin
        image_1_160 <= io_pixelVal_in_1_4;
      end else if (8'ha0 == _T_25[7:0]) begin
        image_1_160 <= io_pixelVal_in_1_3;
      end else if (8'ha0 == _T_22[7:0]) begin
        image_1_160 <= io_pixelVal_in_1_2;
      end else if (8'ha0 == _T_19[7:0]) begin
        image_1_160 <= io_pixelVal_in_1_1;
      end else if (8'ha0 == _T_15[7:0]) begin
        image_1_160 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_161 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha1 == _T_34[7:0]) begin
        image_1_161 <= io_pixelVal_in_1_6;
      end else if (8'ha1 == _T_31[7:0]) begin
        image_1_161 <= io_pixelVal_in_1_5;
      end else if (8'ha1 == _T_28[7:0]) begin
        image_1_161 <= io_pixelVal_in_1_4;
      end else if (8'ha1 == _T_25[7:0]) begin
        image_1_161 <= io_pixelVal_in_1_3;
      end else if (8'ha1 == _T_22[7:0]) begin
        image_1_161 <= io_pixelVal_in_1_2;
      end else if (8'ha1 == _T_19[7:0]) begin
        image_1_161 <= io_pixelVal_in_1_1;
      end else if (8'ha1 == _T_15[7:0]) begin
        image_1_161 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_162 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha2 == _T_34[7:0]) begin
        image_1_162 <= io_pixelVal_in_1_6;
      end else if (8'ha2 == _T_31[7:0]) begin
        image_1_162 <= io_pixelVal_in_1_5;
      end else if (8'ha2 == _T_28[7:0]) begin
        image_1_162 <= io_pixelVal_in_1_4;
      end else if (8'ha2 == _T_25[7:0]) begin
        image_1_162 <= io_pixelVal_in_1_3;
      end else if (8'ha2 == _T_22[7:0]) begin
        image_1_162 <= io_pixelVal_in_1_2;
      end else if (8'ha2 == _T_19[7:0]) begin
        image_1_162 <= io_pixelVal_in_1_1;
      end else if (8'ha2 == _T_15[7:0]) begin
        image_1_162 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_163 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha3 == _T_34[7:0]) begin
        image_1_163 <= io_pixelVal_in_1_6;
      end else if (8'ha3 == _T_31[7:0]) begin
        image_1_163 <= io_pixelVal_in_1_5;
      end else if (8'ha3 == _T_28[7:0]) begin
        image_1_163 <= io_pixelVal_in_1_4;
      end else if (8'ha3 == _T_25[7:0]) begin
        image_1_163 <= io_pixelVal_in_1_3;
      end else if (8'ha3 == _T_22[7:0]) begin
        image_1_163 <= io_pixelVal_in_1_2;
      end else if (8'ha3 == _T_19[7:0]) begin
        image_1_163 <= io_pixelVal_in_1_1;
      end else if (8'ha3 == _T_15[7:0]) begin
        image_1_163 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_164 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha4 == _T_34[7:0]) begin
        image_1_164 <= io_pixelVal_in_1_6;
      end else if (8'ha4 == _T_31[7:0]) begin
        image_1_164 <= io_pixelVal_in_1_5;
      end else if (8'ha4 == _T_28[7:0]) begin
        image_1_164 <= io_pixelVal_in_1_4;
      end else if (8'ha4 == _T_25[7:0]) begin
        image_1_164 <= io_pixelVal_in_1_3;
      end else if (8'ha4 == _T_22[7:0]) begin
        image_1_164 <= io_pixelVal_in_1_2;
      end else if (8'ha4 == _T_19[7:0]) begin
        image_1_164 <= io_pixelVal_in_1_1;
      end else if (8'ha4 == _T_15[7:0]) begin
        image_1_164 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_165 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha5 == _T_34[7:0]) begin
        image_1_165 <= io_pixelVal_in_1_6;
      end else if (8'ha5 == _T_31[7:0]) begin
        image_1_165 <= io_pixelVal_in_1_5;
      end else if (8'ha5 == _T_28[7:0]) begin
        image_1_165 <= io_pixelVal_in_1_4;
      end else if (8'ha5 == _T_25[7:0]) begin
        image_1_165 <= io_pixelVal_in_1_3;
      end else if (8'ha5 == _T_22[7:0]) begin
        image_1_165 <= io_pixelVal_in_1_2;
      end else if (8'ha5 == _T_19[7:0]) begin
        image_1_165 <= io_pixelVal_in_1_1;
      end else if (8'ha5 == _T_15[7:0]) begin
        image_1_165 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_166 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha6 == _T_34[7:0]) begin
        image_1_166 <= io_pixelVal_in_1_6;
      end else if (8'ha6 == _T_31[7:0]) begin
        image_1_166 <= io_pixelVal_in_1_5;
      end else if (8'ha6 == _T_28[7:0]) begin
        image_1_166 <= io_pixelVal_in_1_4;
      end else if (8'ha6 == _T_25[7:0]) begin
        image_1_166 <= io_pixelVal_in_1_3;
      end else if (8'ha6 == _T_22[7:0]) begin
        image_1_166 <= io_pixelVal_in_1_2;
      end else if (8'ha6 == _T_19[7:0]) begin
        image_1_166 <= io_pixelVal_in_1_1;
      end else if (8'ha6 == _T_15[7:0]) begin
        image_1_166 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_167 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha7 == _T_34[7:0]) begin
        image_1_167 <= io_pixelVal_in_1_6;
      end else if (8'ha7 == _T_31[7:0]) begin
        image_1_167 <= io_pixelVal_in_1_5;
      end else if (8'ha7 == _T_28[7:0]) begin
        image_1_167 <= io_pixelVal_in_1_4;
      end else if (8'ha7 == _T_25[7:0]) begin
        image_1_167 <= io_pixelVal_in_1_3;
      end else if (8'ha7 == _T_22[7:0]) begin
        image_1_167 <= io_pixelVal_in_1_2;
      end else if (8'ha7 == _T_19[7:0]) begin
        image_1_167 <= io_pixelVal_in_1_1;
      end else if (8'ha7 == _T_15[7:0]) begin
        image_1_167 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_168 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha8 == _T_34[7:0]) begin
        image_1_168 <= io_pixelVal_in_1_6;
      end else if (8'ha8 == _T_31[7:0]) begin
        image_1_168 <= io_pixelVal_in_1_5;
      end else if (8'ha8 == _T_28[7:0]) begin
        image_1_168 <= io_pixelVal_in_1_4;
      end else if (8'ha8 == _T_25[7:0]) begin
        image_1_168 <= io_pixelVal_in_1_3;
      end else if (8'ha8 == _T_22[7:0]) begin
        image_1_168 <= io_pixelVal_in_1_2;
      end else if (8'ha8 == _T_19[7:0]) begin
        image_1_168 <= io_pixelVal_in_1_1;
      end else if (8'ha8 == _T_15[7:0]) begin
        image_1_168 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_169 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha9 == _T_34[7:0]) begin
        image_1_169 <= io_pixelVal_in_1_6;
      end else if (8'ha9 == _T_31[7:0]) begin
        image_1_169 <= io_pixelVal_in_1_5;
      end else if (8'ha9 == _T_28[7:0]) begin
        image_1_169 <= io_pixelVal_in_1_4;
      end else if (8'ha9 == _T_25[7:0]) begin
        image_1_169 <= io_pixelVal_in_1_3;
      end else if (8'ha9 == _T_22[7:0]) begin
        image_1_169 <= io_pixelVal_in_1_2;
      end else if (8'ha9 == _T_19[7:0]) begin
        image_1_169 <= io_pixelVal_in_1_1;
      end else if (8'ha9 == _T_15[7:0]) begin
        image_1_169 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_170 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'haa == _T_34[7:0]) begin
        image_1_170 <= io_pixelVal_in_1_6;
      end else if (8'haa == _T_31[7:0]) begin
        image_1_170 <= io_pixelVal_in_1_5;
      end else if (8'haa == _T_28[7:0]) begin
        image_1_170 <= io_pixelVal_in_1_4;
      end else if (8'haa == _T_25[7:0]) begin
        image_1_170 <= io_pixelVal_in_1_3;
      end else if (8'haa == _T_22[7:0]) begin
        image_1_170 <= io_pixelVal_in_1_2;
      end else if (8'haa == _T_19[7:0]) begin
        image_1_170 <= io_pixelVal_in_1_1;
      end else if (8'haa == _T_15[7:0]) begin
        image_1_170 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_171 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hab == _T_34[7:0]) begin
        image_1_171 <= io_pixelVal_in_1_6;
      end else if (8'hab == _T_31[7:0]) begin
        image_1_171 <= io_pixelVal_in_1_5;
      end else if (8'hab == _T_28[7:0]) begin
        image_1_171 <= io_pixelVal_in_1_4;
      end else if (8'hab == _T_25[7:0]) begin
        image_1_171 <= io_pixelVal_in_1_3;
      end else if (8'hab == _T_22[7:0]) begin
        image_1_171 <= io_pixelVal_in_1_2;
      end else if (8'hab == _T_19[7:0]) begin
        image_1_171 <= io_pixelVal_in_1_1;
      end else if (8'hab == _T_15[7:0]) begin
        image_1_171 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_172 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hac == _T_34[7:0]) begin
        image_1_172 <= io_pixelVal_in_1_6;
      end else if (8'hac == _T_31[7:0]) begin
        image_1_172 <= io_pixelVal_in_1_5;
      end else if (8'hac == _T_28[7:0]) begin
        image_1_172 <= io_pixelVal_in_1_4;
      end else if (8'hac == _T_25[7:0]) begin
        image_1_172 <= io_pixelVal_in_1_3;
      end else if (8'hac == _T_22[7:0]) begin
        image_1_172 <= io_pixelVal_in_1_2;
      end else if (8'hac == _T_19[7:0]) begin
        image_1_172 <= io_pixelVal_in_1_1;
      end else if (8'hac == _T_15[7:0]) begin
        image_1_172 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_173 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'had == _T_34[7:0]) begin
        image_1_173 <= io_pixelVal_in_1_6;
      end else if (8'had == _T_31[7:0]) begin
        image_1_173 <= io_pixelVal_in_1_5;
      end else if (8'had == _T_28[7:0]) begin
        image_1_173 <= io_pixelVal_in_1_4;
      end else if (8'had == _T_25[7:0]) begin
        image_1_173 <= io_pixelVal_in_1_3;
      end else if (8'had == _T_22[7:0]) begin
        image_1_173 <= io_pixelVal_in_1_2;
      end else if (8'had == _T_19[7:0]) begin
        image_1_173 <= io_pixelVal_in_1_1;
      end else if (8'had == _T_15[7:0]) begin
        image_1_173 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_174 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hae == _T_34[7:0]) begin
        image_1_174 <= io_pixelVal_in_1_6;
      end else if (8'hae == _T_31[7:0]) begin
        image_1_174 <= io_pixelVal_in_1_5;
      end else if (8'hae == _T_28[7:0]) begin
        image_1_174 <= io_pixelVal_in_1_4;
      end else if (8'hae == _T_25[7:0]) begin
        image_1_174 <= io_pixelVal_in_1_3;
      end else if (8'hae == _T_22[7:0]) begin
        image_1_174 <= io_pixelVal_in_1_2;
      end else if (8'hae == _T_19[7:0]) begin
        image_1_174 <= io_pixelVal_in_1_1;
      end else if (8'hae == _T_15[7:0]) begin
        image_1_174 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_175 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'haf == _T_34[7:0]) begin
        image_1_175 <= io_pixelVal_in_1_6;
      end else if (8'haf == _T_31[7:0]) begin
        image_1_175 <= io_pixelVal_in_1_5;
      end else if (8'haf == _T_28[7:0]) begin
        image_1_175 <= io_pixelVal_in_1_4;
      end else if (8'haf == _T_25[7:0]) begin
        image_1_175 <= io_pixelVal_in_1_3;
      end else if (8'haf == _T_22[7:0]) begin
        image_1_175 <= io_pixelVal_in_1_2;
      end else if (8'haf == _T_19[7:0]) begin
        image_1_175 <= io_pixelVal_in_1_1;
      end else if (8'haf == _T_15[7:0]) begin
        image_1_175 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_176 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb0 == _T_34[7:0]) begin
        image_1_176 <= io_pixelVal_in_1_6;
      end else if (8'hb0 == _T_31[7:0]) begin
        image_1_176 <= io_pixelVal_in_1_5;
      end else if (8'hb0 == _T_28[7:0]) begin
        image_1_176 <= io_pixelVal_in_1_4;
      end else if (8'hb0 == _T_25[7:0]) begin
        image_1_176 <= io_pixelVal_in_1_3;
      end else if (8'hb0 == _T_22[7:0]) begin
        image_1_176 <= io_pixelVal_in_1_2;
      end else if (8'hb0 == _T_19[7:0]) begin
        image_1_176 <= io_pixelVal_in_1_1;
      end else if (8'hb0 == _T_15[7:0]) begin
        image_1_176 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_177 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb1 == _T_34[7:0]) begin
        image_1_177 <= io_pixelVal_in_1_6;
      end else if (8'hb1 == _T_31[7:0]) begin
        image_1_177 <= io_pixelVal_in_1_5;
      end else if (8'hb1 == _T_28[7:0]) begin
        image_1_177 <= io_pixelVal_in_1_4;
      end else if (8'hb1 == _T_25[7:0]) begin
        image_1_177 <= io_pixelVal_in_1_3;
      end else if (8'hb1 == _T_22[7:0]) begin
        image_1_177 <= io_pixelVal_in_1_2;
      end else if (8'hb1 == _T_19[7:0]) begin
        image_1_177 <= io_pixelVal_in_1_1;
      end else if (8'hb1 == _T_15[7:0]) begin
        image_1_177 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_178 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb2 == _T_34[7:0]) begin
        image_1_178 <= io_pixelVal_in_1_6;
      end else if (8'hb2 == _T_31[7:0]) begin
        image_1_178 <= io_pixelVal_in_1_5;
      end else if (8'hb2 == _T_28[7:0]) begin
        image_1_178 <= io_pixelVal_in_1_4;
      end else if (8'hb2 == _T_25[7:0]) begin
        image_1_178 <= io_pixelVal_in_1_3;
      end else if (8'hb2 == _T_22[7:0]) begin
        image_1_178 <= io_pixelVal_in_1_2;
      end else if (8'hb2 == _T_19[7:0]) begin
        image_1_178 <= io_pixelVal_in_1_1;
      end else if (8'hb2 == _T_15[7:0]) begin
        image_1_178 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_179 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb3 == _T_34[7:0]) begin
        image_1_179 <= io_pixelVal_in_1_6;
      end else if (8'hb3 == _T_31[7:0]) begin
        image_1_179 <= io_pixelVal_in_1_5;
      end else if (8'hb3 == _T_28[7:0]) begin
        image_1_179 <= io_pixelVal_in_1_4;
      end else if (8'hb3 == _T_25[7:0]) begin
        image_1_179 <= io_pixelVal_in_1_3;
      end else if (8'hb3 == _T_22[7:0]) begin
        image_1_179 <= io_pixelVal_in_1_2;
      end else if (8'hb3 == _T_19[7:0]) begin
        image_1_179 <= io_pixelVal_in_1_1;
      end else if (8'hb3 == _T_15[7:0]) begin
        image_1_179 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_180 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb4 == _T_34[7:0]) begin
        image_1_180 <= io_pixelVal_in_1_6;
      end else if (8'hb4 == _T_31[7:0]) begin
        image_1_180 <= io_pixelVal_in_1_5;
      end else if (8'hb4 == _T_28[7:0]) begin
        image_1_180 <= io_pixelVal_in_1_4;
      end else if (8'hb4 == _T_25[7:0]) begin
        image_1_180 <= io_pixelVal_in_1_3;
      end else if (8'hb4 == _T_22[7:0]) begin
        image_1_180 <= io_pixelVal_in_1_2;
      end else if (8'hb4 == _T_19[7:0]) begin
        image_1_180 <= io_pixelVal_in_1_1;
      end else if (8'hb4 == _T_15[7:0]) begin
        image_1_180 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_181 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb5 == _T_34[7:0]) begin
        image_1_181 <= io_pixelVal_in_1_6;
      end else if (8'hb5 == _T_31[7:0]) begin
        image_1_181 <= io_pixelVal_in_1_5;
      end else if (8'hb5 == _T_28[7:0]) begin
        image_1_181 <= io_pixelVal_in_1_4;
      end else if (8'hb5 == _T_25[7:0]) begin
        image_1_181 <= io_pixelVal_in_1_3;
      end else if (8'hb5 == _T_22[7:0]) begin
        image_1_181 <= io_pixelVal_in_1_2;
      end else if (8'hb5 == _T_19[7:0]) begin
        image_1_181 <= io_pixelVal_in_1_1;
      end else if (8'hb5 == _T_15[7:0]) begin
        image_1_181 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_182 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb6 == _T_34[7:0]) begin
        image_1_182 <= io_pixelVal_in_1_6;
      end else if (8'hb6 == _T_31[7:0]) begin
        image_1_182 <= io_pixelVal_in_1_5;
      end else if (8'hb6 == _T_28[7:0]) begin
        image_1_182 <= io_pixelVal_in_1_4;
      end else if (8'hb6 == _T_25[7:0]) begin
        image_1_182 <= io_pixelVal_in_1_3;
      end else if (8'hb6 == _T_22[7:0]) begin
        image_1_182 <= io_pixelVal_in_1_2;
      end else if (8'hb6 == _T_19[7:0]) begin
        image_1_182 <= io_pixelVal_in_1_1;
      end else if (8'hb6 == _T_15[7:0]) begin
        image_1_182 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_183 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb7 == _T_34[7:0]) begin
        image_1_183 <= io_pixelVal_in_1_6;
      end else if (8'hb7 == _T_31[7:0]) begin
        image_1_183 <= io_pixelVal_in_1_5;
      end else if (8'hb7 == _T_28[7:0]) begin
        image_1_183 <= io_pixelVal_in_1_4;
      end else if (8'hb7 == _T_25[7:0]) begin
        image_1_183 <= io_pixelVal_in_1_3;
      end else if (8'hb7 == _T_22[7:0]) begin
        image_1_183 <= io_pixelVal_in_1_2;
      end else if (8'hb7 == _T_19[7:0]) begin
        image_1_183 <= io_pixelVal_in_1_1;
      end else if (8'hb7 == _T_15[7:0]) begin
        image_1_183 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_184 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb8 == _T_34[7:0]) begin
        image_1_184 <= io_pixelVal_in_1_6;
      end else if (8'hb8 == _T_31[7:0]) begin
        image_1_184 <= io_pixelVal_in_1_5;
      end else if (8'hb8 == _T_28[7:0]) begin
        image_1_184 <= io_pixelVal_in_1_4;
      end else if (8'hb8 == _T_25[7:0]) begin
        image_1_184 <= io_pixelVal_in_1_3;
      end else if (8'hb8 == _T_22[7:0]) begin
        image_1_184 <= io_pixelVal_in_1_2;
      end else if (8'hb8 == _T_19[7:0]) begin
        image_1_184 <= io_pixelVal_in_1_1;
      end else if (8'hb8 == _T_15[7:0]) begin
        image_1_184 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_185 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb9 == _T_34[7:0]) begin
        image_1_185 <= io_pixelVal_in_1_6;
      end else if (8'hb9 == _T_31[7:0]) begin
        image_1_185 <= io_pixelVal_in_1_5;
      end else if (8'hb9 == _T_28[7:0]) begin
        image_1_185 <= io_pixelVal_in_1_4;
      end else if (8'hb9 == _T_25[7:0]) begin
        image_1_185 <= io_pixelVal_in_1_3;
      end else if (8'hb9 == _T_22[7:0]) begin
        image_1_185 <= io_pixelVal_in_1_2;
      end else if (8'hb9 == _T_19[7:0]) begin
        image_1_185 <= io_pixelVal_in_1_1;
      end else if (8'hb9 == _T_15[7:0]) begin
        image_1_185 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_186 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hba == _T_34[7:0]) begin
        image_1_186 <= io_pixelVal_in_1_6;
      end else if (8'hba == _T_31[7:0]) begin
        image_1_186 <= io_pixelVal_in_1_5;
      end else if (8'hba == _T_28[7:0]) begin
        image_1_186 <= io_pixelVal_in_1_4;
      end else if (8'hba == _T_25[7:0]) begin
        image_1_186 <= io_pixelVal_in_1_3;
      end else if (8'hba == _T_22[7:0]) begin
        image_1_186 <= io_pixelVal_in_1_2;
      end else if (8'hba == _T_19[7:0]) begin
        image_1_186 <= io_pixelVal_in_1_1;
      end else if (8'hba == _T_15[7:0]) begin
        image_1_186 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_187 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbb == _T_34[7:0]) begin
        image_1_187 <= io_pixelVal_in_1_6;
      end else if (8'hbb == _T_31[7:0]) begin
        image_1_187 <= io_pixelVal_in_1_5;
      end else if (8'hbb == _T_28[7:0]) begin
        image_1_187 <= io_pixelVal_in_1_4;
      end else if (8'hbb == _T_25[7:0]) begin
        image_1_187 <= io_pixelVal_in_1_3;
      end else if (8'hbb == _T_22[7:0]) begin
        image_1_187 <= io_pixelVal_in_1_2;
      end else if (8'hbb == _T_19[7:0]) begin
        image_1_187 <= io_pixelVal_in_1_1;
      end else if (8'hbb == _T_15[7:0]) begin
        image_1_187 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_188 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbc == _T_34[7:0]) begin
        image_1_188 <= io_pixelVal_in_1_6;
      end else if (8'hbc == _T_31[7:0]) begin
        image_1_188 <= io_pixelVal_in_1_5;
      end else if (8'hbc == _T_28[7:0]) begin
        image_1_188 <= io_pixelVal_in_1_4;
      end else if (8'hbc == _T_25[7:0]) begin
        image_1_188 <= io_pixelVal_in_1_3;
      end else if (8'hbc == _T_22[7:0]) begin
        image_1_188 <= io_pixelVal_in_1_2;
      end else if (8'hbc == _T_19[7:0]) begin
        image_1_188 <= io_pixelVal_in_1_1;
      end else if (8'hbc == _T_15[7:0]) begin
        image_1_188 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_189 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbd == _T_34[7:0]) begin
        image_1_189 <= io_pixelVal_in_1_6;
      end else if (8'hbd == _T_31[7:0]) begin
        image_1_189 <= io_pixelVal_in_1_5;
      end else if (8'hbd == _T_28[7:0]) begin
        image_1_189 <= io_pixelVal_in_1_4;
      end else if (8'hbd == _T_25[7:0]) begin
        image_1_189 <= io_pixelVal_in_1_3;
      end else if (8'hbd == _T_22[7:0]) begin
        image_1_189 <= io_pixelVal_in_1_2;
      end else if (8'hbd == _T_19[7:0]) begin
        image_1_189 <= io_pixelVal_in_1_1;
      end else if (8'hbd == _T_15[7:0]) begin
        image_1_189 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_190 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbe == _T_34[7:0]) begin
        image_1_190 <= io_pixelVal_in_1_6;
      end else if (8'hbe == _T_31[7:0]) begin
        image_1_190 <= io_pixelVal_in_1_5;
      end else if (8'hbe == _T_28[7:0]) begin
        image_1_190 <= io_pixelVal_in_1_4;
      end else if (8'hbe == _T_25[7:0]) begin
        image_1_190 <= io_pixelVal_in_1_3;
      end else if (8'hbe == _T_22[7:0]) begin
        image_1_190 <= io_pixelVal_in_1_2;
      end else if (8'hbe == _T_19[7:0]) begin
        image_1_190 <= io_pixelVal_in_1_1;
      end else if (8'hbe == _T_15[7:0]) begin
        image_1_190 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_191 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbf == _T_34[7:0]) begin
        image_1_191 <= io_pixelVal_in_1_6;
      end else if (8'hbf == _T_31[7:0]) begin
        image_1_191 <= io_pixelVal_in_1_5;
      end else if (8'hbf == _T_28[7:0]) begin
        image_1_191 <= io_pixelVal_in_1_4;
      end else if (8'hbf == _T_25[7:0]) begin
        image_1_191 <= io_pixelVal_in_1_3;
      end else if (8'hbf == _T_22[7:0]) begin
        image_1_191 <= io_pixelVal_in_1_2;
      end else if (8'hbf == _T_19[7:0]) begin
        image_1_191 <= io_pixelVal_in_1_1;
      end else if (8'hbf == _T_15[7:0]) begin
        image_1_191 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_192 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc0 == _T_34[7:0]) begin
        image_1_192 <= io_pixelVal_in_1_6;
      end else if (8'hc0 == _T_31[7:0]) begin
        image_1_192 <= io_pixelVal_in_1_5;
      end else if (8'hc0 == _T_28[7:0]) begin
        image_1_192 <= io_pixelVal_in_1_4;
      end else if (8'hc0 == _T_25[7:0]) begin
        image_1_192 <= io_pixelVal_in_1_3;
      end else if (8'hc0 == _T_22[7:0]) begin
        image_1_192 <= io_pixelVal_in_1_2;
      end else if (8'hc0 == _T_19[7:0]) begin
        image_1_192 <= io_pixelVal_in_1_1;
      end else if (8'hc0 == _T_15[7:0]) begin
        image_1_192 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_193 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc1 == _T_34[7:0]) begin
        image_1_193 <= io_pixelVal_in_1_6;
      end else if (8'hc1 == _T_31[7:0]) begin
        image_1_193 <= io_pixelVal_in_1_5;
      end else if (8'hc1 == _T_28[7:0]) begin
        image_1_193 <= io_pixelVal_in_1_4;
      end else if (8'hc1 == _T_25[7:0]) begin
        image_1_193 <= io_pixelVal_in_1_3;
      end else if (8'hc1 == _T_22[7:0]) begin
        image_1_193 <= io_pixelVal_in_1_2;
      end else if (8'hc1 == _T_19[7:0]) begin
        image_1_193 <= io_pixelVal_in_1_1;
      end else if (8'hc1 == _T_15[7:0]) begin
        image_1_193 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_194 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc2 == _T_34[7:0]) begin
        image_1_194 <= io_pixelVal_in_1_6;
      end else if (8'hc2 == _T_31[7:0]) begin
        image_1_194 <= io_pixelVal_in_1_5;
      end else if (8'hc2 == _T_28[7:0]) begin
        image_1_194 <= io_pixelVal_in_1_4;
      end else if (8'hc2 == _T_25[7:0]) begin
        image_1_194 <= io_pixelVal_in_1_3;
      end else if (8'hc2 == _T_22[7:0]) begin
        image_1_194 <= io_pixelVal_in_1_2;
      end else if (8'hc2 == _T_19[7:0]) begin
        image_1_194 <= io_pixelVal_in_1_1;
      end else if (8'hc2 == _T_15[7:0]) begin
        image_1_194 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_195 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc3 == _T_34[7:0]) begin
        image_1_195 <= io_pixelVal_in_1_6;
      end else if (8'hc3 == _T_31[7:0]) begin
        image_1_195 <= io_pixelVal_in_1_5;
      end else if (8'hc3 == _T_28[7:0]) begin
        image_1_195 <= io_pixelVal_in_1_4;
      end else if (8'hc3 == _T_25[7:0]) begin
        image_1_195 <= io_pixelVal_in_1_3;
      end else if (8'hc3 == _T_22[7:0]) begin
        image_1_195 <= io_pixelVal_in_1_2;
      end else if (8'hc3 == _T_19[7:0]) begin
        image_1_195 <= io_pixelVal_in_1_1;
      end else if (8'hc3 == _T_15[7:0]) begin
        image_1_195 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_196 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc4 == _T_34[7:0]) begin
        image_1_196 <= io_pixelVal_in_1_6;
      end else if (8'hc4 == _T_31[7:0]) begin
        image_1_196 <= io_pixelVal_in_1_5;
      end else if (8'hc4 == _T_28[7:0]) begin
        image_1_196 <= io_pixelVal_in_1_4;
      end else if (8'hc4 == _T_25[7:0]) begin
        image_1_196 <= io_pixelVal_in_1_3;
      end else if (8'hc4 == _T_22[7:0]) begin
        image_1_196 <= io_pixelVal_in_1_2;
      end else if (8'hc4 == _T_19[7:0]) begin
        image_1_196 <= io_pixelVal_in_1_1;
      end else if (8'hc4 == _T_15[7:0]) begin
        image_1_196 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_197 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc5 == _T_34[7:0]) begin
        image_1_197 <= io_pixelVal_in_1_6;
      end else if (8'hc5 == _T_31[7:0]) begin
        image_1_197 <= io_pixelVal_in_1_5;
      end else if (8'hc5 == _T_28[7:0]) begin
        image_1_197 <= io_pixelVal_in_1_4;
      end else if (8'hc5 == _T_25[7:0]) begin
        image_1_197 <= io_pixelVal_in_1_3;
      end else if (8'hc5 == _T_22[7:0]) begin
        image_1_197 <= io_pixelVal_in_1_2;
      end else if (8'hc5 == _T_19[7:0]) begin
        image_1_197 <= io_pixelVal_in_1_1;
      end else if (8'hc5 == _T_15[7:0]) begin
        image_1_197 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_198 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc6 == _T_34[7:0]) begin
        image_1_198 <= io_pixelVal_in_1_6;
      end else if (8'hc6 == _T_31[7:0]) begin
        image_1_198 <= io_pixelVal_in_1_5;
      end else if (8'hc6 == _T_28[7:0]) begin
        image_1_198 <= io_pixelVal_in_1_4;
      end else if (8'hc6 == _T_25[7:0]) begin
        image_1_198 <= io_pixelVal_in_1_3;
      end else if (8'hc6 == _T_22[7:0]) begin
        image_1_198 <= io_pixelVal_in_1_2;
      end else if (8'hc6 == _T_19[7:0]) begin
        image_1_198 <= io_pixelVal_in_1_1;
      end else if (8'hc6 == _T_15[7:0]) begin
        image_1_198 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_199 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc7 == _T_34[7:0]) begin
        image_1_199 <= io_pixelVal_in_1_6;
      end else if (8'hc7 == _T_31[7:0]) begin
        image_1_199 <= io_pixelVal_in_1_5;
      end else if (8'hc7 == _T_28[7:0]) begin
        image_1_199 <= io_pixelVal_in_1_4;
      end else if (8'hc7 == _T_25[7:0]) begin
        image_1_199 <= io_pixelVal_in_1_3;
      end else if (8'hc7 == _T_22[7:0]) begin
        image_1_199 <= io_pixelVal_in_1_2;
      end else if (8'hc7 == _T_19[7:0]) begin
        image_1_199 <= io_pixelVal_in_1_1;
      end else if (8'hc7 == _T_15[7:0]) begin
        image_1_199 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_200 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc8 == _T_34[7:0]) begin
        image_1_200 <= io_pixelVal_in_1_6;
      end else if (8'hc8 == _T_31[7:0]) begin
        image_1_200 <= io_pixelVal_in_1_5;
      end else if (8'hc8 == _T_28[7:0]) begin
        image_1_200 <= io_pixelVal_in_1_4;
      end else if (8'hc8 == _T_25[7:0]) begin
        image_1_200 <= io_pixelVal_in_1_3;
      end else if (8'hc8 == _T_22[7:0]) begin
        image_1_200 <= io_pixelVal_in_1_2;
      end else if (8'hc8 == _T_19[7:0]) begin
        image_1_200 <= io_pixelVal_in_1_1;
      end else if (8'hc8 == _T_15[7:0]) begin
        image_1_200 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_201 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc9 == _T_34[7:0]) begin
        image_1_201 <= io_pixelVal_in_1_6;
      end else if (8'hc9 == _T_31[7:0]) begin
        image_1_201 <= io_pixelVal_in_1_5;
      end else if (8'hc9 == _T_28[7:0]) begin
        image_1_201 <= io_pixelVal_in_1_4;
      end else if (8'hc9 == _T_25[7:0]) begin
        image_1_201 <= io_pixelVal_in_1_3;
      end else if (8'hc9 == _T_22[7:0]) begin
        image_1_201 <= io_pixelVal_in_1_2;
      end else if (8'hc9 == _T_19[7:0]) begin
        image_1_201 <= io_pixelVal_in_1_1;
      end else if (8'hc9 == _T_15[7:0]) begin
        image_1_201 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_202 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hca == _T_34[7:0]) begin
        image_1_202 <= io_pixelVal_in_1_6;
      end else if (8'hca == _T_31[7:0]) begin
        image_1_202 <= io_pixelVal_in_1_5;
      end else if (8'hca == _T_28[7:0]) begin
        image_1_202 <= io_pixelVal_in_1_4;
      end else if (8'hca == _T_25[7:0]) begin
        image_1_202 <= io_pixelVal_in_1_3;
      end else if (8'hca == _T_22[7:0]) begin
        image_1_202 <= io_pixelVal_in_1_2;
      end else if (8'hca == _T_19[7:0]) begin
        image_1_202 <= io_pixelVal_in_1_1;
      end else if (8'hca == _T_15[7:0]) begin
        image_1_202 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_203 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hcb == _T_34[7:0]) begin
        image_1_203 <= io_pixelVal_in_1_6;
      end else if (8'hcb == _T_31[7:0]) begin
        image_1_203 <= io_pixelVal_in_1_5;
      end else if (8'hcb == _T_28[7:0]) begin
        image_1_203 <= io_pixelVal_in_1_4;
      end else if (8'hcb == _T_25[7:0]) begin
        image_1_203 <= io_pixelVal_in_1_3;
      end else if (8'hcb == _T_22[7:0]) begin
        image_1_203 <= io_pixelVal_in_1_2;
      end else if (8'hcb == _T_19[7:0]) begin
        image_1_203 <= io_pixelVal_in_1_1;
      end else if (8'hcb == _T_15[7:0]) begin
        image_1_203 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_204 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hcc == _T_34[7:0]) begin
        image_1_204 <= io_pixelVal_in_1_6;
      end else if (8'hcc == _T_31[7:0]) begin
        image_1_204 <= io_pixelVal_in_1_5;
      end else if (8'hcc == _T_28[7:0]) begin
        image_1_204 <= io_pixelVal_in_1_4;
      end else if (8'hcc == _T_25[7:0]) begin
        image_1_204 <= io_pixelVal_in_1_3;
      end else if (8'hcc == _T_22[7:0]) begin
        image_1_204 <= io_pixelVal_in_1_2;
      end else if (8'hcc == _T_19[7:0]) begin
        image_1_204 <= io_pixelVal_in_1_1;
      end else if (8'hcc == _T_15[7:0]) begin
        image_1_204 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_205 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hcd == _T_34[7:0]) begin
        image_1_205 <= io_pixelVal_in_1_6;
      end else if (8'hcd == _T_31[7:0]) begin
        image_1_205 <= io_pixelVal_in_1_5;
      end else if (8'hcd == _T_28[7:0]) begin
        image_1_205 <= io_pixelVal_in_1_4;
      end else if (8'hcd == _T_25[7:0]) begin
        image_1_205 <= io_pixelVal_in_1_3;
      end else if (8'hcd == _T_22[7:0]) begin
        image_1_205 <= io_pixelVal_in_1_2;
      end else if (8'hcd == _T_19[7:0]) begin
        image_1_205 <= io_pixelVal_in_1_1;
      end else if (8'hcd == _T_15[7:0]) begin
        image_1_205 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_206 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hce == _T_34[7:0]) begin
        image_1_206 <= io_pixelVal_in_1_6;
      end else if (8'hce == _T_31[7:0]) begin
        image_1_206 <= io_pixelVal_in_1_5;
      end else if (8'hce == _T_28[7:0]) begin
        image_1_206 <= io_pixelVal_in_1_4;
      end else if (8'hce == _T_25[7:0]) begin
        image_1_206 <= io_pixelVal_in_1_3;
      end else if (8'hce == _T_22[7:0]) begin
        image_1_206 <= io_pixelVal_in_1_2;
      end else if (8'hce == _T_19[7:0]) begin
        image_1_206 <= io_pixelVal_in_1_1;
      end else if (8'hce == _T_15[7:0]) begin
        image_1_206 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_207 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hcf == _T_34[7:0]) begin
        image_1_207 <= io_pixelVal_in_1_6;
      end else if (8'hcf == _T_31[7:0]) begin
        image_1_207 <= io_pixelVal_in_1_5;
      end else if (8'hcf == _T_28[7:0]) begin
        image_1_207 <= io_pixelVal_in_1_4;
      end else if (8'hcf == _T_25[7:0]) begin
        image_1_207 <= io_pixelVal_in_1_3;
      end else if (8'hcf == _T_22[7:0]) begin
        image_1_207 <= io_pixelVal_in_1_2;
      end else if (8'hcf == _T_19[7:0]) begin
        image_1_207 <= io_pixelVal_in_1_1;
      end else if (8'hcf == _T_15[7:0]) begin
        image_1_207 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_208 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd0 == _T_34[7:0]) begin
        image_1_208 <= io_pixelVal_in_1_6;
      end else if (8'hd0 == _T_31[7:0]) begin
        image_1_208 <= io_pixelVal_in_1_5;
      end else if (8'hd0 == _T_28[7:0]) begin
        image_1_208 <= io_pixelVal_in_1_4;
      end else if (8'hd0 == _T_25[7:0]) begin
        image_1_208 <= io_pixelVal_in_1_3;
      end else if (8'hd0 == _T_22[7:0]) begin
        image_1_208 <= io_pixelVal_in_1_2;
      end else if (8'hd0 == _T_19[7:0]) begin
        image_1_208 <= io_pixelVal_in_1_1;
      end else if (8'hd0 == _T_15[7:0]) begin
        image_1_208 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_209 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd1 == _T_34[7:0]) begin
        image_1_209 <= io_pixelVal_in_1_6;
      end else if (8'hd1 == _T_31[7:0]) begin
        image_1_209 <= io_pixelVal_in_1_5;
      end else if (8'hd1 == _T_28[7:0]) begin
        image_1_209 <= io_pixelVal_in_1_4;
      end else if (8'hd1 == _T_25[7:0]) begin
        image_1_209 <= io_pixelVal_in_1_3;
      end else if (8'hd1 == _T_22[7:0]) begin
        image_1_209 <= io_pixelVal_in_1_2;
      end else if (8'hd1 == _T_19[7:0]) begin
        image_1_209 <= io_pixelVal_in_1_1;
      end else if (8'hd1 == _T_15[7:0]) begin
        image_1_209 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_210 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd2 == _T_34[7:0]) begin
        image_1_210 <= io_pixelVal_in_1_6;
      end else if (8'hd2 == _T_31[7:0]) begin
        image_1_210 <= io_pixelVal_in_1_5;
      end else if (8'hd2 == _T_28[7:0]) begin
        image_1_210 <= io_pixelVal_in_1_4;
      end else if (8'hd2 == _T_25[7:0]) begin
        image_1_210 <= io_pixelVal_in_1_3;
      end else if (8'hd2 == _T_22[7:0]) begin
        image_1_210 <= io_pixelVal_in_1_2;
      end else if (8'hd2 == _T_19[7:0]) begin
        image_1_210 <= io_pixelVal_in_1_1;
      end else if (8'hd2 == _T_15[7:0]) begin
        image_1_210 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_211 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd3 == _T_34[7:0]) begin
        image_1_211 <= io_pixelVal_in_1_6;
      end else if (8'hd3 == _T_31[7:0]) begin
        image_1_211 <= io_pixelVal_in_1_5;
      end else if (8'hd3 == _T_28[7:0]) begin
        image_1_211 <= io_pixelVal_in_1_4;
      end else if (8'hd3 == _T_25[7:0]) begin
        image_1_211 <= io_pixelVal_in_1_3;
      end else if (8'hd3 == _T_22[7:0]) begin
        image_1_211 <= io_pixelVal_in_1_2;
      end else if (8'hd3 == _T_19[7:0]) begin
        image_1_211 <= io_pixelVal_in_1_1;
      end else if (8'hd3 == _T_15[7:0]) begin
        image_1_211 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_212 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd4 == _T_34[7:0]) begin
        image_1_212 <= io_pixelVal_in_1_6;
      end else if (8'hd4 == _T_31[7:0]) begin
        image_1_212 <= io_pixelVal_in_1_5;
      end else if (8'hd4 == _T_28[7:0]) begin
        image_1_212 <= io_pixelVal_in_1_4;
      end else if (8'hd4 == _T_25[7:0]) begin
        image_1_212 <= io_pixelVal_in_1_3;
      end else if (8'hd4 == _T_22[7:0]) begin
        image_1_212 <= io_pixelVal_in_1_2;
      end else if (8'hd4 == _T_19[7:0]) begin
        image_1_212 <= io_pixelVal_in_1_1;
      end else if (8'hd4 == _T_15[7:0]) begin
        image_1_212 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_213 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd5 == _T_34[7:0]) begin
        image_1_213 <= io_pixelVal_in_1_6;
      end else if (8'hd5 == _T_31[7:0]) begin
        image_1_213 <= io_pixelVal_in_1_5;
      end else if (8'hd5 == _T_28[7:0]) begin
        image_1_213 <= io_pixelVal_in_1_4;
      end else if (8'hd5 == _T_25[7:0]) begin
        image_1_213 <= io_pixelVal_in_1_3;
      end else if (8'hd5 == _T_22[7:0]) begin
        image_1_213 <= io_pixelVal_in_1_2;
      end else if (8'hd5 == _T_19[7:0]) begin
        image_1_213 <= io_pixelVal_in_1_1;
      end else if (8'hd5 == _T_15[7:0]) begin
        image_1_213 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_214 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd6 == _T_34[7:0]) begin
        image_1_214 <= io_pixelVal_in_1_6;
      end else if (8'hd6 == _T_31[7:0]) begin
        image_1_214 <= io_pixelVal_in_1_5;
      end else if (8'hd6 == _T_28[7:0]) begin
        image_1_214 <= io_pixelVal_in_1_4;
      end else if (8'hd6 == _T_25[7:0]) begin
        image_1_214 <= io_pixelVal_in_1_3;
      end else if (8'hd6 == _T_22[7:0]) begin
        image_1_214 <= io_pixelVal_in_1_2;
      end else if (8'hd6 == _T_19[7:0]) begin
        image_1_214 <= io_pixelVal_in_1_1;
      end else if (8'hd6 == _T_15[7:0]) begin
        image_1_214 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_215 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd7 == _T_34[7:0]) begin
        image_1_215 <= io_pixelVal_in_1_6;
      end else if (8'hd7 == _T_31[7:0]) begin
        image_1_215 <= io_pixelVal_in_1_5;
      end else if (8'hd7 == _T_28[7:0]) begin
        image_1_215 <= io_pixelVal_in_1_4;
      end else if (8'hd7 == _T_25[7:0]) begin
        image_1_215 <= io_pixelVal_in_1_3;
      end else if (8'hd7 == _T_22[7:0]) begin
        image_1_215 <= io_pixelVal_in_1_2;
      end else if (8'hd7 == _T_19[7:0]) begin
        image_1_215 <= io_pixelVal_in_1_1;
      end else if (8'hd7 == _T_15[7:0]) begin
        image_1_215 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_216 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd8 == _T_34[7:0]) begin
        image_1_216 <= io_pixelVal_in_1_6;
      end else if (8'hd8 == _T_31[7:0]) begin
        image_1_216 <= io_pixelVal_in_1_5;
      end else if (8'hd8 == _T_28[7:0]) begin
        image_1_216 <= io_pixelVal_in_1_4;
      end else if (8'hd8 == _T_25[7:0]) begin
        image_1_216 <= io_pixelVal_in_1_3;
      end else if (8'hd8 == _T_22[7:0]) begin
        image_1_216 <= io_pixelVal_in_1_2;
      end else if (8'hd8 == _T_19[7:0]) begin
        image_1_216 <= io_pixelVal_in_1_1;
      end else if (8'hd8 == _T_15[7:0]) begin
        image_1_216 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_217 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd9 == _T_34[7:0]) begin
        image_1_217 <= io_pixelVal_in_1_6;
      end else if (8'hd9 == _T_31[7:0]) begin
        image_1_217 <= io_pixelVal_in_1_5;
      end else if (8'hd9 == _T_28[7:0]) begin
        image_1_217 <= io_pixelVal_in_1_4;
      end else if (8'hd9 == _T_25[7:0]) begin
        image_1_217 <= io_pixelVal_in_1_3;
      end else if (8'hd9 == _T_22[7:0]) begin
        image_1_217 <= io_pixelVal_in_1_2;
      end else if (8'hd9 == _T_19[7:0]) begin
        image_1_217 <= io_pixelVal_in_1_1;
      end else if (8'hd9 == _T_15[7:0]) begin
        image_1_217 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_218 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hda == _T_34[7:0]) begin
        image_1_218 <= io_pixelVal_in_1_6;
      end else if (8'hda == _T_31[7:0]) begin
        image_1_218 <= io_pixelVal_in_1_5;
      end else if (8'hda == _T_28[7:0]) begin
        image_1_218 <= io_pixelVal_in_1_4;
      end else if (8'hda == _T_25[7:0]) begin
        image_1_218 <= io_pixelVal_in_1_3;
      end else if (8'hda == _T_22[7:0]) begin
        image_1_218 <= io_pixelVal_in_1_2;
      end else if (8'hda == _T_19[7:0]) begin
        image_1_218 <= io_pixelVal_in_1_1;
      end else if (8'hda == _T_15[7:0]) begin
        image_1_218 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_219 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hdb == _T_34[7:0]) begin
        image_1_219 <= io_pixelVal_in_1_6;
      end else if (8'hdb == _T_31[7:0]) begin
        image_1_219 <= io_pixelVal_in_1_5;
      end else if (8'hdb == _T_28[7:0]) begin
        image_1_219 <= io_pixelVal_in_1_4;
      end else if (8'hdb == _T_25[7:0]) begin
        image_1_219 <= io_pixelVal_in_1_3;
      end else if (8'hdb == _T_22[7:0]) begin
        image_1_219 <= io_pixelVal_in_1_2;
      end else if (8'hdb == _T_19[7:0]) begin
        image_1_219 <= io_pixelVal_in_1_1;
      end else if (8'hdb == _T_15[7:0]) begin
        image_1_219 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_220 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hdc == _T_34[7:0]) begin
        image_1_220 <= io_pixelVal_in_1_6;
      end else if (8'hdc == _T_31[7:0]) begin
        image_1_220 <= io_pixelVal_in_1_5;
      end else if (8'hdc == _T_28[7:0]) begin
        image_1_220 <= io_pixelVal_in_1_4;
      end else if (8'hdc == _T_25[7:0]) begin
        image_1_220 <= io_pixelVal_in_1_3;
      end else if (8'hdc == _T_22[7:0]) begin
        image_1_220 <= io_pixelVal_in_1_2;
      end else if (8'hdc == _T_19[7:0]) begin
        image_1_220 <= io_pixelVal_in_1_1;
      end else if (8'hdc == _T_15[7:0]) begin
        image_1_220 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_221 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hdd == _T_34[7:0]) begin
        image_1_221 <= io_pixelVal_in_1_6;
      end else if (8'hdd == _T_31[7:0]) begin
        image_1_221 <= io_pixelVal_in_1_5;
      end else if (8'hdd == _T_28[7:0]) begin
        image_1_221 <= io_pixelVal_in_1_4;
      end else if (8'hdd == _T_25[7:0]) begin
        image_1_221 <= io_pixelVal_in_1_3;
      end else if (8'hdd == _T_22[7:0]) begin
        image_1_221 <= io_pixelVal_in_1_2;
      end else if (8'hdd == _T_19[7:0]) begin
        image_1_221 <= io_pixelVal_in_1_1;
      end else if (8'hdd == _T_15[7:0]) begin
        image_1_221 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_222 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hde == _T_34[7:0]) begin
        image_1_222 <= io_pixelVal_in_1_6;
      end else if (8'hde == _T_31[7:0]) begin
        image_1_222 <= io_pixelVal_in_1_5;
      end else if (8'hde == _T_28[7:0]) begin
        image_1_222 <= io_pixelVal_in_1_4;
      end else if (8'hde == _T_25[7:0]) begin
        image_1_222 <= io_pixelVal_in_1_3;
      end else if (8'hde == _T_22[7:0]) begin
        image_1_222 <= io_pixelVal_in_1_2;
      end else if (8'hde == _T_19[7:0]) begin
        image_1_222 <= io_pixelVal_in_1_1;
      end else if (8'hde == _T_15[7:0]) begin
        image_1_222 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_223 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hdf == _T_34[7:0]) begin
        image_1_223 <= io_pixelVal_in_1_6;
      end else if (8'hdf == _T_31[7:0]) begin
        image_1_223 <= io_pixelVal_in_1_5;
      end else if (8'hdf == _T_28[7:0]) begin
        image_1_223 <= io_pixelVal_in_1_4;
      end else if (8'hdf == _T_25[7:0]) begin
        image_1_223 <= io_pixelVal_in_1_3;
      end else if (8'hdf == _T_22[7:0]) begin
        image_1_223 <= io_pixelVal_in_1_2;
      end else if (8'hdf == _T_19[7:0]) begin
        image_1_223 <= io_pixelVal_in_1_1;
      end else if (8'hdf == _T_15[7:0]) begin
        image_1_223 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_224 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he0 == _T_34[7:0]) begin
        image_1_224 <= io_pixelVal_in_1_6;
      end else if (8'he0 == _T_31[7:0]) begin
        image_1_224 <= io_pixelVal_in_1_5;
      end else if (8'he0 == _T_28[7:0]) begin
        image_1_224 <= io_pixelVal_in_1_4;
      end else if (8'he0 == _T_25[7:0]) begin
        image_1_224 <= io_pixelVal_in_1_3;
      end else if (8'he0 == _T_22[7:0]) begin
        image_1_224 <= io_pixelVal_in_1_2;
      end else if (8'he0 == _T_19[7:0]) begin
        image_1_224 <= io_pixelVal_in_1_1;
      end else if (8'he0 == _T_15[7:0]) begin
        image_1_224 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_225 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he1 == _T_34[7:0]) begin
        image_1_225 <= io_pixelVal_in_1_6;
      end else if (8'he1 == _T_31[7:0]) begin
        image_1_225 <= io_pixelVal_in_1_5;
      end else if (8'he1 == _T_28[7:0]) begin
        image_1_225 <= io_pixelVal_in_1_4;
      end else if (8'he1 == _T_25[7:0]) begin
        image_1_225 <= io_pixelVal_in_1_3;
      end else if (8'he1 == _T_22[7:0]) begin
        image_1_225 <= io_pixelVal_in_1_2;
      end else if (8'he1 == _T_19[7:0]) begin
        image_1_225 <= io_pixelVal_in_1_1;
      end else if (8'he1 == _T_15[7:0]) begin
        image_1_225 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_226 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he2 == _T_34[7:0]) begin
        image_1_226 <= io_pixelVal_in_1_6;
      end else if (8'he2 == _T_31[7:0]) begin
        image_1_226 <= io_pixelVal_in_1_5;
      end else if (8'he2 == _T_28[7:0]) begin
        image_1_226 <= io_pixelVal_in_1_4;
      end else if (8'he2 == _T_25[7:0]) begin
        image_1_226 <= io_pixelVal_in_1_3;
      end else if (8'he2 == _T_22[7:0]) begin
        image_1_226 <= io_pixelVal_in_1_2;
      end else if (8'he2 == _T_19[7:0]) begin
        image_1_226 <= io_pixelVal_in_1_1;
      end else if (8'he2 == _T_15[7:0]) begin
        image_1_226 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_227 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he3 == _T_34[7:0]) begin
        image_1_227 <= io_pixelVal_in_1_6;
      end else if (8'he3 == _T_31[7:0]) begin
        image_1_227 <= io_pixelVal_in_1_5;
      end else if (8'he3 == _T_28[7:0]) begin
        image_1_227 <= io_pixelVal_in_1_4;
      end else if (8'he3 == _T_25[7:0]) begin
        image_1_227 <= io_pixelVal_in_1_3;
      end else if (8'he3 == _T_22[7:0]) begin
        image_1_227 <= io_pixelVal_in_1_2;
      end else if (8'he3 == _T_19[7:0]) begin
        image_1_227 <= io_pixelVal_in_1_1;
      end else if (8'he3 == _T_15[7:0]) begin
        image_1_227 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_228 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he4 == _T_34[7:0]) begin
        image_1_228 <= io_pixelVal_in_1_6;
      end else if (8'he4 == _T_31[7:0]) begin
        image_1_228 <= io_pixelVal_in_1_5;
      end else if (8'he4 == _T_28[7:0]) begin
        image_1_228 <= io_pixelVal_in_1_4;
      end else if (8'he4 == _T_25[7:0]) begin
        image_1_228 <= io_pixelVal_in_1_3;
      end else if (8'he4 == _T_22[7:0]) begin
        image_1_228 <= io_pixelVal_in_1_2;
      end else if (8'he4 == _T_19[7:0]) begin
        image_1_228 <= io_pixelVal_in_1_1;
      end else if (8'he4 == _T_15[7:0]) begin
        image_1_228 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_229 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he5 == _T_34[7:0]) begin
        image_1_229 <= io_pixelVal_in_1_6;
      end else if (8'he5 == _T_31[7:0]) begin
        image_1_229 <= io_pixelVal_in_1_5;
      end else if (8'he5 == _T_28[7:0]) begin
        image_1_229 <= io_pixelVal_in_1_4;
      end else if (8'he5 == _T_25[7:0]) begin
        image_1_229 <= io_pixelVal_in_1_3;
      end else if (8'he5 == _T_22[7:0]) begin
        image_1_229 <= io_pixelVal_in_1_2;
      end else if (8'he5 == _T_19[7:0]) begin
        image_1_229 <= io_pixelVal_in_1_1;
      end else if (8'he5 == _T_15[7:0]) begin
        image_1_229 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_230 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he6 == _T_34[7:0]) begin
        image_1_230 <= io_pixelVal_in_1_6;
      end else if (8'he6 == _T_31[7:0]) begin
        image_1_230 <= io_pixelVal_in_1_5;
      end else if (8'he6 == _T_28[7:0]) begin
        image_1_230 <= io_pixelVal_in_1_4;
      end else if (8'he6 == _T_25[7:0]) begin
        image_1_230 <= io_pixelVal_in_1_3;
      end else if (8'he6 == _T_22[7:0]) begin
        image_1_230 <= io_pixelVal_in_1_2;
      end else if (8'he6 == _T_19[7:0]) begin
        image_1_230 <= io_pixelVal_in_1_1;
      end else if (8'he6 == _T_15[7:0]) begin
        image_1_230 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_231 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he7 == _T_34[7:0]) begin
        image_1_231 <= io_pixelVal_in_1_6;
      end else if (8'he7 == _T_31[7:0]) begin
        image_1_231 <= io_pixelVal_in_1_5;
      end else if (8'he7 == _T_28[7:0]) begin
        image_1_231 <= io_pixelVal_in_1_4;
      end else if (8'he7 == _T_25[7:0]) begin
        image_1_231 <= io_pixelVal_in_1_3;
      end else if (8'he7 == _T_22[7:0]) begin
        image_1_231 <= io_pixelVal_in_1_2;
      end else if (8'he7 == _T_19[7:0]) begin
        image_1_231 <= io_pixelVal_in_1_1;
      end else if (8'he7 == _T_15[7:0]) begin
        image_1_231 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_232 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he8 == _T_34[7:0]) begin
        image_1_232 <= io_pixelVal_in_1_6;
      end else if (8'he8 == _T_31[7:0]) begin
        image_1_232 <= io_pixelVal_in_1_5;
      end else if (8'he8 == _T_28[7:0]) begin
        image_1_232 <= io_pixelVal_in_1_4;
      end else if (8'he8 == _T_25[7:0]) begin
        image_1_232 <= io_pixelVal_in_1_3;
      end else if (8'he8 == _T_22[7:0]) begin
        image_1_232 <= io_pixelVal_in_1_2;
      end else if (8'he8 == _T_19[7:0]) begin
        image_1_232 <= io_pixelVal_in_1_1;
      end else if (8'he8 == _T_15[7:0]) begin
        image_1_232 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_233 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he9 == _T_34[7:0]) begin
        image_1_233 <= io_pixelVal_in_1_6;
      end else if (8'he9 == _T_31[7:0]) begin
        image_1_233 <= io_pixelVal_in_1_5;
      end else if (8'he9 == _T_28[7:0]) begin
        image_1_233 <= io_pixelVal_in_1_4;
      end else if (8'he9 == _T_25[7:0]) begin
        image_1_233 <= io_pixelVal_in_1_3;
      end else if (8'he9 == _T_22[7:0]) begin
        image_1_233 <= io_pixelVal_in_1_2;
      end else if (8'he9 == _T_19[7:0]) begin
        image_1_233 <= io_pixelVal_in_1_1;
      end else if (8'he9 == _T_15[7:0]) begin
        image_1_233 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_234 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hea == _T_34[7:0]) begin
        image_1_234 <= io_pixelVal_in_1_6;
      end else if (8'hea == _T_31[7:0]) begin
        image_1_234 <= io_pixelVal_in_1_5;
      end else if (8'hea == _T_28[7:0]) begin
        image_1_234 <= io_pixelVal_in_1_4;
      end else if (8'hea == _T_25[7:0]) begin
        image_1_234 <= io_pixelVal_in_1_3;
      end else if (8'hea == _T_22[7:0]) begin
        image_1_234 <= io_pixelVal_in_1_2;
      end else if (8'hea == _T_19[7:0]) begin
        image_1_234 <= io_pixelVal_in_1_1;
      end else if (8'hea == _T_15[7:0]) begin
        image_1_234 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_235 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'heb == _T_34[7:0]) begin
        image_1_235 <= io_pixelVal_in_1_6;
      end else if (8'heb == _T_31[7:0]) begin
        image_1_235 <= io_pixelVal_in_1_5;
      end else if (8'heb == _T_28[7:0]) begin
        image_1_235 <= io_pixelVal_in_1_4;
      end else if (8'heb == _T_25[7:0]) begin
        image_1_235 <= io_pixelVal_in_1_3;
      end else if (8'heb == _T_22[7:0]) begin
        image_1_235 <= io_pixelVal_in_1_2;
      end else if (8'heb == _T_19[7:0]) begin
        image_1_235 <= io_pixelVal_in_1_1;
      end else if (8'heb == _T_15[7:0]) begin
        image_1_235 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_236 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hec == _T_34[7:0]) begin
        image_1_236 <= io_pixelVal_in_1_6;
      end else if (8'hec == _T_31[7:0]) begin
        image_1_236 <= io_pixelVal_in_1_5;
      end else if (8'hec == _T_28[7:0]) begin
        image_1_236 <= io_pixelVal_in_1_4;
      end else if (8'hec == _T_25[7:0]) begin
        image_1_236 <= io_pixelVal_in_1_3;
      end else if (8'hec == _T_22[7:0]) begin
        image_1_236 <= io_pixelVal_in_1_2;
      end else if (8'hec == _T_19[7:0]) begin
        image_1_236 <= io_pixelVal_in_1_1;
      end else if (8'hec == _T_15[7:0]) begin
        image_1_236 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_237 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hed == _T_34[7:0]) begin
        image_1_237 <= io_pixelVal_in_1_6;
      end else if (8'hed == _T_31[7:0]) begin
        image_1_237 <= io_pixelVal_in_1_5;
      end else if (8'hed == _T_28[7:0]) begin
        image_1_237 <= io_pixelVal_in_1_4;
      end else if (8'hed == _T_25[7:0]) begin
        image_1_237 <= io_pixelVal_in_1_3;
      end else if (8'hed == _T_22[7:0]) begin
        image_1_237 <= io_pixelVal_in_1_2;
      end else if (8'hed == _T_19[7:0]) begin
        image_1_237 <= io_pixelVal_in_1_1;
      end else if (8'hed == _T_15[7:0]) begin
        image_1_237 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_238 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hee == _T_34[7:0]) begin
        image_1_238 <= io_pixelVal_in_1_6;
      end else if (8'hee == _T_31[7:0]) begin
        image_1_238 <= io_pixelVal_in_1_5;
      end else if (8'hee == _T_28[7:0]) begin
        image_1_238 <= io_pixelVal_in_1_4;
      end else if (8'hee == _T_25[7:0]) begin
        image_1_238 <= io_pixelVal_in_1_3;
      end else if (8'hee == _T_22[7:0]) begin
        image_1_238 <= io_pixelVal_in_1_2;
      end else if (8'hee == _T_19[7:0]) begin
        image_1_238 <= io_pixelVal_in_1_1;
      end else if (8'hee == _T_15[7:0]) begin
        image_1_238 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_239 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hef == _T_34[7:0]) begin
        image_1_239 <= io_pixelVal_in_1_6;
      end else if (8'hef == _T_31[7:0]) begin
        image_1_239 <= io_pixelVal_in_1_5;
      end else if (8'hef == _T_28[7:0]) begin
        image_1_239 <= io_pixelVal_in_1_4;
      end else if (8'hef == _T_25[7:0]) begin
        image_1_239 <= io_pixelVal_in_1_3;
      end else if (8'hef == _T_22[7:0]) begin
        image_1_239 <= io_pixelVal_in_1_2;
      end else if (8'hef == _T_19[7:0]) begin
        image_1_239 <= io_pixelVal_in_1_1;
      end else if (8'hef == _T_15[7:0]) begin
        image_1_239 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_240 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf0 == _T_34[7:0]) begin
        image_1_240 <= io_pixelVal_in_1_6;
      end else if (8'hf0 == _T_31[7:0]) begin
        image_1_240 <= io_pixelVal_in_1_5;
      end else if (8'hf0 == _T_28[7:0]) begin
        image_1_240 <= io_pixelVal_in_1_4;
      end else if (8'hf0 == _T_25[7:0]) begin
        image_1_240 <= io_pixelVal_in_1_3;
      end else if (8'hf0 == _T_22[7:0]) begin
        image_1_240 <= io_pixelVal_in_1_2;
      end else if (8'hf0 == _T_19[7:0]) begin
        image_1_240 <= io_pixelVal_in_1_1;
      end else if (8'hf0 == _T_15[7:0]) begin
        image_1_240 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_241 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf1 == _T_34[7:0]) begin
        image_1_241 <= io_pixelVal_in_1_6;
      end else if (8'hf1 == _T_31[7:0]) begin
        image_1_241 <= io_pixelVal_in_1_5;
      end else if (8'hf1 == _T_28[7:0]) begin
        image_1_241 <= io_pixelVal_in_1_4;
      end else if (8'hf1 == _T_25[7:0]) begin
        image_1_241 <= io_pixelVal_in_1_3;
      end else if (8'hf1 == _T_22[7:0]) begin
        image_1_241 <= io_pixelVal_in_1_2;
      end else if (8'hf1 == _T_19[7:0]) begin
        image_1_241 <= io_pixelVal_in_1_1;
      end else if (8'hf1 == _T_15[7:0]) begin
        image_1_241 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_242 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf2 == _T_34[7:0]) begin
        image_1_242 <= io_pixelVal_in_1_6;
      end else if (8'hf2 == _T_31[7:0]) begin
        image_1_242 <= io_pixelVal_in_1_5;
      end else if (8'hf2 == _T_28[7:0]) begin
        image_1_242 <= io_pixelVal_in_1_4;
      end else if (8'hf2 == _T_25[7:0]) begin
        image_1_242 <= io_pixelVal_in_1_3;
      end else if (8'hf2 == _T_22[7:0]) begin
        image_1_242 <= io_pixelVal_in_1_2;
      end else if (8'hf2 == _T_19[7:0]) begin
        image_1_242 <= io_pixelVal_in_1_1;
      end else if (8'hf2 == _T_15[7:0]) begin
        image_1_242 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_243 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf3 == _T_34[7:0]) begin
        image_1_243 <= io_pixelVal_in_1_6;
      end else if (8'hf3 == _T_31[7:0]) begin
        image_1_243 <= io_pixelVal_in_1_5;
      end else if (8'hf3 == _T_28[7:0]) begin
        image_1_243 <= io_pixelVal_in_1_4;
      end else if (8'hf3 == _T_25[7:0]) begin
        image_1_243 <= io_pixelVal_in_1_3;
      end else if (8'hf3 == _T_22[7:0]) begin
        image_1_243 <= io_pixelVal_in_1_2;
      end else if (8'hf3 == _T_19[7:0]) begin
        image_1_243 <= io_pixelVal_in_1_1;
      end else if (8'hf3 == _T_15[7:0]) begin
        image_1_243 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_244 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf4 == _T_34[7:0]) begin
        image_1_244 <= io_pixelVal_in_1_6;
      end else if (8'hf4 == _T_31[7:0]) begin
        image_1_244 <= io_pixelVal_in_1_5;
      end else if (8'hf4 == _T_28[7:0]) begin
        image_1_244 <= io_pixelVal_in_1_4;
      end else if (8'hf4 == _T_25[7:0]) begin
        image_1_244 <= io_pixelVal_in_1_3;
      end else if (8'hf4 == _T_22[7:0]) begin
        image_1_244 <= io_pixelVal_in_1_2;
      end else if (8'hf4 == _T_19[7:0]) begin
        image_1_244 <= io_pixelVal_in_1_1;
      end else if (8'hf4 == _T_15[7:0]) begin
        image_1_244 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_245 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf5 == _T_34[7:0]) begin
        image_1_245 <= io_pixelVal_in_1_6;
      end else if (8'hf5 == _T_31[7:0]) begin
        image_1_245 <= io_pixelVal_in_1_5;
      end else if (8'hf5 == _T_28[7:0]) begin
        image_1_245 <= io_pixelVal_in_1_4;
      end else if (8'hf5 == _T_25[7:0]) begin
        image_1_245 <= io_pixelVal_in_1_3;
      end else if (8'hf5 == _T_22[7:0]) begin
        image_1_245 <= io_pixelVal_in_1_2;
      end else if (8'hf5 == _T_19[7:0]) begin
        image_1_245 <= io_pixelVal_in_1_1;
      end else if (8'hf5 == _T_15[7:0]) begin
        image_1_245 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_246 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf6 == _T_34[7:0]) begin
        image_1_246 <= io_pixelVal_in_1_6;
      end else if (8'hf6 == _T_31[7:0]) begin
        image_1_246 <= io_pixelVal_in_1_5;
      end else if (8'hf6 == _T_28[7:0]) begin
        image_1_246 <= io_pixelVal_in_1_4;
      end else if (8'hf6 == _T_25[7:0]) begin
        image_1_246 <= io_pixelVal_in_1_3;
      end else if (8'hf6 == _T_22[7:0]) begin
        image_1_246 <= io_pixelVal_in_1_2;
      end else if (8'hf6 == _T_19[7:0]) begin
        image_1_246 <= io_pixelVal_in_1_1;
      end else if (8'hf6 == _T_15[7:0]) begin
        image_1_246 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_247 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf7 == _T_34[7:0]) begin
        image_1_247 <= io_pixelVal_in_1_6;
      end else if (8'hf7 == _T_31[7:0]) begin
        image_1_247 <= io_pixelVal_in_1_5;
      end else if (8'hf7 == _T_28[7:0]) begin
        image_1_247 <= io_pixelVal_in_1_4;
      end else if (8'hf7 == _T_25[7:0]) begin
        image_1_247 <= io_pixelVal_in_1_3;
      end else if (8'hf7 == _T_22[7:0]) begin
        image_1_247 <= io_pixelVal_in_1_2;
      end else if (8'hf7 == _T_19[7:0]) begin
        image_1_247 <= io_pixelVal_in_1_1;
      end else if (8'hf7 == _T_15[7:0]) begin
        image_1_247 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_248 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf8 == _T_34[7:0]) begin
        image_1_248 <= io_pixelVal_in_1_6;
      end else if (8'hf8 == _T_31[7:0]) begin
        image_1_248 <= io_pixelVal_in_1_5;
      end else if (8'hf8 == _T_28[7:0]) begin
        image_1_248 <= io_pixelVal_in_1_4;
      end else if (8'hf8 == _T_25[7:0]) begin
        image_1_248 <= io_pixelVal_in_1_3;
      end else if (8'hf8 == _T_22[7:0]) begin
        image_1_248 <= io_pixelVal_in_1_2;
      end else if (8'hf8 == _T_19[7:0]) begin
        image_1_248 <= io_pixelVal_in_1_1;
      end else if (8'hf8 == _T_15[7:0]) begin
        image_1_248 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_249 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf9 == _T_34[7:0]) begin
        image_1_249 <= io_pixelVal_in_1_6;
      end else if (8'hf9 == _T_31[7:0]) begin
        image_1_249 <= io_pixelVal_in_1_5;
      end else if (8'hf9 == _T_28[7:0]) begin
        image_1_249 <= io_pixelVal_in_1_4;
      end else if (8'hf9 == _T_25[7:0]) begin
        image_1_249 <= io_pixelVal_in_1_3;
      end else if (8'hf9 == _T_22[7:0]) begin
        image_1_249 <= io_pixelVal_in_1_2;
      end else if (8'hf9 == _T_19[7:0]) begin
        image_1_249 <= io_pixelVal_in_1_1;
      end else if (8'hf9 == _T_15[7:0]) begin
        image_1_249 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_250 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hfa == _T_34[7:0]) begin
        image_1_250 <= io_pixelVal_in_1_6;
      end else if (8'hfa == _T_31[7:0]) begin
        image_1_250 <= io_pixelVal_in_1_5;
      end else if (8'hfa == _T_28[7:0]) begin
        image_1_250 <= io_pixelVal_in_1_4;
      end else if (8'hfa == _T_25[7:0]) begin
        image_1_250 <= io_pixelVal_in_1_3;
      end else if (8'hfa == _T_22[7:0]) begin
        image_1_250 <= io_pixelVal_in_1_2;
      end else if (8'hfa == _T_19[7:0]) begin
        image_1_250 <= io_pixelVal_in_1_1;
      end else if (8'hfa == _T_15[7:0]) begin
        image_1_250 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_251 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hfb == _T_34[7:0]) begin
        image_1_251 <= io_pixelVal_in_1_6;
      end else if (8'hfb == _T_31[7:0]) begin
        image_1_251 <= io_pixelVal_in_1_5;
      end else if (8'hfb == _T_28[7:0]) begin
        image_1_251 <= io_pixelVal_in_1_4;
      end else if (8'hfb == _T_25[7:0]) begin
        image_1_251 <= io_pixelVal_in_1_3;
      end else if (8'hfb == _T_22[7:0]) begin
        image_1_251 <= io_pixelVal_in_1_2;
      end else if (8'hfb == _T_19[7:0]) begin
        image_1_251 <= io_pixelVal_in_1_1;
      end else if (8'hfb == _T_15[7:0]) begin
        image_1_251 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_2_0 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h0 == _T_34[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_6;
      end else if (8'h0 == _T_31[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_5;
      end else if (8'h0 == _T_28[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_4;
      end else if (8'h0 == _T_25[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_3;
      end else if (8'h0 == _T_22[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_2;
      end else if (8'h0 == _T_19[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_1;
      end else if (8'h0 == _T_15[7:0]) begin
        image_2_0 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_1 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1 == _T_34[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_6;
      end else if (8'h1 == _T_31[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_5;
      end else if (8'h1 == _T_28[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_4;
      end else if (8'h1 == _T_25[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_3;
      end else if (8'h1 == _T_22[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_2;
      end else if (8'h1 == _T_19[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_1;
      end else if (8'h1 == _T_15[7:0]) begin
        image_2_1 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_2 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2 == _T_34[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_6;
      end else if (8'h2 == _T_31[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_5;
      end else if (8'h2 == _T_28[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_4;
      end else if (8'h2 == _T_25[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_3;
      end else if (8'h2 == _T_22[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_2;
      end else if (8'h2 == _T_19[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_1;
      end else if (8'h2 == _T_15[7:0]) begin
        image_2_2 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_3 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3 == _T_34[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_6;
      end else if (8'h3 == _T_31[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_5;
      end else if (8'h3 == _T_28[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_4;
      end else if (8'h3 == _T_25[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_3;
      end else if (8'h3 == _T_22[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_2;
      end else if (8'h3 == _T_19[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_1;
      end else if (8'h3 == _T_15[7:0]) begin
        image_2_3 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_4 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4 == _T_34[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_6;
      end else if (8'h4 == _T_31[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_5;
      end else if (8'h4 == _T_28[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_4;
      end else if (8'h4 == _T_25[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_3;
      end else if (8'h4 == _T_22[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_2;
      end else if (8'h4 == _T_19[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_1;
      end else if (8'h4 == _T_15[7:0]) begin
        image_2_4 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_5 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5 == _T_34[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_6;
      end else if (8'h5 == _T_31[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_5;
      end else if (8'h5 == _T_28[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_4;
      end else if (8'h5 == _T_25[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_3;
      end else if (8'h5 == _T_22[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_2;
      end else if (8'h5 == _T_19[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_1;
      end else if (8'h5 == _T_15[7:0]) begin
        image_2_5 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_6 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6 == _T_34[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_6;
      end else if (8'h6 == _T_31[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_5;
      end else if (8'h6 == _T_28[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_4;
      end else if (8'h6 == _T_25[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_3;
      end else if (8'h6 == _T_22[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_2;
      end else if (8'h6 == _T_19[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_1;
      end else if (8'h6 == _T_15[7:0]) begin
        image_2_6 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_7 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7 == _T_34[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_6;
      end else if (8'h7 == _T_31[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_5;
      end else if (8'h7 == _T_28[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_4;
      end else if (8'h7 == _T_25[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_3;
      end else if (8'h7 == _T_22[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_2;
      end else if (8'h7 == _T_19[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_1;
      end else if (8'h7 == _T_15[7:0]) begin
        image_2_7 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_8 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8 == _T_34[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_6;
      end else if (8'h8 == _T_31[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_5;
      end else if (8'h8 == _T_28[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_4;
      end else if (8'h8 == _T_25[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_3;
      end else if (8'h8 == _T_22[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_2;
      end else if (8'h8 == _T_19[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_1;
      end else if (8'h8 == _T_15[7:0]) begin
        image_2_8 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_9 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9 == _T_34[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_6;
      end else if (8'h9 == _T_31[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_5;
      end else if (8'h9 == _T_28[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_4;
      end else if (8'h9 == _T_25[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_3;
      end else if (8'h9 == _T_22[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_2;
      end else if (8'h9 == _T_19[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_1;
      end else if (8'h9 == _T_15[7:0]) begin
        image_2_9 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_10 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha == _T_34[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_6;
      end else if (8'ha == _T_31[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_5;
      end else if (8'ha == _T_28[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_4;
      end else if (8'ha == _T_25[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_3;
      end else if (8'ha == _T_22[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_2;
      end else if (8'ha == _T_19[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_1;
      end else if (8'ha == _T_15[7:0]) begin
        image_2_10 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_11 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb == _T_34[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_6;
      end else if (8'hb == _T_31[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_5;
      end else if (8'hb == _T_28[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_4;
      end else if (8'hb == _T_25[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_3;
      end else if (8'hb == _T_22[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_2;
      end else if (8'hb == _T_19[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_1;
      end else if (8'hb == _T_15[7:0]) begin
        image_2_11 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_12 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc == _T_34[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_6;
      end else if (8'hc == _T_31[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_5;
      end else if (8'hc == _T_28[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_4;
      end else if (8'hc == _T_25[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_3;
      end else if (8'hc == _T_22[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_2;
      end else if (8'hc == _T_19[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_1;
      end else if (8'hc == _T_15[7:0]) begin
        image_2_12 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_13 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd == _T_34[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_6;
      end else if (8'hd == _T_31[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_5;
      end else if (8'hd == _T_28[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_4;
      end else if (8'hd == _T_25[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_3;
      end else if (8'hd == _T_22[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_2;
      end else if (8'hd == _T_19[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_1;
      end else if (8'hd == _T_15[7:0]) begin
        image_2_13 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_14 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he == _T_34[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_6;
      end else if (8'he == _T_31[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_5;
      end else if (8'he == _T_28[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_4;
      end else if (8'he == _T_25[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_3;
      end else if (8'he == _T_22[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_2;
      end else if (8'he == _T_19[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_1;
      end else if (8'he == _T_15[7:0]) begin
        image_2_14 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_15 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf == _T_34[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_6;
      end else if (8'hf == _T_31[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_5;
      end else if (8'hf == _T_28[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_4;
      end else if (8'hf == _T_25[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_3;
      end else if (8'hf == _T_22[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_2;
      end else if (8'hf == _T_19[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_1;
      end else if (8'hf == _T_15[7:0]) begin
        image_2_15 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_16 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h10 == _T_34[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_6;
      end else if (8'h10 == _T_31[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_5;
      end else if (8'h10 == _T_28[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_4;
      end else if (8'h10 == _T_25[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_3;
      end else if (8'h10 == _T_22[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_2;
      end else if (8'h10 == _T_19[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_1;
      end else if (8'h10 == _T_15[7:0]) begin
        image_2_16 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_17 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h11 == _T_34[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_6;
      end else if (8'h11 == _T_31[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_5;
      end else if (8'h11 == _T_28[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_4;
      end else if (8'h11 == _T_25[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_3;
      end else if (8'h11 == _T_22[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_2;
      end else if (8'h11 == _T_19[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_1;
      end else if (8'h11 == _T_15[7:0]) begin
        image_2_17 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_18 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h12 == _T_34[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_6;
      end else if (8'h12 == _T_31[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_5;
      end else if (8'h12 == _T_28[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_4;
      end else if (8'h12 == _T_25[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_3;
      end else if (8'h12 == _T_22[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_2;
      end else if (8'h12 == _T_19[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_1;
      end else if (8'h12 == _T_15[7:0]) begin
        image_2_18 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_19 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h13 == _T_34[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_6;
      end else if (8'h13 == _T_31[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_5;
      end else if (8'h13 == _T_28[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_4;
      end else if (8'h13 == _T_25[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_3;
      end else if (8'h13 == _T_22[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_2;
      end else if (8'h13 == _T_19[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_1;
      end else if (8'h13 == _T_15[7:0]) begin
        image_2_19 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_20 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h14 == _T_34[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_6;
      end else if (8'h14 == _T_31[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_5;
      end else if (8'h14 == _T_28[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_4;
      end else if (8'h14 == _T_25[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_3;
      end else if (8'h14 == _T_22[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_2;
      end else if (8'h14 == _T_19[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_1;
      end else if (8'h14 == _T_15[7:0]) begin
        image_2_20 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_21 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h15 == _T_34[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_6;
      end else if (8'h15 == _T_31[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_5;
      end else if (8'h15 == _T_28[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_4;
      end else if (8'h15 == _T_25[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_3;
      end else if (8'h15 == _T_22[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_2;
      end else if (8'h15 == _T_19[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_1;
      end else if (8'h15 == _T_15[7:0]) begin
        image_2_21 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_22 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h16 == _T_34[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_6;
      end else if (8'h16 == _T_31[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_5;
      end else if (8'h16 == _T_28[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_4;
      end else if (8'h16 == _T_25[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_3;
      end else if (8'h16 == _T_22[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_2;
      end else if (8'h16 == _T_19[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_1;
      end else if (8'h16 == _T_15[7:0]) begin
        image_2_22 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_23 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h17 == _T_34[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_6;
      end else if (8'h17 == _T_31[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_5;
      end else if (8'h17 == _T_28[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_4;
      end else if (8'h17 == _T_25[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_3;
      end else if (8'h17 == _T_22[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_2;
      end else if (8'h17 == _T_19[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_1;
      end else if (8'h17 == _T_15[7:0]) begin
        image_2_23 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_24 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h18 == _T_34[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_6;
      end else if (8'h18 == _T_31[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_5;
      end else if (8'h18 == _T_28[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_4;
      end else if (8'h18 == _T_25[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_3;
      end else if (8'h18 == _T_22[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_2;
      end else if (8'h18 == _T_19[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_1;
      end else if (8'h18 == _T_15[7:0]) begin
        image_2_24 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_25 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h19 == _T_34[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_6;
      end else if (8'h19 == _T_31[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_5;
      end else if (8'h19 == _T_28[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_4;
      end else if (8'h19 == _T_25[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_3;
      end else if (8'h19 == _T_22[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_2;
      end else if (8'h19 == _T_19[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_1;
      end else if (8'h19 == _T_15[7:0]) begin
        image_2_25 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_26 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1a == _T_34[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_6;
      end else if (8'h1a == _T_31[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_5;
      end else if (8'h1a == _T_28[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_4;
      end else if (8'h1a == _T_25[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_3;
      end else if (8'h1a == _T_22[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_2;
      end else if (8'h1a == _T_19[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_1;
      end else if (8'h1a == _T_15[7:0]) begin
        image_2_26 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_27 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1b == _T_34[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_6;
      end else if (8'h1b == _T_31[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_5;
      end else if (8'h1b == _T_28[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_4;
      end else if (8'h1b == _T_25[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_3;
      end else if (8'h1b == _T_22[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_2;
      end else if (8'h1b == _T_19[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_1;
      end else if (8'h1b == _T_15[7:0]) begin
        image_2_27 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_28 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1c == _T_34[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_6;
      end else if (8'h1c == _T_31[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_5;
      end else if (8'h1c == _T_28[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_4;
      end else if (8'h1c == _T_25[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_3;
      end else if (8'h1c == _T_22[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_2;
      end else if (8'h1c == _T_19[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_1;
      end else if (8'h1c == _T_15[7:0]) begin
        image_2_28 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_29 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1d == _T_34[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_6;
      end else if (8'h1d == _T_31[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_5;
      end else if (8'h1d == _T_28[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_4;
      end else if (8'h1d == _T_25[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_3;
      end else if (8'h1d == _T_22[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_2;
      end else if (8'h1d == _T_19[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_1;
      end else if (8'h1d == _T_15[7:0]) begin
        image_2_29 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_30 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1e == _T_34[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_6;
      end else if (8'h1e == _T_31[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_5;
      end else if (8'h1e == _T_28[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_4;
      end else if (8'h1e == _T_25[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_3;
      end else if (8'h1e == _T_22[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_2;
      end else if (8'h1e == _T_19[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_1;
      end else if (8'h1e == _T_15[7:0]) begin
        image_2_30 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_31 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h1f == _T_34[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_6;
      end else if (8'h1f == _T_31[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_5;
      end else if (8'h1f == _T_28[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_4;
      end else if (8'h1f == _T_25[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_3;
      end else if (8'h1f == _T_22[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_2;
      end else if (8'h1f == _T_19[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_1;
      end else if (8'h1f == _T_15[7:0]) begin
        image_2_31 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_32 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h20 == _T_34[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_6;
      end else if (8'h20 == _T_31[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_5;
      end else if (8'h20 == _T_28[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_4;
      end else if (8'h20 == _T_25[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_3;
      end else if (8'h20 == _T_22[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_2;
      end else if (8'h20 == _T_19[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_1;
      end else if (8'h20 == _T_15[7:0]) begin
        image_2_32 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_33 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h21 == _T_34[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_6;
      end else if (8'h21 == _T_31[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_5;
      end else if (8'h21 == _T_28[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_4;
      end else if (8'h21 == _T_25[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_3;
      end else if (8'h21 == _T_22[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_2;
      end else if (8'h21 == _T_19[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_1;
      end else if (8'h21 == _T_15[7:0]) begin
        image_2_33 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_34 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h22 == _T_34[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_6;
      end else if (8'h22 == _T_31[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_5;
      end else if (8'h22 == _T_28[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_4;
      end else if (8'h22 == _T_25[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_3;
      end else if (8'h22 == _T_22[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_2;
      end else if (8'h22 == _T_19[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_1;
      end else if (8'h22 == _T_15[7:0]) begin
        image_2_34 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_35 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h23 == _T_34[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_6;
      end else if (8'h23 == _T_31[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_5;
      end else if (8'h23 == _T_28[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_4;
      end else if (8'h23 == _T_25[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_3;
      end else if (8'h23 == _T_22[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_2;
      end else if (8'h23 == _T_19[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_1;
      end else if (8'h23 == _T_15[7:0]) begin
        image_2_35 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_36 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h24 == _T_34[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_6;
      end else if (8'h24 == _T_31[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_5;
      end else if (8'h24 == _T_28[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_4;
      end else if (8'h24 == _T_25[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_3;
      end else if (8'h24 == _T_22[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_2;
      end else if (8'h24 == _T_19[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_1;
      end else if (8'h24 == _T_15[7:0]) begin
        image_2_36 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_37 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h25 == _T_34[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_6;
      end else if (8'h25 == _T_31[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_5;
      end else if (8'h25 == _T_28[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_4;
      end else if (8'h25 == _T_25[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_3;
      end else if (8'h25 == _T_22[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_2;
      end else if (8'h25 == _T_19[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_1;
      end else if (8'h25 == _T_15[7:0]) begin
        image_2_37 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_38 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h26 == _T_34[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_6;
      end else if (8'h26 == _T_31[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_5;
      end else if (8'h26 == _T_28[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_4;
      end else if (8'h26 == _T_25[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_3;
      end else if (8'h26 == _T_22[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_2;
      end else if (8'h26 == _T_19[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_1;
      end else if (8'h26 == _T_15[7:0]) begin
        image_2_38 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_39 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h27 == _T_34[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_6;
      end else if (8'h27 == _T_31[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_5;
      end else if (8'h27 == _T_28[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_4;
      end else if (8'h27 == _T_25[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_3;
      end else if (8'h27 == _T_22[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_2;
      end else if (8'h27 == _T_19[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_1;
      end else if (8'h27 == _T_15[7:0]) begin
        image_2_39 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_40 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h28 == _T_34[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_6;
      end else if (8'h28 == _T_31[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_5;
      end else if (8'h28 == _T_28[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_4;
      end else if (8'h28 == _T_25[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_3;
      end else if (8'h28 == _T_22[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_2;
      end else if (8'h28 == _T_19[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_1;
      end else if (8'h28 == _T_15[7:0]) begin
        image_2_40 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_41 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h29 == _T_34[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_6;
      end else if (8'h29 == _T_31[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_5;
      end else if (8'h29 == _T_28[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_4;
      end else if (8'h29 == _T_25[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_3;
      end else if (8'h29 == _T_22[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_2;
      end else if (8'h29 == _T_19[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_1;
      end else if (8'h29 == _T_15[7:0]) begin
        image_2_41 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_42 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2a == _T_34[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_6;
      end else if (8'h2a == _T_31[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_5;
      end else if (8'h2a == _T_28[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_4;
      end else if (8'h2a == _T_25[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_3;
      end else if (8'h2a == _T_22[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_2;
      end else if (8'h2a == _T_19[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_1;
      end else if (8'h2a == _T_15[7:0]) begin
        image_2_42 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_43 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2b == _T_34[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_6;
      end else if (8'h2b == _T_31[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_5;
      end else if (8'h2b == _T_28[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_4;
      end else if (8'h2b == _T_25[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_3;
      end else if (8'h2b == _T_22[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_2;
      end else if (8'h2b == _T_19[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_1;
      end else if (8'h2b == _T_15[7:0]) begin
        image_2_43 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_44 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2c == _T_34[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_6;
      end else if (8'h2c == _T_31[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_5;
      end else if (8'h2c == _T_28[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_4;
      end else if (8'h2c == _T_25[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_3;
      end else if (8'h2c == _T_22[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_2;
      end else if (8'h2c == _T_19[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_1;
      end else if (8'h2c == _T_15[7:0]) begin
        image_2_44 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_45 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2d == _T_34[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_6;
      end else if (8'h2d == _T_31[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_5;
      end else if (8'h2d == _T_28[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_4;
      end else if (8'h2d == _T_25[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_3;
      end else if (8'h2d == _T_22[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_2;
      end else if (8'h2d == _T_19[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_1;
      end else if (8'h2d == _T_15[7:0]) begin
        image_2_45 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_46 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2e == _T_34[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_6;
      end else if (8'h2e == _T_31[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_5;
      end else if (8'h2e == _T_28[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_4;
      end else if (8'h2e == _T_25[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_3;
      end else if (8'h2e == _T_22[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_2;
      end else if (8'h2e == _T_19[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_1;
      end else if (8'h2e == _T_15[7:0]) begin
        image_2_46 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_47 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h2f == _T_34[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_6;
      end else if (8'h2f == _T_31[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_5;
      end else if (8'h2f == _T_28[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_4;
      end else if (8'h2f == _T_25[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_3;
      end else if (8'h2f == _T_22[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_2;
      end else if (8'h2f == _T_19[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_1;
      end else if (8'h2f == _T_15[7:0]) begin
        image_2_47 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_48 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h30 == _T_34[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_6;
      end else if (8'h30 == _T_31[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_5;
      end else if (8'h30 == _T_28[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_4;
      end else if (8'h30 == _T_25[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_3;
      end else if (8'h30 == _T_22[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_2;
      end else if (8'h30 == _T_19[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_1;
      end else if (8'h30 == _T_15[7:0]) begin
        image_2_48 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_49 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h31 == _T_34[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_6;
      end else if (8'h31 == _T_31[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_5;
      end else if (8'h31 == _T_28[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_4;
      end else if (8'h31 == _T_25[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_3;
      end else if (8'h31 == _T_22[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_2;
      end else if (8'h31 == _T_19[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_1;
      end else if (8'h31 == _T_15[7:0]) begin
        image_2_49 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_50 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h32 == _T_34[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_6;
      end else if (8'h32 == _T_31[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_5;
      end else if (8'h32 == _T_28[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_4;
      end else if (8'h32 == _T_25[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_3;
      end else if (8'h32 == _T_22[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_2;
      end else if (8'h32 == _T_19[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_1;
      end else if (8'h32 == _T_15[7:0]) begin
        image_2_50 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_51 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h33 == _T_34[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_6;
      end else if (8'h33 == _T_31[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_5;
      end else if (8'h33 == _T_28[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_4;
      end else if (8'h33 == _T_25[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_3;
      end else if (8'h33 == _T_22[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_2;
      end else if (8'h33 == _T_19[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_1;
      end else if (8'h33 == _T_15[7:0]) begin
        image_2_51 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_52 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h34 == _T_34[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_6;
      end else if (8'h34 == _T_31[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_5;
      end else if (8'h34 == _T_28[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_4;
      end else if (8'h34 == _T_25[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_3;
      end else if (8'h34 == _T_22[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_2;
      end else if (8'h34 == _T_19[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_1;
      end else if (8'h34 == _T_15[7:0]) begin
        image_2_52 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_53 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h35 == _T_34[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_6;
      end else if (8'h35 == _T_31[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_5;
      end else if (8'h35 == _T_28[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_4;
      end else if (8'h35 == _T_25[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_3;
      end else if (8'h35 == _T_22[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_2;
      end else if (8'h35 == _T_19[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_1;
      end else if (8'h35 == _T_15[7:0]) begin
        image_2_53 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_54 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h36 == _T_34[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_6;
      end else if (8'h36 == _T_31[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_5;
      end else if (8'h36 == _T_28[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_4;
      end else if (8'h36 == _T_25[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_3;
      end else if (8'h36 == _T_22[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_2;
      end else if (8'h36 == _T_19[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_1;
      end else if (8'h36 == _T_15[7:0]) begin
        image_2_54 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_55 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h37 == _T_34[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_6;
      end else if (8'h37 == _T_31[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_5;
      end else if (8'h37 == _T_28[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_4;
      end else if (8'h37 == _T_25[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_3;
      end else if (8'h37 == _T_22[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_2;
      end else if (8'h37 == _T_19[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_1;
      end else if (8'h37 == _T_15[7:0]) begin
        image_2_55 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_56 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h38 == _T_34[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_6;
      end else if (8'h38 == _T_31[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_5;
      end else if (8'h38 == _T_28[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_4;
      end else if (8'h38 == _T_25[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_3;
      end else if (8'h38 == _T_22[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_2;
      end else if (8'h38 == _T_19[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_1;
      end else if (8'h38 == _T_15[7:0]) begin
        image_2_56 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_57 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h39 == _T_34[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_6;
      end else if (8'h39 == _T_31[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_5;
      end else if (8'h39 == _T_28[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_4;
      end else if (8'h39 == _T_25[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_3;
      end else if (8'h39 == _T_22[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_2;
      end else if (8'h39 == _T_19[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_1;
      end else if (8'h39 == _T_15[7:0]) begin
        image_2_57 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_58 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3a == _T_34[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_6;
      end else if (8'h3a == _T_31[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_5;
      end else if (8'h3a == _T_28[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_4;
      end else if (8'h3a == _T_25[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_3;
      end else if (8'h3a == _T_22[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_2;
      end else if (8'h3a == _T_19[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_1;
      end else if (8'h3a == _T_15[7:0]) begin
        image_2_58 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_59 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3b == _T_34[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_6;
      end else if (8'h3b == _T_31[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_5;
      end else if (8'h3b == _T_28[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_4;
      end else if (8'h3b == _T_25[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_3;
      end else if (8'h3b == _T_22[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_2;
      end else if (8'h3b == _T_19[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_1;
      end else if (8'h3b == _T_15[7:0]) begin
        image_2_59 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_60 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3c == _T_34[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_6;
      end else if (8'h3c == _T_31[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_5;
      end else if (8'h3c == _T_28[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_4;
      end else if (8'h3c == _T_25[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_3;
      end else if (8'h3c == _T_22[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_2;
      end else if (8'h3c == _T_19[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_1;
      end else if (8'h3c == _T_15[7:0]) begin
        image_2_60 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_61 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3d == _T_34[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_6;
      end else if (8'h3d == _T_31[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_5;
      end else if (8'h3d == _T_28[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_4;
      end else if (8'h3d == _T_25[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_3;
      end else if (8'h3d == _T_22[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_2;
      end else if (8'h3d == _T_19[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_1;
      end else if (8'h3d == _T_15[7:0]) begin
        image_2_61 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_62 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3e == _T_34[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_6;
      end else if (8'h3e == _T_31[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_5;
      end else if (8'h3e == _T_28[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_4;
      end else if (8'h3e == _T_25[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_3;
      end else if (8'h3e == _T_22[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_2;
      end else if (8'h3e == _T_19[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_1;
      end else if (8'h3e == _T_15[7:0]) begin
        image_2_62 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_63 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h3f == _T_34[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_6;
      end else if (8'h3f == _T_31[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_5;
      end else if (8'h3f == _T_28[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_4;
      end else if (8'h3f == _T_25[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_3;
      end else if (8'h3f == _T_22[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_2;
      end else if (8'h3f == _T_19[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_1;
      end else if (8'h3f == _T_15[7:0]) begin
        image_2_63 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_64 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h40 == _T_34[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_6;
      end else if (8'h40 == _T_31[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_5;
      end else if (8'h40 == _T_28[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_4;
      end else if (8'h40 == _T_25[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_3;
      end else if (8'h40 == _T_22[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_2;
      end else if (8'h40 == _T_19[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_1;
      end else if (8'h40 == _T_15[7:0]) begin
        image_2_64 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_65 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h41 == _T_34[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_6;
      end else if (8'h41 == _T_31[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_5;
      end else if (8'h41 == _T_28[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_4;
      end else if (8'h41 == _T_25[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_3;
      end else if (8'h41 == _T_22[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_2;
      end else if (8'h41 == _T_19[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_1;
      end else if (8'h41 == _T_15[7:0]) begin
        image_2_65 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_66 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h42 == _T_34[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_6;
      end else if (8'h42 == _T_31[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_5;
      end else if (8'h42 == _T_28[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_4;
      end else if (8'h42 == _T_25[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_3;
      end else if (8'h42 == _T_22[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_2;
      end else if (8'h42 == _T_19[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_1;
      end else if (8'h42 == _T_15[7:0]) begin
        image_2_66 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_67 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h43 == _T_34[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_6;
      end else if (8'h43 == _T_31[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_5;
      end else if (8'h43 == _T_28[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_4;
      end else if (8'h43 == _T_25[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_3;
      end else if (8'h43 == _T_22[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_2;
      end else if (8'h43 == _T_19[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_1;
      end else if (8'h43 == _T_15[7:0]) begin
        image_2_67 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_68 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h44 == _T_34[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_6;
      end else if (8'h44 == _T_31[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_5;
      end else if (8'h44 == _T_28[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_4;
      end else if (8'h44 == _T_25[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_3;
      end else if (8'h44 == _T_22[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_2;
      end else if (8'h44 == _T_19[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_1;
      end else if (8'h44 == _T_15[7:0]) begin
        image_2_68 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_69 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h45 == _T_34[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_6;
      end else if (8'h45 == _T_31[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_5;
      end else if (8'h45 == _T_28[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_4;
      end else if (8'h45 == _T_25[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_3;
      end else if (8'h45 == _T_22[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_2;
      end else if (8'h45 == _T_19[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_1;
      end else if (8'h45 == _T_15[7:0]) begin
        image_2_69 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_70 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h46 == _T_34[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_6;
      end else if (8'h46 == _T_31[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_5;
      end else if (8'h46 == _T_28[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_4;
      end else if (8'h46 == _T_25[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_3;
      end else if (8'h46 == _T_22[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_2;
      end else if (8'h46 == _T_19[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_1;
      end else if (8'h46 == _T_15[7:0]) begin
        image_2_70 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_71 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h47 == _T_34[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_6;
      end else if (8'h47 == _T_31[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_5;
      end else if (8'h47 == _T_28[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_4;
      end else if (8'h47 == _T_25[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_3;
      end else if (8'h47 == _T_22[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_2;
      end else if (8'h47 == _T_19[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_1;
      end else if (8'h47 == _T_15[7:0]) begin
        image_2_71 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_72 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h48 == _T_34[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_6;
      end else if (8'h48 == _T_31[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_5;
      end else if (8'h48 == _T_28[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_4;
      end else if (8'h48 == _T_25[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_3;
      end else if (8'h48 == _T_22[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_2;
      end else if (8'h48 == _T_19[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_1;
      end else if (8'h48 == _T_15[7:0]) begin
        image_2_72 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_73 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h49 == _T_34[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_6;
      end else if (8'h49 == _T_31[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_5;
      end else if (8'h49 == _T_28[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_4;
      end else if (8'h49 == _T_25[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_3;
      end else if (8'h49 == _T_22[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_2;
      end else if (8'h49 == _T_19[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_1;
      end else if (8'h49 == _T_15[7:0]) begin
        image_2_73 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_74 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4a == _T_34[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_6;
      end else if (8'h4a == _T_31[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_5;
      end else if (8'h4a == _T_28[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_4;
      end else if (8'h4a == _T_25[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_3;
      end else if (8'h4a == _T_22[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_2;
      end else if (8'h4a == _T_19[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_1;
      end else if (8'h4a == _T_15[7:0]) begin
        image_2_74 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_75 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4b == _T_34[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_6;
      end else if (8'h4b == _T_31[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_5;
      end else if (8'h4b == _T_28[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_4;
      end else if (8'h4b == _T_25[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_3;
      end else if (8'h4b == _T_22[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_2;
      end else if (8'h4b == _T_19[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_1;
      end else if (8'h4b == _T_15[7:0]) begin
        image_2_75 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_76 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4c == _T_34[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_6;
      end else if (8'h4c == _T_31[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_5;
      end else if (8'h4c == _T_28[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_4;
      end else if (8'h4c == _T_25[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_3;
      end else if (8'h4c == _T_22[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_2;
      end else if (8'h4c == _T_19[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_1;
      end else if (8'h4c == _T_15[7:0]) begin
        image_2_76 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_77 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4d == _T_34[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_6;
      end else if (8'h4d == _T_31[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_5;
      end else if (8'h4d == _T_28[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_4;
      end else if (8'h4d == _T_25[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_3;
      end else if (8'h4d == _T_22[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_2;
      end else if (8'h4d == _T_19[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_1;
      end else if (8'h4d == _T_15[7:0]) begin
        image_2_77 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_78 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4e == _T_34[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_6;
      end else if (8'h4e == _T_31[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_5;
      end else if (8'h4e == _T_28[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_4;
      end else if (8'h4e == _T_25[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_3;
      end else if (8'h4e == _T_22[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_2;
      end else if (8'h4e == _T_19[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_1;
      end else if (8'h4e == _T_15[7:0]) begin
        image_2_78 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_79 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h4f == _T_34[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_6;
      end else if (8'h4f == _T_31[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_5;
      end else if (8'h4f == _T_28[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_4;
      end else if (8'h4f == _T_25[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_3;
      end else if (8'h4f == _T_22[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_2;
      end else if (8'h4f == _T_19[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_1;
      end else if (8'h4f == _T_15[7:0]) begin
        image_2_79 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_80 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h50 == _T_34[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_6;
      end else if (8'h50 == _T_31[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_5;
      end else if (8'h50 == _T_28[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_4;
      end else if (8'h50 == _T_25[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_3;
      end else if (8'h50 == _T_22[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_2;
      end else if (8'h50 == _T_19[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_1;
      end else if (8'h50 == _T_15[7:0]) begin
        image_2_80 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_81 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h51 == _T_34[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_6;
      end else if (8'h51 == _T_31[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_5;
      end else if (8'h51 == _T_28[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_4;
      end else if (8'h51 == _T_25[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_3;
      end else if (8'h51 == _T_22[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_2;
      end else if (8'h51 == _T_19[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_1;
      end else if (8'h51 == _T_15[7:0]) begin
        image_2_81 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_82 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h52 == _T_34[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_6;
      end else if (8'h52 == _T_31[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_5;
      end else if (8'h52 == _T_28[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_4;
      end else if (8'h52 == _T_25[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_3;
      end else if (8'h52 == _T_22[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_2;
      end else if (8'h52 == _T_19[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_1;
      end else if (8'h52 == _T_15[7:0]) begin
        image_2_82 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_83 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h53 == _T_34[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_6;
      end else if (8'h53 == _T_31[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_5;
      end else if (8'h53 == _T_28[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_4;
      end else if (8'h53 == _T_25[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_3;
      end else if (8'h53 == _T_22[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_2;
      end else if (8'h53 == _T_19[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_1;
      end else if (8'h53 == _T_15[7:0]) begin
        image_2_83 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_84 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h54 == _T_34[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_6;
      end else if (8'h54 == _T_31[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_5;
      end else if (8'h54 == _T_28[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_4;
      end else if (8'h54 == _T_25[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_3;
      end else if (8'h54 == _T_22[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_2;
      end else if (8'h54 == _T_19[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_1;
      end else if (8'h54 == _T_15[7:0]) begin
        image_2_84 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_85 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h55 == _T_34[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_6;
      end else if (8'h55 == _T_31[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_5;
      end else if (8'h55 == _T_28[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_4;
      end else if (8'h55 == _T_25[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_3;
      end else if (8'h55 == _T_22[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_2;
      end else if (8'h55 == _T_19[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_1;
      end else if (8'h55 == _T_15[7:0]) begin
        image_2_85 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_86 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h56 == _T_34[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_6;
      end else if (8'h56 == _T_31[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_5;
      end else if (8'h56 == _T_28[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_4;
      end else if (8'h56 == _T_25[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_3;
      end else if (8'h56 == _T_22[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_2;
      end else if (8'h56 == _T_19[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_1;
      end else if (8'h56 == _T_15[7:0]) begin
        image_2_86 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_87 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h57 == _T_34[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_6;
      end else if (8'h57 == _T_31[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_5;
      end else if (8'h57 == _T_28[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_4;
      end else if (8'h57 == _T_25[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_3;
      end else if (8'h57 == _T_22[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_2;
      end else if (8'h57 == _T_19[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_1;
      end else if (8'h57 == _T_15[7:0]) begin
        image_2_87 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_88 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h58 == _T_34[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_6;
      end else if (8'h58 == _T_31[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_5;
      end else if (8'h58 == _T_28[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_4;
      end else if (8'h58 == _T_25[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_3;
      end else if (8'h58 == _T_22[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_2;
      end else if (8'h58 == _T_19[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_1;
      end else if (8'h58 == _T_15[7:0]) begin
        image_2_88 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_89 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h59 == _T_34[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_6;
      end else if (8'h59 == _T_31[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_5;
      end else if (8'h59 == _T_28[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_4;
      end else if (8'h59 == _T_25[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_3;
      end else if (8'h59 == _T_22[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_2;
      end else if (8'h59 == _T_19[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_1;
      end else if (8'h59 == _T_15[7:0]) begin
        image_2_89 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_90 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5a == _T_34[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_6;
      end else if (8'h5a == _T_31[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_5;
      end else if (8'h5a == _T_28[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_4;
      end else if (8'h5a == _T_25[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_3;
      end else if (8'h5a == _T_22[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_2;
      end else if (8'h5a == _T_19[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_1;
      end else if (8'h5a == _T_15[7:0]) begin
        image_2_90 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_91 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5b == _T_34[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_6;
      end else if (8'h5b == _T_31[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_5;
      end else if (8'h5b == _T_28[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_4;
      end else if (8'h5b == _T_25[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_3;
      end else if (8'h5b == _T_22[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_2;
      end else if (8'h5b == _T_19[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_1;
      end else if (8'h5b == _T_15[7:0]) begin
        image_2_91 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_92 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5c == _T_34[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_6;
      end else if (8'h5c == _T_31[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_5;
      end else if (8'h5c == _T_28[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_4;
      end else if (8'h5c == _T_25[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_3;
      end else if (8'h5c == _T_22[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_2;
      end else if (8'h5c == _T_19[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_1;
      end else if (8'h5c == _T_15[7:0]) begin
        image_2_92 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_93 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5d == _T_34[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_6;
      end else if (8'h5d == _T_31[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_5;
      end else if (8'h5d == _T_28[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_4;
      end else if (8'h5d == _T_25[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_3;
      end else if (8'h5d == _T_22[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_2;
      end else if (8'h5d == _T_19[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_1;
      end else if (8'h5d == _T_15[7:0]) begin
        image_2_93 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_94 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5e == _T_34[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_6;
      end else if (8'h5e == _T_31[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_5;
      end else if (8'h5e == _T_28[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_4;
      end else if (8'h5e == _T_25[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_3;
      end else if (8'h5e == _T_22[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_2;
      end else if (8'h5e == _T_19[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_1;
      end else if (8'h5e == _T_15[7:0]) begin
        image_2_94 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_95 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h5f == _T_34[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_6;
      end else if (8'h5f == _T_31[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_5;
      end else if (8'h5f == _T_28[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_4;
      end else if (8'h5f == _T_25[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_3;
      end else if (8'h5f == _T_22[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_2;
      end else if (8'h5f == _T_19[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_1;
      end else if (8'h5f == _T_15[7:0]) begin
        image_2_95 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_96 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h60 == _T_34[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_6;
      end else if (8'h60 == _T_31[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_5;
      end else if (8'h60 == _T_28[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_4;
      end else if (8'h60 == _T_25[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_3;
      end else if (8'h60 == _T_22[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_2;
      end else if (8'h60 == _T_19[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_1;
      end else if (8'h60 == _T_15[7:0]) begin
        image_2_96 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_97 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h61 == _T_34[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_6;
      end else if (8'h61 == _T_31[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_5;
      end else if (8'h61 == _T_28[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_4;
      end else if (8'h61 == _T_25[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_3;
      end else if (8'h61 == _T_22[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_2;
      end else if (8'h61 == _T_19[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_1;
      end else if (8'h61 == _T_15[7:0]) begin
        image_2_97 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_98 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h62 == _T_34[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_6;
      end else if (8'h62 == _T_31[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_5;
      end else if (8'h62 == _T_28[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_4;
      end else if (8'h62 == _T_25[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_3;
      end else if (8'h62 == _T_22[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_2;
      end else if (8'h62 == _T_19[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_1;
      end else if (8'h62 == _T_15[7:0]) begin
        image_2_98 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_99 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h63 == _T_34[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_6;
      end else if (8'h63 == _T_31[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_5;
      end else if (8'h63 == _T_28[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_4;
      end else if (8'h63 == _T_25[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_3;
      end else if (8'h63 == _T_22[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_2;
      end else if (8'h63 == _T_19[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_1;
      end else if (8'h63 == _T_15[7:0]) begin
        image_2_99 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_100 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h64 == _T_34[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_6;
      end else if (8'h64 == _T_31[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_5;
      end else if (8'h64 == _T_28[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_4;
      end else if (8'h64 == _T_25[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_3;
      end else if (8'h64 == _T_22[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_2;
      end else if (8'h64 == _T_19[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_1;
      end else if (8'h64 == _T_15[7:0]) begin
        image_2_100 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_101 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h65 == _T_34[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_6;
      end else if (8'h65 == _T_31[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_5;
      end else if (8'h65 == _T_28[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_4;
      end else if (8'h65 == _T_25[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_3;
      end else if (8'h65 == _T_22[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_2;
      end else if (8'h65 == _T_19[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_1;
      end else if (8'h65 == _T_15[7:0]) begin
        image_2_101 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_102 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h66 == _T_34[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_6;
      end else if (8'h66 == _T_31[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_5;
      end else if (8'h66 == _T_28[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_4;
      end else if (8'h66 == _T_25[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_3;
      end else if (8'h66 == _T_22[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_2;
      end else if (8'h66 == _T_19[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_1;
      end else if (8'h66 == _T_15[7:0]) begin
        image_2_102 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_103 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h67 == _T_34[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_6;
      end else if (8'h67 == _T_31[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_5;
      end else if (8'h67 == _T_28[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_4;
      end else if (8'h67 == _T_25[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_3;
      end else if (8'h67 == _T_22[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_2;
      end else if (8'h67 == _T_19[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_1;
      end else if (8'h67 == _T_15[7:0]) begin
        image_2_103 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_104 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h68 == _T_34[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_6;
      end else if (8'h68 == _T_31[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_5;
      end else if (8'h68 == _T_28[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_4;
      end else if (8'h68 == _T_25[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_3;
      end else if (8'h68 == _T_22[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_2;
      end else if (8'h68 == _T_19[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_1;
      end else if (8'h68 == _T_15[7:0]) begin
        image_2_104 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_105 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h69 == _T_34[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_6;
      end else if (8'h69 == _T_31[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_5;
      end else if (8'h69 == _T_28[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_4;
      end else if (8'h69 == _T_25[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_3;
      end else if (8'h69 == _T_22[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_2;
      end else if (8'h69 == _T_19[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_1;
      end else if (8'h69 == _T_15[7:0]) begin
        image_2_105 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_106 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6a == _T_34[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_6;
      end else if (8'h6a == _T_31[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_5;
      end else if (8'h6a == _T_28[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_4;
      end else if (8'h6a == _T_25[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_3;
      end else if (8'h6a == _T_22[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_2;
      end else if (8'h6a == _T_19[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_1;
      end else if (8'h6a == _T_15[7:0]) begin
        image_2_106 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_107 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6b == _T_34[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_6;
      end else if (8'h6b == _T_31[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_5;
      end else if (8'h6b == _T_28[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_4;
      end else if (8'h6b == _T_25[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_3;
      end else if (8'h6b == _T_22[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_2;
      end else if (8'h6b == _T_19[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_1;
      end else if (8'h6b == _T_15[7:0]) begin
        image_2_107 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_108 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6c == _T_34[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_6;
      end else if (8'h6c == _T_31[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_5;
      end else if (8'h6c == _T_28[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_4;
      end else if (8'h6c == _T_25[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_3;
      end else if (8'h6c == _T_22[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_2;
      end else if (8'h6c == _T_19[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_1;
      end else if (8'h6c == _T_15[7:0]) begin
        image_2_108 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_109 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6d == _T_34[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_6;
      end else if (8'h6d == _T_31[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_5;
      end else if (8'h6d == _T_28[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_4;
      end else if (8'h6d == _T_25[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_3;
      end else if (8'h6d == _T_22[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_2;
      end else if (8'h6d == _T_19[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_1;
      end else if (8'h6d == _T_15[7:0]) begin
        image_2_109 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_110 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6e == _T_34[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_6;
      end else if (8'h6e == _T_31[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_5;
      end else if (8'h6e == _T_28[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_4;
      end else if (8'h6e == _T_25[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_3;
      end else if (8'h6e == _T_22[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_2;
      end else if (8'h6e == _T_19[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_1;
      end else if (8'h6e == _T_15[7:0]) begin
        image_2_110 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_111 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h6f == _T_34[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_6;
      end else if (8'h6f == _T_31[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_5;
      end else if (8'h6f == _T_28[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_4;
      end else if (8'h6f == _T_25[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_3;
      end else if (8'h6f == _T_22[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_2;
      end else if (8'h6f == _T_19[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_1;
      end else if (8'h6f == _T_15[7:0]) begin
        image_2_111 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_112 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h70 == _T_34[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_6;
      end else if (8'h70 == _T_31[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_5;
      end else if (8'h70 == _T_28[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_4;
      end else if (8'h70 == _T_25[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_3;
      end else if (8'h70 == _T_22[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_2;
      end else if (8'h70 == _T_19[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_1;
      end else if (8'h70 == _T_15[7:0]) begin
        image_2_112 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_113 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h71 == _T_34[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_6;
      end else if (8'h71 == _T_31[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_5;
      end else if (8'h71 == _T_28[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_4;
      end else if (8'h71 == _T_25[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_3;
      end else if (8'h71 == _T_22[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_2;
      end else if (8'h71 == _T_19[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_1;
      end else if (8'h71 == _T_15[7:0]) begin
        image_2_113 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_114 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h72 == _T_34[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_6;
      end else if (8'h72 == _T_31[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_5;
      end else if (8'h72 == _T_28[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_4;
      end else if (8'h72 == _T_25[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_3;
      end else if (8'h72 == _T_22[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_2;
      end else if (8'h72 == _T_19[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_1;
      end else if (8'h72 == _T_15[7:0]) begin
        image_2_114 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_115 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h73 == _T_34[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_6;
      end else if (8'h73 == _T_31[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_5;
      end else if (8'h73 == _T_28[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_4;
      end else if (8'h73 == _T_25[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_3;
      end else if (8'h73 == _T_22[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_2;
      end else if (8'h73 == _T_19[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_1;
      end else if (8'h73 == _T_15[7:0]) begin
        image_2_115 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_116 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h74 == _T_34[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_6;
      end else if (8'h74 == _T_31[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_5;
      end else if (8'h74 == _T_28[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_4;
      end else if (8'h74 == _T_25[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_3;
      end else if (8'h74 == _T_22[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_2;
      end else if (8'h74 == _T_19[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_1;
      end else if (8'h74 == _T_15[7:0]) begin
        image_2_116 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_117 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h75 == _T_34[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_6;
      end else if (8'h75 == _T_31[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_5;
      end else if (8'h75 == _T_28[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_4;
      end else if (8'h75 == _T_25[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_3;
      end else if (8'h75 == _T_22[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_2;
      end else if (8'h75 == _T_19[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_1;
      end else if (8'h75 == _T_15[7:0]) begin
        image_2_117 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_118 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h76 == _T_34[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_6;
      end else if (8'h76 == _T_31[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_5;
      end else if (8'h76 == _T_28[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_4;
      end else if (8'h76 == _T_25[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_3;
      end else if (8'h76 == _T_22[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_2;
      end else if (8'h76 == _T_19[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_1;
      end else if (8'h76 == _T_15[7:0]) begin
        image_2_118 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_119 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h77 == _T_34[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_6;
      end else if (8'h77 == _T_31[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_5;
      end else if (8'h77 == _T_28[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_4;
      end else if (8'h77 == _T_25[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_3;
      end else if (8'h77 == _T_22[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_2;
      end else if (8'h77 == _T_19[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_1;
      end else if (8'h77 == _T_15[7:0]) begin
        image_2_119 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_120 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h78 == _T_34[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_6;
      end else if (8'h78 == _T_31[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_5;
      end else if (8'h78 == _T_28[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_4;
      end else if (8'h78 == _T_25[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_3;
      end else if (8'h78 == _T_22[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_2;
      end else if (8'h78 == _T_19[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_1;
      end else if (8'h78 == _T_15[7:0]) begin
        image_2_120 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_121 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h79 == _T_34[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_6;
      end else if (8'h79 == _T_31[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_5;
      end else if (8'h79 == _T_28[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_4;
      end else if (8'h79 == _T_25[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_3;
      end else if (8'h79 == _T_22[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_2;
      end else if (8'h79 == _T_19[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_1;
      end else if (8'h79 == _T_15[7:0]) begin
        image_2_121 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_122 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7a == _T_34[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_6;
      end else if (8'h7a == _T_31[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_5;
      end else if (8'h7a == _T_28[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_4;
      end else if (8'h7a == _T_25[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_3;
      end else if (8'h7a == _T_22[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_2;
      end else if (8'h7a == _T_19[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_1;
      end else if (8'h7a == _T_15[7:0]) begin
        image_2_122 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_123 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7b == _T_34[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_6;
      end else if (8'h7b == _T_31[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_5;
      end else if (8'h7b == _T_28[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_4;
      end else if (8'h7b == _T_25[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_3;
      end else if (8'h7b == _T_22[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_2;
      end else if (8'h7b == _T_19[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_1;
      end else if (8'h7b == _T_15[7:0]) begin
        image_2_123 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_124 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7c == _T_34[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_6;
      end else if (8'h7c == _T_31[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_5;
      end else if (8'h7c == _T_28[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_4;
      end else if (8'h7c == _T_25[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_3;
      end else if (8'h7c == _T_22[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_2;
      end else if (8'h7c == _T_19[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_1;
      end else if (8'h7c == _T_15[7:0]) begin
        image_2_124 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_125 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7d == _T_34[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_6;
      end else if (8'h7d == _T_31[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_5;
      end else if (8'h7d == _T_28[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_4;
      end else if (8'h7d == _T_25[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_3;
      end else if (8'h7d == _T_22[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_2;
      end else if (8'h7d == _T_19[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_1;
      end else if (8'h7d == _T_15[7:0]) begin
        image_2_125 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_126 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7e == _T_34[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_6;
      end else if (8'h7e == _T_31[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_5;
      end else if (8'h7e == _T_28[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_4;
      end else if (8'h7e == _T_25[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_3;
      end else if (8'h7e == _T_22[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_2;
      end else if (8'h7e == _T_19[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_1;
      end else if (8'h7e == _T_15[7:0]) begin
        image_2_126 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_127 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h7f == _T_34[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_6;
      end else if (8'h7f == _T_31[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_5;
      end else if (8'h7f == _T_28[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_4;
      end else if (8'h7f == _T_25[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_3;
      end else if (8'h7f == _T_22[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_2;
      end else if (8'h7f == _T_19[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_1;
      end else if (8'h7f == _T_15[7:0]) begin
        image_2_127 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_128 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h80 == _T_34[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_6;
      end else if (8'h80 == _T_31[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_5;
      end else if (8'h80 == _T_28[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_4;
      end else if (8'h80 == _T_25[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_3;
      end else if (8'h80 == _T_22[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_2;
      end else if (8'h80 == _T_19[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_1;
      end else if (8'h80 == _T_15[7:0]) begin
        image_2_128 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_129 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h81 == _T_34[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_6;
      end else if (8'h81 == _T_31[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_5;
      end else if (8'h81 == _T_28[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_4;
      end else if (8'h81 == _T_25[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_3;
      end else if (8'h81 == _T_22[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_2;
      end else if (8'h81 == _T_19[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_1;
      end else if (8'h81 == _T_15[7:0]) begin
        image_2_129 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_130 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h82 == _T_34[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_6;
      end else if (8'h82 == _T_31[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_5;
      end else if (8'h82 == _T_28[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_4;
      end else if (8'h82 == _T_25[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_3;
      end else if (8'h82 == _T_22[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_2;
      end else if (8'h82 == _T_19[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_1;
      end else if (8'h82 == _T_15[7:0]) begin
        image_2_130 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_131 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h83 == _T_34[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_6;
      end else if (8'h83 == _T_31[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_5;
      end else if (8'h83 == _T_28[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_4;
      end else if (8'h83 == _T_25[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_3;
      end else if (8'h83 == _T_22[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_2;
      end else if (8'h83 == _T_19[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_1;
      end else if (8'h83 == _T_15[7:0]) begin
        image_2_131 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_132 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h84 == _T_34[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_6;
      end else if (8'h84 == _T_31[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_5;
      end else if (8'h84 == _T_28[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_4;
      end else if (8'h84 == _T_25[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_3;
      end else if (8'h84 == _T_22[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_2;
      end else if (8'h84 == _T_19[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_1;
      end else if (8'h84 == _T_15[7:0]) begin
        image_2_132 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_133 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h85 == _T_34[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_6;
      end else if (8'h85 == _T_31[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_5;
      end else if (8'h85 == _T_28[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_4;
      end else if (8'h85 == _T_25[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_3;
      end else if (8'h85 == _T_22[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_2;
      end else if (8'h85 == _T_19[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_1;
      end else if (8'h85 == _T_15[7:0]) begin
        image_2_133 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_134 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h86 == _T_34[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_6;
      end else if (8'h86 == _T_31[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_5;
      end else if (8'h86 == _T_28[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_4;
      end else if (8'h86 == _T_25[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_3;
      end else if (8'h86 == _T_22[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_2;
      end else if (8'h86 == _T_19[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_1;
      end else if (8'h86 == _T_15[7:0]) begin
        image_2_134 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_135 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h87 == _T_34[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_6;
      end else if (8'h87 == _T_31[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_5;
      end else if (8'h87 == _T_28[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_4;
      end else if (8'h87 == _T_25[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_3;
      end else if (8'h87 == _T_22[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_2;
      end else if (8'h87 == _T_19[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_1;
      end else if (8'h87 == _T_15[7:0]) begin
        image_2_135 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_136 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h88 == _T_34[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_6;
      end else if (8'h88 == _T_31[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_5;
      end else if (8'h88 == _T_28[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_4;
      end else if (8'h88 == _T_25[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_3;
      end else if (8'h88 == _T_22[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_2;
      end else if (8'h88 == _T_19[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_1;
      end else if (8'h88 == _T_15[7:0]) begin
        image_2_136 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_137 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h89 == _T_34[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_6;
      end else if (8'h89 == _T_31[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_5;
      end else if (8'h89 == _T_28[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_4;
      end else if (8'h89 == _T_25[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_3;
      end else if (8'h89 == _T_22[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_2;
      end else if (8'h89 == _T_19[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_1;
      end else if (8'h89 == _T_15[7:0]) begin
        image_2_137 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_138 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8a == _T_34[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_6;
      end else if (8'h8a == _T_31[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_5;
      end else if (8'h8a == _T_28[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_4;
      end else if (8'h8a == _T_25[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_3;
      end else if (8'h8a == _T_22[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_2;
      end else if (8'h8a == _T_19[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_1;
      end else if (8'h8a == _T_15[7:0]) begin
        image_2_138 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_139 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8b == _T_34[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_6;
      end else if (8'h8b == _T_31[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_5;
      end else if (8'h8b == _T_28[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_4;
      end else if (8'h8b == _T_25[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_3;
      end else if (8'h8b == _T_22[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_2;
      end else if (8'h8b == _T_19[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_1;
      end else if (8'h8b == _T_15[7:0]) begin
        image_2_139 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_140 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8c == _T_34[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_6;
      end else if (8'h8c == _T_31[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_5;
      end else if (8'h8c == _T_28[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_4;
      end else if (8'h8c == _T_25[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_3;
      end else if (8'h8c == _T_22[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_2;
      end else if (8'h8c == _T_19[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_1;
      end else if (8'h8c == _T_15[7:0]) begin
        image_2_140 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_141 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8d == _T_34[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_6;
      end else if (8'h8d == _T_31[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_5;
      end else if (8'h8d == _T_28[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_4;
      end else if (8'h8d == _T_25[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_3;
      end else if (8'h8d == _T_22[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_2;
      end else if (8'h8d == _T_19[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_1;
      end else if (8'h8d == _T_15[7:0]) begin
        image_2_141 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_142 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8e == _T_34[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_6;
      end else if (8'h8e == _T_31[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_5;
      end else if (8'h8e == _T_28[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_4;
      end else if (8'h8e == _T_25[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_3;
      end else if (8'h8e == _T_22[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_2;
      end else if (8'h8e == _T_19[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_1;
      end else if (8'h8e == _T_15[7:0]) begin
        image_2_142 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_143 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h8f == _T_34[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_6;
      end else if (8'h8f == _T_31[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_5;
      end else if (8'h8f == _T_28[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_4;
      end else if (8'h8f == _T_25[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_3;
      end else if (8'h8f == _T_22[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_2;
      end else if (8'h8f == _T_19[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_1;
      end else if (8'h8f == _T_15[7:0]) begin
        image_2_143 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_144 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h90 == _T_34[7:0]) begin
        image_2_144 <= io_pixelVal_in_2_6;
      end else if (8'h90 == _T_31[7:0]) begin
        image_2_144 <= io_pixelVal_in_2_5;
      end else if (8'h90 == _T_28[7:0]) begin
        image_2_144 <= io_pixelVal_in_2_4;
      end else if (8'h90 == _T_25[7:0]) begin
        image_2_144 <= io_pixelVal_in_2_3;
      end else if (8'h90 == _T_22[7:0]) begin
        image_2_144 <= io_pixelVal_in_2_2;
      end else if (8'h90 == _T_19[7:0]) begin
        image_2_144 <= io_pixelVal_in_2_1;
      end else if (8'h90 == _T_15[7:0]) begin
        image_2_144 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_145 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h91 == _T_34[7:0]) begin
        image_2_145 <= io_pixelVal_in_2_6;
      end else if (8'h91 == _T_31[7:0]) begin
        image_2_145 <= io_pixelVal_in_2_5;
      end else if (8'h91 == _T_28[7:0]) begin
        image_2_145 <= io_pixelVal_in_2_4;
      end else if (8'h91 == _T_25[7:0]) begin
        image_2_145 <= io_pixelVal_in_2_3;
      end else if (8'h91 == _T_22[7:0]) begin
        image_2_145 <= io_pixelVal_in_2_2;
      end else if (8'h91 == _T_19[7:0]) begin
        image_2_145 <= io_pixelVal_in_2_1;
      end else if (8'h91 == _T_15[7:0]) begin
        image_2_145 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_146 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h92 == _T_34[7:0]) begin
        image_2_146 <= io_pixelVal_in_2_6;
      end else if (8'h92 == _T_31[7:0]) begin
        image_2_146 <= io_pixelVal_in_2_5;
      end else if (8'h92 == _T_28[7:0]) begin
        image_2_146 <= io_pixelVal_in_2_4;
      end else if (8'h92 == _T_25[7:0]) begin
        image_2_146 <= io_pixelVal_in_2_3;
      end else if (8'h92 == _T_22[7:0]) begin
        image_2_146 <= io_pixelVal_in_2_2;
      end else if (8'h92 == _T_19[7:0]) begin
        image_2_146 <= io_pixelVal_in_2_1;
      end else if (8'h92 == _T_15[7:0]) begin
        image_2_146 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_147 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h93 == _T_34[7:0]) begin
        image_2_147 <= io_pixelVal_in_2_6;
      end else if (8'h93 == _T_31[7:0]) begin
        image_2_147 <= io_pixelVal_in_2_5;
      end else if (8'h93 == _T_28[7:0]) begin
        image_2_147 <= io_pixelVal_in_2_4;
      end else if (8'h93 == _T_25[7:0]) begin
        image_2_147 <= io_pixelVal_in_2_3;
      end else if (8'h93 == _T_22[7:0]) begin
        image_2_147 <= io_pixelVal_in_2_2;
      end else if (8'h93 == _T_19[7:0]) begin
        image_2_147 <= io_pixelVal_in_2_1;
      end else if (8'h93 == _T_15[7:0]) begin
        image_2_147 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_148 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h94 == _T_34[7:0]) begin
        image_2_148 <= io_pixelVal_in_2_6;
      end else if (8'h94 == _T_31[7:0]) begin
        image_2_148 <= io_pixelVal_in_2_5;
      end else if (8'h94 == _T_28[7:0]) begin
        image_2_148 <= io_pixelVal_in_2_4;
      end else if (8'h94 == _T_25[7:0]) begin
        image_2_148 <= io_pixelVal_in_2_3;
      end else if (8'h94 == _T_22[7:0]) begin
        image_2_148 <= io_pixelVal_in_2_2;
      end else if (8'h94 == _T_19[7:0]) begin
        image_2_148 <= io_pixelVal_in_2_1;
      end else if (8'h94 == _T_15[7:0]) begin
        image_2_148 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_149 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h95 == _T_34[7:0]) begin
        image_2_149 <= io_pixelVal_in_2_6;
      end else if (8'h95 == _T_31[7:0]) begin
        image_2_149 <= io_pixelVal_in_2_5;
      end else if (8'h95 == _T_28[7:0]) begin
        image_2_149 <= io_pixelVal_in_2_4;
      end else if (8'h95 == _T_25[7:0]) begin
        image_2_149 <= io_pixelVal_in_2_3;
      end else if (8'h95 == _T_22[7:0]) begin
        image_2_149 <= io_pixelVal_in_2_2;
      end else if (8'h95 == _T_19[7:0]) begin
        image_2_149 <= io_pixelVal_in_2_1;
      end else if (8'h95 == _T_15[7:0]) begin
        image_2_149 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_150 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h96 == _T_34[7:0]) begin
        image_2_150 <= io_pixelVal_in_2_6;
      end else if (8'h96 == _T_31[7:0]) begin
        image_2_150 <= io_pixelVal_in_2_5;
      end else if (8'h96 == _T_28[7:0]) begin
        image_2_150 <= io_pixelVal_in_2_4;
      end else if (8'h96 == _T_25[7:0]) begin
        image_2_150 <= io_pixelVal_in_2_3;
      end else if (8'h96 == _T_22[7:0]) begin
        image_2_150 <= io_pixelVal_in_2_2;
      end else if (8'h96 == _T_19[7:0]) begin
        image_2_150 <= io_pixelVal_in_2_1;
      end else if (8'h96 == _T_15[7:0]) begin
        image_2_150 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_151 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h97 == _T_34[7:0]) begin
        image_2_151 <= io_pixelVal_in_2_6;
      end else if (8'h97 == _T_31[7:0]) begin
        image_2_151 <= io_pixelVal_in_2_5;
      end else if (8'h97 == _T_28[7:0]) begin
        image_2_151 <= io_pixelVal_in_2_4;
      end else if (8'h97 == _T_25[7:0]) begin
        image_2_151 <= io_pixelVal_in_2_3;
      end else if (8'h97 == _T_22[7:0]) begin
        image_2_151 <= io_pixelVal_in_2_2;
      end else if (8'h97 == _T_19[7:0]) begin
        image_2_151 <= io_pixelVal_in_2_1;
      end else if (8'h97 == _T_15[7:0]) begin
        image_2_151 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_152 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h98 == _T_34[7:0]) begin
        image_2_152 <= io_pixelVal_in_2_6;
      end else if (8'h98 == _T_31[7:0]) begin
        image_2_152 <= io_pixelVal_in_2_5;
      end else if (8'h98 == _T_28[7:0]) begin
        image_2_152 <= io_pixelVal_in_2_4;
      end else if (8'h98 == _T_25[7:0]) begin
        image_2_152 <= io_pixelVal_in_2_3;
      end else if (8'h98 == _T_22[7:0]) begin
        image_2_152 <= io_pixelVal_in_2_2;
      end else if (8'h98 == _T_19[7:0]) begin
        image_2_152 <= io_pixelVal_in_2_1;
      end else if (8'h98 == _T_15[7:0]) begin
        image_2_152 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_153 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h99 == _T_34[7:0]) begin
        image_2_153 <= io_pixelVal_in_2_6;
      end else if (8'h99 == _T_31[7:0]) begin
        image_2_153 <= io_pixelVal_in_2_5;
      end else if (8'h99 == _T_28[7:0]) begin
        image_2_153 <= io_pixelVal_in_2_4;
      end else if (8'h99 == _T_25[7:0]) begin
        image_2_153 <= io_pixelVal_in_2_3;
      end else if (8'h99 == _T_22[7:0]) begin
        image_2_153 <= io_pixelVal_in_2_2;
      end else if (8'h99 == _T_19[7:0]) begin
        image_2_153 <= io_pixelVal_in_2_1;
      end else if (8'h99 == _T_15[7:0]) begin
        image_2_153 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_154 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9a == _T_34[7:0]) begin
        image_2_154 <= io_pixelVal_in_2_6;
      end else if (8'h9a == _T_31[7:0]) begin
        image_2_154 <= io_pixelVal_in_2_5;
      end else if (8'h9a == _T_28[7:0]) begin
        image_2_154 <= io_pixelVal_in_2_4;
      end else if (8'h9a == _T_25[7:0]) begin
        image_2_154 <= io_pixelVal_in_2_3;
      end else if (8'h9a == _T_22[7:0]) begin
        image_2_154 <= io_pixelVal_in_2_2;
      end else if (8'h9a == _T_19[7:0]) begin
        image_2_154 <= io_pixelVal_in_2_1;
      end else if (8'h9a == _T_15[7:0]) begin
        image_2_154 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_155 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9b == _T_34[7:0]) begin
        image_2_155 <= io_pixelVal_in_2_6;
      end else if (8'h9b == _T_31[7:0]) begin
        image_2_155 <= io_pixelVal_in_2_5;
      end else if (8'h9b == _T_28[7:0]) begin
        image_2_155 <= io_pixelVal_in_2_4;
      end else if (8'h9b == _T_25[7:0]) begin
        image_2_155 <= io_pixelVal_in_2_3;
      end else if (8'h9b == _T_22[7:0]) begin
        image_2_155 <= io_pixelVal_in_2_2;
      end else if (8'h9b == _T_19[7:0]) begin
        image_2_155 <= io_pixelVal_in_2_1;
      end else if (8'h9b == _T_15[7:0]) begin
        image_2_155 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_156 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9c == _T_34[7:0]) begin
        image_2_156 <= io_pixelVal_in_2_6;
      end else if (8'h9c == _T_31[7:0]) begin
        image_2_156 <= io_pixelVal_in_2_5;
      end else if (8'h9c == _T_28[7:0]) begin
        image_2_156 <= io_pixelVal_in_2_4;
      end else if (8'h9c == _T_25[7:0]) begin
        image_2_156 <= io_pixelVal_in_2_3;
      end else if (8'h9c == _T_22[7:0]) begin
        image_2_156 <= io_pixelVal_in_2_2;
      end else if (8'h9c == _T_19[7:0]) begin
        image_2_156 <= io_pixelVal_in_2_1;
      end else if (8'h9c == _T_15[7:0]) begin
        image_2_156 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_157 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9d == _T_34[7:0]) begin
        image_2_157 <= io_pixelVal_in_2_6;
      end else if (8'h9d == _T_31[7:0]) begin
        image_2_157 <= io_pixelVal_in_2_5;
      end else if (8'h9d == _T_28[7:0]) begin
        image_2_157 <= io_pixelVal_in_2_4;
      end else if (8'h9d == _T_25[7:0]) begin
        image_2_157 <= io_pixelVal_in_2_3;
      end else if (8'h9d == _T_22[7:0]) begin
        image_2_157 <= io_pixelVal_in_2_2;
      end else if (8'h9d == _T_19[7:0]) begin
        image_2_157 <= io_pixelVal_in_2_1;
      end else if (8'h9d == _T_15[7:0]) begin
        image_2_157 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_158 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9e == _T_34[7:0]) begin
        image_2_158 <= io_pixelVal_in_2_6;
      end else if (8'h9e == _T_31[7:0]) begin
        image_2_158 <= io_pixelVal_in_2_5;
      end else if (8'h9e == _T_28[7:0]) begin
        image_2_158 <= io_pixelVal_in_2_4;
      end else if (8'h9e == _T_25[7:0]) begin
        image_2_158 <= io_pixelVal_in_2_3;
      end else if (8'h9e == _T_22[7:0]) begin
        image_2_158 <= io_pixelVal_in_2_2;
      end else if (8'h9e == _T_19[7:0]) begin
        image_2_158 <= io_pixelVal_in_2_1;
      end else if (8'h9e == _T_15[7:0]) begin
        image_2_158 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_159 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'h9f == _T_34[7:0]) begin
        image_2_159 <= io_pixelVal_in_2_6;
      end else if (8'h9f == _T_31[7:0]) begin
        image_2_159 <= io_pixelVal_in_2_5;
      end else if (8'h9f == _T_28[7:0]) begin
        image_2_159 <= io_pixelVal_in_2_4;
      end else if (8'h9f == _T_25[7:0]) begin
        image_2_159 <= io_pixelVal_in_2_3;
      end else if (8'h9f == _T_22[7:0]) begin
        image_2_159 <= io_pixelVal_in_2_2;
      end else if (8'h9f == _T_19[7:0]) begin
        image_2_159 <= io_pixelVal_in_2_1;
      end else if (8'h9f == _T_15[7:0]) begin
        image_2_159 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_160 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha0 == _T_34[7:0]) begin
        image_2_160 <= io_pixelVal_in_2_6;
      end else if (8'ha0 == _T_31[7:0]) begin
        image_2_160 <= io_pixelVal_in_2_5;
      end else if (8'ha0 == _T_28[7:0]) begin
        image_2_160 <= io_pixelVal_in_2_4;
      end else if (8'ha0 == _T_25[7:0]) begin
        image_2_160 <= io_pixelVal_in_2_3;
      end else if (8'ha0 == _T_22[7:0]) begin
        image_2_160 <= io_pixelVal_in_2_2;
      end else if (8'ha0 == _T_19[7:0]) begin
        image_2_160 <= io_pixelVal_in_2_1;
      end else if (8'ha0 == _T_15[7:0]) begin
        image_2_160 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_161 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha1 == _T_34[7:0]) begin
        image_2_161 <= io_pixelVal_in_2_6;
      end else if (8'ha1 == _T_31[7:0]) begin
        image_2_161 <= io_pixelVal_in_2_5;
      end else if (8'ha1 == _T_28[7:0]) begin
        image_2_161 <= io_pixelVal_in_2_4;
      end else if (8'ha1 == _T_25[7:0]) begin
        image_2_161 <= io_pixelVal_in_2_3;
      end else if (8'ha1 == _T_22[7:0]) begin
        image_2_161 <= io_pixelVal_in_2_2;
      end else if (8'ha1 == _T_19[7:0]) begin
        image_2_161 <= io_pixelVal_in_2_1;
      end else if (8'ha1 == _T_15[7:0]) begin
        image_2_161 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_162 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha2 == _T_34[7:0]) begin
        image_2_162 <= io_pixelVal_in_2_6;
      end else if (8'ha2 == _T_31[7:0]) begin
        image_2_162 <= io_pixelVal_in_2_5;
      end else if (8'ha2 == _T_28[7:0]) begin
        image_2_162 <= io_pixelVal_in_2_4;
      end else if (8'ha2 == _T_25[7:0]) begin
        image_2_162 <= io_pixelVal_in_2_3;
      end else if (8'ha2 == _T_22[7:0]) begin
        image_2_162 <= io_pixelVal_in_2_2;
      end else if (8'ha2 == _T_19[7:0]) begin
        image_2_162 <= io_pixelVal_in_2_1;
      end else if (8'ha2 == _T_15[7:0]) begin
        image_2_162 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_163 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha3 == _T_34[7:0]) begin
        image_2_163 <= io_pixelVal_in_2_6;
      end else if (8'ha3 == _T_31[7:0]) begin
        image_2_163 <= io_pixelVal_in_2_5;
      end else if (8'ha3 == _T_28[7:0]) begin
        image_2_163 <= io_pixelVal_in_2_4;
      end else if (8'ha3 == _T_25[7:0]) begin
        image_2_163 <= io_pixelVal_in_2_3;
      end else if (8'ha3 == _T_22[7:0]) begin
        image_2_163 <= io_pixelVal_in_2_2;
      end else if (8'ha3 == _T_19[7:0]) begin
        image_2_163 <= io_pixelVal_in_2_1;
      end else if (8'ha3 == _T_15[7:0]) begin
        image_2_163 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_164 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha4 == _T_34[7:0]) begin
        image_2_164 <= io_pixelVal_in_2_6;
      end else if (8'ha4 == _T_31[7:0]) begin
        image_2_164 <= io_pixelVal_in_2_5;
      end else if (8'ha4 == _T_28[7:0]) begin
        image_2_164 <= io_pixelVal_in_2_4;
      end else if (8'ha4 == _T_25[7:0]) begin
        image_2_164 <= io_pixelVal_in_2_3;
      end else if (8'ha4 == _T_22[7:0]) begin
        image_2_164 <= io_pixelVal_in_2_2;
      end else if (8'ha4 == _T_19[7:0]) begin
        image_2_164 <= io_pixelVal_in_2_1;
      end else if (8'ha4 == _T_15[7:0]) begin
        image_2_164 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_165 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha5 == _T_34[7:0]) begin
        image_2_165 <= io_pixelVal_in_2_6;
      end else if (8'ha5 == _T_31[7:0]) begin
        image_2_165 <= io_pixelVal_in_2_5;
      end else if (8'ha5 == _T_28[7:0]) begin
        image_2_165 <= io_pixelVal_in_2_4;
      end else if (8'ha5 == _T_25[7:0]) begin
        image_2_165 <= io_pixelVal_in_2_3;
      end else if (8'ha5 == _T_22[7:0]) begin
        image_2_165 <= io_pixelVal_in_2_2;
      end else if (8'ha5 == _T_19[7:0]) begin
        image_2_165 <= io_pixelVal_in_2_1;
      end else if (8'ha5 == _T_15[7:0]) begin
        image_2_165 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_166 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha6 == _T_34[7:0]) begin
        image_2_166 <= io_pixelVal_in_2_6;
      end else if (8'ha6 == _T_31[7:0]) begin
        image_2_166 <= io_pixelVal_in_2_5;
      end else if (8'ha6 == _T_28[7:0]) begin
        image_2_166 <= io_pixelVal_in_2_4;
      end else if (8'ha6 == _T_25[7:0]) begin
        image_2_166 <= io_pixelVal_in_2_3;
      end else if (8'ha6 == _T_22[7:0]) begin
        image_2_166 <= io_pixelVal_in_2_2;
      end else if (8'ha6 == _T_19[7:0]) begin
        image_2_166 <= io_pixelVal_in_2_1;
      end else if (8'ha6 == _T_15[7:0]) begin
        image_2_166 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_167 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha7 == _T_34[7:0]) begin
        image_2_167 <= io_pixelVal_in_2_6;
      end else if (8'ha7 == _T_31[7:0]) begin
        image_2_167 <= io_pixelVal_in_2_5;
      end else if (8'ha7 == _T_28[7:0]) begin
        image_2_167 <= io_pixelVal_in_2_4;
      end else if (8'ha7 == _T_25[7:0]) begin
        image_2_167 <= io_pixelVal_in_2_3;
      end else if (8'ha7 == _T_22[7:0]) begin
        image_2_167 <= io_pixelVal_in_2_2;
      end else if (8'ha7 == _T_19[7:0]) begin
        image_2_167 <= io_pixelVal_in_2_1;
      end else if (8'ha7 == _T_15[7:0]) begin
        image_2_167 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_168 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha8 == _T_34[7:0]) begin
        image_2_168 <= io_pixelVal_in_2_6;
      end else if (8'ha8 == _T_31[7:0]) begin
        image_2_168 <= io_pixelVal_in_2_5;
      end else if (8'ha8 == _T_28[7:0]) begin
        image_2_168 <= io_pixelVal_in_2_4;
      end else if (8'ha8 == _T_25[7:0]) begin
        image_2_168 <= io_pixelVal_in_2_3;
      end else if (8'ha8 == _T_22[7:0]) begin
        image_2_168 <= io_pixelVal_in_2_2;
      end else if (8'ha8 == _T_19[7:0]) begin
        image_2_168 <= io_pixelVal_in_2_1;
      end else if (8'ha8 == _T_15[7:0]) begin
        image_2_168 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_169 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'ha9 == _T_34[7:0]) begin
        image_2_169 <= io_pixelVal_in_2_6;
      end else if (8'ha9 == _T_31[7:0]) begin
        image_2_169 <= io_pixelVal_in_2_5;
      end else if (8'ha9 == _T_28[7:0]) begin
        image_2_169 <= io_pixelVal_in_2_4;
      end else if (8'ha9 == _T_25[7:0]) begin
        image_2_169 <= io_pixelVal_in_2_3;
      end else if (8'ha9 == _T_22[7:0]) begin
        image_2_169 <= io_pixelVal_in_2_2;
      end else if (8'ha9 == _T_19[7:0]) begin
        image_2_169 <= io_pixelVal_in_2_1;
      end else if (8'ha9 == _T_15[7:0]) begin
        image_2_169 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_170 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'haa == _T_34[7:0]) begin
        image_2_170 <= io_pixelVal_in_2_6;
      end else if (8'haa == _T_31[7:0]) begin
        image_2_170 <= io_pixelVal_in_2_5;
      end else if (8'haa == _T_28[7:0]) begin
        image_2_170 <= io_pixelVal_in_2_4;
      end else if (8'haa == _T_25[7:0]) begin
        image_2_170 <= io_pixelVal_in_2_3;
      end else if (8'haa == _T_22[7:0]) begin
        image_2_170 <= io_pixelVal_in_2_2;
      end else if (8'haa == _T_19[7:0]) begin
        image_2_170 <= io_pixelVal_in_2_1;
      end else if (8'haa == _T_15[7:0]) begin
        image_2_170 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_171 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hab == _T_34[7:0]) begin
        image_2_171 <= io_pixelVal_in_2_6;
      end else if (8'hab == _T_31[7:0]) begin
        image_2_171 <= io_pixelVal_in_2_5;
      end else if (8'hab == _T_28[7:0]) begin
        image_2_171 <= io_pixelVal_in_2_4;
      end else if (8'hab == _T_25[7:0]) begin
        image_2_171 <= io_pixelVal_in_2_3;
      end else if (8'hab == _T_22[7:0]) begin
        image_2_171 <= io_pixelVal_in_2_2;
      end else if (8'hab == _T_19[7:0]) begin
        image_2_171 <= io_pixelVal_in_2_1;
      end else if (8'hab == _T_15[7:0]) begin
        image_2_171 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_172 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hac == _T_34[7:0]) begin
        image_2_172 <= io_pixelVal_in_2_6;
      end else if (8'hac == _T_31[7:0]) begin
        image_2_172 <= io_pixelVal_in_2_5;
      end else if (8'hac == _T_28[7:0]) begin
        image_2_172 <= io_pixelVal_in_2_4;
      end else if (8'hac == _T_25[7:0]) begin
        image_2_172 <= io_pixelVal_in_2_3;
      end else if (8'hac == _T_22[7:0]) begin
        image_2_172 <= io_pixelVal_in_2_2;
      end else if (8'hac == _T_19[7:0]) begin
        image_2_172 <= io_pixelVal_in_2_1;
      end else if (8'hac == _T_15[7:0]) begin
        image_2_172 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_173 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'had == _T_34[7:0]) begin
        image_2_173 <= io_pixelVal_in_2_6;
      end else if (8'had == _T_31[7:0]) begin
        image_2_173 <= io_pixelVal_in_2_5;
      end else if (8'had == _T_28[7:0]) begin
        image_2_173 <= io_pixelVal_in_2_4;
      end else if (8'had == _T_25[7:0]) begin
        image_2_173 <= io_pixelVal_in_2_3;
      end else if (8'had == _T_22[7:0]) begin
        image_2_173 <= io_pixelVal_in_2_2;
      end else if (8'had == _T_19[7:0]) begin
        image_2_173 <= io_pixelVal_in_2_1;
      end else if (8'had == _T_15[7:0]) begin
        image_2_173 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_174 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hae == _T_34[7:0]) begin
        image_2_174 <= io_pixelVal_in_2_6;
      end else if (8'hae == _T_31[7:0]) begin
        image_2_174 <= io_pixelVal_in_2_5;
      end else if (8'hae == _T_28[7:0]) begin
        image_2_174 <= io_pixelVal_in_2_4;
      end else if (8'hae == _T_25[7:0]) begin
        image_2_174 <= io_pixelVal_in_2_3;
      end else if (8'hae == _T_22[7:0]) begin
        image_2_174 <= io_pixelVal_in_2_2;
      end else if (8'hae == _T_19[7:0]) begin
        image_2_174 <= io_pixelVal_in_2_1;
      end else if (8'hae == _T_15[7:0]) begin
        image_2_174 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_175 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'haf == _T_34[7:0]) begin
        image_2_175 <= io_pixelVal_in_2_6;
      end else if (8'haf == _T_31[7:0]) begin
        image_2_175 <= io_pixelVal_in_2_5;
      end else if (8'haf == _T_28[7:0]) begin
        image_2_175 <= io_pixelVal_in_2_4;
      end else if (8'haf == _T_25[7:0]) begin
        image_2_175 <= io_pixelVal_in_2_3;
      end else if (8'haf == _T_22[7:0]) begin
        image_2_175 <= io_pixelVal_in_2_2;
      end else if (8'haf == _T_19[7:0]) begin
        image_2_175 <= io_pixelVal_in_2_1;
      end else if (8'haf == _T_15[7:0]) begin
        image_2_175 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_176 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb0 == _T_34[7:0]) begin
        image_2_176 <= io_pixelVal_in_2_6;
      end else if (8'hb0 == _T_31[7:0]) begin
        image_2_176 <= io_pixelVal_in_2_5;
      end else if (8'hb0 == _T_28[7:0]) begin
        image_2_176 <= io_pixelVal_in_2_4;
      end else if (8'hb0 == _T_25[7:0]) begin
        image_2_176 <= io_pixelVal_in_2_3;
      end else if (8'hb0 == _T_22[7:0]) begin
        image_2_176 <= io_pixelVal_in_2_2;
      end else if (8'hb0 == _T_19[7:0]) begin
        image_2_176 <= io_pixelVal_in_2_1;
      end else if (8'hb0 == _T_15[7:0]) begin
        image_2_176 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_177 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb1 == _T_34[7:0]) begin
        image_2_177 <= io_pixelVal_in_2_6;
      end else if (8'hb1 == _T_31[7:0]) begin
        image_2_177 <= io_pixelVal_in_2_5;
      end else if (8'hb1 == _T_28[7:0]) begin
        image_2_177 <= io_pixelVal_in_2_4;
      end else if (8'hb1 == _T_25[7:0]) begin
        image_2_177 <= io_pixelVal_in_2_3;
      end else if (8'hb1 == _T_22[7:0]) begin
        image_2_177 <= io_pixelVal_in_2_2;
      end else if (8'hb1 == _T_19[7:0]) begin
        image_2_177 <= io_pixelVal_in_2_1;
      end else if (8'hb1 == _T_15[7:0]) begin
        image_2_177 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_178 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb2 == _T_34[7:0]) begin
        image_2_178 <= io_pixelVal_in_2_6;
      end else if (8'hb2 == _T_31[7:0]) begin
        image_2_178 <= io_pixelVal_in_2_5;
      end else if (8'hb2 == _T_28[7:0]) begin
        image_2_178 <= io_pixelVal_in_2_4;
      end else if (8'hb2 == _T_25[7:0]) begin
        image_2_178 <= io_pixelVal_in_2_3;
      end else if (8'hb2 == _T_22[7:0]) begin
        image_2_178 <= io_pixelVal_in_2_2;
      end else if (8'hb2 == _T_19[7:0]) begin
        image_2_178 <= io_pixelVal_in_2_1;
      end else if (8'hb2 == _T_15[7:0]) begin
        image_2_178 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_179 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb3 == _T_34[7:0]) begin
        image_2_179 <= io_pixelVal_in_2_6;
      end else if (8'hb3 == _T_31[7:0]) begin
        image_2_179 <= io_pixelVal_in_2_5;
      end else if (8'hb3 == _T_28[7:0]) begin
        image_2_179 <= io_pixelVal_in_2_4;
      end else if (8'hb3 == _T_25[7:0]) begin
        image_2_179 <= io_pixelVal_in_2_3;
      end else if (8'hb3 == _T_22[7:0]) begin
        image_2_179 <= io_pixelVal_in_2_2;
      end else if (8'hb3 == _T_19[7:0]) begin
        image_2_179 <= io_pixelVal_in_2_1;
      end else if (8'hb3 == _T_15[7:0]) begin
        image_2_179 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_180 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb4 == _T_34[7:0]) begin
        image_2_180 <= io_pixelVal_in_2_6;
      end else if (8'hb4 == _T_31[7:0]) begin
        image_2_180 <= io_pixelVal_in_2_5;
      end else if (8'hb4 == _T_28[7:0]) begin
        image_2_180 <= io_pixelVal_in_2_4;
      end else if (8'hb4 == _T_25[7:0]) begin
        image_2_180 <= io_pixelVal_in_2_3;
      end else if (8'hb4 == _T_22[7:0]) begin
        image_2_180 <= io_pixelVal_in_2_2;
      end else if (8'hb4 == _T_19[7:0]) begin
        image_2_180 <= io_pixelVal_in_2_1;
      end else if (8'hb4 == _T_15[7:0]) begin
        image_2_180 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_181 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb5 == _T_34[7:0]) begin
        image_2_181 <= io_pixelVal_in_2_6;
      end else if (8'hb5 == _T_31[7:0]) begin
        image_2_181 <= io_pixelVal_in_2_5;
      end else if (8'hb5 == _T_28[7:0]) begin
        image_2_181 <= io_pixelVal_in_2_4;
      end else if (8'hb5 == _T_25[7:0]) begin
        image_2_181 <= io_pixelVal_in_2_3;
      end else if (8'hb5 == _T_22[7:0]) begin
        image_2_181 <= io_pixelVal_in_2_2;
      end else if (8'hb5 == _T_19[7:0]) begin
        image_2_181 <= io_pixelVal_in_2_1;
      end else if (8'hb5 == _T_15[7:0]) begin
        image_2_181 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_182 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb6 == _T_34[7:0]) begin
        image_2_182 <= io_pixelVal_in_2_6;
      end else if (8'hb6 == _T_31[7:0]) begin
        image_2_182 <= io_pixelVal_in_2_5;
      end else if (8'hb6 == _T_28[7:0]) begin
        image_2_182 <= io_pixelVal_in_2_4;
      end else if (8'hb6 == _T_25[7:0]) begin
        image_2_182 <= io_pixelVal_in_2_3;
      end else if (8'hb6 == _T_22[7:0]) begin
        image_2_182 <= io_pixelVal_in_2_2;
      end else if (8'hb6 == _T_19[7:0]) begin
        image_2_182 <= io_pixelVal_in_2_1;
      end else if (8'hb6 == _T_15[7:0]) begin
        image_2_182 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_183 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb7 == _T_34[7:0]) begin
        image_2_183 <= io_pixelVal_in_2_6;
      end else if (8'hb7 == _T_31[7:0]) begin
        image_2_183 <= io_pixelVal_in_2_5;
      end else if (8'hb7 == _T_28[7:0]) begin
        image_2_183 <= io_pixelVal_in_2_4;
      end else if (8'hb7 == _T_25[7:0]) begin
        image_2_183 <= io_pixelVal_in_2_3;
      end else if (8'hb7 == _T_22[7:0]) begin
        image_2_183 <= io_pixelVal_in_2_2;
      end else if (8'hb7 == _T_19[7:0]) begin
        image_2_183 <= io_pixelVal_in_2_1;
      end else if (8'hb7 == _T_15[7:0]) begin
        image_2_183 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_184 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb8 == _T_34[7:0]) begin
        image_2_184 <= io_pixelVal_in_2_6;
      end else if (8'hb8 == _T_31[7:0]) begin
        image_2_184 <= io_pixelVal_in_2_5;
      end else if (8'hb8 == _T_28[7:0]) begin
        image_2_184 <= io_pixelVal_in_2_4;
      end else if (8'hb8 == _T_25[7:0]) begin
        image_2_184 <= io_pixelVal_in_2_3;
      end else if (8'hb8 == _T_22[7:0]) begin
        image_2_184 <= io_pixelVal_in_2_2;
      end else if (8'hb8 == _T_19[7:0]) begin
        image_2_184 <= io_pixelVal_in_2_1;
      end else if (8'hb8 == _T_15[7:0]) begin
        image_2_184 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_185 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hb9 == _T_34[7:0]) begin
        image_2_185 <= io_pixelVal_in_2_6;
      end else if (8'hb9 == _T_31[7:0]) begin
        image_2_185 <= io_pixelVal_in_2_5;
      end else if (8'hb9 == _T_28[7:0]) begin
        image_2_185 <= io_pixelVal_in_2_4;
      end else if (8'hb9 == _T_25[7:0]) begin
        image_2_185 <= io_pixelVal_in_2_3;
      end else if (8'hb9 == _T_22[7:0]) begin
        image_2_185 <= io_pixelVal_in_2_2;
      end else if (8'hb9 == _T_19[7:0]) begin
        image_2_185 <= io_pixelVal_in_2_1;
      end else if (8'hb9 == _T_15[7:0]) begin
        image_2_185 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_186 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hba == _T_34[7:0]) begin
        image_2_186 <= io_pixelVal_in_2_6;
      end else if (8'hba == _T_31[7:0]) begin
        image_2_186 <= io_pixelVal_in_2_5;
      end else if (8'hba == _T_28[7:0]) begin
        image_2_186 <= io_pixelVal_in_2_4;
      end else if (8'hba == _T_25[7:0]) begin
        image_2_186 <= io_pixelVal_in_2_3;
      end else if (8'hba == _T_22[7:0]) begin
        image_2_186 <= io_pixelVal_in_2_2;
      end else if (8'hba == _T_19[7:0]) begin
        image_2_186 <= io_pixelVal_in_2_1;
      end else if (8'hba == _T_15[7:0]) begin
        image_2_186 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_187 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbb == _T_34[7:0]) begin
        image_2_187 <= io_pixelVal_in_2_6;
      end else if (8'hbb == _T_31[7:0]) begin
        image_2_187 <= io_pixelVal_in_2_5;
      end else if (8'hbb == _T_28[7:0]) begin
        image_2_187 <= io_pixelVal_in_2_4;
      end else if (8'hbb == _T_25[7:0]) begin
        image_2_187 <= io_pixelVal_in_2_3;
      end else if (8'hbb == _T_22[7:0]) begin
        image_2_187 <= io_pixelVal_in_2_2;
      end else if (8'hbb == _T_19[7:0]) begin
        image_2_187 <= io_pixelVal_in_2_1;
      end else if (8'hbb == _T_15[7:0]) begin
        image_2_187 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_188 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbc == _T_34[7:0]) begin
        image_2_188 <= io_pixelVal_in_2_6;
      end else if (8'hbc == _T_31[7:0]) begin
        image_2_188 <= io_pixelVal_in_2_5;
      end else if (8'hbc == _T_28[7:0]) begin
        image_2_188 <= io_pixelVal_in_2_4;
      end else if (8'hbc == _T_25[7:0]) begin
        image_2_188 <= io_pixelVal_in_2_3;
      end else if (8'hbc == _T_22[7:0]) begin
        image_2_188 <= io_pixelVal_in_2_2;
      end else if (8'hbc == _T_19[7:0]) begin
        image_2_188 <= io_pixelVal_in_2_1;
      end else if (8'hbc == _T_15[7:0]) begin
        image_2_188 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_189 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbd == _T_34[7:0]) begin
        image_2_189 <= io_pixelVal_in_2_6;
      end else if (8'hbd == _T_31[7:0]) begin
        image_2_189 <= io_pixelVal_in_2_5;
      end else if (8'hbd == _T_28[7:0]) begin
        image_2_189 <= io_pixelVal_in_2_4;
      end else if (8'hbd == _T_25[7:0]) begin
        image_2_189 <= io_pixelVal_in_2_3;
      end else if (8'hbd == _T_22[7:0]) begin
        image_2_189 <= io_pixelVal_in_2_2;
      end else if (8'hbd == _T_19[7:0]) begin
        image_2_189 <= io_pixelVal_in_2_1;
      end else if (8'hbd == _T_15[7:0]) begin
        image_2_189 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_190 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbe == _T_34[7:0]) begin
        image_2_190 <= io_pixelVal_in_2_6;
      end else if (8'hbe == _T_31[7:0]) begin
        image_2_190 <= io_pixelVal_in_2_5;
      end else if (8'hbe == _T_28[7:0]) begin
        image_2_190 <= io_pixelVal_in_2_4;
      end else if (8'hbe == _T_25[7:0]) begin
        image_2_190 <= io_pixelVal_in_2_3;
      end else if (8'hbe == _T_22[7:0]) begin
        image_2_190 <= io_pixelVal_in_2_2;
      end else if (8'hbe == _T_19[7:0]) begin
        image_2_190 <= io_pixelVal_in_2_1;
      end else if (8'hbe == _T_15[7:0]) begin
        image_2_190 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_191 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hbf == _T_34[7:0]) begin
        image_2_191 <= io_pixelVal_in_2_6;
      end else if (8'hbf == _T_31[7:0]) begin
        image_2_191 <= io_pixelVal_in_2_5;
      end else if (8'hbf == _T_28[7:0]) begin
        image_2_191 <= io_pixelVal_in_2_4;
      end else if (8'hbf == _T_25[7:0]) begin
        image_2_191 <= io_pixelVal_in_2_3;
      end else if (8'hbf == _T_22[7:0]) begin
        image_2_191 <= io_pixelVal_in_2_2;
      end else if (8'hbf == _T_19[7:0]) begin
        image_2_191 <= io_pixelVal_in_2_1;
      end else if (8'hbf == _T_15[7:0]) begin
        image_2_191 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_192 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc0 == _T_34[7:0]) begin
        image_2_192 <= io_pixelVal_in_2_6;
      end else if (8'hc0 == _T_31[7:0]) begin
        image_2_192 <= io_pixelVal_in_2_5;
      end else if (8'hc0 == _T_28[7:0]) begin
        image_2_192 <= io_pixelVal_in_2_4;
      end else if (8'hc0 == _T_25[7:0]) begin
        image_2_192 <= io_pixelVal_in_2_3;
      end else if (8'hc0 == _T_22[7:0]) begin
        image_2_192 <= io_pixelVal_in_2_2;
      end else if (8'hc0 == _T_19[7:0]) begin
        image_2_192 <= io_pixelVal_in_2_1;
      end else if (8'hc0 == _T_15[7:0]) begin
        image_2_192 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_193 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc1 == _T_34[7:0]) begin
        image_2_193 <= io_pixelVal_in_2_6;
      end else if (8'hc1 == _T_31[7:0]) begin
        image_2_193 <= io_pixelVal_in_2_5;
      end else if (8'hc1 == _T_28[7:0]) begin
        image_2_193 <= io_pixelVal_in_2_4;
      end else if (8'hc1 == _T_25[7:0]) begin
        image_2_193 <= io_pixelVal_in_2_3;
      end else if (8'hc1 == _T_22[7:0]) begin
        image_2_193 <= io_pixelVal_in_2_2;
      end else if (8'hc1 == _T_19[7:0]) begin
        image_2_193 <= io_pixelVal_in_2_1;
      end else if (8'hc1 == _T_15[7:0]) begin
        image_2_193 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_194 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc2 == _T_34[7:0]) begin
        image_2_194 <= io_pixelVal_in_2_6;
      end else if (8'hc2 == _T_31[7:0]) begin
        image_2_194 <= io_pixelVal_in_2_5;
      end else if (8'hc2 == _T_28[7:0]) begin
        image_2_194 <= io_pixelVal_in_2_4;
      end else if (8'hc2 == _T_25[7:0]) begin
        image_2_194 <= io_pixelVal_in_2_3;
      end else if (8'hc2 == _T_22[7:0]) begin
        image_2_194 <= io_pixelVal_in_2_2;
      end else if (8'hc2 == _T_19[7:0]) begin
        image_2_194 <= io_pixelVal_in_2_1;
      end else if (8'hc2 == _T_15[7:0]) begin
        image_2_194 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_195 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc3 == _T_34[7:0]) begin
        image_2_195 <= io_pixelVal_in_2_6;
      end else if (8'hc3 == _T_31[7:0]) begin
        image_2_195 <= io_pixelVal_in_2_5;
      end else if (8'hc3 == _T_28[7:0]) begin
        image_2_195 <= io_pixelVal_in_2_4;
      end else if (8'hc3 == _T_25[7:0]) begin
        image_2_195 <= io_pixelVal_in_2_3;
      end else if (8'hc3 == _T_22[7:0]) begin
        image_2_195 <= io_pixelVal_in_2_2;
      end else if (8'hc3 == _T_19[7:0]) begin
        image_2_195 <= io_pixelVal_in_2_1;
      end else if (8'hc3 == _T_15[7:0]) begin
        image_2_195 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_196 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc4 == _T_34[7:0]) begin
        image_2_196 <= io_pixelVal_in_2_6;
      end else if (8'hc4 == _T_31[7:0]) begin
        image_2_196 <= io_pixelVal_in_2_5;
      end else if (8'hc4 == _T_28[7:0]) begin
        image_2_196 <= io_pixelVal_in_2_4;
      end else if (8'hc4 == _T_25[7:0]) begin
        image_2_196 <= io_pixelVal_in_2_3;
      end else if (8'hc4 == _T_22[7:0]) begin
        image_2_196 <= io_pixelVal_in_2_2;
      end else if (8'hc4 == _T_19[7:0]) begin
        image_2_196 <= io_pixelVal_in_2_1;
      end else if (8'hc4 == _T_15[7:0]) begin
        image_2_196 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_197 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc5 == _T_34[7:0]) begin
        image_2_197 <= io_pixelVal_in_2_6;
      end else if (8'hc5 == _T_31[7:0]) begin
        image_2_197 <= io_pixelVal_in_2_5;
      end else if (8'hc5 == _T_28[7:0]) begin
        image_2_197 <= io_pixelVal_in_2_4;
      end else if (8'hc5 == _T_25[7:0]) begin
        image_2_197 <= io_pixelVal_in_2_3;
      end else if (8'hc5 == _T_22[7:0]) begin
        image_2_197 <= io_pixelVal_in_2_2;
      end else if (8'hc5 == _T_19[7:0]) begin
        image_2_197 <= io_pixelVal_in_2_1;
      end else if (8'hc5 == _T_15[7:0]) begin
        image_2_197 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_198 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc6 == _T_34[7:0]) begin
        image_2_198 <= io_pixelVal_in_2_6;
      end else if (8'hc6 == _T_31[7:0]) begin
        image_2_198 <= io_pixelVal_in_2_5;
      end else if (8'hc6 == _T_28[7:0]) begin
        image_2_198 <= io_pixelVal_in_2_4;
      end else if (8'hc6 == _T_25[7:0]) begin
        image_2_198 <= io_pixelVal_in_2_3;
      end else if (8'hc6 == _T_22[7:0]) begin
        image_2_198 <= io_pixelVal_in_2_2;
      end else if (8'hc6 == _T_19[7:0]) begin
        image_2_198 <= io_pixelVal_in_2_1;
      end else if (8'hc6 == _T_15[7:0]) begin
        image_2_198 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_199 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc7 == _T_34[7:0]) begin
        image_2_199 <= io_pixelVal_in_2_6;
      end else if (8'hc7 == _T_31[7:0]) begin
        image_2_199 <= io_pixelVal_in_2_5;
      end else if (8'hc7 == _T_28[7:0]) begin
        image_2_199 <= io_pixelVal_in_2_4;
      end else if (8'hc7 == _T_25[7:0]) begin
        image_2_199 <= io_pixelVal_in_2_3;
      end else if (8'hc7 == _T_22[7:0]) begin
        image_2_199 <= io_pixelVal_in_2_2;
      end else if (8'hc7 == _T_19[7:0]) begin
        image_2_199 <= io_pixelVal_in_2_1;
      end else if (8'hc7 == _T_15[7:0]) begin
        image_2_199 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_200 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc8 == _T_34[7:0]) begin
        image_2_200 <= io_pixelVal_in_2_6;
      end else if (8'hc8 == _T_31[7:0]) begin
        image_2_200 <= io_pixelVal_in_2_5;
      end else if (8'hc8 == _T_28[7:0]) begin
        image_2_200 <= io_pixelVal_in_2_4;
      end else if (8'hc8 == _T_25[7:0]) begin
        image_2_200 <= io_pixelVal_in_2_3;
      end else if (8'hc8 == _T_22[7:0]) begin
        image_2_200 <= io_pixelVal_in_2_2;
      end else if (8'hc8 == _T_19[7:0]) begin
        image_2_200 <= io_pixelVal_in_2_1;
      end else if (8'hc8 == _T_15[7:0]) begin
        image_2_200 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_201 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hc9 == _T_34[7:0]) begin
        image_2_201 <= io_pixelVal_in_2_6;
      end else if (8'hc9 == _T_31[7:0]) begin
        image_2_201 <= io_pixelVal_in_2_5;
      end else if (8'hc9 == _T_28[7:0]) begin
        image_2_201 <= io_pixelVal_in_2_4;
      end else if (8'hc9 == _T_25[7:0]) begin
        image_2_201 <= io_pixelVal_in_2_3;
      end else if (8'hc9 == _T_22[7:0]) begin
        image_2_201 <= io_pixelVal_in_2_2;
      end else if (8'hc9 == _T_19[7:0]) begin
        image_2_201 <= io_pixelVal_in_2_1;
      end else if (8'hc9 == _T_15[7:0]) begin
        image_2_201 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_202 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hca == _T_34[7:0]) begin
        image_2_202 <= io_pixelVal_in_2_6;
      end else if (8'hca == _T_31[7:0]) begin
        image_2_202 <= io_pixelVal_in_2_5;
      end else if (8'hca == _T_28[7:0]) begin
        image_2_202 <= io_pixelVal_in_2_4;
      end else if (8'hca == _T_25[7:0]) begin
        image_2_202 <= io_pixelVal_in_2_3;
      end else if (8'hca == _T_22[7:0]) begin
        image_2_202 <= io_pixelVal_in_2_2;
      end else if (8'hca == _T_19[7:0]) begin
        image_2_202 <= io_pixelVal_in_2_1;
      end else if (8'hca == _T_15[7:0]) begin
        image_2_202 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_203 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hcb == _T_34[7:0]) begin
        image_2_203 <= io_pixelVal_in_2_6;
      end else if (8'hcb == _T_31[7:0]) begin
        image_2_203 <= io_pixelVal_in_2_5;
      end else if (8'hcb == _T_28[7:0]) begin
        image_2_203 <= io_pixelVal_in_2_4;
      end else if (8'hcb == _T_25[7:0]) begin
        image_2_203 <= io_pixelVal_in_2_3;
      end else if (8'hcb == _T_22[7:0]) begin
        image_2_203 <= io_pixelVal_in_2_2;
      end else if (8'hcb == _T_19[7:0]) begin
        image_2_203 <= io_pixelVal_in_2_1;
      end else if (8'hcb == _T_15[7:0]) begin
        image_2_203 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_204 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hcc == _T_34[7:0]) begin
        image_2_204 <= io_pixelVal_in_2_6;
      end else if (8'hcc == _T_31[7:0]) begin
        image_2_204 <= io_pixelVal_in_2_5;
      end else if (8'hcc == _T_28[7:0]) begin
        image_2_204 <= io_pixelVal_in_2_4;
      end else if (8'hcc == _T_25[7:0]) begin
        image_2_204 <= io_pixelVal_in_2_3;
      end else if (8'hcc == _T_22[7:0]) begin
        image_2_204 <= io_pixelVal_in_2_2;
      end else if (8'hcc == _T_19[7:0]) begin
        image_2_204 <= io_pixelVal_in_2_1;
      end else if (8'hcc == _T_15[7:0]) begin
        image_2_204 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_205 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hcd == _T_34[7:0]) begin
        image_2_205 <= io_pixelVal_in_2_6;
      end else if (8'hcd == _T_31[7:0]) begin
        image_2_205 <= io_pixelVal_in_2_5;
      end else if (8'hcd == _T_28[7:0]) begin
        image_2_205 <= io_pixelVal_in_2_4;
      end else if (8'hcd == _T_25[7:0]) begin
        image_2_205 <= io_pixelVal_in_2_3;
      end else if (8'hcd == _T_22[7:0]) begin
        image_2_205 <= io_pixelVal_in_2_2;
      end else if (8'hcd == _T_19[7:0]) begin
        image_2_205 <= io_pixelVal_in_2_1;
      end else if (8'hcd == _T_15[7:0]) begin
        image_2_205 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_206 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hce == _T_34[7:0]) begin
        image_2_206 <= io_pixelVal_in_2_6;
      end else if (8'hce == _T_31[7:0]) begin
        image_2_206 <= io_pixelVal_in_2_5;
      end else if (8'hce == _T_28[7:0]) begin
        image_2_206 <= io_pixelVal_in_2_4;
      end else if (8'hce == _T_25[7:0]) begin
        image_2_206 <= io_pixelVal_in_2_3;
      end else if (8'hce == _T_22[7:0]) begin
        image_2_206 <= io_pixelVal_in_2_2;
      end else if (8'hce == _T_19[7:0]) begin
        image_2_206 <= io_pixelVal_in_2_1;
      end else if (8'hce == _T_15[7:0]) begin
        image_2_206 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_207 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hcf == _T_34[7:0]) begin
        image_2_207 <= io_pixelVal_in_2_6;
      end else if (8'hcf == _T_31[7:0]) begin
        image_2_207 <= io_pixelVal_in_2_5;
      end else if (8'hcf == _T_28[7:0]) begin
        image_2_207 <= io_pixelVal_in_2_4;
      end else if (8'hcf == _T_25[7:0]) begin
        image_2_207 <= io_pixelVal_in_2_3;
      end else if (8'hcf == _T_22[7:0]) begin
        image_2_207 <= io_pixelVal_in_2_2;
      end else if (8'hcf == _T_19[7:0]) begin
        image_2_207 <= io_pixelVal_in_2_1;
      end else if (8'hcf == _T_15[7:0]) begin
        image_2_207 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_208 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd0 == _T_34[7:0]) begin
        image_2_208 <= io_pixelVal_in_2_6;
      end else if (8'hd0 == _T_31[7:0]) begin
        image_2_208 <= io_pixelVal_in_2_5;
      end else if (8'hd0 == _T_28[7:0]) begin
        image_2_208 <= io_pixelVal_in_2_4;
      end else if (8'hd0 == _T_25[7:0]) begin
        image_2_208 <= io_pixelVal_in_2_3;
      end else if (8'hd0 == _T_22[7:0]) begin
        image_2_208 <= io_pixelVal_in_2_2;
      end else if (8'hd0 == _T_19[7:0]) begin
        image_2_208 <= io_pixelVal_in_2_1;
      end else if (8'hd0 == _T_15[7:0]) begin
        image_2_208 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_209 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd1 == _T_34[7:0]) begin
        image_2_209 <= io_pixelVal_in_2_6;
      end else if (8'hd1 == _T_31[7:0]) begin
        image_2_209 <= io_pixelVal_in_2_5;
      end else if (8'hd1 == _T_28[7:0]) begin
        image_2_209 <= io_pixelVal_in_2_4;
      end else if (8'hd1 == _T_25[7:0]) begin
        image_2_209 <= io_pixelVal_in_2_3;
      end else if (8'hd1 == _T_22[7:0]) begin
        image_2_209 <= io_pixelVal_in_2_2;
      end else if (8'hd1 == _T_19[7:0]) begin
        image_2_209 <= io_pixelVal_in_2_1;
      end else if (8'hd1 == _T_15[7:0]) begin
        image_2_209 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_210 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd2 == _T_34[7:0]) begin
        image_2_210 <= io_pixelVal_in_2_6;
      end else if (8'hd2 == _T_31[7:0]) begin
        image_2_210 <= io_pixelVal_in_2_5;
      end else if (8'hd2 == _T_28[7:0]) begin
        image_2_210 <= io_pixelVal_in_2_4;
      end else if (8'hd2 == _T_25[7:0]) begin
        image_2_210 <= io_pixelVal_in_2_3;
      end else if (8'hd2 == _T_22[7:0]) begin
        image_2_210 <= io_pixelVal_in_2_2;
      end else if (8'hd2 == _T_19[7:0]) begin
        image_2_210 <= io_pixelVal_in_2_1;
      end else if (8'hd2 == _T_15[7:0]) begin
        image_2_210 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_211 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd3 == _T_34[7:0]) begin
        image_2_211 <= io_pixelVal_in_2_6;
      end else if (8'hd3 == _T_31[7:0]) begin
        image_2_211 <= io_pixelVal_in_2_5;
      end else if (8'hd3 == _T_28[7:0]) begin
        image_2_211 <= io_pixelVal_in_2_4;
      end else if (8'hd3 == _T_25[7:0]) begin
        image_2_211 <= io_pixelVal_in_2_3;
      end else if (8'hd3 == _T_22[7:0]) begin
        image_2_211 <= io_pixelVal_in_2_2;
      end else if (8'hd3 == _T_19[7:0]) begin
        image_2_211 <= io_pixelVal_in_2_1;
      end else if (8'hd3 == _T_15[7:0]) begin
        image_2_211 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_212 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd4 == _T_34[7:0]) begin
        image_2_212 <= io_pixelVal_in_2_6;
      end else if (8'hd4 == _T_31[7:0]) begin
        image_2_212 <= io_pixelVal_in_2_5;
      end else if (8'hd4 == _T_28[7:0]) begin
        image_2_212 <= io_pixelVal_in_2_4;
      end else if (8'hd4 == _T_25[7:0]) begin
        image_2_212 <= io_pixelVal_in_2_3;
      end else if (8'hd4 == _T_22[7:0]) begin
        image_2_212 <= io_pixelVal_in_2_2;
      end else if (8'hd4 == _T_19[7:0]) begin
        image_2_212 <= io_pixelVal_in_2_1;
      end else if (8'hd4 == _T_15[7:0]) begin
        image_2_212 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_213 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd5 == _T_34[7:0]) begin
        image_2_213 <= io_pixelVal_in_2_6;
      end else if (8'hd5 == _T_31[7:0]) begin
        image_2_213 <= io_pixelVal_in_2_5;
      end else if (8'hd5 == _T_28[7:0]) begin
        image_2_213 <= io_pixelVal_in_2_4;
      end else if (8'hd5 == _T_25[7:0]) begin
        image_2_213 <= io_pixelVal_in_2_3;
      end else if (8'hd5 == _T_22[7:0]) begin
        image_2_213 <= io_pixelVal_in_2_2;
      end else if (8'hd5 == _T_19[7:0]) begin
        image_2_213 <= io_pixelVal_in_2_1;
      end else if (8'hd5 == _T_15[7:0]) begin
        image_2_213 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_214 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd6 == _T_34[7:0]) begin
        image_2_214 <= io_pixelVal_in_2_6;
      end else if (8'hd6 == _T_31[7:0]) begin
        image_2_214 <= io_pixelVal_in_2_5;
      end else if (8'hd6 == _T_28[7:0]) begin
        image_2_214 <= io_pixelVal_in_2_4;
      end else if (8'hd6 == _T_25[7:0]) begin
        image_2_214 <= io_pixelVal_in_2_3;
      end else if (8'hd6 == _T_22[7:0]) begin
        image_2_214 <= io_pixelVal_in_2_2;
      end else if (8'hd6 == _T_19[7:0]) begin
        image_2_214 <= io_pixelVal_in_2_1;
      end else if (8'hd6 == _T_15[7:0]) begin
        image_2_214 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_215 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd7 == _T_34[7:0]) begin
        image_2_215 <= io_pixelVal_in_2_6;
      end else if (8'hd7 == _T_31[7:0]) begin
        image_2_215 <= io_pixelVal_in_2_5;
      end else if (8'hd7 == _T_28[7:0]) begin
        image_2_215 <= io_pixelVal_in_2_4;
      end else if (8'hd7 == _T_25[7:0]) begin
        image_2_215 <= io_pixelVal_in_2_3;
      end else if (8'hd7 == _T_22[7:0]) begin
        image_2_215 <= io_pixelVal_in_2_2;
      end else if (8'hd7 == _T_19[7:0]) begin
        image_2_215 <= io_pixelVal_in_2_1;
      end else if (8'hd7 == _T_15[7:0]) begin
        image_2_215 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_216 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd8 == _T_34[7:0]) begin
        image_2_216 <= io_pixelVal_in_2_6;
      end else if (8'hd8 == _T_31[7:0]) begin
        image_2_216 <= io_pixelVal_in_2_5;
      end else if (8'hd8 == _T_28[7:0]) begin
        image_2_216 <= io_pixelVal_in_2_4;
      end else if (8'hd8 == _T_25[7:0]) begin
        image_2_216 <= io_pixelVal_in_2_3;
      end else if (8'hd8 == _T_22[7:0]) begin
        image_2_216 <= io_pixelVal_in_2_2;
      end else if (8'hd8 == _T_19[7:0]) begin
        image_2_216 <= io_pixelVal_in_2_1;
      end else if (8'hd8 == _T_15[7:0]) begin
        image_2_216 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_217 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hd9 == _T_34[7:0]) begin
        image_2_217 <= io_pixelVal_in_2_6;
      end else if (8'hd9 == _T_31[7:0]) begin
        image_2_217 <= io_pixelVal_in_2_5;
      end else if (8'hd9 == _T_28[7:0]) begin
        image_2_217 <= io_pixelVal_in_2_4;
      end else if (8'hd9 == _T_25[7:0]) begin
        image_2_217 <= io_pixelVal_in_2_3;
      end else if (8'hd9 == _T_22[7:0]) begin
        image_2_217 <= io_pixelVal_in_2_2;
      end else if (8'hd9 == _T_19[7:0]) begin
        image_2_217 <= io_pixelVal_in_2_1;
      end else if (8'hd9 == _T_15[7:0]) begin
        image_2_217 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_218 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hda == _T_34[7:0]) begin
        image_2_218 <= io_pixelVal_in_2_6;
      end else if (8'hda == _T_31[7:0]) begin
        image_2_218 <= io_pixelVal_in_2_5;
      end else if (8'hda == _T_28[7:0]) begin
        image_2_218 <= io_pixelVal_in_2_4;
      end else if (8'hda == _T_25[7:0]) begin
        image_2_218 <= io_pixelVal_in_2_3;
      end else if (8'hda == _T_22[7:0]) begin
        image_2_218 <= io_pixelVal_in_2_2;
      end else if (8'hda == _T_19[7:0]) begin
        image_2_218 <= io_pixelVal_in_2_1;
      end else if (8'hda == _T_15[7:0]) begin
        image_2_218 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_219 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hdb == _T_34[7:0]) begin
        image_2_219 <= io_pixelVal_in_2_6;
      end else if (8'hdb == _T_31[7:0]) begin
        image_2_219 <= io_pixelVal_in_2_5;
      end else if (8'hdb == _T_28[7:0]) begin
        image_2_219 <= io_pixelVal_in_2_4;
      end else if (8'hdb == _T_25[7:0]) begin
        image_2_219 <= io_pixelVal_in_2_3;
      end else if (8'hdb == _T_22[7:0]) begin
        image_2_219 <= io_pixelVal_in_2_2;
      end else if (8'hdb == _T_19[7:0]) begin
        image_2_219 <= io_pixelVal_in_2_1;
      end else if (8'hdb == _T_15[7:0]) begin
        image_2_219 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_220 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hdc == _T_34[7:0]) begin
        image_2_220 <= io_pixelVal_in_2_6;
      end else if (8'hdc == _T_31[7:0]) begin
        image_2_220 <= io_pixelVal_in_2_5;
      end else if (8'hdc == _T_28[7:0]) begin
        image_2_220 <= io_pixelVal_in_2_4;
      end else if (8'hdc == _T_25[7:0]) begin
        image_2_220 <= io_pixelVal_in_2_3;
      end else if (8'hdc == _T_22[7:0]) begin
        image_2_220 <= io_pixelVal_in_2_2;
      end else if (8'hdc == _T_19[7:0]) begin
        image_2_220 <= io_pixelVal_in_2_1;
      end else if (8'hdc == _T_15[7:0]) begin
        image_2_220 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_221 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hdd == _T_34[7:0]) begin
        image_2_221 <= io_pixelVal_in_2_6;
      end else if (8'hdd == _T_31[7:0]) begin
        image_2_221 <= io_pixelVal_in_2_5;
      end else if (8'hdd == _T_28[7:0]) begin
        image_2_221 <= io_pixelVal_in_2_4;
      end else if (8'hdd == _T_25[7:0]) begin
        image_2_221 <= io_pixelVal_in_2_3;
      end else if (8'hdd == _T_22[7:0]) begin
        image_2_221 <= io_pixelVal_in_2_2;
      end else if (8'hdd == _T_19[7:0]) begin
        image_2_221 <= io_pixelVal_in_2_1;
      end else if (8'hdd == _T_15[7:0]) begin
        image_2_221 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_222 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hde == _T_34[7:0]) begin
        image_2_222 <= io_pixelVal_in_2_6;
      end else if (8'hde == _T_31[7:0]) begin
        image_2_222 <= io_pixelVal_in_2_5;
      end else if (8'hde == _T_28[7:0]) begin
        image_2_222 <= io_pixelVal_in_2_4;
      end else if (8'hde == _T_25[7:0]) begin
        image_2_222 <= io_pixelVal_in_2_3;
      end else if (8'hde == _T_22[7:0]) begin
        image_2_222 <= io_pixelVal_in_2_2;
      end else if (8'hde == _T_19[7:0]) begin
        image_2_222 <= io_pixelVal_in_2_1;
      end else if (8'hde == _T_15[7:0]) begin
        image_2_222 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_223 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hdf == _T_34[7:0]) begin
        image_2_223 <= io_pixelVal_in_2_6;
      end else if (8'hdf == _T_31[7:0]) begin
        image_2_223 <= io_pixelVal_in_2_5;
      end else if (8'hdf == _T_28[7:0]) begin
        image_2_223 <= io_pixelVal_in_2_4;
      end else if (8'hdf == _T_25[7:0]) begin
        image_2_223 <= io_pixelVal_in_2_3;
      end else if (8'hdf == _T_22[7:0]) begin
        image_2_223 <= io_pixelVal_in_2_2;
      end else if (8'hdf == _T_19[7:0]) begin
        image_2_223 <= io_pixelVal_in_2_1;
      end else if (8'hdf == _T_15[7:0]) begin
        image_2_223 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_224 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he0 == _T_34[7:0]) begin
        image_2_224 <= io_pixelVal_in_2_6;
      end else if (8'he0 == _T_31[7:0]) begin
        image_2_224 <= io_pixelVal_in_2_5;
      end else if (8'he0 == _T_28[7:0]) begin
        image_2_224 <= io_pixelVal_in_2_4;
      end else if (8'he0 == _T_25[7:0]) begin
        image_2_224 <= io_pixelVal_in_2_3;
      end else if (8'he0 == _T_22[7:0]) begin
        image_2_224 <= io_pixelVal_in_2_2;
      end else if (8'he0 == _T_19[7:0]) begin
        image_2_224 <= io_pixelVal_in_2_1;
      end else if (8'he0 == _T_15[7:0]) begin
        image_2_224 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_225 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he1 == _T_34[7:0]) begin
        image_2_225 <= io_pixelVal_in_2_6;
      end else if (8'he1 == _T_31[7:0]) begin
        image_2_225 <= io_pixelVal_in_2_5;
      end else if (8'he1 == _T_28[7:0]) begin
        image_2_225 <= io_pixelVal_in_2_4;
      end else if (8'he1 == _T_25[7:0]) begin
        image_2_225 <= io_pixelVal_in_2_3;
      end else if (8'he1 == _T_22[7:0]) begin
        image_2_225 <= io_pixelVal_in_2_2;
      end else if (8'he1 == _T_19[7:0]) begin
        image_2_225 <= io_pixelVal_in_2_1;
      end else if (8'he1 == _T_15[7:0]) begin
        image_2_225 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_226 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he2 == _T_34[7:0]) begin
        image_2_226 <= io_pixelVal_in_2_6;
      end else if (8'he2 == _T_31[7:0]) begin
        image_2_226 <= io_pixelVal_in_2_5;
      end else if (8'he2 == _T_28[7:0]) begin
        image_2_226 <= io_pixelVal_in_2_4;
      end else if (8'he2 == _T_25[7:0]) begin
        image_2_226 <= io_pixelVal_in_2_3;
      end else if (8'he2 == _T_22[7:0]) begin
        image_2_226 <= io_pixelVal_in_2_2;
      end else if (8'he2 == _T_19[7:0]) begin
        image_2_226 <= io_pixelVal_in_2_1;
      end else if (8'he2 == _T_15[7:0]) begin
        image_2_226 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_227 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he3 == _T_34[7:0]) begin
        image_2_227 <= io_pixelVal_in_2_6;
      end else if (8'he3 == _T_31[7:0]) begin
        image_2_227 <= io_pixelVal_in_2_5;
      end else if (8'he3 == _T_28[7:0]) begin
        image_2_227 <= io_pixelVal_in_2_4;
      end else if (8'he3 == _T_25[7:0]) begin
        image_2_227 <= io_pixelVal_in_2_3;
      end else if (8'he3 == _T_22[7:0]) begin
        image_2_227 <= io_pixelVal_in_2_2;
      end else if (8'he3 == _T_19[7:0]) begin
        image_2_227 <= io_pixelVal_in_2_1;
      end else if (8'he3 == _T_15[7:0]) begin
        image_2_227 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_228 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he4 == _T_34[7:0]) begin
        image_2_228 <= io_pixelVal_in_2_6;
      end else if (8'he4 == _T_31[7:0]) begin
        image_2_228 <= io_pixelVal_in_2_5;
      end else if (8'he4 == _T_28[7:0]) begin
        image_2_228 <= io_pixelVal_in_2_4;
      end else if (8'he4 == _T_25[7:0]) begin
        image_2_228 <= io_pixelVal_in_2_3;
      end else if (8'he4 == _T_22[7:0]) begin
        image_2_228 <= io_pixelVal_in_2_2;
      end else if (8'he4 == _T_19[7:0]) begin
        image_2_228 <= io_pixelVal_in_2_1;
      end else if (8'he4 == _T_15[7:0]) begin
        image_2_228 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_229 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he5 == _T_34[7:0]) begin
        image_2_229 <= io_pixelVal_in_2_6;
      end else if (8'he5 == _T_31[7:0]) begin
        image_2_229 <= io_pixelVal_in_2_5;
      end else if (8'he5 == _T_28[7:0]) begin
        image_2_229 <= io_pixelVal_in_2_4;
      end else if (8'he5 == _T_25[7:0]) begin
        image_2_229 <= io_pixelVal_in_2_3;
      end else if (8'he5 == _T_22[7:0]) begin
        image_2_229 <= io_pixelVal_in_2_2;
      end else if (8'he5 == _T_19[7:0]) begin
        image_2_229 <= io_pixelVal_in_2_1;
      end else if (8'he5 == _T_15[7:0]) begin
        image_2_229 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_230 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he6 == _T_34[7:0]) begin
        image_2_230 <= io_pixelVal_in_2_6;
      end else if (8'he6 == _T_31[7:0]) begin
        image_2_230 <= io_pixelVal_in_2_5;
      end else if (8'he6 == _T_28[7:0]) begin
        image_2_230 <= io_pixelVal_in_2_4;
      end else if (8'he6 == _T_25[7:0]) begin
        image_2_230 <= io_pixelVal_in_2_3;
      end else if (8'he6 == _T_22[7:0]) begin
        image_2_230 <= io_pixelVal_in_2_2;
      end else if (8'he6 == _T_19[7:0]) begin
        image_2_230 <= io_pixelVal_in_2_1;
      end else if (8'he6 == _T_15[7:0]) begin
        image_2_230 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_231 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he7 == _T_34[7:0]) begin
        image_2_231 <= io_pixelVal_in_2_6;
      end else if (8'he7 == _T_31[7:0]) begin
        image_2_231 <= io_pixelVal_in_2_5;
      end else if (8'he7 == _T_28[7:0]) begin
        image_2_231 <= io_pixelVal_in_2_4;
      end else if (8'he7 == _T_25[7:0]) begin
        image_2_231 <= io_pixelVal_in_2_3;
      end else if (8'he7 == _T_22[7:0]) begin
        image_2_231 <= io_pixelVal_in_2_2;
      end else if (8'he7 == _T_19[7:0]) begin
        image_2_231 <= io_pixelVal_in_2_1;
      end else if (8'he7 == _T_15[7:0]) begin
        image_2_231 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_232 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he8 == _T_34[7:0]) begin
        image_2_232 <= io_pixelVal_in_2_6;
      end else if (8'he8 == _T_31[7:0]) begin
        image_2_232 <= io_pixelVal_in_2_5;
      end else if (8'he8 == _T_28[7:0]) begin
        image_2_232 <= io_pixelVal_in_2_4;
      end else if (8'he8 == _T_25[7:0]) begin
        image_2_232 <= io_pixelVal_in_2_3;
      end else if (8'he8 == _T_22[7:0]) begin
        image_2_232 <= io_pixelVal_in_2_2;
      end else if (8'he8 == _T_19[7:0]) begin
        image_2_232 <= io_pixelVal_in_2_1;
      end else if (8'he8 == _T_15[7:0]) begin
        image_2_232 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_233 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'he9 == _T_34[7:0]) begin
        image_2_233 <= io_pixelVal_in_2_6;
      end else if (8'he9 == _T_31[7:0]) begin
        image_2_233 <= io_pixelVal_in_2_5;
      end else if (8'he9 == _T_28[7:0]) begin
        image_2_233 <= io_pixelVal_in_2_4;
      end else if (8'he9 == _T_25[7:0]) begin
        image_2_233 <= io_pixelVal_in_2_3;
      end else if (8'he9 == _T_22[7:0]) begin
        image_2_233 <= io_pixelVal_in_2_2;
      end else if (8'he9 == _T_19[7:0]) begin
        image_2_233 <= io_pixelVal_in_2_1;
      end else if (8'he9 == _T_15[7:0]) begin
        image_2_233 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_234 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hea == _T_34[7:0]) begin
        image_2_234 <= io_pixelVal_in_2_6;
      end else if (8'hea == _T_31[7:0]) begin
        image_2_234 <= io_pixelVal_in_2_5;
      end else if (8'hea == _T_28[7:0]) begin
        image_2_234 <= io_pixelVal_in_2_4;
      end else if (8'hea == _T_25[7:0]) begin
        image_2_234 <= io_pixelVal_in_2_3;
      end else if (8'hea == _T_22[7:0]) begin
        image_2_234 <= io_pixelVal_in_2_2;
      end else if (8'hea == _T_19[7:0]) begin
        image_2_234 <= io_pixelVal_in_2_1;
      end else if (8'hea == _T_15[7:0]) begin
        image_2_234 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_235 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'heb == _T_34[7:0]) begin
        image_2_235 <= io_pixelVal_in_2_6;
      end else if (8'heb == _T_31[7:0]) begin
        image_2_235 <= io_pixelVal_in_2_5;
      end else if (8'heb == _T_28[7:0]) begin
        image_2_235 <= io_pixelVal_in_2_4;
      end else if (8'heb == _T_25[7:0]) begin
        image_2_235 <= io_pixelVal_in_2_3;
      end else if (8'heb == _T_22[7:0]) begin
        image_2_235 <= io_pixelVal_in_2_2;
      end else if (8'heb == _T_19[7:0]) begin
        image_2_235 <= io_pixelVal_in_2_1;
      end else if (8'heb == _T_15[7:0]) begin
        image_2_235 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_236 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hec == _T_34[7:0]) begin
        image_2_236 <= io_pixelVal_in_2_6;
      end else if (8'hec == _T_31[7:0]) begin
        image_2_236 <= io_pixelVal_in_2_5;
      end else if (8'hec == _T_28[7:0]) begin
        image_2_236 <= io_pixelVal_in_2_4;
      end else if (8'hec == _T_25[7:0]) begin
        image_2_236 <= io_pixelVal_in_2_3;
      end else if (8'hec == _T_22[7:0]) begin
        image_2_236 <= io_pixelVal_in_2_2;
      end else if (8'hec == _T_19[7:0]) begin
        image_2_236 <= io_pixelVal_in_2_1;
      end else if (8'hec == _T_15[7:0]) begin
        image_2_236 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_237 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hed == _T_34[7:0]) begin
        image_2_237 <= io_pixelVal_in_2_6;
      end else if (8'hed == _T_31[7:0]) begin
        image_2_237 <= io_pixelVal_in_2_5;
      end else if (8'hed == _T_28[7:0]) begin
        image_2_237 <= io_pixelVal_in_2_4;
      end else if (8'hed == _T_25[7:0]) begin
        image_2_237 <= io_pixelVal_in_2_3;
      end else if (8'hed == _T_22[7:0]) begin
        image_2_237 <= io_pixelVal_in_2_2;
      end else if (8'hed == _T_19[7:0]) begin
        image_2_237 <= io_pixelVal_in_2_1;
      end else if (8'hed == _T_15[7:0]) begin
        image_2_237 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_238 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hee == _T_34[7:0]) begin
        image_2_238 <= io_pixelVal_in_2_6;
      end else if (8'hee == _T_31[7:0]) begin
        image_2_238 <= io_pixelVal_in_2_5;
      end else if (8'hee == _T_28[7:0]) begin
        image_2_238 <= io_pixelVal_in_2_4;
      end else if (8'hee == _T_25[7:0]) begin
        image_2_238 <= io_pixelVal_in_2_3;
      end else if (8'hee == _T_22[7:0]) begin
        image_2_238 <= io_pixelVal_in_2_2;
      end else if (8'hee == _T_19[7:0]) begin
        image_2_238 <= io_pixelVal_in_2_1;
      end else if (8'hee == _T_15[7:0]) begin
        image_2_238 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_239 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hef == _T_34[7:0]) begin
        image_2_239 <= io_pixelVal_in_2_6;
      end else if (8'hef == _T_31[7:0]) begin
        image_2_239 <= io_pixelVal_in_2_5;
      end else if (8'hef == _T_28[7:0]) begin
        image_2_239 <= io_pixelVal_in_2_4;
      end else if (8'hef == _T_25[7:0]) begin
        image_2_239 <= io_pixelVal_in_2_3;
      end else if (8'hef == _T_22[7:0]) begin
        image_2_239 <= io_pixelVal_in_2_2;
      end else if (8'hef == _T_19[7:0]) begin
        image_2_239 <= io_pixelVal_in_2_1;
      end else if (8'hef == _T_15[7:0]) begin
        image_2_239 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_240 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf0 == _T_34[7:0]) begin
        image_2_240 <= io_pixelVal_in_2_6;
      end else if (8'hf0 == _T_31[7:0]) begin
        image_2_240 <= io_pixelVal_in_2_5;
      end else if (8'hf0 == _T_28[7:0]) begin
        image_2_240 <= io_pixelVal_in_2_4;
      end else if (8'hf0 == _T_25[7:0]) begin
        image_2_240 <= io_pixelVal_in_2_3;
      end else if (8'hf0 == _T_22[7:0]) begin
        image_2_240 <= io_pixelVal_in_2_2;
      end else if (8'hf0 == _T_19[7:0]) begin
        image_2_240 <= io_pixelVal_in_2_1;
      end else if (8'hf0 == _T_15[7:0]) begin
        image_2_240 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_241 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf1 == _T_34[7:0]) begin
        image_2_241 <= io_pixelVal_in_2_6;
      end else if (8'hf1 == _T_31[7:0]) begin
        image_2_241 <= io_pixelVal_in_2_5;
      end else if (8'hf1 == _T_28[7:0]) begin
        image_2_241 <= io_pixelVal_in_2_4;
      end else if (8'hf1 == _T_25[7:0]) begin
        image_2_241 <= io_pixelVal_in_2_3;
      end else if (8'hf1 == _T_22[7:0]) begin
        image_2_241 <= io_pixelVal_in_2_2;
      end else if (8'hf1 == _T_19[7:0]) begin
        image_2_241 <= io_pixelVal_in_2_1;
      end else if (8'hf1 == _T_15[7:0]) begin
        image_2_241 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_242 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf2 == _T_34[7:0]) begin
        image_2_242 <= io_pixelVal_in_2_6;
      end else if (8'hf2 == _T_31[7:0]) begin
        image_2_242 <= io_pixelVal_in_2_5;
      end else if (8'hf2 == _T_28[7:0]) begin
        image_2_242 <= io_pixelVal_in_2_4;
      end else if (8'hf2 == _T_25[7:0]) begin
        image_2_242 <= io_pixelVal_in_2_3;
      end else if (8'hf2 == _T_22[7:0]) begin
        image_2_242 <= io_pixelVal_in_2_2;
      end else if (8'hf2 == _T_19[7:0]) begin
        image_2_242 <= io_pixelVal_in_2_1;
      end else if (8'hf2 == _T_15[7:0]) begin
        image_2_242 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_243 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf3 == _T_34[7:0]) begin
        image_2_243 <= io_pixelVal_in_2_6;
      end else if (8'hf3 == _T_31[7:0]) begin
        image_2_243 <= io_pixelVal_in_2_5;
      end else if (8'hf3 == _T_28[7:0]) begin
        image_2_243 <= io_pixelVal_in_2_4;
      end else if (8'hf3 == _T_25[7:0]) begin
        image_2_243 <= io_pixelVal_in_2_3;
      end else if (8'hf3 == _T_22[7:0]) begin
        image_2_243 <= io_pixelVal_in_2_2;
      end else if (8'hf3 == _T_19[7:0]) begin
        image_2_243 <= io_pixelVal_in_2_1;
      end else if (8'hf3 == _T_15[7:0]) begin
        image_2_243 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_244 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf4 == _T_34[7:0]) begin
        image_2_244 <= io_pixelVal_in_2_6;
      end else if (8'hf4 == _T_31[7:0]) begin
        image_2_244 <= io_pixelVal_in_2_5;
      end else if (8'hf4 == _T_28[7:0]) begin
        image_2_244 <= io_pixelVal_in_2_4;
      end else if (8'hf4 == _T_25[7:0]) begin
        image_2_244 <= io_pixelVal_in_2_3;
      end else if (8'hf4 == _T_22[7:0]) begin
        image_2_244 <= io_pixelVal_in_2_2;
      end else if (8'hf4 == _T_19[7:0]) begin
        image_2_244 <= io_pixelVal_in_2_1;
      end else if (8'hf4 == _T_15[7:0]) begin
        image_2_244 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_245 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf5 == _T_34[7:0]) begin
        image_2_245 <= io_pixelVal_in_2_6;
      end else if (8'hf5 == _T_31[7:0]) begin
        image_2_245 <= io_pixelVal_in_2_5;
      end else if (8'hf5 == _T_28[7:0]) begin
        image_2_245 <= io_pixelVal_in_2_4;
      end else if (8'hf5 == _T_25[7:0]) begin
        image_2_245 <= io_pixelVal_in_2_3;
      end else if (8'hf5 == _T_22[7:0]) begin
        image_2_245 <= io_pixelVal_in_2_2;
      end else if (8'hf5 == _T_19[7:0]) begin
        image_2_245 <= io_pixelVal_in_2_1;
      end else if (8'hf5 == _T_15[7:0]) begin
        image_2_245 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_246 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf6 == _T_34[7:0]) begin
        image_2_246 <= io_pixelVal_in_2_6;
      end else if (8'hf6 == _T_31[7:0]) begin
        image_2_246 <= io_pixelVal_in_2_5;
      end else if (8'hf6 == _T_28[7:0]) begin
        image_2_246 <= io_pixelVal_in_2_4;
      end else if (8'hf6 == _T_25[7:0]) begin
        image_2_246 <= io_pixelVal_in_2_3;
      end else if (8'hf6 == _T_22[7:0]) begin
        image_2_246 <= io_pixelVal_in_2_2;
      end else if (8'hf6 == _T_19[7:0]) begin
        image_2_246 <= io_pixelVal_in_2_1;
      end else if (8'hf6 == _T_15[7:0]) begin
        image_2_246 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_247 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf7 == _T_34[7:0]) begin
        image_2_247 <= io_pixelVal_in_2_6;
      end else if (8'hf7 == _T_31[7:0]) begin
        image_2_247 <= io_pixelVal_in_2_5;
      end else if (8'hf7 == _T_28[7:0]) begin
        image_2_247 <= io_pixelVal_in_2_4;
      end else if (8'hf7 == _T_25[7:0]) begin
        image_2_247 <= io_pixelVal_in_2_3;
      end else if (8'hf7 == _T_22[7:0]) begin
        image_2_247 <= io_pixelVal_in_2_2;
      end else if (8'hf7 == _T_19[7:0]) begin
        image_2_247 <= io_pixelVal_in_2_1;
      end else if (8'hf7 == _T_15[7:0]) begin
        image_2_247 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_248 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf8 == _T_34[7:0]) begin
        image_2_248 <= io_pixelVal_in_2_6;
      end else if (8'hf8 == _T_31[7:0]) begin
        image_2_248 <= io_pixelVal_in_2_5;
      end else if (8'hf8 == _T_28[7:0]) begin
        image_2_248 <= io_pixelVal_in_2_4;
      end else if (8'hf8 == _T_25[7:0]) begin
        image_2_248 <= io_pixelVal_in_2_3;
      end else if (8'hf8 == _T_22[7:0]) begin
        image_2_248 <= io_pixelVal_in_2_2;
      end else if (8'hf8 == _T_19[7:0]) begin
        image_2_248 <= io_pixelVal_in_2_1;
      end else if (8'hf8 == _T_15[7:0]) begin
        image_2_248 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_249 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hf9 == _T_34[7:0]) begin
        image_2_249 <= io_pixelVal_in_2_6;
      end else if (8'hf9 == _T_31[7:0]) begin
        image_2_249 <= io_pixelVal_in_2_5;
      end else if (8'hf9 == _T_28[7:0]) begin
        image_2_249 <= io_pixelVal_in_2_4;
      end else if (8'hf9 == _T_25[7:0]) begin
        image_2_249 <= io_pixelVal_in_2_3;
      end else if (8'hf9 == _T_22[7:0]) begin
        image_2_249 <= io_pixelVal_in_2_2;
      end else if (8'hf9 == _T_19[7:0]) begin
        image_2_249 <= io_pixelVal_in_2_1;
      end else if (8'hf9 == _T_15[7:0]) begin
        image_2_249 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_250 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hfa == _T_34[7:0]) begin
        image_2_250 <= io_pixelVal_in_2_6;
      end else if (8'hfa == _T_31[7:0]) begin
        image_2_250 <= io_pixelVal_in_2_5;
      end else if (8'hfa == _T_28[7:0]) begin
        image_2_250 <= io_pixelVal_in_2_4;
      end else if (8'hfa == _T_25[7:0]) begin
        image_2_250 <= io_pixelVal_in_2_3;
      end else if (8'hfa == _T_22[7:0]) begin
        image_2_250 <= io_pixelVal_in_2_2;
      end else if (8'hfa == _T_19[7:0]) begin
        image_2_250 <= io_pixelVal_in_2_1;
      end else if (8'hfa == _T_15[7:0]) begin
        image_2_250 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_251 <= 4'h0;
    end else if (io_valid_in) begin
      if (8'hfb == _T_34[7:0]) begin
        image_2_251 <= io_pixelVal_in_2_6;
      end else if (8'hfb == _T_31[7:0]) begin
        image_2_251 <= io_pixelVal_in_2_5;
      end else if (8'hfb == _T_28[7:0]) begin
        image_2_251 <= io_pixelVal_in_2_4;
      end else if (8'hfb == _T_25[7:0]) begin
        image_2_251 <= io_pixelVal_in_2_3;
      end else if (8'hfb == _T_22[7:0]) begin
        image_2_251 <= io_pixelVal_in_2_2;
      end else if (8'hfb == _T_19[7:0]) begin
        image_2_251 <= io_pixelVal_in_2_1;
      end else if (8'hfb == _T_15[7:0]) begin
        image_2_251 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      pixelIndex <= 32'h0;
    end else if (io_valid_in) begin
      if (_T_81) begin
        pixelIndex <= 32'h0;
      end else begin
        pixelIndex <= _T_79;
      end
    end
  end
endmodule
module ImageProcessing(
  input         clock,
  input         reset,
  input  [5:0]  io_SPI_filterIndex,
  input         io_SPI_invert,
  input         io_SPI_distort,
  input  [10:0] io_rowIndex,
  input  [10:0] io_colIndex,
  output [3:0]  io_pixelVal_out_0,
  output [3:0]  io_pixelVal_out_1,
  output [3:0]  io_pixelVal_out_2
);
  wire  filter_clock; // @[ImageProcessing.scala 23:22]
  wire  filter_reset; // @[ImageProcessing.scala 23:22]
  wire [5:0] filter_io_SPI_filterIndex; // @[ImageProcessing.scala 23:22]
  wire  filter_io_SPI_invert; // @[ImageProcessing.scala 23:22]
  wire  filter_io_SPI_distort; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_0; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_1; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_2; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_3; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_4; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_5; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_6; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_0; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_1; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_2; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_3; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_4; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_5; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_6; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_0; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_1; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_2; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_3; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_4; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_5; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_6; // @[ImageProcessing.scala 23:22]
  wire  filter_io_valid_out; // @[ImageProcessing.scala 23:22]
  wire  videoBuffer_clock; // @[ImageProcessing.scala 24:27]
  wire  videoBuffer_reset; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_0; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_1; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_2; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_3; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_4; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_5; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_6; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_0; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_1; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_2; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_3; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_4; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_5; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_6; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_0; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_1; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_2; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_3; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_4; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_5; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_6; // @[ImageProcessing.scala 24:27]
  wire  videoBuffer_io_valid_in; // @[ImageProcessing.scala 24:27]
  wire [10:0] videoBuffer_io_rowIndex; // @[ImageProcessing.scala 24:27]
  wire [10:0] videoBuffer_io_colIndex; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_out_0; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_out_1; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_out_2; // @[ImageProcessing.scala 24:27]
  Filter filter ( // @[ImageProcessing.scala 23:22]
    .clock(filter_clock),
    .reset(filter_reset),
    .io_SPI_filterIndex(filter_io_SPI_filterIndex),
    .io_SPI_invert(filter_io_SPI_invert),
    .io_SPI_distort(filter_io_SPI_distort),
    .io_pixelVal_out_0_0(filter_io_pixelVal_out_0_0),
    .io_pixelVal_out_0_1(filter_io_pixelVal_out_0_1),
    .io_pixelVal_out_0_2(filter_io_pixelVal_out_0_2),
    .io_pixelVal_out_0_3(filter_io_pixelVal_out_0_3),
    .io_pixelVal_out_0_4(filter_io_pixelVal_out_0_4),
    .io_pixelVal_out_0_5(filter_io_pixelVal_out_0_5),
    .io_pixelVal_out_0_6(filter_io_pixelVal_out_0_6),
    .io_pixelVal_out_1_0(filter_io_pixelVal_out_1_0),
    .io_pixelVal_out_1_1(filter_io_pixelVal_out_1_1),
    .io_pixelVal_out_1_2(filter_io_pixelVal_out_1_2),
    .io_pixelVal_out_1_3(filter_io_pixelVal_out_1_3),
    .io_pixelVal_out_1_4(filter_io_pixelVal_out_1_4),
    .io_pixelVal_out_1_5(filter_io_pixelVal_out_1_5),
    .io_pixelVal_out_1_6(filter_io_pixelVal_out_1_6),
    .io_pixelVal_out_2_0(filter_io_pixelVal_out_2_0),
    .io_pixelVal_out_2_1(filter_io_pixelVal_out_2_1),
    .io_pixelVal_out_2_2(filter_io_pixelVal_out_2_2),
    .io_pixelVal_out_2_3(filter_io_pixelVal_out_2_3),
    .io_pixelVal_out_2_4(filter_io_pixelVal_out_2_4),
    .io_pixelVal_out_2_5(filter_io_pixelVal_out_2_5),
    .io_pixelVal_out_2_6(filter_io_pixelVal_out_2_6),
    .io_valid_out(filter_io_valid_out)
  );
  VideoBuffer videoBuffer ( // @[ImageProcessing.scala 24:27]
    .clock(videoBuffer_clock),
    .reset(videoBuffer_reset),
    .io_pixelVal_in_0_0(videoBuffer_io_pixelVal_in_0_0),
    .io_pixelVal_in_0_1(videoBuffer_io_pixelVal_in_0_1),
    .io_pixelVal_in_0_2(videoBuffer_io_pixelVal_in_0_2),
    .io_pixelVal_in_0_3(videoBuffer_io_pixelVal_in_0_3),
    .io_pixelVal_in_0_4(videoBuffer_io_pixelVal_in_0_4),
    .io_pixelVal_in_0_5(videoBuffer_io_pixelVal_in_0_5),
    .io_pixelVal_in_0_6(videoBuffer_io_pixelVal_in_0_6),
    .io_pixelVal_in_1_0(videoBuffer_io_pixelVal_in_1_0),
    .io_pixelVal_in_1_1(videoBuffer_io_pixelVal_in_1_1),
    .io_pixelVal_in_1_2(videoBuffer_io_pixelVal_in_1_2),
    .io_pixelVal_in_1_3(videoBuffer_io_pixelVal_in_1_3),
    .io_pixelVal_in_1_4(videoBuffer_io_pixelVal_in_1_4),
    .io_pixelVal_in_1_5(videoBuffer_io_pixelVal_in_1_5),
    .io_pixelVal_in_1_6(videoBuffer_io_pixelVal_in_1_6),
    .io_pixelVal_in_2_0(videoBuffer_io_pixelVal_in_2_0),
    .io_pixelVal_in_2_1(videoBuffer_io_pixelVal_in_2_1),
    .io_pixelVal_in_2_2(videoBuffer_io_pixelVal_in_2_2),
    .io_pixelVal_in_2_3(videoBuffer_io_pixelVal_in_2_3),
    .io_pixelVal_in_2_4(videoBuffer_io_pixelVal_in_2_4),
    .io_pixelVal_in_2_5(videoBuffer_io_pixelVal_in_2_5),
    .io_pixelVal_in_2_6(videoBuffer_io_pixelVal_in_2_6),
    .io_valid_in(videoBuffer_io_valid_in),
    .io_rowIndex(videoBuffer_io_rowIndex),
    .io_colIndex(videoBuffer_io_colIndex),
    .io_pixelVal_out_0(videoBuffer_io_pixelVal_out_0),
    .io_pixelVal_out_1(videoBuffer_io_pixelVal_out_1),
    .io_pixelVal_out_2(videoBuffer_io_pixelVal_out_2)
  );
  assign io_pixelVal_out_0 = videoBuffer_io_pixelVal_out_0; // @[ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25]
  assign io_pixelVal_out_1 = videoBuffer_io_pixelVal_out_1; // @[ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25]
  assign io_pixelVal_out_2 = videoBuffer_io_pixelVal_out_2; // @[ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25]
  assign filter_clock = clock;
  assign filter_reset = reset;
  assign filter_io_SPI_filterIndex = io_SPI_filterIndex; // @[ImageProcessing.scala 29:29]
  assign filter_io_SPI_invert = io_SPI_invert; // @[ImageProcessing.scala 30:29]
  assign filter_io_SPI_distort = io_SPI_distort; // @[ImageProcessing.scala 31:29]
  assign videoBuffer_clock = clock;
  assign videoBuffer_reset = reset;
  assign videoBuffer_io_pixelVal_in_0_0 = filter_io_pixelVal_out_0_0; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_1 = filter_io_pixelVal_out_0_1; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_2 = filter_io_pixelVal_out_0_2; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_3 = filter_io_pixelVal_out_0_3; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_4 = filter_io_pixelVal_out_0_4; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_5 = filter_io_pixelVal_out_0_5; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_6 = filter_io_pixelVal_out_0_6; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_0 = filter_io_pixelVal_out_1_0; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_1 = filter_io_pixelVal_out_1_1; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_2 = filter_io_pixelVal_out_1_2; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_3 = filter_io_pixelVal_out_1_3; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_4 = filter_io_pixelVal_out_1_4; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_5 = filter_io_pixelVal_out_1_5; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_6 = filter_io_pixelVal_out_1_6; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_0 = filter_io_pixelVal_out_2_0; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_1 = filter_io_pixelVal_out_2_1; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_2 = filter_io_pixelVal_out_2_2; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_3 = filter_io_pixelVal_out_2_3; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_4 = filter_io_pixelVal_out_2_4; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_5 = filter_io_pixelVal_out_2_5; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_6 = filter_io_pixelVal_out_2_6; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_valid_in = filter_io_valid_out; // @[ImageProcessing.scala 39:27]
  assign videoBuffer_io_rowIndex = io_rowIndex; // @[ImageProcessing.scala 26:27]
  assign videoBuffer_io_colIndex = io_colIndex; // @[ImageProcessing.scala 27:27]
endmodule
